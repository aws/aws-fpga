`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Zsg04eHsmrkwhG9zvpgQQjeSUORE/CUo9y+/mnGaFaA+nno9VQsbp4wCIDbHJIVGAAg68bwmoF52
cbITPRKrr5bS6AiVeu1l3p/StVKrPy8i/6BQBmKq9aK5gAP3SPmIzPivrcOM+tqC9v/5+rzMCWN9
JO7Q5PnUpd2e7W0VSbWz262oUmZMGjtAAH3WmTF5g+Z67qt3JzHMInfdtpkVcPcPQ5zsV8M1GuAi
InD+lN1vn0HDQL89+YNrSKko01Dz9LV77y25Hr2xwJcX2++xz9YDB3LcpPC7W4iyvrCH00bNMhGS
A8pftQ1UP5KqP9PVn4/51K+TKygJ6EPQ4HcVKw==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
EP3E7tBPo4ovxgYew4KGB2yhxyLbOg0kMRJ6EM4DWXsT8cCyafiZpR+pkpktccU0F32YjxILKghD
c4aMEdHdWxCfpuxQzBfvmVfHWJY/6ef/bX9LDGLo8O0BUEjVG0ai0aS7ydsi2IBEaQaga4esZQvw
YcY5v/AK25A4YXkVVJM=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
Pjq/f0nec7jI/jj2HUo1mZGaBuvb4B9BxB51fRlxPuE3WU0lFmWcLZRF+5ildKjWaWAOHmcd4X9p
Kf2PIua3+NpMMjPg1b5CQfQ/5Y/4PjOp21KPyI4/dR91G6tR6vsz6cXne7nIySH7c2GS7PM7RnCh
kjljIN0/68XwW3AAiq8=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2160)
`pragma protect data_block
eMDyyfThTI7SqCuKeLjpa/wDC0WMXwuT1Iwj5B5vIuNAAej9PKBqa1JavKctpuvU45Im+3m0/ek/
afTTjuJkgNfQBvf8X2R5NMLzqnWeXzip2WzvlEXHN5EE2+0wVeHKB85R/5YI/d7hKg8CwVHdos9L
3BJwcKq6qOc9wW1WTcBXASQ0nq6QUTRyEvfFxAs3F6ay22G1HVKfvP2CiZP9iaP35qKBBxgj2Jij
0ipdsFgPQuzEMdS7hJ52CvekFkNeIv7G7zhjGkJ83PIbPpjknpLZYJl/dk/DgBBIz+f6YscSKJFp
PqLrDtkMdrmKmCJVdmgZC9RbbujDa7MkGahogTAny9o7QJnWUaCVFl/CjMyYKSStw0sC6SkZXHMs
BR3GLqNsNuXItOc3cXL++jCtD7/U5UJQKLfCmLvPZK2x1T53gU+cf1reY1/+EujiBjYN7w/HpmhA
EH5xerC3e6hNvOuL3oJh3LMAEcfAMuD+0qF4bhN/VERmxuy9KWJz0rJDX0mEGdE8Jirlol7cR91z
+kspXS1FhlQVKvdOVilyqtaHPkkqlanX11IaNfcZYb1LN2kx8xFj9eYPeMi2/MZZDdaCPvaaxajY
dgSsQtl298wCJMPgLNys0wqTEABwXiZj7qTPFi1Ubwpm1INeolrZKx9h5vSpj4xYcrpyd4COS1dX
dGglk86+LsGVoQCO5+zSx/Lp5CI4wqCPhvmCNqrRxsmL5bTFXYEtIN9jUMLdB1ABrmyGZMg08htc
Qio7jHEKsfN1JDNOtxMEi1yIaT2UP5Noiau6qata0w3Rb0pLQdOMIBglVYxZV1y+3pOU/ayhlbgM
5ZvQhpb1xIR4eU2rlNNvh9K+Ag56RZDmf29SfCL5DXGt45yxWcnEK2taItzdA+9doHiyHpC6clSH
BHoBDSA9TiV+7CnL3/EZH1xN2C/wUIjZkF/EVxXXI8r8xD1qDTt2HvmIVlycLig/4sJHKDBuAjQR
riS9VxvbJWYlssJgTcO8p4NP6h7YW3euudLNWg5pYSxezEpXboq1jiZQm427OKs7oay7Uzt3cxKc
seboYyj91uhlRsiblzvb6tGnkq+r5GOPQSYcGK1bROuYZiL4pNJ4ljU5N1sRi2a19zIuFy+R8JAO
IIZLhJzQ5RG1GJXTUPzlte7FwyhKCP+7NrbAbVlgFiWjM5Xa/jccyGKhpbwNeIJQZGojW7LPLAb3
oVoLNXDLJRJic0yDATWSM/vqJPrF31mCpdFioCPOtr0jzGRGTcNX859NQzgvpvbtMWNqtVRz3G/H
trWpHCu58dOiq//hOxVuBtWYsB3Sbt/w+ydhD7oooA3KbnfiR02ExKSV6T94Y81xdy4jSyBnTCdE
KuBhGhiPjmdED6fu13hxgef/I+0LpJo/yckOqqsO1A3R4eOoxpF16TGZfaxfE+cAGeQi7AmdTsBv
NjU51SHGTOsZXmPRYszqh0d71zpCidA/urQ76/F4lGDSPRqmLlq0C7qaDY6u6BA8suJXunY5SW18
clN+LRtEPNrytgnacagEe5p76qxLfMxbYpK6f9/xWaC+OvY/ik9+r8Eh4qIoADd3Qr9ElOMGdG2Q
Bd3wwTVdpbOeFMNLUtCcx5/zZSxrEhLFLiHZcO7TOnuLIZNF9T6R7ei/liY3vTICEzyWnfz91+L6
DkX+ZtMFrBYdF1YCfcrIpjgAR6H6R04FzLZazARuDAFFdEQ3ghhXQ7xvAC/ZWdL3Nyw+xlzk9/x+
VB1xTerMuOkIRtF2fXaU0u/VVmVOGVfUX69Ap8yB9b8rj4XDcHJuGKdnQ97o3mkU3PmXI5bZkhIn
vDdM2d3DNYSJfjrBjvmBppxRXJsb12YcUywFQDU9ZhG0TmASEp4G1CVsQsX+WdIVFBCW8eCmsQRT
VXUPRqdpxKdXfcyS1w9D83jusVWQJOtQu10CoFVwJvvJsqck/Tp5aUrpqRnWoYjS/TXSh2j21+K+
C297+XkL5/XHXuxD2cZE0IfV+k2boLT/VHIBy7Zwulb1iijMyCYB+CRZC17YeYBRP61BwL/lSp1r
aflXpU/gd/BxW9bdpH3aPSC+hdqhX0Kp7PdUu7kmT+q/MXlSqBqfZEcu6HQecYVUx/fGx8ICqjhR
+bvFBh8S6MX/zV7j1av0OVjRFjPEWLQkxUn1+jH2yjUbH+mfim0+RguKN3Kw68MuEsLokcF/bp/j
SKn4ohLRErnTzAiGtd4sVH1xdFu3EDp6Nb/Z/+rshXZ5jf/La3V5XgLHJ55ZyMYuegZCmCC5wGdo
S9w4t+n09vNPyEjacGN7INlIQ0utnFZ1KW7fZ01iOSqvTHB/ws9THe7q+T9RZ+PTKM7VJaAQ1Hkd
ZXP7cs7FyI9muKV3xrXIYwgmCYLM/GUVbMrD+P8VxtD+pUn2C/f1A0H4LkUhUCygDUu4YBfnn1vY
MJRBSg49hxo9i78bVhTAveSskOKSfXjO4vhlMdE09TOPheWG870t42sUWDQhMCjpI/bbfWYI4KGm
Vw+Ie50SoVNvPw4gpY40FZCjpnhgvxHdsxdXWcBKyRMnu95f3bk3DLI6WCvfuUCljAhEksI0/UR2
LnJOhLxwAHbGya3imPqwXf4WYsnf0WL6Ogo9e0m3YKm1NdRdMwKl5z/disisqCp9uN8tdHcn4jan
9jtlFBmMyan/Q9ORNinXXxZUnxvY2JEjIFqAk/nosGVIpwCtAdA42KuFze94GAQAzTEDGvjSLWVN
oO4kiHs444LpUopMuC+DXgmCLDwsTVECyZKxgPffFn7mcxvQMkjEVjQgb0T+hR1jk09ySw+Oj5+4
Wdt/EBvU2Mlpi/cPgB2sIrPzceM08JKQfHeLSMpdatk+bx24NFxouklYb1F3Pj0X8p2v
`pragma protect end_protected
