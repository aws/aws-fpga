`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
nXTphsbaHLT3vjv1XQxUZ0Ifl+FAGceIo1BmNg8/DSRn3UpsF63ewaQBDwhlbVwhr0jmXDbNcs/u
YkOJeVe2UQZ+s97R8troomPkMDu4WnToiHy3Vbui4RMBnkG5BKy8eWruoTb/mMLfshrdK4hpkegX
pq8PhUQ+CQAverO/tO8KFhwu/A/KjW8PRy710md43+KI+2DoKTcXx6FF9o/H/6ZXlpsF1V9s2UmP
BhkpNNt390ooVHPjNjwZ4pDnQsI7GTOsfe6TID2pjLehGK9tQuvpS9TBOteau2X6bmfxz0wI/nv3
GOm+6sf+mpnnaO+MN+3v8xHWaORzdTj8ZfboLw==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
moXH1PeIV0A51aUWU9q+cEHxr/sYgU7/g7ODnTsVDpND/SUVF9tlZRxgPM1Jdq4wzmoWmHNx5r/h
qePRIao4cbwYKQFRSm5WoFCHguUazwqYverLwciFP+gkngVMuwBMaHhZxtVdlBnzT2H5H9FDqUOs
9tVMHxatv8ERpO5EVfo=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
XjzD3FQCvyS5P1ZkhPdFo93ukMpy8GaUJtTwl2JK+vUdDA8Ab1kbvNe//djVwmulpHvWbQv5fxbm
JOwoGeDeI+evIyIjPdumlwR5MgOWaTuzMzIqNKE6rfQ5kL48iLJXvnINbXPbJ+KgehVo1Bg9sqSJ
HWpI+EdbjhPmkZXeOfM=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3056)
`pragma protect data_block
dSqopU9NdDDcsU1p4GfkFdGJP4O1Czqbb26B7uxio3BP6X7jlNfYB8AcHFyz1DP7ip4kZzmxkW3Q
u3OdMNV7razIVIvExpvs7n8UKA0TaBU0ZtMXtG+1hEkuCGScRPCNZlKJhrnHnyxQZwvbpT+FoQKt
hRSWhy8oC2/1djBqkgcfUF7Kz+L5hIkR/Pil2oqfF7uog0D8sTQU1o5Xgf0vU8w4jPkKvGEL33Ut
9IZgFkOIH0E1XN+73p2fWs9ID2axBfsS6LlQZcSJEx8KjlP/tsmJD2Q5TynmDYFN08CRH49EiFPq
7U49H1WZde2RnF7E0mh1m97pwuoy1Ce9jPpacyeBQnnSYKHTNbL0yD3UlfjQduTBFqgq82gxjDIB
Muz+aYiu51wYA9YY0ZrAqD+HWJ8z9aPV3h8QO2jiKm030oSsesArnmccPwD5vxE04j6YI7KsbZnK
Q3SbhlvvXGWmxjABZVT5+Jy1lRzVCS9MyiROLxAyaO9tjsLCSorVJtbm/1vcHBWdo/eQFg/eobN6
6/afMDmKSwTEaMi0ze6xSkhd2z6B7ImEu8YTrVKQC9uFSWt4kXuIu7D6BOGNhIpCkz+qDbrDfdgu
mM2kaaVudAx21nMJgBXvvNh3S1YDrExucCdQoPTe0ZCcskzeMwXEIJoo37Fo6QNkxfAaIrmQ4Jm5
pobsBLZa+30OdQwiRI479wza/pTeJpTMT28JwWCi9rwbvw86zie+v8gEkXceRKYb0Wj9Dmc6mFxv
DeH0DsTE+7iqPagt6DUDN5m+jK1zlgyDdRgPqjWymmr/PNuQrwb50o5ZHeKi4s9sPJtBr5XEdU/h
j5+VIrjxXU90u1qTR2qRY7cQphN9wTR/CeUpkqwWb7wyVjR1eN0G2hqB6UM37bppzxX6sf7hsSyl
AWsLFfrrV2AT48S117EllpUIsJ0wVKsU6MFHnJUwapqnz1Z8kjT81yMy2HVOMDbf4gQMFt90gJfK
XvtJqNmxhPFzBteG0B0E9gcKHcywANby8z5//NWzihoNpPhXWopcPJ32U+Ek9F16c/XM23ccVNj1
V9sfxAGfIvdKv56t68WcYOKJyFyOUwzoN6OhP1oJyQU6xmUP4xOOWv288OvAAqG5E5Pi7DyIUxr6
I5me29Oi5kztrkANaU+WDKYF9vwbHFMb//f9vgnkARhSf70qjg9WhYU1eT0u0sKTI6/S6SnGKJxZ
nX+oY6oqZn6BmsKznEJw/HsSN5y1UP0Sh1V1yVitDx4e19LdKjeKf9AgDyJ5M4e31QbfxMgLWv63
6avGe4oWiglF8dnsJLi8SVENW9ofh3eakl21qEso7lADeBq9kNB8Q7R9zyGPCmxSFIk28H5EBJio
ApipBfxL8kbHdzi/ECPvjsmLdEIjgASXEs4O3ulHcT8TeFj2VlvC8t8siwRs8cakJ46R8c/l0IPi
Ob4gXISlnTTMA3x/9Cm/EsWBELCEQuZ/XDeNVob8btF40wc5XFxDK5r3X7HaTjovf0fnupViNHFD
W+2IpmI2yGxR97Lm/Q/RGec3lNlSegFEkSEuflA6lYCBG0v1m7QGTuJGoTHPu32rEUfRC0NgT1WA
pDdq8OTWAMLu60oJke7dOUOVb04Acg8YM09e429BaGrl7ERoq2UkJ8QlOIVvYcbYFicWlLaK7rm+
1septRa2paqQA+vfy+J2nXVN+NfKRoYxuRIme6WXtde7jMBFptugd/EruvRkAxMd2V2iH/bxU4gQ
PpRMeYqsJAFjXVejWi1Uku6tvV4QhCYSxPS92TN3UJ9SFpTEyA0LKqjHr24oUYgN8t3V/DBKExoM
fyE7JQurVVs3hchzrOU8NYmjmXRM09vYQJgD17FGz7Rjd6TDRYPzjqAPRByFIu4IaQmBIYTu5lrc
kGYKMBEVkRcTmwZZ9jy3G6OgZ++bD0G/OqtDpOoDOy81ch6daLaSgMnBIChowTzslZ3nVDquIot9
1jYO+zUtkB3PqliRT3jmsorW0b7hY5n+f8s6E/aw3MHjKPuGoggdFfjGHU9QS1jC37DySa0fVof0
V7HmbQCHMAv8EjZqzzJZGa+U4bQlraq8V11CC4E8B6gm8zQRvlVuJYd3qmGVcmcQpSxeVIHPMmQK
xWWzpfEM9sZVZ1ftq3bW5OhDtbI5efuz7jxH+j5B8K/INj+jQ0Nm47HJhdtsqUC78O6webxljm7V
zHkDppN39wfxIycLrQ4Z6EwZKEMv4tJO0mIR0hRMdKd4neinSU9jvwT5JII5I86qpetbsx7ryFJB
pN8tUQvVHRhYe+r/3cb5XFGc2MI0QC1UyOHFMnPYR1Goc09r45PNbo4NXNkj0vJjPGuAoSz15icg
Y2oo/9RyzEl5CmiewDZOHH3WH/vNTEehiWj9qG54JQ6XpaHv+YAn02pE1skYpEv2cOI1y2JLV+Ew
XQMnULYiMdv+FoMXqjWnYhN7IuvPwCJW6bh/0vl2V6SHUlJ7e7AhyNKLMrv/xcvB6HB057GJrllh
dGDrmEid1DsfM5TunYOiJ8EaO2RXik9hiTaEy0zrkNRCPhwDaMB9e1OV+nNc6bK/ysZD6l2x7uQ0
PAVw7SMo0MliqubOZ9PVKxCjO2mwPOls7DEujNp3bEL5eeO2c/tlbfqb8kkhnYe62LgTUgOoWVRI
N/4+R9XhzPyyRFHrJxicV0v6epd5BJ+3H9AjA9XsLIh/FK5MCmdiAmUdFSO3GO0g4PrA8cnB/yXr
aioc8RxEs6OMlQk52zr7Pq/ZoCoXwhFUS2iJIXbD5wwczW4oAp3iVV+r6f4aLt0824CECqUHNd3e
Cg9HY62CT6KCtNvYttCgQEHhIfXEQFEK4hAVkGm7CRHTKVW2qHidUroI0cV5NS7xzAgzcJk6Yibb
x+DEG5hl9ojcGxKml13UYkXglB24LZ2u/py6SVeWOehrqnYYPaK9Y9/ZH6qHiywpiWtizodgTFja
u8IYV+gzep55bPVDcj9UunNVyedUWIeESLrqMpyHDI3WcvdeKHCEHNV+ZRfjLX/oNCoHtO9U3RC7
IT4zFhgfaht3oWa16RyJueKoQ65Jpr4ZbQbIz4pTt+wuyvWrR9skhmNsWHiss2xDuLpnTOVARs0l
GWaYLs+cmoFy3CsB4lOOaQExJCayI66AQgMaNenzfskY5fazXdekIATwv6n13Dzrea4LHcRZ4BzE
cYGMBoR00kbZoYVzJ3YYPDkTJIGNi+qUiaQLSCh2pkUkFXdHLJnhC6jgms70FCiifTCdwv5OGbG9
T84bPADNiVD8VMZIA9hZDQ61K6RVlMf3HycKj3BV1ChJjuQ2hdk3Xym4hzlEcqNZq8oyiMRbTSRZ
JIUCShKiUEVPckncl4n4f8Zr0P6bFuGG/HS+yHjrrxG71Nv39D/zm0VMXNCv6nOOzoqsCkMih2Jj
hNxN/fv0SdZFjyxNZqU9RondE9ozT9cEhLDcmndPL9aIm4zShT7W41uNDhW5dPXTsEkrnYR+eUwB
NTfU3gx3gXOuGoZftMUyhAmlibOIJVV1wYv2Kexu1L9Qve7sBrIIOKTgKoqL6izEPBQ2fs3kX/7l
NRKSWJqxeWCt9CEcGyyEOtI5usALQ+PnsTQ/x3BPZ6tBQIIZqA2c4aHCpaHE8Cod7hXSJSY6pAKy
8rNsoJv4moniLpB6SyGBx2/6zDlrEW6008lgUVEnW98YUmMuSHkiS6fZ1l01MwMlD12p7N1WUf+H
LAshvYpP/3oRJQPzXiDN1go1N9xf0FSxjYury3t3x1xso3mokDfyiXCHF34bopYGP7YnfryO+XKg
jMqtWRfpT50WNmRt2BDY8VI52SpxJzT1n8nB7z4O800fcJPo1EqHRfZukIRW0FkEnlJxqwg7x9aU
sewYmFDY8xyeYO5jWiFGUY61ri6Gl7TndHOUk1NKNHyItfz3KOhWQzmCTUNfKJ70W5NkYZbyDDOW
JJvgGf3lpUKZkC9EkLEQy96ds7lB+J/5BFB6d8Y8sD9X4A+Eec/2PJyPE7BaQC195dTSSoM4CKof
1ndmrs+zNNF2S26s+vmSw0+uYCe0ibk+Joo370CnsMfsEFc=
`pragma protect end_protected
