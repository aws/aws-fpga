// Amazon FPGA Hardware Development Kit
//
// Copyright 2016 Amazon.com, Inc. or its affiliates. All Rights Reserved.
//
// Licensed under the Amazon Software License (the "License"). You may not use
// this file except in compliance with the License. A copy of the License is
// located at
//
//    http://aws.amazon.com/asl/
//
// or in the "license" file accompanying this file. This file is distributed on
// an "AS IS" BASIS, WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, express or
// implied. See the License for the specific language governing permissions and
// limitations under the License.

// SHA: bddf8457046b3a64e63d28d7e334020b6f1d09ee
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
rJ0c6LBVhJ+AJJ7HccLBgTlffpb6jJPb7887SuP2KIVHLpATOUYOmJQ/Mb6Vvgw2o6lAP5xMUxWE
CbqKAe4vVVhd6etoG022MtX+uHcMwS77uaQODDYE+MDqtfS3HHqyVLekalu5ExjcnlDVZ8lqC9JC
BDr3OItAf+H9SNxTiC5BH1L7mwnnV12HVfWPoIPaYhrHRnrtQIu3hEh/EUw4StT5i8buhWRzLxgV
Y047fvOZ4vvD+CwhybFB99mx2H1WD2Wp7xlLfG6cMx1J0851zjY7Qb898z+GIp26c/+B/En3iSAu
1t9ZBrdL/9jfr78LNtjJ83dfkp7EVr3WbUZc6g==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
eOH+uFgVxGzzjHMABF+P6OdJ42M9yVIU80xR++BJGVXQLLZmS8/u458ZftvDm/oY0ALFh8zqfsbV
j143/ghaBiVa0NcX7f2aqtCaraznLHg21i9Yejnk+zyGBRLQcU4wT7KmXltGuHQWgEbOWqoO+I5S
RT97pWbKQFk7GDSKhUg=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
XVVo2RWK84SRsMk8WdLZztGrmVeHTbpo/J9eJb00cuQW/x9EFVQatfWiRXPdZIxJmRuV5WCQnb38
jPkNgf9Wqg4F5+ncuIkA/1yfOOYEXAAECSToxApo011KSrl3Yk0DGeCncFkV8/qYVXw/w+KwvcHK
boU+jLCgJt0rFmcD/H4=

`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
d+ScrqijwH9M4fdYj0c0O8Oui0ZZzjjAlKkExw6AvTEkZuLcnKnoR8UMK2q84Rce/6uBgZtAs3IO
3+/bEniOSA==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3136)
`pragma protect data_block
H6TJs59wtckL8dRHSi7zZg1IExnc+CUfBxiTe+dLcexfccABAdqgqb8U3cR0e8GaU40j4zwzhGOF
BmeLWmBnmNw4XwYJwQ/bcTkfvAFl/kgtDLCyMfHdDfuJFGOY2W3xAm/4X6OCFr3Ti+s2gWCQtnhi
78A/wJshwfDFy3uJgiaXFWIPecwJ7sfYmv8WoLFut7m5ZeRHONlSHpwW51F8dfBmEymJH+MXLwyH
VIOoYueSOqW0x2STH5eDnmuJpoBP7Pvm/euit8sxHg0QoF6oyxDEcUmm7vGp200p5sr+pILZbbQ0
6rvQ+QEfwgCHgLslpocfkEC+iAdcTL6HCtNc5ujTDz7yUkmR3ZyNeujvGwNvbL0BVR2h6AtMa3YU
Miyg3PAlrOffzRl4RPxSnNMZ6ByFQl9rwmPRGZ+B7QB0bSUWxQRWBMiteT/RkSxjzPeyMDPf9Zva
+Q43fW/Uos9p4ehszkJSc9mfHzeAWOVt6flIYdQ0QcEb0u/to7ZR0b6W6oKxjg5V4ctduMySb51Q
1f5HvtXULFkP4gxQzRGRLDwVvTRVQfl/3uG9iwqI6qSIKj54vHTpxXL1AtAWnFG+Dayk209MfZN8
Rdp6swBHgzWYA9UE03YD3RL1kjLy4uNhzIvz+vgG0QLn92H/FbxK1xcF46t3QsBnlxNpHqf8laqN
R/4PpC8OIfiowa/yLZBjDt4+BZXqs8ZYbRgxnei3nS9ksWR+4OFshcf38JB34zzcgXXILyBzvuEv
9+xzRtMLdcnc5Lpsvb35IEvjQYZs0l+XLrngp6PyQhRzA7+N+rHRo2Hrg5Z1VaBPt80b6bTh0CeN
UnS24lsie6AD/v3RRbp1R4t9hj0UPziVG35+/xjlL9xGKHWJIvVTwg2hDvSEzegt+1cZ38CXONKj
ZRt7hEpt6XB1mLoHrftsd6HZqg9k2KXaf2xH/SVuOknfQPIM8jaB5uLyrvzmN1Fk/mqbUlwCSZXI
6pYKIcjs/dcdmmawNm/88LlMuAebNAPMdlsab+rscoEzvWDzP1t06TWF/pGAdxdLDqxcibqnRGWs
O1nXxI889qXhTd74w4lyf3epRzJ+vokxycWwRYdQnwtPRFDV9SpYlLIJtllnUBsvm5IDGaTkX/t5
N8FtZWbRzSY/ps7moZGXizL8AQcHGfffUjw3iIvZSMNoPS7ZozIP2UD4UvCviDbCgAmPZloJMP9H
l59x8vc14W7oF23F3rR58lMnWZYg0mQyeBLbh5Qb1Mcw0VZ+f6pqbeZdUMDrqi9vODRsPW4db4Cs
5zxYw0xULID7f/sP1XKPT+0tD7bv5oA0ZYH6ZBqgG0/pkBMaFai57EqHztu9RekLYad1DhRUVMtx
ZNI+JtlY17bSIyrFqf2F6fi46Yia+Fy9eDkRosfW1b6pXQdfbnilEehy6QgnKFW0zQw28WbII8vB
UztSoZP0MqsbUPPqJ34IvPs74X8SYGSL9yLppnCK7dER70JPv6s+NJ0WsAAnJpUSHSUDpB5CgZAT
PGL4B949g+8xG+d5D48y4Q0vJAJNKbqxN1jz3jfclqjvwRCDx8M+PiOTN1IQCfRuf1g6oalPQKRS
C0svf8a/qgKycAVqQEMJqQ5bnUXk7aJAaIZQXaxjR6U7NImzK5xTLTimj3rJZbkTg6tToJadYOH8
Jb/C6+6k+L2DQuGyM2awO6ZFWKWL7bV1qqREFoRHiA/RTak0syoCGXAnozurFswrKbfFgWfQnwK4
4pgIxp4KrxUb8L1akSZjqGp8c3e6HV1sJmop67+tuHKuX+QWWeygJjvLunMZ9R5B+pq03mxX2VBB
Lg3U9B+Q+AsvlfYBdNKIEx1yaMGu1G8kB08L+bwSYgbchvHqOhjrEugcR+iaGHgOYZoqq7x+nm4l
qzXu/i831oEhng+jVZtrWy5FzrZpfrP+OQXj98xEhTh1pNZu2tuIa8gn7go1uJtTKX5pKfea8CUd
5gBVsyOaYdLtQ8K1LfK45R7nsODsbwlqkp0DBIBISSJ+jKLDXAQhItErDqCN54xf0KF0VNvsG+Jb
/qVzVXHmtFVC4vrEZ9jw820O9qgnI9nlvlpXC8OV/YwP1Cqf/rx2aQPUlTHDZHkS1f9J+/xw6PPV
zuSjzVOOrUN3uSGMEH+PBqPSDrKME3u6YeGwhvSaqLAq+Pja8We/krqfpud+D0808uzrHXjqd69g
unZQ/qGw9U+ZXGLiOk/tqKIIimXPgTX6wEGps0E3UTxbjEPowRH1OsKI5yMXoZe63mFADcoez4vI
zURZ3Lol9b+RYBUgrR5ns5pwTh1VnMu+DI1eoJAXbHZgY+31nsEjr4sZiHX8vZ+HwYwOAB4gBojj
DEFTJcRPS2x54UkgNFcv77qL6UQk/7b2YKmC9bmZWgzElnUS9pjZOQcZa31y/MseOrbh8CCkZ+Xo
0yH1sXIXdQSf3U5yEDWBJaHHfRss/hibDJiQOXE0708HHNtsK9djTRmCJC5cQELqjmFqoaYdfaPC
drUaHfiTlFWcgGmQD37EIvITufnAfu1ExhnMCuaR/rDvu2QYHxVF5mGxxtnfg/YpIxIs2u7eQ5sz
cwqO37n31NT2ydepejZlgwJjbUM6LSxvWdFsgmsw4/Qe5u5IWT9zRrgTe08iFtf1jL1NTpDr9ZLZ
POesO70shM9g7ZLAM6wdxwHvKzjnDFj8471RcGR1LgBHddsj/QEyd9tYuyfNpCICNz1cmyvIFa3t
iPT4NjDHU6mihh6eoYz3nYnx6HU5e+OWA3v5Zj69PDp2lM5z1HkrxhGIBHU7uxj3FjXI+YhRvZax
AYKbRPqjOqP6p/hG8tgLTK6bPm3f2ky2TJHGyyOIjsmry0rHh2QLe2Kpi8E8GIUywu1jYfmeh5Hu
esjEx4sZ8Smb3n2dWE6TuE7YO2uy3WVVd1rV5LjlAGr+35CQIIBYNz0qNgaQQT99Pz15eCmZQcE5
VgDYC8az/ny67+6x6QVZo3faC/teVwGZaxeqnnlrOXMK/owSs7+kZ8CsHGouxsn21Bam66oixqb4
DzsGieSRcsNaCeDfe0ZBCBlHYnpLYuGau07hadKVhyaJvBH/9fpJtWE0uik6CFfCvk6mcoCAWtdL
fjXSDXQ0rS5piI3psRIeMyRKENXYs5Qu9Z9zAfwo2SJN7jh4v7rVQg0zkwNzWBsYuqeWNQzL7TIK
RWtZb8YXJ+qvyKtPBhcUdWKdTShWneKlJPH6F1Fg+JwVR164/XpBuAbS+JIYf0iXW5UGgwZTd8qT
TKJP4Wr46CX+6REhBAVNbU73/9vHDThaY+edRjE04kZL/95XkCHzg884sLr4TbS3ily9CeCDyHqa
MjdSdLHJ2/JFbIA6IjN2axCxKkNfxDkZ9D7z6Tnsx06AzS4LNxeqM9zNvWuU07U1alNMIdhWuB4W
fbdrYJX+Az6hHbEQV+KkNEODuRoYt8Qjdy9AYZSgzX30CZIUE1mVsPeiUVwlpHmpL3BiS6667R2K
IdZ5B7avrxzsgBHWLB6BAr4OSXTbgEEhXpbb5qLTdqQ4YmDXh2Piz35oOxKpUgifMtB9ui+kGsL0
Bmi9LBHLUpCaVylWRdG2ndU7mqdWg2AKFyAflCPT7POzdYfCjcL3khhgKBtHs0L56PMyRYY1X3M2
TOWKlrTHwq8v0kGKtVr41SyxFGklQjEXHP2rEFUkdP+YJ2dejeGHYuoxmyupO4Guc9ZDghKkSZVV
uUkj5LqOuhSrZ5JbFff4o2zsKSFV0bjOgYWdNByROtevNoXR0oJmqHCdsxYAs7mI12J0A6eG9WJH
eC1CiemtVtdFYJxZHYqmIdPH28kx3Sp2zuASst780kQVPa+siibFfAa4dWFNCAdsCE9bV4s88ZsZ
pqnLsj5ErTQmyKj2h3ggU7OKUAEpYUj5qfCu2HkAR5Rfp7ELuDqVCzGVE3+Bs3/mcX4aLac+EaWQ
/sRD2m0phD1UzvFYBsmKHShdzIkv/VTMn635NmYPwVYoPRAVoS8LB1g7CHLBd1u9qQoX9WSwn3yl
M5BnrAENpxg91cA5jK8du2wIsZc9YwLg1n49VDmA8F/Pz8Koi6OjBDWF7Aoed3TCg5o2lh9s4G2B
YtzENjn/j5g94dMtuwLZfuys0acnUnOhAQJQPPVWe8jjeny3BKva3gKAN4RGFxbXKkrj0kEfddP3
Gw==
`pragma protect end_protected
