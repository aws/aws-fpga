// Amazon FPGA Hardware Development Kit
//
// Copyright 2016 Amazon.com, Inc. or its affiliates. All Rights Reserved.
//
// Licensed under the Amazon Software License (the "License"). You may not use
// this file except in compliance with the License. A copy of the License is
// located at
//
// http://aws.amazon.com/asl/
//
// or in the "license" file accompanying this file. This file is distributed on
// an "AS IS" BASIS, WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, express or
// implied. See the License for the specific language governing permissions and
// limitations under the License.


`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
EHLq/BFuT/D47Wdttwfql23h3EUI0dQK1d1Pw5yx9FfFDFbo9Wa1ocUgixra+aNICZFmZECRlZCB
7MofS89c02Ci/uXlbebwvaEWH95ZYCrAB5lkS6rGE/tU3IYnRyBSk5iBvobyevOCamNQ1wrDgZx4
7KSd8nehtEDbOsljAg00que5+GCc5kv6WkHdi2ZCJAgtFj5ZUa/ECo+nxn/gJj2qgF4DvnD+ZBTD
KIMxof1rPu0kdjHXc+v60jliZDOmDLeFJybU+ub7wB6nL59pqxhWhAn54H2w8jLigXISTwRPwxTX
T03CQqkix9NIhWSm1vte76ijOCLtUFnw79IT/w==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
ddYYxOrqkNeyTmkWK6fdt7aNngfChDGdCiQ0Se02L+vJu8+ooT5VhMe7uCHFTZP+GRySntOowP2u
po2MReHtv1U6TkUXd6oZhYKilRK9oVXvikezuYbaQZ+3I8b0WT7TiNTmfz6KTovJfulxHzd2A50e
RBSl0fGJmVaTy4ZgM5o=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
kU569mtvJIff0Cdy0ubv7R8Ev7el9mUu/BDn5i6CguaPENaFGp/yPgJbwbtRPDP/zoPsNRcCAOw/
g5JycUonGa1afe5/DtJHOtqTMYyGujGlXMfx2i8gwny44aDHZU6jO0plGk3WbrhgoPmCetXZuVPy
m2fVrKRTRJTDbjIbd7M=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3696)
`pragma protect data_block
c2eGtsg9O340CVf5E8RH035v/1mD1ycVGMS0KJ4gMufLgtdL/cPZ0wbqBfKao25yTjMfbB+8OyAo
40Tb6vyfAMDt5CM2QBQkE7jN07GRkThqdY98hCRaMDUc+CnCh2lMdrwKVCfWojxdOvudOxD9IDrH
HbQRtRfgUdA9GV0z8ignm7I3SzaseTZmZPbjIWavftfo6AL+cdtdJQ0JWbX7GpZFycD45guUwk42
kWs5VERjvsecJsoDzjXy1gLrvliPDK3wuuTBiejt281/NNljVH8yc5GfzzsY1W33kAnSs+MUHnZr
8PMzEwUZjMSUHGm2HZE2EM6Rkjwvn2dx1LfAW+8LjQ5DoCq2yNpU8A6ZZfTomrfSLTeEfNb2uHwo
mBxt+sktooBAa+UHN3mFLBP3ubfxpTZ89wx5n8P5yVzhiuB8dcvMJ1TerxwBIRZAs2YeCOJHYGst
oPDace3Yf01uu+eoyRqtShYCwq2EicRfTcOUJpuyC5eTkWmw73yue/E37Zz82+D1aP9AIj2L7a5j
rDanHp9L4W8PqgFX0bpANfTfFRvOpRSyVST3cETt6nflwvzy/yNBLO06dFiKF0yMWz8r+WeeAmTY
qn1m9FDiVTyAhc1kd1tusJ4QzoD8mx5G4Pln3M6j5CGgBHtMf7EvCSsJSVWA6cMu66ExKHnF62GM
Ehv0SBtHVucwBlKqI2oIKz2fDPlRmHgsMujzrw3FuURxXQBsApn5JVK1xZ5XC7xZB6gnWl5pXtDT
M/FAjwqORJq5YOA+qtQ3pGHPTdteVIuu/6PuVoMZBCEO7kWF33W4iDWq1vADOqGVT4z+jIjP4wE8
4bf0zqoJ8Y8koML6gveqt3xz2E2MLAyRX3szhmcJa47sqIek3ZAgoxTE6bTQnczJpnYIullxGkHh
ZXlVaWSVgIEPwwbc14TlgAkwqdvS3VkHaFYWakCfU59QO7Pj9lBUMg6k4nCbrS4PI78jga7LNPJJ
gS5+idIeks2jQIN4r8gnNpROCprd1gOWfWyfv5uTg+sId54b3xV8JsTbM+f1Fc1d+p50thOL0unA
Aw/Mvv3Iukiz80H3DR/zkOxxPzXFZPzyt+mGGjUttFuO44VYJOSl811P0BmGku7FKjWPSQqdOIhn
JgakzLWxNxv/YOAGzhqzdo6Do9iTqUV8Opl/KPmlI1hgrRtoERzmMABmfloORo+XxAazJJpwcxib
oFnXpJoV+DRiXAT5S59q2hi+MsSGlsYVpvUtyJiALE9UtaBdxz3Xk60hw6zXWjAmVDIZY24NBXFh
AVuftE9sb4ik17ZRRFKS3OAJIOxIAq/4dzNhmm0XJFQbczYFOxTSfyR520DHdlvCppW8gWrmfgtQ
kpey1I6g+F3G16MNRX0bIFNHNNy10zT14GG2b98yF+MiyYDzM6Na0t6J/jVtCCBjL9lsZQCoH+3I
yVRKisxVWoimYleGPmyCuFgzCEG+m83UPOJZz1Lo9jaeuf9+XkjIUg4Zd05p+NK5xCJN5zBUrQpK
c7kSb/BrcBLm+uTwbJJuJaz+36Ujfb8A4vbmZAyknafIeeW6tRdiKDusM0U0lsbMzpsqNQk5xvsn
VKqGRD2rviXpSanVOVH0nCkFFMv32rM+AlfiLTODxubXxlWSW5nvp0+A0ZztnKiVhR7Ynu8kpf4X
BDH0gg/GlsJjCnMMdUaUA/2XN3V3RZVYn/QrSX0ynO5gJb6qapiA6vn67RmI3WBUUG7gFJyVBmA7
oMMsaEPYwlKoUB14ZBYeOl7FFvqJg/OgNzZ8K6SWun1JGeiwAn3hUzpDFUsmLg+xF+fu6/ittGAb
dH3FMubs1fohtc5WOKsd0lMQteCqj9FMFLHZnSGLf4di5EKFGk41wWyPPlUgTlS8Y2oL8kDxonbe
Scy2S8625anW1WElGcgVWVo2L58BI+aS+dnUyawlWnwzrdZq2XhLyq08aVK6sf5wRTL1cAjgBbEE
zAG21TwboZEskj3NT8JdaTTj/v9HDfxcuNiLu6hs3DRqqO3eDQ1mwf8RqSrEZdZCblf3oYsjnTGe
6DnJlgtsaa2iRMHSw6uZMtZwkOTX4vvYFnh4uTVyUiyJfxRmULiOjlcW1MHgSjk1bUmGUhzjuhoB
xcTh6w4J79GWUYx9wUFb6gOR30q/spnDlVfpK+GYUrVJBO3oUOjkRepdQ4rvtu6QrbsgjbOoCRKH
sg+bL0JuLyvb10Jq0gqemh+BtkZ2PxmqsQ41GgOGMgQuLgMjsU1v3gDQQv0sSxxFx8Zx8Qd6wFJA
b2kMY1RerzPXD2L5EdnES9YEoKuzVkuCJu4F+JPHxOy58fHiGhtRAFR4mFxg3ufu0RIUZkT1DiHi
4uAE6+Pna6OC21H5VQdhCE4prL4arX/4u4gDOSwYUNvT5Zs3SyusUgww6fj54oq0iBKNP9RthNRp
9W/XW78HQb0R8A2HFqvG0m834g6E8F5zyY5WV91zFVU0iQXCxXaZVqKrbndUFTzICdfV2xuPkO/i
V36Rgyt/bu2uJc/47NdfSYi1LuAT8Q3pjsE59N+Pg69mdF9MKs3FF+cXc8U5OGE/cYstKpec+8Ef
1VCQzdgtGg0ENWMZEsEutMxd1vU3anFOHotrKlUUGhE1lLw+AUzVAgNJlRXNBs07C1/n7/EtFIpc
LQjHE1Pz3BgeNNKlS0nmP1y/RjxehThv+jSgz8yeuvVrVI6YH7jmMETaMk9Bg+TRD7mw8sqVAyZ2
kG5juq3VKlf6Jsg4eZzDLYzKv5G1SvGefyd/wt2/Ub3xGG7ZFQJIxkQWFQxbKp4DiLOSxLw7Clrp
ON0WPBz0fNaL00mOKTgczV5T1R8MfXU2/C8pBEhdZlW0u55gEzNXT4H2SuosISOkgVHl0RGuC5R0
bALtsCplnM0M+98dURrtbKxZ5cvsWdE+PsF/AFk8Fk8YUfGBaEucoWaRjBug/mGW65WqLv0uI+RH
ZBuWMUPVlYSyEIfDbKIIXVIPQrcvVGF7YqdhJY6+QwtiW1McQW4cBhcBmzwQVzVavQDl4LpIl0IP
osq/SJn5A7Yq6X9UcHw7JX5PAH+ljyPVZAAHo8tMQk9IdSnpWt2BWHaOCrKL7raLbrYQ+wlxp4aG
njtXFdepgvT7+WiCBJ+dpNneEadHpF73is6gxR+O0Z/5XOn6XW4xkk2VJZ8QE7G05wfrVo4FBwUu
Ykxf/dFav32X3N+dEb26csMEQTkzo4w+nEyalNLo6S9plF9Z4V88G6lW/WznDMb2lAREYjIVPRte
uC2cMBnuF9PQ8Mc6HETF9GzcPSQ2FnBHi6djAMj1JcHMEA8agqIYgloma5FxLSdPBMVEKMBUma2v
aIjZnLjU4k2Fcz5n6rSojFheu6Y5mhoDlCjtGnb2k4wKKIvK4rMZS+eS25HFUh0XwiD4HjSsDAgW
mOO0wUGKuGBt1Mxgz17I3jZJogQOxkS/2FF+isq9r5RA/xfJ8A6IQ3JDLHYrBRbLZiWDdijKS0Yj
lNggKjslIDQKP49L2nDjXMEV09DPYtV3y8sX6eVKu8eLp/LB+GdF4cucAQ0vQ4a4nxtsyS20ZmZ0
L7HjEnGA8gzOsYYsuEYLUVyb90s8yWeSlMqI9b5jO2SvkSry5FrjIP1NbwlsOtodqUtl90ozkp+u
bq8DkUCw/s4dwgrSG2qtclP8otlEUxa0u6NGE3nKtJopIiyJL7O5a+i1OJeisMT2LI24qyO6chbl
SaQcYFqsYcgNCkjPesNpWkVXINXpy1HRUl6O8N/LZUyLKvoe8VbKnunKVbFXLh+toBTawXwTYrQA
NINBmQBNWTqjIKGFgQ7+PNmhrmAwzyJdMBQFh8l5xqmmkBT2Vz4BNJawJ7Kh0itjwX5ciKpqm+/s
aHIG38Rs2oyeX9m+cP5p1c2wGRobwBoNmvMxStncICIzlr5hclVOnpeJXMHCIRl6Ct+aHGjgGI9d
JChMQ5hA52rF1xnWNMI8e4WMvngclkT9jHzruLNn4PikE4WsFHpy79jCImYFn3Wv9u9Rlfz4LWr+
P5wzmPeXxw49cfRR3Hky8PYzbKgyugtQNgcqtaorvMOtckf957cstxItEeQ5A2FaVYWIskVYOkzu
AbZ1h7dNy8s0diDySENynd6y39yZBU/MYcu+Q4jj0tifjmSkulTn9LZS/CNxyhJU90er0XTCxUK5
+NE5IhTlkbUKEtLE4DEJ1umeHI9kjrLw/BMTH84FK53DnPC5eNBGSzAKDNTCDxigMJa6HfA0eSB7
MT3A3KuL0FL+NXOzw2EiRion1dfwqzdCW2OLCl06Mq2ZvMcX2RA199tgazlZ8CWhLBwove4yUxP5
I4rOJ8S56DzMc6kTG78wADVAEjP6Whfrd437kHVlKD0GZBz3UxOtMfRIrAw2ZX382VDaozt+MXfY
zY/sbnjeeP5iTgEst3XxfK4kTCT9kgFcWqMgjM+wuGUt+4eBzATX7IDHRcSwq3K/2KYty6U6udPR
9tp9ZvD6FDY/Ww3oq1nISXO2Led7kpIo1Bnm/uRsqr8KSrE7gMItptCD7evpDE6mfRiFygI2vgC1
tqbxTzhPWTzkndAgW/e0nXA6QEh2/GmR427NItMhwvMB5AbI7r25URupXk3VL52uPN+L2msoIhfE
xaFbjHY6IOfTWIeU3YJB7j1cOyktTDWQbCmryeA+MWGn8OU7tRNGWlTh//HJEopfzeA7bnxYqgVS
gczUKvi0WvTJEvSjXjHZdkoiDaytGTr45Ch9DHfq/cfqz5OmcbC+r2UyecUZRjcF5rGM1f0B9+xh
OFQORjPyxmtU7rOW8L9ccgUmxzLprqFMGkqAlhN6UwJt61QpdyGo+1Alv/cPCO1C5q/OTbVji1+E
fWSDOCNM6QmniTtluIrJSIRdGb/arpe3yaeIRq31Zj3nHLOMJzY06LnbroDvsTnP
`pragma protect end_protected
