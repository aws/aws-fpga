`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
KozAwAUN8Y1BAEleBFIqlAFGYmHGzOQQOLa1wEGMALoo3LQfSf3HI+kYH6K0DLmOLMexr/0jI1c0
RjHVOmdMmVJQXO6y7+2mBmsKoCXS/0hnNayg1K8QBPa1r/dNbwyjNA8sC85+ZOG3t0jVaEeoocuF
T8uTIEZfsqOpmOM6m0SCciWSljskqhgHiqDPPotFJ6AToYZAf9JG8Wj/Y1eyN+HtWPCfONV9ni/H
Hj7R3cYAJqwno5FrzJJ4GLUsnKXTzB8Bc2cQDYyuANNlDBuNJ4VPzQFiWBJ9BYe9mHey2GKj+YjK
MgIRWgGJ4qOHtgSw46y5t+AzkEhBzDZqtab6FA==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
UBrDSrgifvmpQRCQnPGW6Iz7NiOBRE0/TiEfc9H9jITR1z7wiwo6BQHwMheU8/RkR9FDhY7YkHgu
G5v1jiUjIe9/qCCtkABIkk0sV4EkaTIxaHE3J882JdPm58VkHTOPFs4wmVw0S1uMQiq2M+ad4zNZ
2wimbmmPV8Mr2YD0gNg=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
Wog99WPzsxCwKH2Mwe5Vqk5iCMnV4HoK2dnxk7LShzzmR4Y7qIJ6HCFM9cSKy+Eju49SwjnoHI/f
Ov48Zo6PGxr1N3P8kO9J35J5uXn2hzyeVLHC4GJRe3LYb8JWE7k20csAd/zjZnhnY7+OukGf0Kyv
laFel2rSDaPOnuIr+KM=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 45184)
`pragma protect data_block
pl+ZgnQUhhDpT7Pk7zqOnfXtnoxJQuk0is3N9PlyUAQrDmRxiId+byzdyLGJpQ4qjq8JLQEZm7P1
yR4EepKrcBOQukp46P/xMuJq/I2Tjrs4R1u49pBFVuLXb7t1LyHwKhYcFUfr3GiGaGxmpF4GQUSS
NQf1/+0VTEi5WiQuiRaRYQVx9XfOhnE7aLMkN8v2OBgVtFkAt3fPz8OWQd8NNUiGzaXaRfca6E/9
yy0tJAG/ARmOLV/sjMYo3Ay3u9TsL4xvwXOmn+qNQhd6hruNayTcINtAW0lZqjgkPiMX0/ibyzJU
q2sgM0roDraHIp5k8hGGMLFXPIUyN1Dx+0ZBAaUNUjZinfVhyegWk01RTPyKvJ5m0lJfKyA1SoeQ
pZW52GNO8RyiQMclUghh8FxDPVF8q8Q84B3wxVBxNtACWzP3vmRVAscPui9mMRfxijua7wojtwGy
t7M8U/QHo4i8F0BkbIOcu/AFLd4B50BaBk1luZB5dmc2NV8f6u521d+wRg4ZoEE9N7COXWgq0oKg
ThtOxihZcqEWsPzROeKbFFxOThJMoO8z/LtZ3L3YXpHUyPZgcPrquNmZQaL9Qstry/T7oscKfpfz
GQTqzD/dfSKyKEl3sc97I60i8vgK4R2/10x8eHOvQLt27q7XnOLrJFPlw7zJnBqS1gNDTUm/n0Gu
zxd1m7TxpEdUDb3RP4wT/WlpLRet3m5tmOaW6OAeGv/w6EgK+Kbz+8ufOoeCYVPxYPrDvEuuZOk+
rxG3DKu8K/E5/Sg/6dlnQQJtXC3CV82/p3cThrmzeGj/adp42810CGRHWEiyDyZG1T06xMHgeFiL
ZvQGXYmFtWcatP0xekXqDzF2b0RFKlsPhM/4C0Wo8ZWjBSWGsPzEeDs3020QQL+azidQQuyC4mQh
5MFkhWKvy+TrKs1x/GRyGwEiwS0YlUICZnjTz/zSBvM6vuKZNQTstree3lYiGGvKmPh4YNmK3S/g
PexGLZqSPX/ulXbGpQ7iJzsfYlMwlPj59BvcSygE6GaF2k5RFSbUM7rWwbj23ASwjopOwDulY8hr
VWXwjG6+7X8nrqaAE2WzAihoBcX9jR+cxbRoAxzayK3jRXdG7BBCw6ZiSIKbD+HbYD/FyDkzadiV
0tf3oWF/3eZyCQ3jOKESFd+Y3LH2XO37NkJrp5x74DNrT4yr3aFrAzOexkBKFC+mv1iiOZyCNGFE
kwDJa31iWMvcb6WH1qVBihqXFamdULtPvEggPVCAMGx0AIOL1z6JnBAO3u6bV3o2Z4RhKbRpCDyt
gvN9zkxfg+2srU0Jd4pFGMnsTC0nXEKo5Ss4LX+tZVFCT+UTNO5lMQbPQSbRLdOCHxvzudZdBe/g
r0aL+9RJZEAm+1rIqxwD3KTGkhoTtX06qr/CSgwFNQbADOkk0LN7OtCtXiFbVO41i4MjWcr8ep60
NrD+8CK/UUbcQl4TgC2HwE9Ig1vhjEQIE9nfqIfGgIMV2lwlBYucIAofT8r7l2ZWT7QgnGkdPmmS
vVJPuJVGNj7vSfG3vdEgxQKUKa8qBjKjqHWZBqAMqKXrm/RTW8NuGB/OGVCW0KrHBQw5SICjfuBd
z+QfjXfn3HlbVkYNY7YxywqnD6FnhKAwsH3nCWgMQVg7p3MwJeqkX4wJis/+osEakXe+dwoh61r0
p3kqsojQ+XkhFZ7wchc0b55uJYbvzR+gX6kzT4mw2bT+M/MmkwF9ccK3hbwWpRBI5kYttQ9Ze64Q
bo2gJ7V8NMbTolhJr0wcRIRn6u0yUiOCHcOmwTNZqbkRpbPoOmrpiSRmd3sCPmtFm+O/VbPwJrny
x5ehLJ76fnwDsl+pXZVDev1ZOfKnVfcp29OQYQcoq/PyjoB7CLgT7vmUHPA89O6ccBZ5eNki14bM
DSILpce1iq8GOYIbLPPyk036lBhDlomRfHVMe697Skt+GkJYx40fYbaA4ug26Tzgb/hsGazTgg0H
TRGrQKpw3PN8M/mbRrolsqcu39IlAyJwPvDeK6it+XZM/RoLDHfsF9swb9c3v26/eEryIZ+XKO61
lmBqGxOcFXQKHs99RZY+ga+9DGk8q+sM29M7wbPiz21iLHs2HWsbPesA8GwzF17S8IX1BTBhTfeq
58bSLEJtRKBhzM9ZO57TkyfQacmRKBgvECErgHLnkT264uxzju4bEkMG4W2081Mj8RG9jqe4ZwDn
Uv+f7uvyIXS0L19079Vtf6SJwru+ZKJVdxwLJrBc45Io29YSERpat0BxoZCcG43S/1iBpvR5JS2k
9jbGxpO9pjWYs19bv9e24XPO3VEv9jq2RxNVcm4CAQPESV0apBwMLF9vn1VFf0rLCan5w8RjaOXr
t+y5odzpfvn4UndUPQI+EA9+c3gnM2j/dnP5nBJz1LMnstO44Rly0nd+4VJogznrCoTRm+4mtJvL
ZHTBD+XP5m5YeDqtyu8H6bUuPT51F/hG7fzG0CAhGi2osF1JiDpYLcBUHTUbODXd5ZJvXmYVcdQb
A2vss3U628XtIsPWpzGHTcFy3QbQK1eabaEVWRJdOAJKA7V06yfnNHHHJRNHVXMS+RuiqCyIYIqr
LQpkjAt17xBkH3SVe77hSHHyZ4UIPDDVKGrn68iC0yaIajOiBYURKzjt+VNgxKKqDYESrYEFaZPQ
7jNNH4C2Tw/quIqcwHhPD452jYZanL3dkySelHdaW4qGUBMjeoTxRzoak6ltggNxjSKOCz1vRNT1
vd+qKuKuuKUnGw/esBTagQLsJzLo30qpjyfiQx3hKQfec2fQbQRn0Aue87gePUwiaZ5tRy88AQbu
WkWoMK6ZKc9VF5uB6zCU8kLApkcId8D5T/o/Y5DCE6/pBCCvGTdXBrmc6edUaeWxAo0xtp/2yZ+s
l/KVo0z9nM23Y/W1CvpEbUqIUsZujqufgN9aPHygMcxylZ4QMfZd+Bgiej1AaAkYI0bKhGyVOIGw
Rn8SYG2zU1ZEAEMkiaRsakyHccUOzkF+g8BLnSwEdXJfE92fx78ZtT1JRIqHe3reQpxEfbNqi6EI
3pItUOmKWApq7mFbA1tqsN7L5cSShw/8i9QSGZtdjo3XWijudHV5YqbLW43NYTQhHo9AOwfZyI5h
fRoASlgCMANJ9PRqWbeX52G/A91aLLhZthF5GjwZNkZ4Ob5+qsY2Mj+IBEdOUDU1WKt4qYIl+l3f
jRV8sst6m4RTGLAnBdTzomGM1VYu0iS15/Au2J0Ba1fboNm3t7dGpd0r+j/Xv4K/6ZPSGFKiQsD2
O6NrkR+d/z1ZlA5LEmSItWcmNBHA8wFv7vmCWZpntlnQdLxoF2vPBJjwQvFE6ZTrx16tDOKJrxXf
XO/2XhDwTaZtBo2OLPAm3skLivO4b5IdkuyNBA91c19kfpCblNyAXf5l1UvcdzGvYuEdOkFtJZDV
o9udTuKMEGa4d7ZR3OQyC9urttVK2+nDt5geEN7VFAE+RKje2fDTh+hC9hkvFPyRyKukR364zcCr
h7pc4n8h14sgebxixL3IMfHSjyp2lmgJpH1t1phSGI4wUUv6lwjzq1MnrlFyBl0twmGPoQLJ8qFN
IuOKatLyq08pPzhCpPsnuH9nIL3WHDpYd4xl744MCr4N8FM0qNIPmhiRM94JQJ1D6W4t55NCVTsU
4y84mJ/ZIrMpUR3j1lAX9V3VPqB/honSm+FBkq7dUpj0j648IfBR2DRj8YNoXhGzo+sNcku4fj5Y
Ts2OWTM70YD78Pg1RpdNkUbEjlchzWhifS3v9vgVQpOSKYh1m0zLL62614n8i42Q5Y5k62CAQWJg
l6EVO5im5hme/TpX1FHoMt1o+M8HKwIJAQ+Hys30PdD81omTQy06KxdyUOGZ9V1ZLDLa3Qb8VSXw
rJMLzxTe8KF4DCNdVYg7nsKXw2Tys0lm+iYuHcRGWRrmak4C89FSJCpNGAvviBqTWX/VkFVG9Os9
THI/ZBJ1VxEDLzWUQFHXu4e+WXIlEOKtX7gx2nEZwdQVEjZ2mzLY4qN3scyKIUPhxAKnuVvgWjVO
gJyVCouSwUC08tr9GC8LvvLX9HRkjiPCvdkQfdMMrw+N85tVfoQFOJ97Dtc+FykoJjDAKEWs/N09
QiZBVzhvNiL46jln7lq9Oea4lLXimg9efl4nWtMQ2Ow0AJtj7dt0Jqkj1hmac7BE6G4vC62x2ZWc
BhYS6euk6OmLYDYkjz819a2EcqH+Reo2f2GrN/H39aiwPkP7RBH0xCjhQ0HAGeVHxSkiKMmaRybg
XB031YV/ltq+BP/uWLs/xHII4lzO2o3uxbpTLJVDoMOC5CLC1mwpdanZwwWE3UPkKQSpxXWS9r0f
GfdCixZVHlTBcEeJ8+QMP3AQww6cnNaXUVpVt/xhDzVuCVOTGYrF1d/JnuHbltViuZIUKxsv1ckG
ry2ByBC34mJW1os7RKsTyjvvS84vQAjpMiExes4yuUtynotxE+/m41Y/NM7xbH8Kk71xVUTT2ZBn
eajY9JNEBTJtkV8X7ZzgZw4Dz5xHrNbS8hhNxzkxBVyWrAHMzT7lUWeU6mc+2Wjzu6RVKx2Dyvp2
Edk1LMOOj1FUzowiOtndkiK9Zg9kT+8QGLKWrDFR1Oq0/PrTZzbNUeeVtwfgzX1jvouMeGCcMuHk
74MVD/WTQpxAj3jsJd2wE6DaHZeMW/8/Ho+Z1ZwLRCcGqynfLdZuEH8R0uFMU04TuVQRz3eXiEiY
JKXH8Dvf0oRj2AZjulhSmq/hCXdHY1TbQ/rDSyvI+1rR7U8t4BAk5H6/D2zoNz3rKnX0g+nrKG5H
cz4BgVSjDyvJMEtd1wfcJNnUsxgXDRZXbZH3tHQrcfuFta93bdKzwNLmI4YpQObyqJjJ0OrhR99a
L/yxWn+nYOTb9EnqXmj9d0aI7aM3aFHAhDK3VzGvs/IAkOHsaQusY0PMAWSjb+l0ptd/O9C56Jrd
D/K7YMHkLdlgoJ9WOdAXbdbKioK794MZsP64w3nH1K1T/qqXoud14zko+4WAKnywrPsInJ2NDmTI
EqcwSFgmeCwmQuAIpCDvak1INyM6QTbm/yIPRds0fT+SHuvpSDlhr1RFCTiAdBcJfit4V2SiAYtQ
dbKG80SVxytHd1CLQHiSCDkB9/pRchx4o63fdc7rWSo6yvRv8VUlX/xhNsbi9XNFLIf1Z52oNLDX
aSfArcHlTJX/iWKyGiVnHZemQh0s9IyHri3fttPmr2JKpMXdcQL+RnBDHxFcdRK1fwnnsTBjeYrv
MNXHWRb8E6S9udzsDToIikxRNw7RM81QB6Nt5KKkekxOroROipV62y81JQhD4e9DueZwkV1mb/AP
qaHu0HB2eEd2vSxUvD/zIp8JD5oeSgpigaUaizRtT8hlh9viB54IBWgMUZ2CXr4F0a/t+SJHnruS
HXuMFmstUMccSTlyfWqdinTGu9bCR9NXsOGeatI3XTQ8VsyCvsiPLmcWbIyFltYEAaARZcUKzPO0
aYq1lX/R08SkodgpMtr9z7anbrGTnnvJssRsZx5UCPSUupUA6lBXwYHy3LInyjlUDNIu9XiuqKtV
8nFpmnsgdd3RP+jUF6LtPcBtljCP4YdfzVcTC58jGBPADRVePWcD2eybKzXT01uUcORUj92uGxRx
1rAvmwic1tl5s5NjcPeC9yezNicK2wClWQk48gOpMOBozWRB6/B9APUegtEvMva0Qqce2eV/MV45
xtu8ygW5Ea1Nt5f+01nBxNVQP7FeZ1gCDyyObfvmfbTMKKmeoV8efYkKy7jYuOxpJ1PSDXwmyvmq
KW/9+IrkxNgU9JjInVzUMcCcJJ5n7lYS/va2a7e532pNqB135zHdBkoszM/34YB090u0WeE/T/2N
Z8ty0IXqrxnxxdX1w4OAKctxCpfH6eWY2IbGSEi7hWwOmLWX7K9Y8TrjTIY7hSEFcDJj8IrYYmO8
A+tbNaY/q7LM6N9IntzoVtJ0EA/KRefjohxQRFzTNAVe8yaDST4LThyIjzXzFrYu8ZdxFT3vD+EG
7WMH3lmMnHvtVAjWw+Junevte7pmLNGK9dMzKG4AWAm+VpEfjjsFXe7I3PiVq6yxUrEQ3J2UXtEi
LAKKmE3kAYP8CgxCzmBIPZYPJ+J4R9u+conFld7wY7DAxumO3SEDudfMkV29IX80SmFykS0bmfsN
3tIBNdZ3KYC1zV/MNOeZ9pMaVGDlz4WQHxLekkgfi6XdEKLgeAYzoRaO9RWuEme6/sneAVOEmm9h
ROqFx1zS4QliJ94peM+mpsDk5sL6tBMNv/Kg3dtF5b/D2wGgdpf9M9W4UI/GV/GSRbAZRgRrASf4
PUYhsFvW0NAQlXzTSq7pVQIfXrQH/mpJ9sOzpZdBz2awBYY3G5ABibJ6Xojski7JjJGBa7Z+qY0x
yvDrefdgkeIksNxQ5V41gPCvJsR6+WMZkVcmXSO5lAenn8mmvD/9qWNVDjAk8O8dCXqoAJVmb+2o
8AiGF0b6yrlbjiUUtoe4h8K9qGl3ba1V4YqRwkGC5rUn62j4AUkI8OlJkvgklADO6PsjnPBALuJM
ceYS3m3jKnihSFEc4FAAZXZZ2z64nwX+0RFxBItWIG+bIyQb1+wvxsiLP6Vq6ihU12mqZMFG6RrZ
WZyMk9y2bemE3yJrp0ZTATx84wxuuqvz2BuWVyGN+mQa/1C3TP+fRCKNVgczbbgfFvnlVxj82CPs
Z2j/qKe/FgnEPcoHONRa9+bdl8RLu94AcyXzuQbsS6q3zE4LARzRluHa/v+2V1yFQ1VgULh8DH+L
EO7NrSRoqVCjR8yqCiW/58k9YsX9gyhimVDPiWr6AmPTI28nPKgiK42gkDbEEp5Ljj/xZvF4afk2
o924kTxxvpsvZDZBnGrie3vmoMJyLMMPIpXOQ/MuM4bIzW9v1AKQEfw/epD1/EhO+wbvU0kozI/1
XaQGRk1zkWbG5JYYycYzdemGOC8IVfgtc1p+kpLu6PJB3FuLvGCvXwD7st7PKPyGbMnv3CnZFQ0s
7T4dMcRYKVqoc3InMI9HHLkxB/zIMuZfP+eh0HHk6ueKowu/lgOIyvl/KHFd+k7kRIW8IAQq7NRa
1QaNuNW7Ams22qxgh7BiLCRlyqGI0PLqm1tO/wh4cF8hqwZE3F446Zkx1tJ+WKT27FlCs1Fq3VDV
TeqNaHSZzlMl2cgHUVv/i4NYXSXx+ONRwNWOtFdNAQqyiceWCApVxt9gQbW6JLlMkpjm0a9TGJN5
9044ml/oc+7NW5upkOgLgjIv8OxRNnWK+4U75d6yM2DU0IkdsyEYDz5FtDdDd8eB5J2FR3O/ihWF
Kb6uXH/NN167wL47ebBUhdUvXQ+seTjGstg6o7vCiBSUwpwZ9OjtKoujQ58A/cygNf4F43zJGTLs
Den1GRmJ4s1wvPIV2O5nCUTtASteiIqKmrpjDqfzJbea8Xc8Iw1WVVOg1npogx/RVA6D2apC/BTv
G824uMM41H+oFBOWj+pKV1b5dCRgZ4Uodw3ilZvgsl4j8xRsp/JuxcvZZuh6zlz7+k678cQE6IoT
6qNG6rwGKOsO1Hne7rXrfI5KYXZcXoy/XtvdRka1cECfo3l/1ljO9rgHwJEcJv7pu1Ud5Z1BECtB
JEP/DFTh6GN4WnUd7r9L5R493PC1knftCPch6KKD5bFifitmUfEfPAUmq4gmpUkYXzZ8Ozx8/Wlu
tb/O6D89AqqglXQLtktxBcDj9jMSF/B31ekis8ce6L+zZ9JzL/+NEI/drEMH/+58yJTJOI49krJL
BmuqBzQmmt4pTbT4ojLWwDIk7Xlbm1HT7GGyVC0pHW47S2fh1tdjtCQdHYEjy5ciBtZVcHjc9ANU
l8nzzyUYwryplQsFEUYA6LSxqvjJ4/Jcx7fF1KPNpKeC0u3Gitk8WkyOTz8zyiV/b1tiM2gnQann
TEVwcOEkSWT7eZnpewUOyZdJg3bi0itvqrHTnffrwydhLp4AZv/hrYNiTfEcO2ATMKfPbUG/E/U1
5fnSFSKrU8AMma2tuKcTyIQ6lSFrGpTB7lob8GRmypkQYk05onVocZy6JpD8bi0hGyzFOmbDg8Gp
mAvrqHKVoan/vDCq5EyZrJ+EhMsBsZq0J6mkVWiqLp+WHOJWTE7TVyJMYJ5fcTVi5FUgtuKaODqo
29ky/fgENOmgWNXiEkIlH4pPeKWnFpDKSK4j8KQFzc+PO1p9Tj2FYNsL8Gq7tOV/Dz6Wms9P7/Y7
uButy/B6GOGiw8W+WUm5NTrL5NrpYg+uMqI0kb+qZQV+LFOlLLGjJgB3pxgyATc2QpB8jGtz25xW
ICRoXxuWPQ+Lp1jYwsl5dgdhOmsDWHCxxCZA5lgGOn6ta0Xdz4DLCy1qviY0C8YBoyJAHVb9UCAk
HG7F+vZXHumVsA8yFLxUi/qJhEm8PPxcB4DnXXSOeBL78jG9aqRdM9harP/DuTGgSTd5rlNl2zfP
CHnuWVWpjf54M2oXs6OFHGbUx7JC0MSV4+e8PNGaXv1D04orIlv3UBfnyyATIxyRD6tdOVd22Tq2
vcRwy+Jr95xwkLC2oP3eca1dNlKcz7+0rI+bxkj3rxv4n8yhL95G3BfD4u4aF3yCntmohTpKuCT2
bPwl9WAP2UHJ0qki0z/FMj7fXC9G77Jq8eDJX0kgK3Meat+Xd040m/5HFU0Gn2jw/P+lNQB4JLGM
tJvbWc0h1x8tHbks6ols7klbhqstTR0+klIXdhSrYn+OikFI0v5TCTmdXn9fHz0MPbm7zdff91UG
jSd7iiE73GnQSTKV6/lIL7Km95PkhNoH1CPTsEpvD3DuG6PtppXi93myeyKZzZKKdtMydJTY8fXR
i+6MkHr09GOa/oJdizCTQiCS+YWQNEKhaX8ywjRpCQpmTmzCU1GRn28noKM+9XemLlu1qCDJXh+v
fjch2DdTsunu9miknmn1yiHs17hKQfWHcY/KYvSub1QcRFJ9bf2cE+eFDmym7Dp0YudaEbgYenQ4
UBPAlFd++MrZZ6N0ItOWwaHKmfyjkIo+op2VJlJe6SOLZwtz7161hLKsFdps80lwOfB/Z77oGOmG
pH3VER5TeHD1TL2L4XiEz170WjYjoUTnYas7BBRiw/INDNIogb5FlUsNQhe9epBXhbJ6ZW4LLtnz
N9+Pl/K91tocSjMBLjN7cJyPP3mRP7G7s7Iz7My8vuRcbaF8EmvZdjVxyOQwKK0FPCSTw9GS/VFr
O45jslqgH0DldnBqQckMpHHg+Pdnswrc5HTIOs4r5c7moRDirJF8fZ7As+0Hhsvp2hQh9jQ/vVdu
WpVmwnVlzZghMenb8FAIGT5+Ag8H93VlI5s+m349Gad28OC3lF9WbIDPOC3+fSca/LDBRrnjUO+W
Wse1a5NKQzi2ZvRV2xeO4GeKGATaWQ1Gd2NF7J9sWpzeDcCFw3o0xIoR0jCRXbP0Ll2e1mjvRihC
UoNYik07en+KK6ron+J4uOnqFriQbPwcLH8i94Y6lynea+sFBzPI0LEZsFMfRXDjUOWk0JsIxLSA
z+BfvE1P6LWZv48G7YsH/HHXRxjsp1ShxkyxlqNpqyjDKFqJL0lilh6FStDFYes7DmO1UZRdPnSi
iz2n/VBodrDC2XDsovCY6iJzseWRRvG6+hsg8hQin0V+viWviQU5hcRAmVs79+nUGyjwNoq+TDMC
WIwAtpOTuQ0O5yLoJb5L8fPLnhU1Ib+qvjcJXTPGipX3DX6PGM/aUhod1InNyRGU7Tgg/ZNAASHg
yO9EZfMC5k52qe1TKoZ4gDRQvGkLuSVwv8oClVbqZPPR2FW0yzgOi6SEZp09nA8nQksq8yR8JAn/
8iLvsJWvY3HEqrYO7V3BiCixy/3CmCy+GmvTPz4HeNf3oPjZbpO/lX2v851jmiOOkUe/G3dksHx8
jkutmAp9dVXxRqqjXZUvA9L6JF8DZtrHgGvKpkzidz/EBzE8+xRZIbREJ1DtIABPt+JqaktPbGtL
i4tcH5Yfofv7oGtI2c2V6Ue+PEYwxITaD/wsKicxkj2z+TEiD6ynXSnEJwO2fKFu5JxFytI339df
BnFhMS+XYv30D5pQ3yUE80mOmg9yaXjHIk4Lepu/l4nRIQIoi20QFLzyckhrfnYWX3XBXdUxF98l
dec4t6v3Jx0RZX3hlFCHn+Qz3aM/7CrYtkQHZGdknufeUdI9DFgzviWMPfdhI+iuXXTzXn9ptxET
IzWefnWj06OAziSZ89zzWOW5i3vwRHseE2y2f8zZqbFruGY5lNUcoAv+G79TmhHlyz08T8UhQrBf
BOBxwSulJGi9kDxAAWYPpbvq5bNqiA+GA1+dFuPAUJlSKlG+AWCg94Gg1PP4U+vPois3OuSYqcsf
0xuOf0bDMPZHys3mR4beNvpPa/mYNr6Da6CUNiHcqIvwYleG0p3zoF+EoqY23OhkHDsygjCO19q2
QSQbhOA9lIN6pLye9f8HiX+6U8X/PpiyYaCRR8Fq8xFK8+c7omiWvVLsXSGI9qjCn+jqRCXv7Mcs
MSXe0uxedsCBbpj0enESeWu2bJjsrDOq0ZJt6tc5tkjIpQRg3S1/0kX0LSX2GowFwLOz8FgMy2LQ
cowFytRlK6OaX6xg3oIW/NUE33fz+JTqkcO1QxtsicDEmhoD0LWLXAbNCibumgPvb4nwXj0FZXVR
cw+wEeguwEa46PWP/uqio6Ojztd9xRHxks81+RfRgLqtnaxKpeaEBbj/OPKLs4feHIu9OolZ/pU+
VrD4paxFElMDJKPIbgDlmo9e5+mSpkCrY+/VEsbsjG+3yGWhogs7W1PzIqQlGdyOwxbNdA51I4NS
FNlOTIePH+TPM0vUMKqZ1HfMqc7uR0c/enAXAXMz7GeKjgm+tQq7ENnu2LgvNWdiHVAMaYmtHupC
LMq3mdo2kevSy/IVGK86Izh4ULTiVwGliyisfgOdC3j8ZImfwmURGZJeqWXSuTV0bqp3XC3mfkl7
/DVe8Q9emtGNFf2BHHqsB9rFwpqhETiwfM5mPlnJY6HL+lk1XrWcH5yO0lzSno1jt1w3rq/JRwKG
SmEY8gLrYP2mUDzy6sn+vfchSMLYGJu5T7gJnIMFOIyIUXVFSuGvHPmVLfdDv237jj0/pBDu0BPO
tS9U4TwAPIO79sW2UtmD5YudObTQSWbLw0M0qOFYvSPws92W8Um2dQrkaFY2pqxbu76COOeU+BSC
73iCdTLXXbXFWOTozoieDgdi7M+odmWGkpgJxfy8bd3k/FKxWidCo2BSbil4PUO/Jgm8/+o9XA+R
lBLcRHk4OkIF5UEr3+ieMe8EG6MF6fyBo5NG71O/qvVBsF66TAUFwPOTVS4d1zZKkjYTY51/OfLS
WD/BT/oZFzGPGtAttrcIWqC8yLCEe2QIje4cBSB4Muj8fqH20ZIgpYxYlL07c/0SE099fbAiNcw7
xDFALaoF7F578H5lWrNWapvJKLMmkru+0aUF31kHIImg49UscFfElroa1inqQjBum9fiXRY97tQo
2ZOaHxSzY7yhoFBsmBzTn3Slqy/EY1WKfXWFx58s2R9KuICGUMKWIor64VI1PBYtlUHlbJbtwlr5
Rhx7hjJfgPnBNh/PNixfDdYz7XNwgOgWQcL0nARruDich/CjBLmzafoDt0YPBpaarxtAvEhPICkX
nHeDwCh///BQWh2D6QJN5hXQ3KwYHjz8ANvfUQuWvRVIsbsrSR2l00NegkhodKNWoQ8YlSZQpilR
zGK/EZJ8VBVIr3ISssYfEEpn6xfd0lQnP9XriTogcueF/7M50/gzzOGhLRv6WacoeLiuAeaRVZcT
6EjMtdAO6egO4r7xh6F1rt9PsXmzFSiIavsesoTT5fAbavpJfCQqwIWxSBSW2B0EoOPEA7MSGm/l
juNFr+eig7xicQSZjVv5YF1XVpA3XNTNhgSDMaIeHbJCSy0K8rzO4Evi2YRX8aTyIzfTLCUmFoHK
lbUfzFY2S9mOOdjHadV+XtOANXpW6qleKsuGamhWtptOHqes/VOuH8CYE/fI3zfeHEhagicWKDUN
mVj+dwKL5Z5a2YUDkajCHjsAEh1q0/TyBIHu4IlcKSvn7wi/ObSThTXTyv6RnqwpzFUs2Xxv4XY1
UnbYkf1kEAnqpQnmB5YvK1oCyfylgXGFDJF+xtE01eNOPSjdOPwVkV3kK3TFJY6ZdL/d0zGe0cQ+
y0B6lTDw2e9QTR9mULRfS+v4sQh47ZqfUsQxQxWJFME6T5QejAao2h4tadlG/9xw8HBNBU/gJlLs
MqL/fkHWmW1R0BzPzxZTSFEkPcGQGoatlaw+eYBNFflk7SgiWrtgDcc0iK7N9wH575KStcgT/2bu
j5U/av/z2llnkiJQzae/ynzDetXB2qYa4mS089+DUdrqF2lO+eaQfK1xradT+o8E/c12T9jg7QAc
8Oa93fSHRedthpTFPfOU8PbsNxm37K7Gv5G8KI03u6yP6JWngpCqHTGiZDrUEDm9R/vwyyjB3K/v
EwzOr8q5TBvXb5DjuZzg06xCGnK8OqjiCEDwITqEDn65L7L2VtHQYahr90WYu/pN068kctXB/w7t
8qPHizKIxN2+uG1d+JrMpoo7hzdTbq7uOyWeuCPSc1jIBJBDT7E2Gc/ccpqzAR3NpfOLcdn+agxJ
E/yExJkAEpqnTCnPpNQVzSwnyR+jcEZND/mE8B5PWwMrMOQESsAGIVLAPj0gVlf/9J4yd+VioMyd
KvXF3vLu8/Q8B0ZAlpU2fp/ckLFIM9gKZ8O9L+b+lCIJGiULav5UvLQmsbdFvCT2Lbh8lVatWvOG
ZWJ/hjwdxp5YO9n48RbqQA7Qoe4QN7MugITee7Xoy72G0uzoh7IIXQm72klrPl/Mnap5uBWdwubU
k7FmY2sk8J4HKnr0ofYXYZVdJ3bEnjn8neBmPpJeg5OEzizvo7pKk5KcthatFA3wPK6TEB88GxER
3veaJnGUR9dNFoRjuuznKFUpCK4pH11gWDjd5jH9GxBmPp8td32LCyGURyM9q/9F5jBhngZQX0fF
ri/yQ0T3RzlmH+x7E36GU3E9E8dMqP/sGhbCb5I1Jvurb5PtqNTIK5VU7pj0f8ZKThQ8zfvblzph
qKbeCfcNOFjLIr13/Sl1xlIKoLVNR7/BzscdfKEkh28zPR56BFWLi4vXGrkizSNSeiHFNfeS1Sue
3fHC0oKEZT1wHn+k82nAYeVRjNb2g6nV9UIXLqsZfp4ipbqnTJie2sjRW2BV0nAd6OnWgURSqHvm
WxcP0c169E8vb6QEBR9RObepYJ8YBAOsH4zLaoF61O79aHTc+wujxCw3CcSp1vARUfS9OseqD0bU
4pl0CVes7C5+oxY9TLZPrdt5V2HWxrSt08VXHFSIG+Xweupyb7SpKSOo8g1dWNHWxOXi6zoisghx
4a7Nry91Tx3BdLQnbM+GmEvzbRUeRl2UAY8XIW741vtxj6mxaBVasg+rpuGhPntjTrXlh2ZY7unw
qI+YyY5HF9ve370rvUW+HPeYagouRbeFqRAfVVEFENvMvwvhCnJl0CH7Oc2d09IhAVAAdf7Jdhxd
bJu8Hvsc3ly6Otyr48JXvtB4yJ/S7DXmrMzYDxGi7HRxUS0kS7XODsmXUt+17VxdH8KwXM27d9Lc
gdze6Y+5nHDAGEWsRBkAvyd9AvWbqF5rAC1V4yjEfI6JtA7430R8V5SkJ6aWz4FkkVAoZuhFOFyo
9GkY9VG1q6wWeQrRCl2iPa7j7rou5+nb0F8iGM/yUY/ygKnILbMk6/AdT63rqE7VsLwNl4OZn7Sw
dAecK8JiLmDTV2o8AKazcw+SP+7JtTOt0Pdg5/lfBROT0/YFpWPGx41XDFF30J0Hi17RhhqR8Eul
4KXCNR4Yl+O1YN9yVD5z5l0KdInUM6ox+oju9hSbiaX1f6TxCgu7FmU5DiKeAK6JH/0HwYeuMAwB
t5SNG3JC7rslAHuCnAMx7Q2zIuvPAXi2iPF33411t4lZEX4w4cETfcb1mQJmkveyidVWqrqlIaSh
DENnZ280qfURXb/B9NO+LEOFUa0uJcysteuYeTLAMeE3rID5TRFZMNxC4UNdBpj2OVje2tLaS6Eb
NFZwOngE+zgcCWjju6HWbw+7nwi7eD76jV61w6T6GP8Lk7eQFNV+nULk7k3iDkt+rIsRJW4NevDE
M6Y9Jje20a3rCP3T0ZoIc6P0H5lUPIk5XLNlv0fH4xKY1saMye4Vq/LFt7O7+pGPTjqAHPtGXUqt
qoOV4QtIN9CPlNe8eIArmbT00pVGDdgQk1RETEuOuhVT2uHjkAK+GoIrSu5mvoXZGwJOTYdLdJEd
NNpPJjfMIbRb9Ae4gDLoIuw6WZGvpnpXVJDwhOEjDrPVqGOsO8fGHtYl8/vpkBQpBhdsa1/O9aEr
JtEhjMMgO/W2PrjUSo8d3D6Gq5qaCyPwS6BctnySL26XhPWd3CP4x0spfy+33YM2HrJtm2rZkAeR
+odP/eyiKbG62UWxnny4NJukXpcJc8WDZtZ+NmhlD69tDIERUxXQ2KDhL2nMr+VvvY01wHQXfukL
ORpqJAUMHqSe0yRVBIgf84KhNHre2wrww04iD8t6MMrefQitDYEP/vpqiErm7NzHRYPgC2/nXk2D
+C1Y4/c44JkbDTvjxCpFyg/SdusUJjaKx5L0s7ERPg/YdqwnfwkpiECxruWlTY08z6nQIU+9AIo/
a2JFEsGDZqbacC6FEsRL6B9mVyExIFh42aQXuomRazbupdCYaYhaFnSHHpTMuEI/zcVFA6Om9hLL
m7TS1AyNyfGPSwi2b+pcd68a1YkVaMCLQpco/MspirgTyqOU32EML9nwMr+ew4S6k0xRgwWiYk0v
BhB0b6UjY2w3uN3HvPdjJjgkSiog2AL3ngxoLafenpz5uoxPDEKLalnB0vNZ1rCyxSdJoU7/T+/r
Eg4eCMHC33lq/uDpvukGRIuw+VFNQC7bx33CCawUYwFSERslIFrWfQpdhqfCoM55QeR7anUNWb+N
IYDRJyeFSznz5ASe/Iye0Ur5BOwbEc9ygiwjPSsBx8BLFpaUaNc/wrXHKSafqCHP7o5VWqxmpVHb
OUTLG3HmKz3DG92J3sJ2kU0ogAreVZJcULZJ5uP46CWRaLEhknmRfZHIMzUq4dkgiIyPunjhGarM
lM+5Ym0p20AyFCG1mH+dm27hN779e1qvZFbUXugIbHsWFHDHDlu7htkbSzOdO0XwRlCF+SHivF/Z
NEE7g738UyeHlpdCP91FsQcTe2D0cnX4MfLdwWa/jVko3fpDHaRYiS7bY9VxQx0vzDwTju5W7cvD
mubGsd0WWh6xoZEQvYJW2AkzHoXXs4w4hxn+2Aj3pJI9ONMYBUNfq4jg8DPAKhqCij8OA4xOZ6aT
xcC3ssiaLoAX/m5EdNr+Qz0keqDoKzXGiMepiVRg//uYV56bXDONr6CMyZ2gjl4uot5GiQoh0E9V
yoL7aA4S1+CQq/boD3GoxNIeacc9HWFTFFctUeiA3quFdvpttaf6GmKYgAjYEY9sesrtuTaTJdjt
OxsqKLeRmPN5PrkEldS7kCfFeiRVm8RrI4tbbQ3sV43sYe7Q9mS8GxBfUci5XOd16GxLpzKaEX0D
K1e/1S+cCZTxdV0PIXDyyWVFWD8lu42HVh+T4wgaHTBl7wYhKT6u/1KsanNySty3jmcoVP7tBIkt
UgoTRS4HkPVSnPhm+gbs8LJdnDjN9ZtgZr/XfT9B4n1EIDsXHUtRWDayJOe7hWTlca1SOkkvlzgH
M5lIOSXIq9ewbCLcXP+GFHTA47w4mDKCezw3l3ntRqpT2z/eaxNYgeU0O7cqRpShPIn1AYGppBiP
ywNKSVQdJmBxLN9zy/n/+XE9H3wyX5FwoHXjkGb3LmqxTVYivX69faXnAIuJpISYZ+vWAV7BMFjl
4LWmcgOv0PkgKB4dUJeWBfEV5O9GfU+M1FzYYfyAeAz/JT0nPmq9RklWx4yKB/n73WC5aeumPfmy
deK7r4WQjNPkEZMAaXeqts5QPEyPeLojncOO+uUV7VvKIO1t0n+pCQ6ue/TNvNpUnrYsj/iDxE8s
jZMK0znruN51ST/NGTW4p4VvbOtHmRSpY+Gz/MUH9JybU2eI85GJA7vj62I5OeAnhOuUS8of9UzW
Z52hKezjevTSHaHkmAQXeKAabh/MIzaFjxMM1e+TZKnFzx6CjeLcroVBn9VfKMb8CkvglSagCGT8
WEWVTDA22nLe85H03TgjtcEnx2W018z2NuVJEpJK9hPQfHVfpXzyX45HlQqXcSzzbaDLj+CtNjnf
3EkZ+IKgbKt55T1QZrl1iCeEeUeGVehDxOWPTtW3nYFyUtNK5bbYXdp5F/IpJE4vMIqLD9NennY0
YBFHnIdw3IrQJy+ywBNg3Qh+VBoVCqHkZWVCNfbLlBvjew4HcWdI1TuGDFuDl5FFit0D0uNiaosJ
Xzao34iIEz0HlPY0yVaNe5emLaXvIV0o9qgdlWRtcPAqaIO5HKzDBs4vmavGplByZgSzhkwkUFyU
ytH3ijHux+/EGo2VpW2taxqinpEjbEaVHd6Pm9bHazqpOshbop2fgxYB+8ZlkFFTmehBdZAhdm31
Q8Xugq36mGS5r/04X/rMxzlIlBlEhWRI904jBTH+19EXyzgChUyeD0U9Ae/kZ+B/vQMZEXsWSZAv
NcdoUdKlJ94JLG2tXzbsVmX62rbbhXlSmBtHeEeYxodo6wSpdJm6lVYc1F0O5KLeA4f1co4ic4y9
YmX9aX48HaF9xA3YNacz4Br6QPn0TjG+v1inBkrm92tQd9TpPirNcN/4odz88GGxDL48cGOpsMtU
3Gr+EoHlXL2Jpv/hEoHFG++Bn3x4VqJ/eyjvo30f32h/qgA45qT8cpdHI1rXYP+s4Jtwra/A9Dtn
Kr906MJVOmiR5DS+XyHEu9PUixSC++TEFsacF0ezw4ZZanySo75ahUv3QiM2csGghz4VIhM68sgG
iaGewo/ECh5g+JP36LVA3LX8Z2a7xybkXrET4Vslrjln6utC+qOViqAZiiaSr7DMQkxKdlB55bru
2m9hRKwTyuOVEQHCEA2QZOq9xlsoV2UpTnr9bJy2v2ouy19ZDJaq8cRG0LMCBFMwPz0h1tDmASFw
YNsJXtrpCCeQ8ZdN8z2wUrF8nIZFUKkgCvebZ3pfdr7fJt/g8xdkqesnegd080tPQWZQsvuJvuDl
3pxZSTJJJe162DAvrFblbqk2vZrO8rT7utTpPhsCGzBDJoiZmY3p/9LgNNrcAK06zQtbIw0RN7bV
JKqEx+M2eFYaOzSUYWZYq5WXncmcALuGSwv8VBVi15Cs8dPiTrkx62KubQVZ5LtXehOsgPDDBBf5
H7iwNJXWdUTcM/8lpQWupDabOwL2YioncoV+169tIoPDfZk/O5uoBD6heZQseMnX2dl6rFQxhFem
N62b0AecP+2txIN8dD/gDmITeXN26x86RiuTWhnPQjIgPhL//vLGUB04W8bQoHsY1kgQ1wv/QeR2
ROSIerT2G7F0rDsPfEGn6LIctg9vEdT0fb878kvhENaAj4UyjMFEc2neTXfToMHfT2O7Odvu7vHH
CaIl1FPwFjTDYWZhfnWwpobxj5SV0IM1OUA3xxVkZeUDPwOTXMx5G76LV1QfFsVqHNBWI2eZNfLx
hsSQqVNc9gIZq9kDfjOdQxSTBK1C6MpFGCWUgptaQ9+BJo0OhY6DL0xwSkpm/XrTOgUcGHC8gCxw
suPK3NYVysIrdxj3z0DXecnpdfLfnKGVR4lWTpako4FKEWPPCUvVvY9N3WjJwjyEPHLd1bRdScB7
rRHASDv97Kp0TMQO4PnQBa1HzbQdD8wUmbjxWmeJxjr9N6KbHsloAaUz5tRnzHD3Ck9DHJluTbBr
uh1jiITWnMb6ri7CwQFFiq8Kwn6gwnFCbhUJAB+CC0PE+32tKJKeQjHL/7P1SXIfQmpNMFo8l6xp
scgUpErlzKf6EQywzBlRnp0EVkh68vZb5ESArpz+WxkgKG221r9uhY6GsMR50gh0UbPdYHqK/US2
GDqE3D7z1gcCjJzYiYC8Lr2eq/DyvD1qtX4nKdnpN0RcoGKaOdjCvYgMe0j3tPtRe5vFWemlyxRD
Yp7rv6qCWUPLx5RRvAYkrkTH1uIecP1mhSwhdPAmEq8UnCqQTugLj7HiQ7NbhyhufqEQDfJgZZxz
+62/DsA8gBjSkWOL1taPHwRlRW+kcDSDAOhdkb2b5FwBVaTyfrzwpOHCUoIowJjXqdgHPQaJy+j9
OskWWjA2WFmvA8AgDR8/TU5pJYNPLG/ymFdEkFiz8+GgbDsctXAMCbw2Wf5nhQTwYI/SCUeFrgP4
zLrW79WGVPxhqlNBt1kvPgaggwv6JNw7bxbw9eXpagGXTBqd8vMGU0mr+xRm2morLrfnztolG6Gn
E4iesIHjNo/V43OLAl2UNLHYR8aPlIMRYzygrxSpw1/1JIFlDG+d/xVt83S7sDzGjsswhu5NXDbp
NUd/kqLH9mk2nygxGe6ts4VIX89MWBo1NgVs/Ex3EB3ryqjFAHhxUe8WY/xZtmJ+oxBF//Eoqni8
NsFVl/hdo9r6GDKB8NF+eeKtciF92LpUUtWJf83oT0LplijARnzoYSVu6llLEqDUDxk8QBONqnVK
s+4ZbAW8/fcUeu9MF1ZhN/HPg2B5xPvu/XTb4re0AWby7rC0GE6yDjHtoHkDK6xRLDyfi4/M2oMP
xPr0735lGL27d1KCZeV5AMy8m/e73kugvxxbGxuEVdyYq8Jhm7926hiFtXlIOMesID2Oil6tmfat
XYudty1ON3hT1cDIiN4SmgM/dNIVKxydlejB9q39xXBwV4VyAmjPpwpEv1ocZYSNo70m/odr3CU7
6Uh+8C/OBR/9+vbCIFs86eGo1CdpseXfg0GZmlRVC7ixzuHMGuC/W3Sp974XBcbeIlysmNYu7GyG
YCl1W/uxfN9L6agYrY99dB81imrXmgZMnjLZb+1wI8vi64hSAnbzgeEEXCj1tXoDOirKSgraqYIE
CLKn/b773DwXS6t5fsN9u8UMJpmX2S5w7X48fYfk3bCon3u91CpK6A4t6mswRLfeTEPMgXVzyZ3r
c13eBZ1XB5dyWHw6aTaO2I7+bMx2H82qHEEjm+LLNyTa22acbYBEzj6DzDLeHciNYkXFwZrVvO5L
cKp0p8SOgk5JQ3e6X6WbnPPEuAwQZ8XaWr35Na/tG9BHWIG1uhGf3Z9w7e9prswLYmlzusGc3AIs
dSkq8Mwu+I4ScbD7Yu+JdskfLg/QOJEpah7NbrBjbAoFi9QP4A/7B3BjbW7L2JTOGKzZfboBS9xT
jnEUb4BY9t/qhCzV/cl0WDvaW9lQ6IR2fjvTcxllU0XwL8xPQyNmLaxissQWqtvnbmvT5B4TUh71
1sIbJ+2I+iY6Ez7xqqA/TLP+7CmY5HxWoVdggjS8k+83xwWnKdcTvDQUL+MHxjkPIC5lEgICfz/T
E7vyJk95RGodmp9m/wgIWoMXl0di3gb/SZVLgs9jQOmBbS59dY2UIzNXzZkKomGxJ+QnRJK/nQwN
TPAIOZNYplMvqCZ6P2Eny0MjGFkp5OV2RzhHe+xF0MA/kn5iKON76y47Gy4uBjz5nqpFd6DinCch
4gGJhNYmG4jorlaZ2BhCPQEcNgi/ZQFZefqPSvIkwp2kuVrhmuWekbM2ATW7EH7l/U+T8vJi0Et/
G/Y82A1byO52sm5fIoYhU7guHzB7PlOUp2WLcBeLjam3LjmxOo7U+LEFGJDnxoF8Nbuk7MS0/ohN
CkACP/7P/Ha1L+wY1vHS6oefDSP16mn7IVGxwdvEFxvlm0c5S6YSfo6kkesbFUOu74SdA6SyxrRc
In8hSLLfbdxAWmU2CdNRGJeg+IO/ouV8A7DDNXAvZ0eRnlHSgjvSDbLb1uAXxFUX71FBDbJYMZwN
Y/6D/2YGA9nS7Lj7OsOa0ERQbm1po7RsuyI4x3qCfk/zQ51ea6Pgo/RDyVtvXmikeev9V8ITJb39
Ai9N/FoPTHmf3aePuNpXqEdJeTMT0SjKtLHFwafSPNIVaynNj6OKgu2ctgc0cvbr4G6SJXHYlQGI
REHL/8Zil3s6XfiabQk0dSdzO4J7yFGCgKKh3H8m9FDp+Rca9hV8j3+WLVhvDeUtYNOVfRHwjlwN
x5R4vqbXFUws13wbf+kOC3rKacrpkxP26BMbeKmRzRQiKmnmvh3usRJvC5aCjBoBDeF8wvUMbQ4J
1y4E0I4dLx8XXQbQY1ZbmOHdV1OmaYihfUcbDv3ayaAFQlv1bPBWIU47f1nrSmTkcvGgjNKu857m
BHf2UPgvESRVZW8eWOX8Wu1WZ9Fba7F3+NH9jLXly2h55uOQ+np3YMPEnVK6anVTkb4hmc+KROAt
NFgIcBMV/POO1l6/KBxwmN/Xlhg4N+5x64+Baea6+ZsqqvXXfarMwLy0LGWU3xdlJCRIO9QoMCSw
DCclTGmkoNRctCm6xTPtDn3HdosmpY+VNSQLUTVVpxCzXjMB2s2SzLpmEgdXPFmPKEw7iGAnrVjj
TfJgAzWBxLeB6IU4I8iKUIiju5a3IOyNa+qXaX1FVwnsh8E5d4Q0lTag+Qhw2wFSryGnb2aznV+w
/eKuPQI2llafUc1VnPlr/OG0ncs5hFrGtL/jU1nxOVOXW0VMf8A/DIurn3GZ3Zld289vm4tlhjtN
TOJYdAJcHFpf0kxqAhCDHlm03xeWeJ8wd1BRhcc+ZramVnrJZSH73j5/DMH0rXIitGZ2zrwprMV/
3qVpn0akban0uEasC95JOE29CIHeNcf1Ytaqq2EZPJ3SZLH+Sh7k8pH5c0wKlDTD1/uOxUrbNmCG
4708rwLflCQuX/7sKTRhme2+hwz8gKQxGTYbAqEQXJ7z9hIZlS1kpqCJgUtSoR/AMxfMa/ixHngL
yP/ytxhm9FyuilB1345vIQ9ufOr0jgpQvbla+Ii7w9Wq7sqGpbDJl6K9tJvWBa9J9qkVcLYJgQR7
/bvEoqzwEn8lQeMShW3UfrKpJ2gJqPCTzYG7DPOXZxMh1wljt1epr1uxYHQ7+ovLYe0pMhs10ZD2
+xbdbL0PO3LicUq+4hV7uz/btoVNoe9tQTT6Q6HXFf/B8rwD19dEwNeYid1dK+lWvPvu3Ng/LUbm
1bcL2FpvLJpj3xTcGXXUcvQe8W4wKIZTsv7wAHOb0b2GBHBVunPEEytWK/oB8lTvLZk9eaXZiXYN
7jMZgizg1YzN/lTCAQqh4GINZUN9RkZeBEP0VupvOk5UVEv3vebVuYo1y9yzdbx8UFgHkCVipFh/
d947W11xQvSE60XHKq0hNZHNYwX8j9V1Fm8KTGzImdSPQ8zrauq0+Cq56WDaacTVxBAYPeJNSDmb
jt4LYCWhV90QUm+909BVNy2FYviD0rit4W2hqt7gzvJ1FROY4ZVLs/2+aSeTnGylRC6ijjmKVZsc
HY+JynsNUBltGDNc/0tp/j5Ue1US1+AcRy4JNE1GgD2TfXYf1inKyDDBOs5JTHBhNATWiOpnBnaH
1vRifQ2g+zzpSKwhLRhpOBO+R+MJI1hc2PaWiPks0FERlsDc+fh3wZZAf/+ADAFuctK/wq5sDkKi
7nXrP2dpaRNdsB2PFPZLipvIT87ZoQEP7ukCZrQflaKobll+4WxHJyiIzCWYunfTqeX9ecfHX2bL
T/sJXJvv+Q+zfXXfUIjp7R3VhLPpbRX9pWIEAvGlZShDTyOE7pioYCcrsAGNdAZl8068iifEXQM3
kxLTtFAzV517kCq/FAlwbofCi6N+d+Py7SaWx0DhHybm8nLCPTtKsA2AuP9eAWJzJfXG0F51FjuP
+EEz2GeT+kUaP7iIa0t/Z/t5ZiN8IyWJ2FYssHzqYCd78H6sGQqQv0zRY80eCqgBplfNhxSLDROI
DwVPsEnfgvCEiFnc+YIi+hSh0iiJ9qJ+tdbsWQDRWQe6Ay1ORftifvFQz+G+LXY+6MPXdjrTCmvz
QBpTUYmzkm4tqxGuguOUjb9dxBCqXemxdxOq31BEfovMV6aqQbrINxcakdWUQ3KXV/cF3OqriqWG
l5cr9bRojxozK31b7R7ajmMFHKekuwM6fY9BOnQ6N3Pl65yQgmCf8IFr4skix3zFVkKw1ONuy9pu
xKH30qR/u+9OvBSh+KDtw2oX1SMIcEQTc8vDgEvJ1F5znNIyOtUTjSa2MfEdynH+ibPMR8GXSRbA
kOJww3/wcEz7lQPOy3ZSQSaotTiMqDroMDHQI19BjJwCY37R+6xtqPu7yu3kTYg8TEeawNGXdJKQ
dJkI5s6LQQ4wn5fk8XVB0eATxuYgRmelYOgmiv7HjZkcJOFhTIRe0R4G/V7nXJNJ53Jas0FwED1Z
BzY3TRsa5mA4oPxi9fNmtrG1BlQyF//SkYRhQenWzCbKJ4AmIBrjkrYzZ0tH7WeWcf8r1owg3LVY
dWh4JTNmPWvnHXlmbpFdmiHwb0Iv8EcXzNpuX1djiSs+mLChWKErezrb93HcSqSa7/thePwULh8o
zqU9qZK8pQu65Ltw97/OqFCx8FJJ1xXC00vkq/4hQrIETIQAr5gRGJRSyZIuL2CRpdpA/FWGMeut
n5xQdCyitNnPbU0r402vpk64eNRcdFJm41jp+yeZ8q0VZTGJAIoHp5uBHqVyVUBF1o7lnLTUqt6R
RwB3+oLbBcqWVhSxP4I8CUMDwF8UYLbuFAjsYYcb1wI9dD1Tg12EBQOdyrSvBscLUz8Jgm1jHgSG
mHnilWgmeaKCCONlyu4kgGBAvnKZOhBBFedBGxPARYcA+DkJ+31upxhBpnPvonB0cv3JjtfymqEb
hyOZyNigUlXa5IaS4l+DOoMSbHtS8yp1eIsw7sH4Q+jUC4+THbTmbH8BjMTPxqoWu8+9DwFkl6KK
3KtGPQBQPtGjxoNc/lM6MVYa4u5vFxjTSbzm2AZEeeN+xQDGpy0xQUY70mJjqaCNyT7VroTVaOYG
Xp/pUqpU+atjTxaIl/fhOJLtw3k9x6wbCFRon7qVvD7shZABLNnRWe8r8qRiRhpr9p1BW0LUdcc3
whphPjQSzLX52pCfPQY4QrxaCzqBCB9AO1KGKmMG174KOIJKL+NYLvB0GgO8eX+c0zaaD7n3/JfU
jQTwpHXf9AstoZteYJ8EqppX0LaoOFM7ZhEzTnKUnoWQluev8HEzXiHGVr+Yff7B0lVH5W+rKvDe
FnstAyFd1B/v2T4ufLCzmtQrevLSDcg8FLCumwzxwUl7qT13mvlYI74/S6rzvekApRCheK2uBT9T
x+fqBA/njI6bZmASpD53DuuNWTObXh6a4QoL0LXj6CSRHhygUgMqYx3NycZEmMmTRolrWP8SYxTZ
NBQ4c75vbWQ3fNbd1PBbanEp9wLf/sfnUoTfMSai7vxkNv0aL6MsZLlS6jiLQVLjq1AABZ2/dS5K
P3btamgHON0YwLDlAoSPn0fUcg4TF+jS5/nrd46m0K6FZvTN78yhy4UBvFZyxiYrbm/vz7TMB06Y
RA6ukf96HEi4w48DZJ5QSseBgdDIduAowyn56BeZ8JUl4wnCJVi5E28PnztsSn2U2Ojb3Z665F22
GWTbu4dYzWP/FMHUoEjUe4RWzird9F+D1NHawWiUnbISIJThVw4QHclbMUy7K4BDyHVrOyGhVgjX
QpQ7V1KWugn5LdwUz46mZGx0EelEX1/gq+cAjcnFO5i6fRCt9PEBWiG3JhxNbiXYV/0IbDwTlK2w
Mp6GMy3kz7ypS2gIHIir6HqY/bVncctRL8gSwv/jCtIVxPJOzz4e4bdW/ZuXinvouSsFZTcPbB2/
mmGseUlyww57AAQl3pcySW5gtWbat90AQh7UbKrhA+0vMvPDoPkU8VzVU7JwpBOSQTJ9zn6NKIB8
i/Y+eg0pI1I6DO4Rl9/jiWZf0jezM9pkQPjtwla8xjIzm01gbneDp3XperfSrD/124lZVhp7K3a7
PoGLWNCGp+0Cx/WRuygDMpMkphwckfPZot4HL5c0HlrbG251JHJrHW/79N9mjxgybTbZajvHwX1t
0ecohUpHofkVhcgeA04KWrb7ky5ExQIn9TCC2AqTKyZY9vKN+x0dAwAdnDQmbfTeUU/gP9Mq7hLr
1aG8w3xyXEcPe+MQik9dDXX0ROtKmYP2uNm20uh/FoEdOAKuWKWXc29Cdk52IhuTEdOMzH1l3zUz
NGt2fg7IsEiDRu3jj8HylIWNbP53Ks4RLVGk87n1RjHixPeCdzmCv6yTKnXOuLG5f13niabEYcXj
M5ZmmtPkRkpuqbeGY98Zxa7jWUDLflmNUeEBNqG6M4pPGuM9JV1BcG6l4UAcwOMHgecWiOI2PV/i
fJNXdox1Zr7SBKfAICL6otuIfJqfUfH+yO2uD0ACS8Gxtc/0/T6kDOoSi201s6W+xWMCS8rkid4a
wk+NuIyByUgnsbcqADEEDtWxSKWF2EFhhyS0Kcir36tqIqA9kQBHYPIsbEDHlJieppnpqpYyQE5f
4X9Pe0RdvkQ1COrcNr5V/Dxokm/cqJ7LpywxYBBpRiAAF/aLFUAF82uj+IW3HVtnMYwyYZDf5FvE
me4GW+GuugRLcBKODNkI5zkvI13KSJ6Q0HNtdMvIFP3oBw+bnnZQk9ECfHF2ouRP3okyV/RdXLlj
Lb4a4mTURs/m5XIrafUiJbmOZbAAbqq3zNieEkRuF4iiRMhB5XPwKwjMRMwqCfgTDVp9DrpsLFKa
il04UUOB2nHFbspK+1YJNnClAx54UL53cQmw2nUmsStCvDQ3IYJv5NgYyywfzgEBEUYOBjI6wm0M
AkxLOeIzTLj4TkJYN/9/rZAY0QWrvBddoOr2h5j85vbli9amvbW3bt/82nPpT2X20BljReAqUNKV
Ee7nqoxMoTNJtv+OVc/80SgWjnVzhC3I46fNiU9LrXm4TCF3iwuI6jw3ANd8+2i0qE7xVMdRd7hc
E6De7NuD721Pl5kzYPdcMbkEbHgJ7/YK2rf/6D8sqMPdMNxoT2Y3xencWgLunpIbm4aUFz07RG/y
NGWiw7fv/TneLwv6GbXy6G7jlZhSov9Jt4gX8/hK9SsO+0QSestO7eDdVkZz0MRSUuMFuMpVoEuo
cRccrxk6lMDdPbSCIl2QAleLUSUzRS3J6rCZzIF41Joij7VXYIjSeM7fK2Z9qEW6TGap1fREO6+t
DmCTGXBAJLyca9BeBGFz3JBUyW7PWG7A67CNck7Risr5H1Ng/t+pxa/Gsa/Z1JGkUU1Oh+WopqSV
Osc3Crfu9tlex4nfCSvtTv0RBV7marB1tsVPTKKnIBP2VO8n93Up+xutRmjSygGgN4+AgA01wYNf
q8aQ37r8KWGzPzXTTESaT+YCb9chHGRln6U/XGPLawzDJEXEim15hlC9DwiDcwYX8RwrS+azXRSz
M+APDxpXzpKcmLdkNEyJMISqhfcYMecommoio/RlANrFSFNpwiEr4gmmkmVrKIwh1xk9HfNcHHYV
WpM71QyIGt0aakOf7cS8Ur9RJ2VKFGyMbqUICfGWWjp7EoaUaAsKtOPtW/zuwWGx4JobrSnkZCsY
g1Yz5juUnBKJzqz+RbJ6dNUdP/bGvQuUvp79yD5cigptirm5XVzEXp7lnf3EE5CpW2ZgIDvZWp8r
2umZs2yvWria9NnEWXGpHyj1xwX2tmnixv5hhKtYoSxOn0CQSdmjXRy4Gs6Gn8Y6l1aFlfjIizyO
kv1GYwdjx75+5eNlaizftXwAT3L+sI9NYExJUPf9hcIPEOS0IoGCI06FzXPBM69Os80ERwbMq/dQ
mwuWiSIhlUEI8xwqUxNiw37EZSrjDUD8GNG27+jAfyWSnzckI2mZW2afXWk1JivI9SNMSmeecF+3
sS+qQhVR4N+6jBxFqytMc38t/tTb0ezOHcfxswoowyqH7zOM5RcsSRWw1HVKORp/eBTs5ihuBz+v
I83PFYoEXn+agbJPChEPkyn6u64Yys1OhAhv4zjHGwt7Pq2KrqkfLiYJ8DCtyi1+rpKdRyfCRz6h
l/m6NkMhUrnaOh+Ydrtp2/JZgK252Z0U2mVSfBljhCP7Lh/hTyzXDmljj6cD+GF/1MhOzV/gj837
TGDqInP41Mf0S8Dn3xA7Y2sBvMfIcGxXIIMO7rV9wwUpLD6ijJ2nDW+zcJfFpRet7YyXDuSwE9im
3iB/THTMRjRjOM4sZdYMCSN5cDN8Or+Z8vKczYGM8Ol5ZnsDP81JZC1MX4QXzWo6/PzSWaSekEdy
c23OYVf2HUYDmzsT7dAVEhkXLAW/BPP78QwFgIAWI8ey2T6NiIzRlTLrvIpCZXNQYRSSTwGGtvhW
EP/gjRzxY/u+HIDIS4FSLGoj+ZCOyyIp5r8Sc5fckuN9mnxgzK/BqHoEqdmEp30rHcu8inriLUZ7
aSDu/FYvoohQtBDsSnfQPWKGwU5blvH7wF4PXj/JuMjhVVzsztYeufQRIa/cH1CxNikIXzfweBQh
HfedTX2LL8heVfmAN3nQ18aZqgZG9D67AosZ5DKJ3NXg5b3pzpiRodmbi+3dYp7FTFDkds9pE4w7
tV+2NmUVZ8wbWpe3QPgQJKNvyJV2t80gVPj9MZ1NwUdhWD5/ZF1v8i8HvnYZ1myRM4aOKblX8bUq
CgjuYw0qeuJvqO9bgTFvcqT4TgArKuYZ4VmDH5ONXW5ogy3CYC3Ew99kX6y8m2hRcxXRxcV2Lam8
ajtf9iLllgPKxARZ2xCZ/Orz2oybSpcj6izJUg/2tuz0vh7kIE+u2yayPOFkkcnWt06Pe+fxwaJf
QP8SI7p3VhD1Mq4Z5vplYbWkUMpoSKSRrXKvMXqicLJpmuSg38ziwxBa0JV5wTFGckHUr77vWg6A
gWFaKoawJvIqAitI9uv9eP19K08yIrt7VyHPqaNJWT1xgDnstiGexO3ajMyHxG/bskzZiwL0jXvv
aOBOl2Qk/5NXvKpg25UdhYU12axa0VyRVUQ6qUDeABo0k88NEcr/ruINOGD4TubCAnsprmb5wqay
1qLW1vSC/i0X9a/yEV0UP7rGa1LePDILAyqEgk0U67t92H7VTHF0dnVFvBHYxaleYn30u4yJ5fm0
o/rNzfezSJCvOELe/JWwMfE3xRLZsc0XdYeg0QnBZFIhKX+4SJ8rHze9RKt8P3ml0KFFgLVwXWji
YA+YOEkKPgt50po91LH1xBcQhIUw5kXVFfZNHqwGP1dh8yD3GsBAltob2jXANyriuyqZc7KPF5oB
YXjXgplJXFH47VONrb/pzK4k2B+fInMLDnVct/im2bDBbghvogMOV4Y+qvflQb0ulC5gcUDbnreR
HKG7I9SpxzpxDh9E8mr/BKaoOH8J6wB2boKatmFscRDadmp1rV6KlmVJimqHzLQwgYtOgIG1ZJU+
MImveNhdFgXIj8FhuwsCHqdjfSkciVgDlfYazR85xkZmCjaRKLZYFCWU/zyWKenZkSyrH6Tohpi1
rKD4CQetaeKzzyVEyPIwKQc3ep5HBudsjTPW5NqYqvtX21xFYnX3z6GtJb3RPBZI6EfHxfFwEicJ
pL/5UmZ7f8V/Xsj/t8i/k6v7/Zi4wrJAT18F2uMr0WYrzSzvRcCX/YOpsGTEV6LZW5rCoiFBVti/
fF10zT1Iwri8NhMwG1vZhnL5L86DLxNcQqXztLClFBqxZlBKYC8tDZGPUvB1ImU6mZQVlUdvAxRQ
8B3tIIvyPXy5jqppoP3YnT18JvYMGsePJZO0wtCfWWTl1TsoPogqjdeA9LWcnoqru/c7ybTp5KOL
uBhGP+G+hdczm/p2237DUMHG6+dptRQ+Dd+aSEM7OvctbK0bbjtkg2G2i8X6WzebYUWNIWBgGew4
W0FTbRsjhpMtFtTNucIpQ65nQf44jOUeEkTy/zElYx4gTijZLdVtADTuPj39EeHcqEfy5UsXCOAC
Nx0tpeXVkTEHkTcR50k2kKJmsfjB/RJm/ZCfymLz6cb4cR67BlQRRvqupQEVX0jEGfvdOz/4pWLA
r3NiFLabh1Bu/Ec3ZLL3MgDCCQR7tw7o9qQJTUEmkRxVaEt1dFXsHg9A4JWCCxMKOWENOHbr6422
yAZVxdZs2L8pm6s+jRaw/fyzA8Ech/wixUphegAkESW0PHKvBg0L7wgzR0Ey86VgZUZKH16YeVW9
eH60Z7nq80eLvJHUkscgXTse0WjsHlwa9MGuoqSuIweSjrXRe7dPMwoeZiZBGtdKLwLxAzD1p9qQ
pgxaNWGCi4DCYEwQJA4JP4qfHpDz/NyqYCTNYgMtlygVJ0Vkcbo07eyFIHMkMhuz97RRMkDyfEh1
1iWuCwxJx25V/CKWJ0jP6KfmA5DPXfCZYFb/Wog6QKsMS4vx9rWBb2JfKP9yUT7KjLAQP2MwNB9a
/d61uIiXOJ33FXi7jaxxiHDskf11sWwUeUYIICcZR+DASH5a2L5ZQtU53/EN7SOpFVMf7NKFkI/C
0azGn65YEvzLnS9attKAg40wubAmWlIPZoSu000mNf3EIoLnykF3nFgLEBMHllNBWGgpSpyGTESV
QEvkEDORDFKqXmWNRoF0Nru2cXIXXMIghS4nuQMOxlOjGC+ZO1h2pmlJYzvRiIdDMOykx4sJQr1E
KlWUMrZE9mPkFVXtg0gzppGQvQ/lTqqne9K7WLh5Kr3XG3lvT/atL7/UC61oMHHApYbuDx4AWqNV
HksLl4JU8pEh8qHBC40bsj6l9o0xFfaviMHqhGh0JDC1uVZWZzj+9F+Lix0zzk6/E7h0000HtLKy
CrgkxBRSyPoGO9jUr5B6/Lo6+Nh7v1vVGjougscKtANpJ1q37gsxrcz0me7g27k47IxVxokNJURY
7vgXRqxog1XawYQ10bvMCBQOwNK0FmQPpGuk2iojKBcKvbS0DC2sniXFTru1Y9WoQpSEZjqx22Pl
O/8EZyrbdWqHT/yvgC+J9/SCZs6bXPBbG0Sr19pXLvTNKZVsYL614/+XdVey2JsQ/Zuyv1MAvK1a
Cq4Gx+krRzxnOzEnopdCwqrMrC77WelfBZzlbhnVQkTsaA6WCp2nVyejGbK64xQQEy0rgZjQMpHA
c6uiEo7kyLDF49svpjPwbJ3V1hd9VmiqePAmEJuNoArU8rNGsQcgFtwIPIlwz+/i685+YUPnsR6W
vScffeVKpsp1i6/nYRDJKLMqETa+LxaBZFzK16nwnOi3nGfFEzb5K0pF4bwUakKt9EaTd4b0tgYq
v3ltG5rmyIOagagULMY31a7iue262ZnOinmS2iHbUgwqlLzwCS0+THpHPmmqkxoKyI4Yz78ho1Pc
GRQ0dlgWt+6RHOoSwJ1YCQ6jGJoE6Erm2h1YaWKA3tT5Rgm4m7qTYF658zIr5lAba9vfF8en8Tge
Bi7g2ze/izehLDU2zdBFOX0LCpDYrnqNZdlXd0Li7MW8nQef0xOslZXL5ep9tA3eLeQseFahgrRf
NdKgT3zFWliwiIpNFBkG5d1ptPgNvWlLV5Qhn3nS+LItDpH70sexB3g9kN6aYIjWhN63xw8DPR33
M3eJku5lG/BJpzIznZmUsC7Ep3mbXX9yG12k1CNvDmWZKYs8uGby80AAw8XwcXF/9HJhzLynLfV6
bCy3NK5evQI8aKzDWemUS9MVwKz8eAODnfG7Wv5Nv2j88zvG0gxYybum2Rahn23doLx0ruFeTTmY
sCTVAa5oVeaWRzQ/AHdsaVOpXZQN6MUH8euHlFw9CiFwQmZMZaWddg2NW861O6lt8sN05ZxA8sA8
gfvLd9AH8nuukhxdWlTDE/yb80ba9myv+gUceBB/vsi1M4rQIafxe0jwxVOhC+LvOcz8jxbEFAfR
l5+eePaDobTFIj0SmSkMAoawYN5c5SDePxNxGlOi8NlL16307WP6TTVgCbkgmw5ifSCrHRQzGIf3
rMAmg4ORp1nK6TrlmDbVPkbwj6R5iBxrU+FFFRo/RY5JfxDj1QvrdiY6EtvFdRknnXESF+1+hmxS
gMnLUv8rYg1vEg+2wpjiYzRY5NJbkqQ1Qs3rQkYkGfWiQvGSQKczn5oZ8HpFHFNN0f2q4mQUDNXc
k2+WtM2AKNWh+xglKO1y8eOAZ3BTVByxMeUw8WNqL+AwwCHJNmoU+AEjH3uNTNMB4p83EKFJGLgE
zcG4iojeusp0Op+vGfIla920RnqZ9HetK0FgZx08+Z/HK2d5+EY+yVq2mvq2PsvRebWrzR747BpH
xQ6fpwJyLUSo1fG5mOrfL/RGz62Hu56kWljVdvDQRsJPZZGsaiCrEU8d0swM8NXc1Mq8gtYji2K2
+51hSu17FtBuG9e4G0tlTsVsV0obDpK/B3rvXhw57k0P9zmw+behguAjAVnB+Ev1h1/USlIx1GYm
3nf75IwpLRop39TloM1kPTZcJP2O2FQTfSsQx0C2WzCJmqCOW/QfeaaJwOI4CKkv+oSVyXwn+76J
Xvzxs1op96hacsOX2Xl150JUU27y3rD3wgR4zgwkGseFb9D5NVGIDB5qkJprBJqYyHoYBVEc7qxC
hHPSg+mJYnnu11wCbJGRZsG5V0FTHI3bEXIgmlTwEvaDeUFlzHQQYRVIKII/XkEIEBhSRlZ4UlOm
7+PfU3QeDAbZXX38p2J80y5cyLX4Y+2N2xmoTf9PUNGCBRe9Zku4od5XpfkMBrJTSwv4tBq2RC83
EcBv6nAQih+L+VtyMVTndQm45h2qwYWv7U6G96oNZFZurUtayZ4kxOVha4NMGAvN1F4jhbJUEeu5
T0JXx84yVwbxWaBRm5VNktnQOkxCya0alv/sqfkBExUHoj7fUM+CjAKrVxgrSu6Sm+LF03T4asTS
N9PDtEgWhp5E090nBXIfxeE0TQacZI2Ua0zpRdfqSyBhQuh7Dx41uhbnism3UmTzRkyp+gAOd29n
c9oRjIUdG3gfdnoHAy23u3iq/2NTDoMmIhWVRw8Ftp+89Xw1wTfydjX3cEYTyVdlPyKBhvbSl7ZC
LfOp6uuduE+hqUf6RLyVRDNc/2MfulUmqz2c96m0Vc3O3NhC2hcj0zlwEmI/aqKtrAI5In7nYxnY
gFxX0dqOgj3bRZGnaKfr9IYEXvgWA+GPoLw6JTD4Qv5LpGkdHoTarcAy7tAniwbpNPem9vYCdmaZ
MReZSIAh0+37lzXqYWqGjTdAd1V8DuVrmlytHgcBz2v9Nb9ZAgQMHZ+e2K5VtgZbLXWDouSnZjHT
EEOuGbCsSu6KaaoX1QstWvsAL/dr+VrwJi7XlHLEbSNGtfN3TDZ4pSPIC2H4YyDQdi/zVyGJCycU
ZZyxYWWIRlxk6eeUZA8/30FSjQBlzsql3G2t3bUH0lOFlaqu1hO9e3RXBeMUcKY1GdslKXXVi5HR
MkO5FcmOiMMuJgj3Snz1rABt7w+zuHUfDKvolbeOMfjIf/NYQ1VHXWXJXq/7RQYegLQb+NkKHxgP
yBuRtIxdLLgEIXBVUuVn3Sv6yd/UMiEhGdo4uKxTeysatWdiefPIxlZLgFp6E1SmZFWz0SHa5m4t
WsCt1fd29n1tvE+JbkiT/qx2fulegzvXr82Osfw0W30aBFdi+/laFMsvhBZUlxMt8e9eqoTDlvav
zgMNuqZlbqZ+cGhd8tbBn4DTkRbfHxDwGHFLC9knXeQ2piTBLYIbNOBaKDIN9M4SAn1FsN51uEB5
20HG6nqGN979WjkLWCxLdzwG0JsFS/uaZcPI13ohKpJijdsH4dWdrLDWkkb916diV/plKiGKkRq6
LAaf09QQ9oebO7qXcYsiTcFMI9OULCW9qN9k+NKBd5s07ClegEbs6Waugq8xlQTpr8p9B9OgZ6pD
oQLrpcGcDdvvU3VvIlJ1H8E3ScCWA7oMe5JUYJyGBaML/0AyJmuPwPbb0s8Rj/E/XlWk3Vo/HZNH
g0DNtxmMKg4PzCjeWVKtq9XcUBI978BXqesg7PiPJqjmnvsC9nZ/WCUms13yg9w5oxVCGPx886hX
OXzVi4XrZeKvBKypFWl9afGPio8pMc4Pr3/kg22Rzt3ceC61k0sQQfjPjH9Uf7FN0P+Uz70HFzW9
pJ4+05QfVxFoDF2Vagr0gQD/FyqUGz8KYt+VhWcwyS+J0IVFQaJplISuF2XIXQhBVhllDS4GvysR
tSRBFsgf6I4wrPr6KA0cq9H125fRTrJDkPSK2dzRcxUV/3AvJnNNYeUDWUkFVjFwWH4LIRy2PGrf
qIRdv8i2qpDyYRI+/eae0SYLeuQKMrIpkm9PwrT3AZib6YGvtqvZinhsJ7Cjlf2RImKh0auA5aSB
buCPUun3nfMqtoBEgygJjyGPW563GJj60fv6ipral8Nz6eDfoMZhTt68HnkMi7dcRPnjtl68t3k+
5v64tvtkU1eqW29eIhEM5xbUS2KScSDUe2sWKT9hIHJMlTsdT1506KEZWCvUMsUOgudrnd7xtOOh
GIoFmLLYnvi2tDPOSlHBOMNqd6Hqkf2LFEH1HVgD+aCAJ+UvAPU2Sxf0JsAQtExlqmO0Ud5kGeMx
UK8JMuG94vbUIeV0/A1S2PI7hUrQc+5AsnfhxZLkvtoSkmrzBsLhri38RqXDNuHXQpjw1RygFl/W
UAUYgGNOonWyemfdfVuJNwxNwxNmFqnpviY1gUJFQKd9DlBS4JlJjLJZaeZvWcuhPOQgBbyMx/ai
dQB1fqH/tlYURz81iZfS+I6166uT7w09MUOQbWM9k0Yg28GN2K+U2e4eDCmnlzMWXnBL75yWBcAM
N6clI6Uv3/iHVTrqm/xC/2IWk7A2WlfoocABcBysSwQGmmypVhVXFpIHcMvih+GiOGGLZMV+wlq+
kPt49gxXPCgpyhCxi2Q0d/aAXfYR0JpOzxOojJGgb6tu0pfZ5AuvqCqmX5V4hyoNacZDSOBdunSp
LKWbD2FiyMNAk/1aYL9/MBMhwngSoVIsaCmk+90nttUlJMgxPsdKA1xMhXtMgf/7s87aJnC3dpNb
5+wWtmvacJjzqcFtUAgxWwSUTvRiIeMEtCuR1jk35Cq98O02ouTrmyUsCXh1pbnvJtqZjcqH+B/S
+uPkZIvdEolzvdyXsqvguN6xpwQtnAANyLjzoHv1IX1Xy6HMcvF5o+dglxd+8KJWjpV4BFggjyTM
rxegKomRS8qz/7sePNEVR/M8J08gvX6EhUqkw+PUQhrpwMjAAlmtFbS5cOkJTLF9vg3rWGOvx/B+
0XnCaDmuum+fAGoCbDNsGmlypJYHGyX9unIouEnWQaH4TlREFbn2lJDJ7tsjSvaATn96gtJ1hHC6
85bcMQ+E6zrQUYJn78y7v82u8wvFDoDVaZfMG0pGJauCQ71pjfOPCRllUKd0Id3CzhKf1eLofAcm
cftjk00ZPsoXVFO/wXKPAGp6oLUwNwFsbIOMYRo0HaYAw8DM0hSyfmCArVhZ/9+9LXV9lQNhTPNK
RxafSU4p6OsZbu/eeXun+lcm7zNqOh2mD4p28UXmN17fYJGW7mhhq7SyzrLtssgKnQS14y+UAMkl
AN74mteNrr5lGQpsEhgZ+QzeHm5IADD7ZiBE/FpzISzCgx+No9IKClRS6RiotSU14L7UsomDeOFD
3Mdof8gAWvmPEQPKWVWrLVYyWGSF2lAmcrOK3Yc8QB4L+NTYTtzfRbDJMknCM14/avNgBmiPP58z
w1jvzgZDLSrhAPwRVhEhCOFyqnc2xNvDE2BkukcfBViHzPh6fnI5nsWV/roW45+4sPa1JRxuY4wN
R07JYNYd4LcvmePmciyUgoGYbstdaO2EmliDReElUfU4a+5ig05u58cBeAjC+miaQdj4McPz3Dq9
sVjsK8joGAGwedUbDIKm3z8hFWkdFItCcF+NOh2kchUup1g4RPy4/wRSZ6wu1PiAzSuY+KSZ+U9c
P9Txn9aO/qYVAt0UTdfobxMoKft7js+EH3ex4mt6rCH3AssHQtqM+hW9vEAMwScMRBbU8E/stA2t
KS9t4LbR5KvKy6/Hrzi5a00rsH3KIaYKPoRU68CTcRtYMXrX/LLGu27/STd64SVXYn1R1y7w4NOu
miO0Exz1HEzQs4rV+caUNMOKjzv6KJVY7ZmbtHLcwJmxEMAnSEAeJ1bHa8fOsHGajYWZ6frtfx+E
G3wDFzt8Mzzskbvd4XElH43nfrvYn8DRancND0dUn+rnHLHj5yhRP/dzMhrXbpWQ+FXbFh96hYgI
WkPWlZTisjK+h37ZfiFHKIG7vHE9QNEii1MMRtrbXPhgWt+Y/RJdhRgYIdnj36DGC5wdrDuinhRB
FcmfMcfes0KIFj6VvLNdZeWvqCJZPC9ceiYMwQKp5EnEksI8OWrkdu6QWCVMQu/AhGZ0bTSWV6AP
IpxUCeJoGG8W+3kpv9tutXbusPgsEWnwbncwsrg6eLe2uOjw70wXoyHH1XWHZIKVNuANRegYrwo3
o6RJ05PK+7gT1ezgs+UiyTsv7wiR1ZiozJsb49seGxHoUKU2vtr0I0Ie97XuN2tMWJaHao6eYQNF
C0478Y6lflFak4cVIx4HHyby2rr8mMK3n6hm2Y8sJNof+T6MqdQQWAX5aZ0SYBwgWAMgKDQNh2MI
bXCMosMl26Krsm/kduUQw1ptWPyBnMEdfqpjWgQS3/fpJMZrzKt7rHU6A4P3+/L1+msB6znMOdSH
3D+5/QAjzY9Z0oKRyyymkJ7LWC/kkzBq65C1WjVc+ODQgl2nzZV3ACg4ONd3QCkbSWHFIyKY1iyq
83pvyyYetwzHA2OWNdCssk9mRVyedHLc7Q4GgKSlCY7Or9N8hjvyzZ4NSZV2oeKS9KUqD5U7DaOx
0dvqHDlJsCpDLnhg+bp8LqZnMW26KW9J/gRNgdWcmDHoESx3N6aJZGUH9Skg3R7DKiB/CO77Mwud
8LyvwUQAq+/HtJDijiBGf54cNjUSYgbCXi/fZW/2VWSg6R+8wMnR19EQjCbA0SfgssNAD3RlC3Qs
uefw7x176AA/E4Hh55J9ziel8WFP0kaLGMFUFhIyZCGyKeVnU3NFwZCjo7njywW1NrAad/SzmRsb
y34dVpRoegFfLOmUlCSdChmjJsTyh8FTlysO3l8auhpRUpP88W/71licFC3Ebri5FKuFuvSd3d1X
16OKv0taHiWn3tif5NEdvoAOjONkGvSobkgkspyTguEn0bdAUGPnGNhTUOtAWk/GiRgEaXylqplf
QIzjidlrr8wEGep7CImcFwkwqJNM9ojybKQyx791lyG7sddTN0NPV+byeRX5ukKiCAZZyt3HQMQW
6nnugJ59SRumzyGTw1aU1o53dDYsquv3fSeEuuNU5SH4kzI8mYnPMAmj43bPiz3um+fZRGWcv70K
A2Vf4U9Vf+aXbWEYQBQzFjNdHgIsrFNVvpxvHFBf+oO5KtmhiM91IU196SQRzrdjCcskYqkS3ZUq
+Xj6ZfDKEXrGftdc4B6suSdyjZw2K4b9lI0xgxZzwKTC7ipJsgY2XxAXShY3lerh1piCz9K97rWv
EEJnK+V1RSDY0VJwb5sroUHN2yZPjOrvwKxa5YYWcNy3iXHrh2R4NXPgjxeCxCOGpOPfEthfclPn
tjMWys1aOGkKKX8IRdA/XZhQvkF1PGoRurIRg1ltFt9gnO2+zzOYePUkFHb08ZZvExcBaj83PR1w
Wb6pI+kCxbh6JFHV1ylzn9HpOvufofAnuZFmDqwb1VceVaMsTuV4Z/+dF6x/0YVE4Omm/9oRcv02
2NRs8hriA8IbLxFLKgYVG6NzXFaPlTfnK0ONCJw3Yy+eapWMZqaJXHROrs9Bqr0jMHzG9oyCexDE
amjOI535veNQ/BcWSNSCay3REBlmIDUXkZlQOSwmL9zSQRLVkMx7LFGU0b8Nv2Prfva6C2szxx2Q
UyqwP0YsYWwuSPqwIr0l032Sz5Ij7nmYoAINm95frExBDqTkHB4XSrC+suCGzIOK13SBbQQCSL0j
kR9scSoOVMlRlsNPsnRwivK2+0OEko0W5R0syp8kL99KJ6Q1ueGZSSQkDaTg3a3Cagd3STiVKesV
iByWaMsNhIrY+qRFkEF7fVvuP9y7qT/RzP/C4HgLIRJnf5g2RqiKKyMgK398DzStXr42oyMa4lOq
sBrhaZS54W7NLjnTlpTSCjtqci6xkjVzk+0jiFfXgCs7wBTrO/BGWiAy7AF8JSTt/dKbADwiz/yT
cO2mEWhLaYetYOur5eeuwz8fh0Q7psToDLnv+ZOjIB86+mNC3t/q21Vx1sqSAn2u7gv39jPoDqfD
WoafGS67KMtPu3/tc9Jf6VEfDanIWKiVQ8XphWqTv6IRW3H7QJT2/yq0UA/dMHBvQPPRLv8rHKvC
F2As59nwVzF4pHVB8LFCG2UT0kTp9BvTAtSszDtyAS0TP3HwAQMUQZSMyP+9iUgVIen3qhFJkihY
yB7G7lFXxp2QftfElI05boktc5YwDVOYjM+IFnpWsXLBuOuuqQwDGj8o+sARamjdRRrojLQnpjdD
w6QK2RFDQsTVeKFCqTGscul1IKMuqf7KPek7CByEvW6woN2mETA3ejwtyBSSRk7TBFJiEm3Q4nLa
eVmwDMWWNo5rWOMWCRqXiR/vIyEyqEjfhYnh8rJbNSdsTxhicFWlINYLcpedvpK8pfwwVMDMpxY9
cZ1aBZPdatSR2NCtr55zfQrse6fahjp/Sjih91uUGQqOresozYMTTZxcwaP2DAoMqAxcO4W5OoMV
kI1WE6mGDnF8rC6sBafBW2etzTcT/ruAeJ2i8vuf3Bg0juLJgZVtDRt/pkSrYxWtRwKaUlBofiUw
b/pjl0MwIpluevfoXcQpq+dtOLlnSy75TgFT5rrIHVc1gm41feODtoZKJoXx0TQBMM7Nz7ufdas/
XXT/+9vy76aHc7UafENGTSmm1QSeBujnlm25Zws2R0guKiX3G6HicRKAtkHnVASYn5w5hYo7BWqM
cBDOd4yB66ooHNatIhCQMMDvg3G5m2rt0v6ZgNCQ08XyUEg/+uTIX0Ge8PNm1vCNxhautwaybOrn
WRsLvf3X9ZDsjFrCJa6NSSQW57ahbMx6Kzl2uvQED/+Xf8F68yFaZZxU53Ed874uP6vQLnQNUm/g
KHM/Z7u3gw+a4IMcm4J15Fhp47rheN5vLQum4j9irBzC3uQoYMGYofVW+I4TLq12LmEliFPw8Pgt
quYYzdhIj+c68bLC8GPqAVcN2VQY1YGuIjVemUDTcKg6kxN6MfZC/4WKEZsM6rUXaQHqgIZyDgUb
rfsc6lRpCvDx9HLiBc1n5TR0YKXMIHcdUSY7rkx+KVQHJsdv7mI7mBPlqHHyCP5tMCiHvAsiBtyM
6dJLDkd+3KN9YwybV6K2tRkZzAkgG7XLrGXKqc+92R/qLJhc1T85ZvyzQDW8+/xH4V9daH7pzLcO
RWc97tv3M2UzgZkE17Rm5eYGs2k12JtAo4x/O1ucmxKMJK1glDcaD9WMJ9g56BZo+R1A8/wh8+jK
5AlK86fwzZtx9L/yXzULQo+Lb+2nfjsgBLfE6KWW8TQqigfTYtxU5h21DgzCEKY2Abcu0Ae24CG0
gC4SAGm+L9Z4KAXXj+rle4KyggDiXCWguWo876jzlAz+iUXTU7j4uh05igjOUm53NizY7EwEGPwJ
ijWEMx+iCQ0mnJZmJP42uBWVv7Bf8JNdtXfdbpXmkHHJTxvH7k068vF26UFx62ymiWWzNwFfTWI+
AJ2EcBbc0XwVn2N5BapXHvP3a0BrTBxrzmlN1nrBHpD8/JimZiCOQOdcAVWavdm47wMuz/cI8/0Z
0b+lHpjrgMmY8zxMWK075W0ohYEY+lCuvzQcYRT5lCPrPv5IFVtUkf7Q2MoxqPS36ASsi7hDLt+V
RhN3vHk1t7gP/ZMYt6mEe0JGDDwgnpHMajTg4ktSl6f0gFmKasTGSlM2unOAOYERAhLfAebYhbg2
ZymSI8Qunhd4DrPhmKC7tvN3DzHZNKsxXpAf5HGydBl7WmphYidy0Im9nIpQ+zapgxc5shZ6M0hx
oyj998h1eXo5FYxmhRCR5ui+xfMd0y8lw1XYcJU819RI6mRlG/2wdwyay/VuU4AZgZXtZV02k2qZ
qHwU9N5C7KxchpBkb9r4o4+6tXprisV73ecKL/MPBc+wBJm2CGchzPrPLwAr/uRpqNyYr7bp7Wr+
LtXNIkpJi/T5kbW3sSOVVTGYf+nInxK0nCtlMKXfqGN1Gi4dKFCMExvROL2G8+RtSCJW0BDNDlWs
rKLcXhKGQg7XTdI1V+gPG0OZyEp/7gsQ160vrPuqC5IDQXBWS3XEBd0I6HVROOg1qo4WqzdOKKOK
0lvzSwqsksn9X9AVaqYqdgISDS0Rv+utOkkxdkMQ94P6MGnZmrExVsPUqSP5Hd/3rqESbszM8CH0
/JykBQEmefCWuVZ3wBrjmTpfF+oDdks38XRAknFSf5TzLbOe5z4+CUTPe91K4nTdN1p/+GGyXALQ
3LI0Slwmc5i/BONzxKjjm/ZGcev/wAVhqm3/gCnA/RejURip7QscIVF+zOslOae7djzuDnpUq/dJ
pZIpm6qgakfGtLBDymg9VV+DFq6um3qStbzwjEnCZK3p9H9o5rmbOhs/cj9FFyyMgO7Hd/AiADl9
jt32cA6VR2YxwXiemfdE0WTeGipJPa5e/n/w0kakh35bkdkeoutuYcfCqHwSwKU97V5/oWdcNO9e
O1YFtUZ3/oSz08o8vZK19e+cGQbEjtFnIMP6GFMwBmE02CFNG722JcrF10K4ibjL4EuCP3WV/6Sh
feAfMfflqO+orODOKBbUpmFFXEzBtm1UIz20SizATWTol97M3+wjekJ1jNMCRs8y62QnnwBTfkxk
Yb7ChHrVqaBgTjPgVOQbgMALKHUCyGZ4kuNMGGlxGUClXsvZDejbOQ8/CZuGDur/xQf3d5RQgZqS
SHkBIl09l9PQHpDv8YDxCePoNldOdcxkUy8Ap1Z2cTzkMJhjtgqITUyNUCA/91nkXAnmnilZR/n1
Xk5jtlHu/gR7U12JJHNmWEElGXYvbSQ3dLPHH4CMfHHn76rYiSMZwf9DENS1Aia152GCjzwT7vOK
+QLs+4xlMX0ViT3G3FhTwZXQdQzi9tENz/lzyEAU8oIriGfOkMEzdcGmNXymCh1c6RcogCDNfJQU
9hvMR3SmzLGN2wp1eRC0AZQB1Ol0PMF7VXVU69YnfPkXOp7g9I/0h2147NvDMdUK+1tiFCbYvGCy
vyEa5QW5I7dD6m6mOavJJRJJxaqmcc80HCws7id5dFkGAIQwkCYORYWFNpnkxXpeM1Rp761SRdIX
qv9jftb0g3CQ7rY2wjzMb6zqMi9gV4GMF7DuJS3rWwkR/V79wOxZteLwvHJxjdt/Bu1VVELrov72
kjPHxC1/Omf1CO7y7w9fSqPjeSD1eE65ZGhAaz2NMqXFYSfhItVTas5frPzv5P1qo8XRYvHGAXOq
H39QRAY5bsmVQKDFRlP35nJ1OniCw5d03jdCk/Ws7Oc4oYo6XikogtVJ/7iKfOrFaqI3UWJQXax9
l90+BhAgqMJuR1aGuNWEraUO1O//DAP57jvx+Uj20YjXgxzIId/M/vZijlJ+fR/+CNX83eUZJa0b
aueL1abVcsdl84NMoQpmOJq+I2iy1qai4ow83F0P4pydDau6emqGYn301/xRUI5L2l51B7QnxuAg
8ZG5Y140nZOK9yzhSauhRObhlc7Z/HzyI9uAenozq2MUXpoNXSAKsfhbvGikYFT/RFYwiugf8DU5
MsSKrZgv3MCoiW8CfsPw8sGM/QdSHpqi9UbIq6r9q0E8eYw+qbp+iAecZASTNP1L/oJ1EjMcMGJu
j5WArRrAOxR6m5clzjp+UV2C6MdbjihPZfjIX1MjvkRl/sePvN1Uu+oHdHw5CSLO6wRS5UmPxN2l
pxIQamBNy0fC/JIv6vueW5sqCJSh/02PXyCXS6j/u2o0SzmyLzAMJzfMpSd8L9skpb1Vy3ZkoOqx
GQIZpvXcQydLS8zO9WGZ3KZVeDoqDRgEC7/FJ6rxp4/FF9iAY+PMJdWfwgkI/bLgKwzdfgELO0mP
AZakf4eDXy1QeGZ+gIO4wNDd27kHF++ucH6U/CLgyDM5GgkzStnV4z1xrHP8SUmZ0p7k3+f1s+/O
n6WHOmnsTfYBTyKxoPb8INmodpJctiekWJssQANMa+3aBvCAA/ListYAPMJHcqvopowf4l2MerGK
gBXclzm8M91EQ2ECdj8yb+gjdSP/6MQXKaNwHzgX/PD6n0sFo7iITwdz1xM60F18MB2pZGIDKnmk
6wlUemkz2+RPPCUBkPZVIl7JWxEnig3LLnUJxisa5gQUfpWc+B7eboLBOT6rzzMCvTBtDG6Gwf/W
ib/o3JgazbggHrKm5QHbfPwJVdB37FipRcATpK481z1LnyJLlzXbKruPP8XfyDDA8EiZQnE+wGZV
OFEinlRAv8o2JzoriAJEQUALxhcnn3LYcf/NJHfRrM0vMqc8S999nBTLwcejdCJ8SbMbwrJ5OxHM
sKLNqxLqJWyPqm4EYbgyYpa+U6eAIq1zkeQd2L5qPi1/INYYWWzUxlV2D4OO/bN+TIIxk6C4PCc9
cWIZ7VotwvmqZmduTBBJKyUCH5+SkbvBHkuHoU/e7xlL2k67vb9M60DVDFH50dkI+H7DqkW7dvvA
AjsSzQyYNxiUliGRuy9XSthXheG/w/GXRZVpBzHbJlDTwowNbOQzaBGG2ET/yTJMcGgFQOo3fq2J
DNHgArazTn2jEjeLhJmUD8C82TnK2RLwtU8Tih9oot16wGmip1nbJliQJDr9YQzaOXQrSqhgNEvn
6XeqEANu7bWAnZDT5PmXHc3kHTBqYXSPntFss1DCctHIRqnorTSEHkBF3MPHifnmWuxoybw4Lvt9
zISIUJCSyBOjcbUMQvcdlDLLwVDtu6CJ866nwcvJGtww43SlKFwmNwDQcuL55HAf4n4t+0TYL1qO
sfVN0dRVBIgfA/L5cWAfY/01WHdLFnbkSzyVP9UmilLYvJFU7ixFiLs3NXeBjKCTh7DE0ULfMiVn
/A5DMBAW67+nIXapfQpAmzZM4XTykEHzXRQhJFv6EyVbwdanJYyXSlZl68aKmC2NveeZLfiOaeu0
G+i355LFMb1OTQdlU4eFPjx2bDI4lI0XXj4RfjpdtgKqg51dLRU33QScKF2cwqBbU7rbVDOIjhQx
ugOvSSN/IT28o8Cg2xBdq6VoF57ZQvGEArWxrCC0o9kbxgEv7kXBZYqKOUGtuLImYwjObfS2jb1n
PDJOeV75j6k7rJhsRkDgYImJ/jP/hK1EPYwv0wH90YMhy7KrvtCjhBGzROhTzQqhNr5J9nAcrYDk
gbxSl25rxGq2fHvMbt+5TmpjjBOtBLjQeN+7BNKjSsnwdoUvldfIS+LpmBzEvfjo+0V/0pHdyseZ
EHZPQuIH8DLlgGihwEdHnrmX3arng9nwcPyG8RolRLmqwU9qlnEWvk4Ajug2mMI9bBDcCfEy4aBO
P/wBaNkUHLxnvae0Trnqll9gAw9r0CETh7eM3ebmHWXumpWCy9LfMQaQr9UWJmqxYcZGmm4G1/jj
lyZjL8/yH9d8ZJ5E/MufajHuoFcfRMaLITp4UP0niUlBLTdtLfPYwO0Gyatjmq8N+FTmx4PMX/Ha
lHrzN3GOqsodspwWTNdzjU9rph5ZWtFglhLh0VbovzIoJDaaddcNFsqYuTVatQZ4SJMZsfr9qn87
X/VskummqAAineJUiBs87LQw3t4JRkZZVWA5NwPMJ+4tNdORAgTkPCdskD5P3TrT0Du3E5uiqe+N
qCYgdzg7AtuoUFRJ0ojO+qVF7UJ5ARKMvbwfWoGrE1PjFhaIL8BM7p335LFN1X2s3ksd6A3BMcUX
9jbhsEwWT+5+qjMneq/1kz9fMrXVuk4RuL9+FoNHEX1BbJiBUtgBbfLZv3mvlRJeQdMZ6iF8uX2B
DO9p/IJ6SxHWz+yCoY+DlDbEnL+Gg0O3E+1B6X14Sr3oM8rGufueM43aT6kKG2IBuhm2OnZtYUBv
UTps39el/b3jj3TRPjwRljyyLLrXQ1ydjbeYlfpZZ79xqW2ZubI2Q7addFgVRrgVlX6WW6qF428m
/r0trNbOMmzu/yWHso90lul/+SQrSHk5edzzS4f6q5n+++XhQGZfNvK7AcIlEViy605RMEihbrDm
vy2iqiEw/20tLoq7QYORu0wvTekONOxmu0IAZRDCVMTG1nPhB0oYC8HVGiQ3MgkNG3mGcMwP5mPR
plPnn7MmIrtf90zmNKefzWtsaeG7+R/K2bd8Su6A5+V3CSFuZ/A8EdaN6m2ep6Nhm7Y9q8y/rRQ9
/i4f0Ukr3vn4OlyNoLRQ1QtWR35S/t+nykZPeDGj3FNNt2fERDn+xpU22kCuBDSYIlLCQOWfP1QH
tjBaj4eHPpJGHc3kL30naxfo/aTo68+Y8bZOnDfzupLZbPtEL78JcsAtYrSnNTW5pzXHcUdePlUO
TrDqRZPbCjUk6o7Jf171JdW/bs2plqj56spp6AKWCCmgUD9YDJOC8+NXYCU15+GsqTYfC4DaQAuw
awEY9mJXoX/TZnEFACEJHoUOFQ//JoIXcpeAR1oBPs+yPJ8KpYM6lOxCIRvvm1jyg/pKgcnjK3VT
dh5U5HlMnNn74X/vBk90t5WvqW0NZ3P4BhTCrSpwFevYRnrUohqdwaPEJMQUS8S/sC4JJPyqU3cZ
cF/ysZP478K1wunVT1YvRJIuOPftGima809VUE7VDU8wbYr7y6R7WsqcWfKqbFL+j0frEEMvAVAb
t+dNrO2ByXyefNdYlRd7xgdgvEQ9guMNFy44vBqPBErblZq65YNyN8Ug0SMV+ko1W4sPkGikcm4/
dg3W/VxpXLXJifkoMuXBWi46YQ9ShrqNdf9DNnuRK84/jWxE/a4eMKqxW3ErEzzkn+MxFWhoLJ5v
wQn0xnQ28CwEBEoaVBKSoEujrvNTOIVNpfbg8u1NvRrHhpcsFRhGii7CLb+7DGwplD5jPTd9qN1T
aphAnnY8gLySuWqbhELcwrgR3UgkNWvLaydc8VY0CgaFq/21YWDF0v4ONxO6V6iLIBjcAJl1l3E/
opqnVvg9216fdeh5+nmlW0v0aeC3HHoMwr0edBNXgQFSWMvfZJnbgRLawwiihd+c8tajJ9gIBAnX
oPULhsnwzALYBxfBKiwZTN27ycDjFTrtuuU2pap73JqdISZSwbjcMJAzPtZ/LnrV8VYlgzI2g7dK
nJKx0NJhDr+r5UFBWYiu0f3hXntIuiSWbmnFrOEfDCUlj0B2b3LRy2qg99ybQ6EhKFAJvJP3egJS
H+xCAmQnG2oLM4chs9t7fl/b5PmjLe5sZUx/2tnPBs0RjWJYwcPek0lewDlOwXmrBzJ+kIvW3ULK
yIVS6/iON76NX281VmPG99iC+Wu+Hekb4p45toTL4ojTfk7ti2qwxFEimwVzcsAHaJWEtLZZajtS
XUJwI9T/c3fIJFav8ihvehO18zme0whbvXH+b8L0BQuhQpOy0+5cVATyAB1TCLp6yHMS4jdwz0Ic
Kyqo/Zw6eHbwbb9mpj7zuKqlE7XBZmEQ/oIuGvE3j4h/JqSOLLci/DBgxfFZ4Mhq35ceHGvJ0XeQ
0/+45PgonuI974Vr+m4B4ZtftPdeHT7ERzZ2F3uIzhyBT3M8WWhg9lc3GGNzWeUmECBdjZ2F8IME
EQfumxr5Tpf0VMmqeVWrB3pQU53bxIugJKBieqlxJVg0ALw2Wz0vfMhVq6sgx7iK991C2Zc8wWjP
tu5odqEsR9T2jADAg7bWKV0JWvhJZ7ZnF41y8XzCo4rr9SOngFpJFg4+MO03TfwzRVAzoUBFV8Ef
a68Oy/l5hU95rqo6hPEmL2Mr2bNRQQ+Lmzl2eOm09pGrx/jlvA58FZ+YL696q+/uJzwT1Xh3Czi7
3HZUeSFcnZ38bIgRp9EDGxcPJ13Rs9NyN2QMATchTV6ztE9jkml1FVkuI8Tbfe/G5c2wVcXP9/H9
lXjBqSGw8wdhB+rY8yQ7Yz7Bm36t3s1GS0Uz6xh7KjcptaobAH/whENht9aAHRybL2PEgJCxBDoH
AWpxGTZizYhSqghL1zNM4gR+gzAiGqLALS7cay5LTZXH0oYXCtLJKcC4tZjjyof3+oGPK+skvGfy
SXS7jE348p2uwaRU4/UBi01VJA0G7iAM7/K9N25JkdeVkGqxJ8crdKeYPmflYDuDJA0Ln/8kZyRG
Ii8ueGRePETdkwq1oDbuhwdJX9MFsGA0UUZurDfSoVk19xlKw+s2XtOcp8fIaPunrOIcjjsx15sv
CtoGYfmzkpCBKZaAQ+OCdzBXAmcYZun619eZ37P8wGdASwMkUgjIrKNMd6NKmghysbv+LpiIdVhq
FdIkigw6GuTqo33gnU/3+yMob1k4f/JshAbiXoo77XaFqhtggZJDVETZ9KtU36vGUi6TQBqa0Idb
Vw/OT7jVi4qS/vUREr9C4uV+DSw0j7r5QF27Buq82Ma+2MsfdHw4Sa+36SsIr/lxW9ojAuIFz/eF
Meq7iXst/pYlE1B9UBm6ybpO7INk/PfmkLUJf+khk2sajqsofl4cw8Twx89vv+fTU2+YMTOSseDf
KMgw2U2SmgAdrpuCgS6Z+f2bXIEyX1D1HZJwik0jPKbzGWITk2bdoIIEKT0WQAWEaUKenqzfNBta
EhYD0h/RxdrtNNS9yOZUJoJRUqVRH9D2t2HyOr/38OO4OFPVWQ2dwZ6PI3sSu1jWqEaqshZRXv37
JuaT7iD0p4K5KwaoYPEMe9WM+LlL5+OQucJHL2zHVnLCm1VXkOmdlmGeiE2VWNjQY2XjCi3pDub/
PLsetN3wrmI8fdyXqY/Qt43NTwcFOusqxYI30bm7SPLlJ85IytVdLu08G4Wa13EVBy1rReKpBVhv
X9JGBfRpG8l8Rn4xgOIVCB7a9OVc/mlvTbdp2CsX6mcUQMuVb0cyw+9Syoim5gAgy1sCMNUyKCE8
3uh12d2XbH2JQkKUKiBXQsOMZkI9v1TygJYm4myKeWxs114iI0eIC1wNDX8Q4lML/GaB6YFFCDAj
TQ8smOiKpFTtDR0tdytTaeX4imAmOUIjmEr/0w28m7kha5Pu3h3LkQFRHPTsl2pVmRaSBC7IgEr0
FKjaZta7SNYuTGnnj2WgmObuHSKk9FJrjFi06i6YHb8wG3HR6S3ZY8pdGzRJ26SaqTkbUnH/NjRp
2jcZtxfLVVnPJx8U6Wnv+AE6MyWpX1hw3lp0VI/gqiP1knCZ1Q6um2Gjow1SFwNJ4LADux3XaPFz
nzzeKJOO+uaOZTOp3JOLD9IJDaLd0LWIyeXVA2NNnVAXhG6u/ZwWSCLznhJFLS7W/aEk/lWmEWj7
w6Htfc2P8mpas3SNnQqtbFGWUSEu71yZQW+wZlO/VbN4lTSP6VHOCw6AdoebwZJzZzs51k8fdRRq
SclzUPyOfCqfMUg9hvnJ1BFgDrvtwb51KF6RlVvyeXcHSxk3C44uNmrlrB1NhlbZH2HkJ4fQBt5r
n0wU3X7F4sjmosbWW5Xx9PAXVg2ub8JVGe5CbPxdp5d7sOjmcttHF9hxriZdHhiNsIcEPXo6BRqr
e2fDR1gMG3PSKv8MIl/6vz2wlq0Zq5atoI1LZUohLHfb+qcQdevleWU44b2lqLeyQbDXkiIYBYe/
vruXY8kzhc8wGBelhXrCBQC68bNVcuIOQoa1S8bRFOkxZkc+zUFmdNShunDVIyQrdbkWjbUO60zZ
t/qcKCATEAwyzRc0Xt9riWRGiIUbdNcR5/ptl7Ugs4i/s/TnniK9sPgbuE3Eaw7uQfVY8tbOrcfk
E2qokQZcgyIyEr80Wba6SxtextW6b0dlZ6KbYbNXS/9Bv/GLQjb8uNU2tWJbhDYrk2Y0jjmk2uue
XDYpkRtbaxAKkR0PrDGiCSP+Yx34xyIiEDFcNT/CQcNkjUHZ8OScu30QYx9wP7rJnins8sNklq4u
lR/itptoDqvjB2YsjnlMtXi3B91JHFZD0c5nkW6oDTv59cKqFmIhUPLkaxnde7GkK9apm1GuO+E9
5OFunYIjWD/IcdXshxLzxorjvlXErpnytDoxncVyOmlxvQ+qdNd6kdEWYnAZ8oGxA1+OB0kJUqAA
Rn+H9OMFhA6fvCLwSSsPAioO1xCVHqEKvz5ApdiF7jrYFwwSRqWnwdekO63z6W3dEnUiQUBSFFZG
y6OIK/JzJtHoDuhLYIgRLZYUmr8TaZiajUagXuOPl1HRNwyHD/Q0ZXhgCHo3ZeYcAvZn/iOBQFVw
aK/hfCRDkDAZsh5n0hWaoUHaL5lpaGy8mO3lv2YNF0ctlF6fI/xalJXvsz9D8NTom0lKnU+SAvpQ
1URACrfe4CqEk0vsPSB/nqF/diCcfiWs5dBnGqifl6bTNzbjnnDlih6HtxLq0lWQ/7RLBKadt7Nv
11fyFNNWl9mw6c/bzCCdqBr0zrCYs0wiS2wnsLFTJ6ZZAXDbYYd1q61ePcUbcwIxVYIL6XpTInsn
zwbFT9E6CUvdGVC2m3Zd50a/Ygpk2IbQCIyUH2M7HXIFGlB+FkOmjLN8bd6DyK8Fd8CqwIwxwpTC
3hb4bQIUf+eihCwVvqY4XOWSFzZhDU7jTJlggyKhcPuDPMVj/2GIezxxCb0jlOa1kxfT3bs3gBIo
tQRLkmEReVA79XjeACfnRSVlFXm/jIpI4Ru6Ec1+HQsUpKbg9kUtJdX2TQWrXt0QdHP9v4CVt60u
nz+oWdwk4uhROGaLBg9qUm66FcIiy+37HU87hz5dndxd/2iaC2mVyAaqQtmWivxKAVbeabXS4tWq
aNgkKfL52Nzww+a2IDHnAHfc8zmm62OS0f56S/V2Aw02qHF63IW3Bd55z7pUNPCHCQ2sOC7Acj63
chiyHED01PSocP3iEG3wnr9udiFOEcxZptZd6cK7RiddkW5Q3HHqu6gT/erY/m4lKGykVsBwsE5H
6paOid/2xRymzGxcZyKMmun9TreBeGgHthY3p9bBKgBAk4OcLaIOVBgVvzPtSXF/vn5vpi9+eVnE
50PDjQcQKG/N28R6DXjHGBpLCrqsv+nvDCNEdouK9KXnkJ24y1k/Ksk8qQkdFV/Yx4ibUXESdGR8
iOqww5AB4H0et+G1MbhjdCSYhPKgiDRbRflJUEqGLnKSW68DcmB2O8XwJan1XOXD2mTCQPYbxu68
ax5QwCInF3zRL39W2A3GqoKuQjV3IL/wcrL2WkTiUwPw5dLYsJVcKFPe8JOKPVh57mN4gBZfs7RD
Z3G6Fz7ahtKRFE5RA1CJ5vO3/fZEUIHFAaTjeDhfjEIz+y0cbuP29ownIaqGaN7Gd3VIukf3T4I9
wPo2VDJoSRobXY60/eU0Rf6W6Rnfig4MtoEnIrkTC6Rhov1jXzv2C+ecnfVvFn1TcCJ2utQD/n9N
d8nQTIW/HCEv53MogRI9OhSxssmhXlI8loL4Lmc0c4oHR3Renu+IDl7r45ngvfk87YqoKW6YrjYp
Afwqhm6M1l7ZM9/KcfpyNKT9yaTmekfG+ZE4+Je7K7aOBiCGqN+OJnJ28AGWmZSOoxPgJZmJg0c4
GacgTH0jNA9EYd5v40a/nNobI9XOincY4etdeUzUiIdufgLgXFZK7wKrNxm3wBjxSGP6sEaE+4wO
cb8kfo0OVE4tTpk/hqdEi1mF//TPN1fIPSQtkixqv5FmwRevDhvPP8rWPdMOIRK0n7YgVOVgd4bD
O6pjS7PZWv+19S3SmF8VO650cUrPhjZHgq+RJRq+FHeq1VGLGN6uDABpYpOkQyuJ5vdsG6JjEeJj
mS7e3VVMkx/XVbcBnoJcfKe1ji6NZorESuPMIBXMqo7ViBrxoS/T8Jh/8Fp/P4l17d4uoBY6ufAo
ZHycfxjsEBjrPKC9jzibccnX4NAHdf7cJRQO4hhBrOLaDTCNR2itWxjRRlX4CwkXFQLbGDM5PsWN
KGWVREYt5uFzP1qyJPIDwIXPOlmCDF50ImAL2FrcVvaXJ8rYscOFKtTHWk0+gELUemqcYZfnzmP8
jTB3Tp74FNg1uLOF/Q+lFJh17CHAcIbcTlHjx8sXmE6tA4qkc0YyXktkMtKFmYMfOFQRfwckOfGU
FbySCDigzZMLjU1Ah5mYjFhYNEhA9bBVrPq3bPDW6M9/EG5XprrKOHJsyMxcrt0kfTZLjQ3gC3gn
Rp5sJSTz6iJL0QnitQL3BNgJCHvCnZUq44ZooO9Gt1uhU0zmO8w14LAGdrNnfhs68bNnXWUq8zxd
o9jGZ4KdpFh7pOK/Rgqq0TZJUjoiqS4C4uTvdxEMKp19fClDj9+FOoiREpm0n6O5z8zO+RLX01nj
ZTtd+E773BF3ZrP/P810aEiC2aRM4izaLxplSI5u2TRkk1ReHOlbaOhKsaPiQ3SSdKmQ9dZbsrjE
T2QbI9oqVmOHA/3kZegwa+fkESRegzIOtiFBswitbNsBxpcx8jv29GlfExoun2Ldn6qoyK9rrHnl
4o/mPV4al95eQBymxONMKWvPCxVYgjzIAxdD3/3xLjsSNK4gmdT3Pl/42847caBlufI6pju+6dg1
VhSgjcwBytDLZGTrPyx3mz/45ciNZTy5bGDnebyAtrfsTCKFKcUCgCL5vb2eJC7uuEmkVJPFeIvE
UsRNK7nGYqwdTw7lMDaDA9vlNA4pW/fDDD0UTIIrTmKh7GQJ+s8wXfSpRYpRfM3Sbi1xb1LAbRZ9
0ze+7fdqtxsdlSjR7OwcoxZGaDIhBV4P4zKaROd3PbnZu7gkTNfezKXk3UPHpwxFifJ/q0CcoWug
ZWIGuVpRu8NpWrNAL4PLVY2wDIh/vmq04/fmTK8BOhEuZ7ZURRcSCGjYAeQX/CxmnEly6sE4WOOO
2RBdcwlQUOm5rqLPvOJ4+K9Za5ih3pVdL7bBBjvTW46NIyad/O16OkKSuGdMAXqio/w9yUaVB9PB
15UHjptVwgKWuCy5yAeJeta4S7h/ZRadh6ZhZDGexJr55zttC00aMj+q6GcW8TUxWnSZnWWHnF0F
HRqqo8jc8kQNiDe/BM9WaMyeEe8FY5IoKhXtHcl6vqpM1kLe8xuJPW0Wg8gIYYmqwHKxuoOaRPAT
SyAvVifUaMD6VZ14yQnahFnTy0bWXaahwB5TczMW8Yae+X6HmawkeR1XZ7XVEs42abtK7lYsuacK
w4DeUqHN2mQS+w3pHqM1zNane/MXMbhvjp0g5Wvwmmoi8bH1WyYXWT6ud5gTVwUwiQoZlwBzyO85
h50RjXK4yOGEEfaVeDpeOpnsJQFh1piJ36ViAoCSU2b7fZ2PFpiLg3YnygmDbaxMN1LO/83kpAx1
b1OEx70tL0EReL6EWxqrvSbO1PR1wThJ9X0bOnWNwwDxhq1Vg7lUV2XkYbgXLtip2CyIrh3i6Cyp
s7RqAtH7Twd2w+jq24mECYL4HuVZiXfi6kf3mk1wdNJlfW99PrbNYedZfN5wkI8UfiB90N2nrka4
NsLTKJ4QpVdmrfS4MFkyX6dicjcR7wPI02tdNQGVwoAtzUdwpOK0N5h8qqwkrjj+AiONzvkZafdF
El6gbVv2Gahiq1aD6qDx5isZTcsB6Aew61WPUuXdfnp6BN2QnYtvEExM6YxkDFtuFTVOU1myM13p
+QMIxZLA2sPFipI6iVwn19+Gcg+wNE7fM/9r19/7BtpSO/f8GdDLtRcj2Cs6J6klc3PiAocBetqJ
tCNvBTtjNmVs+dSXml/5b4SVePwQzedT5qUhHQk89YZO9kUFhu8Mkz/TTxL2e1VCpPccS+1kq8Zl
37XC7UpC/VCuTNvklGWfi5NsSNOowJ0xNWKm+N8oyShvX20P0JEIrG8RRX2mEToYnWFqTeYbjhY+
13/ZtaDC2GUNUOZjxR3Z7BX3yiHlY2U6MArvNjQ2a5Ovwyr5/h42vC7vOA2LH5uYTupnNcFQfkre
Qt23FTgZhx6T7YMHfYUb5BwLbnkBazB1g4VbgDfttfaeOf6/8WfoNAg0feQY9Vvf+ntI6DXlgkBA
vS7q63Z9ZZpwq6tdEccpuFqianAQemESyVqSAQ8YSEsxjvccIBFstww/4jrVDIWfRiGTWpoF3v+P
M9VePq1anbdqO4/Z44wDGkBsTKrooePf73szXeKfKtu10nWkP4ReXGpU6nhnqWinXKDPNBEljL6w
5bsKm8ooxswGj3YETZFlVFh5OI6Dy63DtWT9DZfnZcD9s7ROJf/EpEqrjd4tvDG/VAZ1avHYLmeB
qzUhrG8l5pcrCXWsm3eQM2vyvYD9i2ozpuKm6DMYWJAJXmUCmxarHtDfOK0x2K9ag1wvFezoDkoe
lh59PKbDnlBIT+CBsHq07rDY5TS2NyD64ejtOdB2MbHo2HfoN6jOw3uP2pA4jp4gf3fDYeZbryG6
CmCR81dHZQ0lOEQ6XkNACzEZh5c1caKTM1pPy7xFHcyj9q7aXwURIWSrW5Qcj8Waot62ZDGAL1+x
MBPOJ0EM1VAAxQ9vg3lrApkYitg+BCDZruxVkOaKQZRyp0Us/TMfekJ5vmEMbCxuvsyPHbJXqgyF
lhlZlzcZlObcVADzq4OiMB8WLw7C8GmbhHLZ7LxGcB7GVIoIN4dSgUewnmO6oERKAjgjcYVnNe3w
205rMXVqnI7EJSDc3iVnqUoolZEnnoMyWJ8B7Lndu4cg45YT0pJYQK5yA1nv5H5bJt3UeqbFnRYN
i7/Mg/Z5d43Qn1NUBhVHD/0ypYCYX8yBY7nH6rdhmkwQIYNEP1MymSSnCc2A+zkM0+oysFOO5kNC
xN5P6ag2/ZU0yKiuEJgzW2nCBD5js7fWteGF9BkTifv0palRSMBQJY5fl0gptMPCoz25iKLg6Wdf
Xntv5yKPMoPeoruwF6voXyCrckBcxeoWxnTDObFmCtT4Q62nWPsT9aS6dG1FBDN9scmZ5JkljqMv
KNSQpZqgL7XtuvGAYz38eYeYDaPShG3Y5sego1xRVM5vTk70Y+j+hZK4KCJvx9R2Agwh9XfmzIUH
2RJBQSCMI3GE/t/YfnNhVTRThmggv4eWLI+/7QG8iWcMh9p0E2Q3KsiIku4Pxj52KnXRB/9trvjE
XmsCCvJqSZdd0m1jPYlf+fzMQ2tcpQyGhsT+zKpMDEe7+WjiGZMwzD9hFtfmdTBMx8zyJZbwd/tk
WaPZU0BVFMjvRli+vUSamb/O8Ezne32J9mTjG3fk658CfHjNOs7r+S+dlUp3fUE6HaHZV13T0KOM
ES9xMAmj8XCBJzCcqW7sgdC0VffxoYeGx4czrOTYETxexw4TnSRIH72+P6XjIICanARTg0TSgcsx
Qy+RSe5WTkMrGEs6ZKISGa+mvpecTLb9bu6CAkTQ1DFBagvh5N9Fo76A2kzOVj5XtH74QmZSO1s0
ojCIUgyw6qT7EoafqWhYoiWHlWHGDjY6DwAMjzUaJVoB+kxQGtOM0xDzSm2oOoz3RydYwyMUmpk4
uxGj0OLqSCQGysrZxTlJjN5rnB1rmSU2MLwjRLGF8P5NF7Z6OLkjQz8iXCUMnpciSwjbQ1INnk72
kiKTRmXrbQkWrQ0oFXUX4EXflybNdef8ZryIcwoj6AWDwUjBpYrMV0LcIhJMUM0sqZVc+uScZzLU
upS2zBUjicgCjOROljnlnw9kPuTT/KNzI/UNQ3m6PIe0PXMMwlmqqeYp84zgnkDyHsm8hN4FH7+f
+FLwtVF12rQI/amjtWZe+B9T11fsST+34UzojZAnBcqRP5BufG905TGka+LsDNdL8TWfNKdb0ijN
2vm6hAz6O/hiJFoCLDQbCICixPVV2mjmQj1Nbs8/x1ZXiGkRTgp1Iq8AxiQ8+lJUwetH5if3wDu+
KsM5pby+EXWF5mk15wit3sAToBowObNmgpajNXFXzLI6+uGThVsERigu8F38Ul9UOcLhmbO7Lu3C
FwVjlL2857gz75euOd+GpDkyGS61XuuNP/ifUUyOOn0edVc9zx/wg3Ib/grZLuYj29hr8A2MVczC
oCx6UDVGFV1U67GrYIBOwUnNzSxc2LncuBkUD6dcvIXVM/LGHX5An6iMzdZC2C12CDwvZi2Q2xlu
DfMjTApNFaGvhD0uPJYyOFoUO0cGRK2lewx6ZozTVCZboDJxrH6h0bsW+SnxyB08noRUHaTIFkDN
ywQE/rzPX83vQZeGlgm86zHDRH6mU5Dh3H3HdQJFHlvTLOPqIfR4P/LsmaS0CKtEET56qRZg0/uS
ydI21Vddpq/R3flb72oGw+WZ/M+/SatOM/PADP5NlhbIyRhb8n/mVtvSh7Is2mT9epAcijJy2LUk
NMZJYyo/m0ELFS4rNsN7WPEKapCSJuPAjEuqvDtVRf50B+VxBq/70s8VtvZfSnznAAlYtSkMAu8B
keMDUDeXnY7cBUUjPzQ/b8WUJAChWP1A9o41Hf2b/CnSzAWDNjRxA48aUq0xkFsqEkspITl5jx1I
nS2TxJq5mLuX6aRPn0PoV2Bl2UEa4v7exrpSBnDqP0yZ1Dbcos8DSpTwEHNndR2cc4rn4+iFlWaP
EGJEHw3cUY4e1upxFhaYd6P5EBILC+D+FX3obEKxyLClGPYn6hbiZh/Dlj80iv+Wsak27HLxVKE2
Z9WlP/uQL1QDPave18aDyUGavbT2HLOtNbUGG1CyrsSKIxTMulbcWKZue0pQJRcKM9m0EGFwy2xV
Uvz+XUZwYapN8uz3FPwRpWdGB3kw2YqJN09nOGfbdE4aV5M72wFf8mDZQdIp5PFZu3yO5DqAeWjG
bRhxQ48txyoKrzfiS86L1amKWxrZe6OH+SaqbcBuhFG1OxPKD9P2P9hJM8veQE9UtYUcgSD3alQj
FtJb/10X7Ay7KGOrIxyBlREmsKboiH+QjTl/cKkumThKQyolFMvzu/6nCp+7hGUhMXsNu2FCBoi1
sQsFRaExdDgQIvY1u2roBaMI54zpLqvwpEU0LDpOtZ3n89oRhafRTgH12b8yu4TYt2zIpAd7c6Tg
be0Hch/oDGFzOeJaSqeMfQs4mZwSgsyNWxmUj/ALfveig3WA+acJDkUcGVAOvOIacCR862NybV1q
bbAQtkwiJspP+OeEK/ARhkOWuzvlWqgXlYxsHdYQlIEColILDaT0F0VpdquoIQE4m7OobQje1vnh
CHKNdjAYjN/4BXikoZ5L69Jokv/JORLjZitXFYzmtcMF07txNYg4UW57uful1mk1Z8O5bpkKkkCM
xX+ZJrdlNpGbyPPiqjqihyNQEPOoYujYJW8B7LEd2MNNtGk3mQkYS7WOcgNBONEXzjVz9T/fHmT1
7Sp8qr6cBOIfb0ZogT4+W8orfM7o/tjwdgjs1o3bwEQhnbNRTdqxJOQVDgLHtVtQ8QBj0BON7UFi
BNrkbvYIKYYe91XMcWQSjgrqbaytlBMfVG5GaYfJEbBUqd+ZK/XLt7naFJDJcxmO8mL0KtuEhGyz
f4ber3OgCkLjotQcPYKV/tBLZifK5Tfkg+auA6/u+I4AlBK+YzCXKFfB8GKxFMzmzi6pm+MZYVSm
8DctXXrdtKwKonGeYluR5FEsiKOYwH5vgcZbDp/Hwv3dd4Rg/krCycteNcr550ZhsnEmdRBZVjQm
Q6DAvPcwMdkRH34WcZfYWAI6DcIBCoWXQRG2Tiy2pIvJFinY7CtGO30BGHlOYMUx2C8QDbYuka+/
1ZKS1pgQZOr0u5lh1MGYaORGz0HFItSFThLYo+x4t/pVybYxDELZQFT6xijwmXvCNBqgxSEW1HDC
VaAkK5GIcFIIVNNvJzlGWhSseKEMnrcraSXX2KlZpBw5rzNRB5RfnLhMXGxWEhILS3zRfAVp8CgH
qPC2WPjVtDHKRx1mv1mXcwB9vxlfARs2f46BugnGqWW3UTBMEaCTTav0q28DoG0S10pNAAOfbP40
DKO3bsL1mwqAiuVpMAIKXXgQ3RQkv35eQ1fsO06NCmsqwRZgWMj8PmX5msNFu/phnbS0YF8pcaw0
g4Z3mMQnbDASQ7VsUjALOzyVGHNcMXoHQweCRez50Ms/9BbDlqnBpvMEIBfX6Aj3kXKRUETmmAOc
aDGZ8C9+o6g5ylRVCD30DDH5jWpfwQIorMKp4taiEjV/hunhv0T97K5Tk8JItbERVBNBjTL0Z3x2
esVvAsQiPUVFlEXMoDABiWXIWzJECArc2PTljqfmKTsLoGcwn9GSUASHRRpD9Hn5tkymDkHPFjHU
X4tl286gFE2JjPJv/lqUwk5sZR3J/PvZ5rYwbKLxR6p5p0YGGwLGudFIcoippfsnHxo/aZbTSwr0
e7G772mqyPZhDT8RqMlEtppwhhXNJujQwHCQ3K4xadRWTg2zJpUW+Jak1i+o6gL/PFZ9Ucv689lb
0AghpbB6R5I6ySKp4GjvQ2v7zWKZgtr05oNIAM9rGJ1qqebDha4ijiOK3zFdS+NvtmN/IE3uns6Z
vJTkCKK8MVC0YLzvi6qH2cEzoo+laldfdbfbbtrWTpNriyo7DI2EtMz7zyRE/d6VRQrZgeMgrSDI
nU6qvdclWyZ4g7rXGpaobRJFXjLpJ2MZT9h02YcUXAqbNKqzoxHlct9g6XxJKBGBXZJ1IT+zfJkm
fQydzEqr2OQcMGOCs4TO3Gc4a44flUKl03tm3J/n1DlY+3PlIaO91RdhTns6wOePCTYHMNeyeFGw
KvCFYb+1duIsMFuULTlYj+hJ44W7Rd0ldVUxbP+eCjY6CdZuZYminEy8jnu5uRR/D6pVQDMjKaHb
9tLFjpwjMpZEgTa/HndVmobhUPDuViKHTak+2JcFAANkSXsklq1DOtGDk1FFHTcIwpS/L4aT90ip
ePxGzXDqtFvjgx4J7rvmWBxnKXptiah5cwmccZhERM0l0b8O0GXnsHm7ECmiaccc6mlrPyKD51J8
wZIjjLun8GiHh+Okjw0IZT1BMB5qSeS2oK7bG/haXx2aqnlmY9q6hHqbTsHV0vDvOnkFCWdkeZzh
JWVFnSXGV/weZmLwPQr7evKrcTcBBcQASLUyPCwOZvqU5f4LEvoRyH/EzbgcjMEfI3bpkiFfPWF4
IvA7z23g1oTXP6sx4/xOkwYWXlx8ul/zrmcHJCDOgqZgt8VsirywNDBfQSKibZnblC8SNtj9jEKQ
FKfCKihiYBthLjjT3QIYCGCwqKsOWZGMPHwF372+VtbGiYQVxJFRy4pgIJOCPpi/x3DcNMlHRHF8
Fbx9j0LOIZp+Sr0BkTJcDL5siIIRaaArfZ+JJ+WoTEqJMWBPvlikwkQu0Moj+gphqjhS0Y+Rgxeu
RbdS5sitofjXt4XJFpI8pxC63pdRgmA1Xu1IJ6Il7ChIRrtBNSvoTdnv0GK124wcbMgsxOMP1agT
292r1kmmSna6XeJBFvzNUxhpGrwkndO80VDJOEmIlvgdylZ1iJaR4p+gIf58AWsP1Uc4LC59GAK1
0XABoOha203sWhYx/GVPi5CPiuF08sS/zrmCHRB/rPK3GnZc2Pm1WxpF1gugYkeKcjltPdQ03Pgg
DHpNSjlY94BxgtQ7EeA2GQB/lc5RXX0ES+rZaH08NClZ9TvC/xGI9XxbicczWPyaIvm2AIJhIbtv
+jXD8ln/R+MHxe93Zxcw9OSieq7HyqpuJHiu40SshE8ico/w8I8aNWyFDnr5+ThSBYogLP6Stlhd
vROTEOY2WEcSBlCTbUmvwqdeQCv5aRlgnlHg78Sk8Pc4H0Eqi803dkwgtQxf+QIST0/2wPMTShDw
ZDEuXNoIiiPtOiQhXDn7Y17NDDN9qWDUxigSc8W0Ww/zoPgYM5ZSfjlOEN373WutWwg3MpmDjKxU
g75UMOmYuiW4Wk34P8BIYGxUfA8YDzmEPocK4xxByMEJPwdOBLJZojVBGkhjmy0kyVvnYC08R1Mi
+CZ24kUaF2r7sz3hIDJbKKgzRmYkW9zEIEK/FNpQtt7+J2dql36qARChwdBpV0ymyckwg3EyW5Fi
g62KCNaPAQItq9DWhGRL/RX7fnLvRxyb5WC/yK3SujsajSOpcys31s2YQGjagXq/G2Sq4LgVhWFi
d+W6/nbXp8X1GajPD04PPz2IycXzL3Bqpplq0rZ58kqOUF9JG6HPlwtqXz+rjZNHWTbgAuti/4Ky
NZp0e89APUCj10Cl7HXBfZjJif+t8osdSXWaFucsFQOXSXaZ292nTeGiOCBY6kFhW/iMn482u6e0
lnqpco7FccQ182tFoGdzlijOTWXsEamlYnTfPnJ+FdyupfcgJ3v03wFvS49O/RthTZBhJKhGsodx
JFQYWEww/sBD3pBkBQh++G6xt7LXgNfz5Mn0W2hk1BHdr7alYVOlh5TAEfoD2InXmUWXFgIK6ZxN
jaBCOTSEU8xsXKkfMzDAn1Rt6tpUnL9RnADgOT04OD+oHdNyG7n3IB3p4YlDY/yTLCnv81pzvcAt
/1KFFCPGxEggzrIwxBZIptTYWC4CBeRLtGGOQcVETdMWF7KKBdRtLqbqofHGNas/2gRcfi/hA0tb
6XZMX9ndCoFZQsRyVHzxr5WU8A2ZjMHhHcmou/9dm9M/C5nB/yJWl52HRM1ZVP87Y1Y++sKWWmTr
efurOQrMM7Yp0/K384e7Ejdm0I0XpAa0QXG0i+2kGv+DJyndKw4lCIb2W/qoUMItY9MlBMXCU2hT
JbqI4EG/xdUZ4RETCG+g99en7+bsDx7XMhtZLUwYYJ07M6QqJkqID8VMRoDtwkp+KUrBs5fk4ON7
goecjF9Eu28jfs8x6XfXu76lIEZTnq1lODr70EtqjhuGeXOcMOHH6r7NKUdLruQz500M5PQDVsLF
YRY5asks/rqCwdNj18VQ3wH765yL4I/WqeTHyyfy9eGFHrL7YthiJCdAN3q5gTgvjKAY8alvcmq2
aNIzCtTfKPET18mVzDxvdV8fsvJVfq22A3Td/vGtIxYU5HWphLoD80j/wdIRUlB5zvueDzjdpxR+
8fXnWwQ2uoqGCvNtyvr5+VLSTjFDJaNZo2N7W6YLJDD4IgiKwpnp3W2lF8+ZkDuoI09jMeUv1w/6
00vhLAjtoRjwl2um3e6KXGmye2cvqIft+uNJIJMiOfA3STHoKNQzwaQxf4ywNq4lFJ9mk6KCPRlh
ai5qKxxMZ945UOV7tXMAhS7oi63SVyWlbnDg1MWypDBsho6Lu4LBTu01me0uiGoJDuBRvfmhdTog
w3QJSi63YNFd1bY5sTW8M0NixYRdBUS6wNnULgdzokt6j/e/M6uWiLS8fZshDzhEgxn3bQpySyT7
CPp52K+VOBu21FQ/P2A4sww8u+niWLkTEASRTRllDTbu15P3PsObxz5LTrNFJ4jhEvVCG872N+T7
irf7PjJup4sS+6RfjO6qseQL/eDlLjkesKrre19acjqtlHsjiBpuWzXy8jXeJa1cmWCRMeCOCUx4
xAJmI0Jv3xwojXWUtYpvkCgzZBrJ+n/Fn/yj0qefy0/CUkmrE00oi4qQjGdksAAdXMw3Br/oHOqS
veJVxdKvTnG/xim6o/nCqX4sYbfksIh8/Chn4u1+9SxX11diY67pbi4upmkSX0HHCVViqQyKtHJ6
72emqA6LvHZyk6xGFVFvxErUAqirvMd6mlb4+reJOroshvmOGLCWUgsCE5WNqJCQLdtE0GdCF2sd
J6B4E2r5H3eaJzC5HWrZLdzl12nocz7UCUzAPEv00BbFFRnTLRFS/u7pSq2wt78cgM9eoR/vv3Co
bjjPy6kAWo1kWOHs+9hljpk/i+JbWt4VXNWL/RIWChllMZVXpXXdFxDO1fgwBBdCa5HlKoLFit5g
1pu3mPj0oNUAX9681XkfyxzYQnbqTEBE6mtX9UYigI4jkrHsx573eW1zvLdVyhWteBL9/FvrEDSG
CdeNC+T4ES/CqgM/WdPXC9RU5MiwMm+o5/kwnm2V1rkdsu1QxP6TrcxWi0fxbYYh2BjnMc965VvA
mZMJvnegWjGNXd2IFg2j1c/9hkHc+NqkFQdq0vG/z9eK3vVwOitY76wx5CAKEBdhQjk47R8feRYP
oD6W4zPFmjfonIvbseOG8lG41n1oJBC5tCmT6v5SCvPc39vQsRiiR1kr+bLxQDN0S29iAc+Bo6hq
aePk4YopiCcc72fHxvtHAVJ5ZCnZfkWCMem50rckr8zlD9oE59r4A/ZlR3JsZcE+MvaHRv5l1i2l
f86kFQ+Dobd5Qy0HtKTPJNEOq94CVqfe6aE9iZNLIaKGuRLO65aEnVQ0blONCmKNxKOYO3vJ8vpQ
HSyuZxHWDBkw+5e3qcmEi0D3zSeOdwLIej3fSDMdB5hYEBBdwkn63sYbQ3z+LkOSrnEW7/z0W1HE
/29q0p70fYlG05t8h0BmAsvvw7wjCwDERRYP7N5lBF/5WJXPO8RHBAWnYf334Y4NS1KXPGGajtyS
V/daxIvJsME4VbFXMV4CMGg4/QwBYo0+7zfEnVx15Ed3v9mwYt1vt5c1A6R3e8DMF/j6JYjxlogF
jBfkgORudKwSp9bDEgDFOF7j0YZnZE3MUL5mwmBpS3uFvz2XbQSPIn3ReKuH0WlUvIGRNapY24MO
cOIQ5nBSwbswsrXpBHvflPbauqp229lCvLAnEDIcedD8T7Thm/JVt0PmOVOeTXyWJCVIiLRlbK2b
tqVJ1lOS77TJlyJwyvoeURDM+H+H9UqD+pIw1rWjz+/iTT9QAsQPbAx51h1Fv3NTPrwvyL8yiSoI
zn351ESPlvAGm/dy9FuCtKBGmuee2wkVW6+TOrQZfH3q24B8NxpvlX+vM2YQ3i1UB1v1eOMPoOKY
56cNrdWQRHazBqNi9jij/YCtqGcp7RWvnLbZipyIqMT4mazyj5nfw5x8PDap0NgDrqz4lRndwCow
WUqcbn/QDo3/l/9JX+bOoKQVO5n2wSt7Zi97qAoUJGcma0hp7Te+Qzycr5yKnYBdbAWQ2Vmz97Q/
O+Heh+BRaNhFywxj/D4osZXmU96kJnCMJ7qdSnOBFo1U42zD1bdI0QB8VvglYiu/N1Ic1GBw39PK
aeKbWElqGrDTsTAQLWSo7YjJ2QeHs8JbSHEeqNIDVrS2pO8L/tJez89+VJmvSsEk871j1ClzLS7Z
N7tBEWNJ0iULiLa8FtPrK7onTWbT87fLjWNO1h84keFJfNvs6SfWBUL0E7tlMpl9A3Ie9aAmB6Fw
5a+EtvC4VgQR4cVQ5tA7IcAXBobLg8tw6TPIEqWrcTlupq4oMwADIMiT5ez2oz6SxxfVipavoxSL
RmIr5D064yfe1ix9jzgvYK7py90OvlrXHzy98EFudLXG5z6PqRnZEIhMx1kQhxEgXjW08uD9o45+
CIqa52ihJq9IskfCZKSq7iarGNdsRAvn5XVniG2CwPjRmjjFKSKErtTkR8yGpSo3RWX7qHBbN80P
Dh4CiH373BSMimX3+Ezpg+5v9ug+/LZxHp3HSLzhWMIB2zyd+SMNIl7+wWCiPOT1BBstSoxVzsyI
TZhSaMGdOeWDE4rmzfit88PtNbUygvgBZi4GD4SsWiKQkGbRtVENVWMNhe1o3yboaJWSmRC5365o
HOlXaerM/rPa/tWe1IBBoGYloDE1m9JeRuRz67aL7tuLAhIrZSxCuuNVR1GaQ7ZNSOuHVNmRTBwO
kKwam4sqMzVgiDdvPYU5rWSQRO8vV4JDs5SginrSk98AStLPWP+EoGS46MkaJexhE6yDNWmm+u0v
wJRoT2CB+Vi7ppatmMvX3zUAUO/+qnd5IVJ3NqFA5yMG6mRMZPzPdg1onTtH+Je4qmqFUIaNuQE7
WYsYNHILRrBdwraRPEIGfBpvObQWiGnpEHXUD35zDr9OLXQm7XiB+RbxaiBbIBQ6WEwU7ugHaiDR
5MjCoq9ioSn2f4WKe0cd8iNMFOMSMY/5qHArmgnzrVsppREOLcBWzlvbpCE9Je7L1dGXCMNqyQ4n
dyBnJg4fILDSGw3LP4Q8EHfq8U8uqfX296/oMKd8pPFie9cUO+zh/KaKTBpMM8ztlK56XxE4L21j
CCXTyCmxlpdCEyBXvy1Zow5KpmNIIJZLbd97y6X0aqboV8TNzSZ0Z3fB9vW89/JcIiIYqv8WppIx
Euh5K9HoYqQNgyM1nPxrU1C3JWGumu1GSxY6zuzXwivR3pTVAkdTDV0BCBJf1PAujD2nE0prWPE+
m2VvfSoYbWDAkIUIHKjCY7KYrR1NSltsl4XRfxiGobHBT6cKHT3Fs36MasP4AHUQSU1t7/ye/kca
9H+g1JT0xndildTIp22JAxl+vYyMH23/SNLJXPDq5UWgNraCnDp14lrgmYIX7hHnpwqbbiLGKrGw
ncdZrAUGC9EX92zW+x3jnM82TodbVoGMbtqbcD72I0zVvH7c3R//IQ==
`pragma protect end_protected
