// Amazon FPGA Hardware Development Kit
//
// Copyright 2016 Amazon.com, Inc. or its affiliates. All Rights Reserved.
//
// Licensed under the Amazon Software License (the "License"). You may not use
// this file except in compliance with the License. A copy of the License is
// located at
//
//    http://aws.amazon.com/asl/
//
// or in the "license" file accompanying this file. This file is distributed on
// an "AS IS" BASIS, WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, express or
// implied. See the License for the specific language governing permissions and
// limitations under the License.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
KkxEMvkzGr7TWvgb+DdrxziVEO40SqBS+n4ISOO474lTZ3gCsx532R6xfk1G0aRP5iJlKbfQwhyq
Z8IGnsq4A5sF8SkIywH6a1J3m359q0h5aKoNqjAsnx40oLBB0oNl7so+09yNBJhiIFHGxX2QUNGZ
gxyXZobloMDJcWZadvfoaTBIlFBMJvU9dPpsVLnrkV9VVooKQPy3UZHP1U9rt24SUDZw0ivYZJn8
qoIPyA7G+nLAHpv4MhJ+X4Zif0Cer3i1kzeovIaK44a/iUroecQijLjg1/P9P+roYSM3pZxLTpRs
crcc1qNZ8u1hWY0v03Ra4tFy0UcNxsaZZmLUzA==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
mQnPC80m1yjlMgU+XKJ7eH3iJpFUSRMIheQhree+rm4/VAyodjiwzc6ViY5+CCoFAzwfUTuzYDOn
sMCRmow4kuqnD/uCZtlABYjk5669MnJQccs2/u8lRqhIBRb4cgGn0Iv4rXZhiI0Ze7afM1W687ok
C9n5GCYCTr929izfZO8=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
SXAXvM+hez0pqTLP/Lnhglb0NIdaCJs0MMnk5P+kM9gmjghSTgqcusbB5TbdXWaBQMd1jRD8Sbyf
CZXZODnFBKdYH3UVyDjrlvVw7AvCt4HP0EJ/GAo6mIkO9ToXQ1fkU+DEe1wSf8M6EhvBpG0LQHq7
IU6wzCibQyxUXemUMKk=

`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
dZKhXPqB2VNqilvBxdUZ9MunW52mDULkkgS/vdz+N3G3l8SMatbfoOVpiP+Z8tJPP9T38l4VRIYl
Uoa5/20VGQ==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6304)
`pragma protect data_block
q5Km+rZAsjhuUqEqgTW35o8CEutXpaCUCc7eKCimy/PjgaF0E8LJkVK9+H7YpAf9s206ymi7QqOZ
W/FaZHw0YakUyAFLUQxj4zXb+3IffZpM+C77Krb2JDh/Y6L6npyghnGL+D+E2HSluuJads9zm7Pd
tF0m2nAgA5MU+LPTy55H09JmbuudQdES4w3iuKJ9vyTermlYtdzeA3MUC5LaNKwJxWPxK20oKDKe
Yk6xARe+k9/B0dY127QsK009LoUhlhDjiAYoO4V5N0/37LdiINyvjeNcRu8v+KXxrrWnGpQ+4EhR
Pak9yKM1EXC517FwiyzWvEMLQp7pLOtDVb2DpxYU1O5fPVEzYhg+owRjxWQMDJvCd93aQyIqv2lL
204YCEMmmeeudcadwzvVxZ81T2tG8OQFhsyAHZLfFetEnoCAUdKdT2rn7gCFOBLzht9/GeS6cghI
rQ9DmMv03jX+SekzIVcLRDulZkIkyqcR5fXbyEmwjf9FQYDa9nRDBzQsRFB7FyTjVVurw1x/lzDm
HIrdgL+zsVp0X03wH5jRz3pWKNU8xHabXlp84bhq/jX9LHQhbd7i26IxQngofym2MXdHPuic+40F
Aen65y+GCQe/Uh7HqKILknSUmvil3X4eaOEiiLNDtgEw813W38s6BkT0Q/T19bJ7Pqdw/xGN6cnH
eombPxpJl1qndi5cNO6j0N1Xfq+0QkYKrBsRAEVap9WVF3j+AH6AsNbzZBC/ZrMaF5gvQwK+O0Sw
c7g+rPj+d9pHlDV+UICXtKltVSa7eNsNctbp9Fe392AH0B/GHMN6JVLh9i6GG+UJP3aYgXj92Xeo
uo3xjhEOxClW8WmG93Q4MFwGp7Hw0jkhUoFWYWMlFnps2szWxCrqOVahtb92I/OaMaGWuhBlaARD
sZQ9Rgy5fPCZrqBXzb8z5Qd+L0F2Jsi42KywSu4XnJ0HjqBl/spUAa8jT2eK57EQ43AfscF8K449
TxGNqyoaXJJUn9mJgmyKRTkxwpz2UOsfdcGitbV/JYkPPjZqBYA0Dun/AVeT8Pn2y+sPsDb+nUu4
/UlGHCnEV9JtJaZID8wmrjlLEB3xGlx98KaRmliopb342whZbSsGltQ4RmizeMMqxpWl+nqzgc0d
z0Lz3bzNtxGEWCSNK212+Q/4E2vjCfwS63vkfg4s2s6dGDMcF2Hwck9WugO9TCS85FLk1pws8LA6
NMreH9YIhcqS/CVreNsYFSwSxZ/AxBSVAnSVcEaBg3Gsr2IfJgCzq+xu1ORp6ccj666hY8ngmgSc
2Awvp3sLmvoyA4d0n/+5qvfoc5gwnGDLOf6ITxQjdW9Ern0j3I/xwvauuNuF6IGDC2JspZxlfRnW
dDeNPThtjTnZDtiyN1abIBSuQoTF9D4JHNE2cn1f0UAVob6RZ508hnDtu2ZpV7dUaHvYvHCmCZLG
JvwooYWc1jSD7u9+T2o622akLAD0RiORXin41scCh8sGDU0w5gnS9et6Vko64VyTv81NdZ99meDN
9R2zuWb6+mGp6L+ntBeqcJx59NiNVAoApXikGFJx5CRvBdp1NnBarj/epcWOYZYNKK/JJ6nA8kO8
cO6++7IIEYcbR5C+Dx0hwDLYAOMBUW9YNfjnsiFJidEjyoWXcXYeguVJzCq3RN0K002NmWh4ac6R
PmeW1s+zRJyBgC4T6mLvTTaVxGxB/3jKervOlH+NIS9OwjRp5TxrweNEFVMYmnLVm+fKGRj7jsHN
9WNDGqdPCCeANLFVp/DkR6Wqaqsn7uEdUbSRljMpKZ8tp4H3F6ognKvjKUXPWltfzCkXT6SmUilk
vpt6a/kaAfsRrPz8q+LqpS5cdcCfEIDpb/1jnMkwNpwxcQvq4J/qZnxEpGn5PZ0NRFY1YWzecgod
App+3Z8TAbge0wQIQ4E2G80qJ1dkMXWD4vpe4AALXOK44zuAVIa4hip2ZvgpeEshmkhDW2qb66+h
p0NxUym5s7d+Vxs8kOx3XYpbqpzS1NbQFD5d/WszjAlIkl707sAs+JYNFKFXIr7VNLIWh68CzEeU
umk6hGXJr1RnXcpNJEfj25VuJPFfmOTY2zh+Rqp+p72g//mfQMeylYVsHQyZ1TSh6SXLwT41VXXj
xZJQlRTTwePgx1R57aKwyMhPiy2U0JG/1s3xg62DkbttWjNKX9DJ3R2zSszqjGnc1XVpxRsh22SG
F5WvlFdSnlkPs5iBQxvNAwK3R3OFwEE/WQjKOmgXb1zac0fVpOfkL4plNJl3kIqf4MUL7/mitTKh
nXSeE6hauozCKmJpSp2h7MSyHeBdV/HQLlnmIviDAaz30JukudmYLfx7gaf61LlTjWpfbbFFCEK+
SOkISxKTeVuFlnHhrGCKWxkcA648SRMYUpvGgQiLiMueiq2+weig8iuTGsE9F1j78RMEtFeeQx9j
7KZ5Cn2LaDnLycif+GrupZkpvFsyyvNnXL9dfjJMXARKp2NfIeEDX0axf0/oWXmibH4aMMUozoAh
o4Ja4Qq/TAtt4hrXwGfpR10HwyOZ6DliTqQUN7bMacxamHiNnVMElyv5jT0eH/s2LUQ5hTXMEFme
e9PesLl+TNVGwkmArv+fwTtb5V6DjTmUjBrSm7msL45WvxmffeVNtSicIW10nOMOIF5uad+gDtiC
CoAfmlAf8JIYH4v4JijTnpAtsbgAZX2Mp5hO6+Kw4UZZpTuMIwcmrOI8i1WCl1Y5zRDG2uc9H1XU
e5ZxcDbZpbLIQHK6dDM+eME8xgh+vLLRuxPcYIL7ml8zMeAvCC/uupTjs+Uivu6/9eqySpruTjAU
SGU/hLdOS6QTn9nEJQZ6KLKRya16GwzaNrYsh85X9swGPjCc9AHX1m+pOF0ocFyuQYR2Qo0HLA8d
8tvxvF5CSRKy4JGxBQmfVvxTiEmdgavAlf38Lp9oNgi0Z46JQ1i/RXmhagaLAyrWUUXTUxPZDUnG
heShdj032gnf7Jk5dIlGg44KljGkrl3S66sh4uf8Ty9/rcVkuDQSYuVq5JosxTvZr4KQGcupVYuQ
WRP7fEMuDezzCObCuicen7fsiMffR5OuN1R05L8xMtO1H5FwaREofRJ4WVYipi0E9HMKyfhby1OJ
gGVPqKAx2dqWnMx6DP+usgWhTt9MC/nwdDTzoJErxoxw9zfpUUmpHdeAghBVB4gBle3nyEhS80n2
M2/HK7FYBw2SwP3gCoM26ImvRtusKekywEWU6B3ChJt6jgMp0VCWc7kCmKndMGDZ0xytS/qbvVfY
Qkx03CuP3dc59kdVjXLbI5aGO8eSwyUmv3sFMR/jbd+3DnozcwIL58o/H3vvBDgpvgvUKrUgbICz
cgodj71Tl/bV5EHBwKdIOZZ+441cu6KypYeeUKwq+enLB2ZEssbJHx+d3xCfzCOWBsmySSlJ5H7g
bb8mf/pONxGvng3njznBCWA1O/SoewtZtu5jQlvB8FljwgPBT9BzyzOp3COCCV9fHWD1xbC7yOGB
Thyl43IYkxEXNn5cVo3tsME3omTsXmLn5HFroyUcVO/UmD84ctJE0/nVffYyY9FYngfea7xNEMgV
Sg00QFXqGt+pH+KTVnzFsAUgiVfw3+F/xRhqQ5uiF3fqh55vvByVIPJb9nQ1LKIby31EmD3fjCCO
ZMpdg07lLF159shxm6iorasGHrt/sEaTTqrdRIQh1FS2PuTcqSiwcEG44plkwpBo5uJby11/jevp
kTUZSQB5DRYR90zDGSl4h0yh0Fe/FxKSJAcqo/XCULJZ/BWLTN2z7piKyvx4Y7aYwy4NqEhVaatX
VpWrHOUJB8AY7jwu0kyRDQl7W4o0sZKHlQL9MpTEm+q7zhUyfy0t6NP0igVk8H4vu7FEfDJmulnv
hiT5SLQJmGlEyCsctiekgdUAISarxLn2V5UJDQF/U/BEWVu56h+KpYevUIem4CfD1Xgijbdldq5N
PWIvw/UUdkMlDmZkIhzlLvgs8/M3bxaPp/ypCJ+y5u2PJSzS2WIyounuqCdBAPdNdVZKdiuXcUty
pfGAAErpbxbQejfZSIO0CxOxxYw/loqJ0MQUYekKxpW7ES8EwfuiCPh6xP6ZfLF+IwVHEyaZXWZN
zB6SRRdPEgfR2lDV9Av7GiHDEyyUJ6EW9FF9u1l/5T6COlmSHogAIVP9M+wZW927KcXdde8E9gOe
PU6SEOPBSrwY0uuEYVV2WUFLV/nZXGy924uGyNVPqiRWR4BPCdm/w3yDML4mXGAlU+u90Wh2qNWl
gENPmlwi4RiLpzwhCJ+TN/pNEd7bRE/8SBYJoHfGdf3HG9p5sE8tM0GK020TYvY6HQTQJtkB/OqJ
2Q28KtTM+pQ+7LuUsHBzk8TefnZXdzLa3DRL79Kf5EzIA4USX6UVim4aoFg+J8L3Z5d4OZU7JdrC
P2tmDW+BpU/NmpNit3RNbxdFT5zYSVsDy89SWPZYh/T9UNv18L9DPsrfpu54KtkvQI7KzSLqDHko
iF+IflyJdaPHw9D1Rcwss8X3zrHhx7WvXtzchSI7xIyETWyN3uojdtJfCjP6BsRyPl70JqLgXkkA
Edzpm0XaWEV5GEEnnzdphmpsYdT9H3L2F5O1218LaOMzON2sq1FCSwcm66BhEMDgJk2qQqM6b7RA
ccW2zxiBbWdzxZwjXiY+WVW9+xXG8K9cX1n6MqkKefEII06ugJ/txfetWwNZkPQbOG3ly1sqM68Y
NwDkDFid1ztdB5qjIm1fS96K0fLg3gc5oi7vSkXr2py5wrOz9+TmxhS/omANdWcouZvKOEthe6XT
xI0mafZISN0xBiifBHkydU+Xki1HHbFyBHv84NdmIV4sAkNzyq7FIlYvtpDdOnu8vgavwR/Ca2Lb
tvGlPNM7AUhDVZpJ4L6vr9y6r1CRju/gGMvbjPoePzyYd3rjVRkHo9ot1AedhT893JwQkZSrRgee
8JC4nPaopK5SnMyHBwIgK1tp6DrFv3vre5uTgB6CLDToLiB9HEmce32dvtmxim/X+Fs7JDCUfa1q
dUgujMg57GJENSD1e2j7a85ilwWtZ4Il+YZ+fD/GZ9yBr8fjctlDjY9r00POItFew0LXeaZdXXWb
3OUcJQUJY4aD5yh/geouBhgI/DgT0k4Pp0KPqCaYT9awcKB8usv5GQBUt7fNeoCQsObwe/8ImnGo
szUSD4P7RQDDClLeuMIpG1d4N6LbZ+nKJEWfwa5+Pu0cQwNQPvM2g7tP3MLgH4NW5eEI+Rk75txW
mRQvPce5unb397wx4WlZjSUl4als2Q1ppxFMxStrjr3krYK/pHZWcz9rT1Wvb2ggb3Gfb2rOaapm
ZGBoIpMKcg3EPfcKQc6l4vy23LYNcM6R4S6Hnsbfwn+Kvzs6DUbEM0h/GvZZAJeuGRSjwyOq7qVb
2SraW1OYhdgKdFslB/Vy+a+NrUzmoMpTDK+3GW/HEZKnwJ2tTegYr5nbFiHp5dipKUVbubwd5gr7
vB02RX9vUmgnAKlK6dmlf3pnxtWhUpmZdswVHiyyfkJJPWrFtRNHo/dzZd1FFp/KoVmRyEtWLOb+
ofp4C2QzAnLFaQxiOaKGtrHOX0SksBJj05+lyn25AMmcBevEbTRMqrNwNxXsYou1WkFCW6iyKtsl
mdSTzQGImsvvE+EUuJ0C7aXwLnEQF3U19oXkwYUyX3H6YXbu4Lrfi/4HQNCIwkuJZUl3pCLPCT7p
w7MiEVgwdhyGscpb0Rp9rcr4GuTpDtLWm9eyceFUGlz1z82Kq8LszlxnDiUQXXMwcaG4bXI0CiIf
QSs9uYmm9fVcLVmWRmX3VSJjp8lw9+RNMeTafX2iNzsC3CFUU9hkKxgzGBT1Awvk4OYAO+9dmncs
djiKPa7yc8HvyCm/HgyRvkbt/wyHoW6btcclAUkTuUW1wDJEmnmD9NjvuDanTtYmWsPNbljyGh29
/pHVaUCF6xA0CxvCZ/9767QcXDe9eCc0RPDTjG6zBH1B3IFlL6uQrt0jY7Uek62+kxQHEE7/nK9K
buMxgs+gVYSgjKMI+hGOy9QK4iE9C9t0cShZwabeiCTH4tJI1UoJmXmKOu7jQIwta64zOSxPzftx
Dpex8cAvGZMNkY7Qa1oSEfi472rDnGKtnr581aTH6VJHFk5sTk3F61KHWKSbfXwfn+kW3RN+6DVq
sOmk2G9A1nbSbp11dCGuqKOz5Img/ctSMfoXtGbVgW55duKvxmI/TcFvubFUGpYH8RVFXN0smFtj
quf+JST1LRmWawdYQtSQw5OE6MmCkr9Chk51KtY80ERmuatEEdv3HU4+O+IUtyNSR+CaEXVftLva
oGH9vRW2uhbqzS5kSIeF1hn3PpouHWcXFDWz00WE4R1T5lzq/ULhg8mUzchqyDU1ZgxLkxbGES1U
8Mw0ruDdLcxXQAs/ov4JbfKTZ9uJiYhTHjAu78ZLQPzRsownJO0RRgk+d2kHgAxIIscE2shMawsG
CsuZiIEkQJVcVZJp4ziVQHKlwWZGO5FzHaKNGIfiCyUJy0EadugmHklNRF0b6R3ZxsLTdrB4mnxe
bzwvF26+12PcPmw9SrFkY1xbOzDEJF5SmDiF0aLByxGisMJ+c6VhJObfMG/6Glc2WW6TcbDtUhOo
pU9SWBZ9jIlFkkh1IdeNCQVo9G2BxtwwbqBJOMOfR+UFXzEekPfQ8cZkcjPTJTHQZlGnOna0tdyN
54kEJlbCi5VV3T4EoeNrot8OfG5pd4F7UHLVntBZNeVurASePetYspxJbFI9gJlrjVa+NMJRUt1V
we2QIvmvjk5N4Q7NK+yxd9cQ1GWBXDhXFW2hF3sJZihui7vm1bZaoSZA1DBfbtfHmhchk2pY+VVg
jsMaBx6Aw1DgQ78HJwm24EgA8jlvOEQMDYFkjdBmru+x7xeiTxr5y16EQWeeBb3TDdGMdNWVtjOr
O+XQH8T+B2mXPQBsqDstK5vZ7K4VIgY7iAgP+K/loXwTyMmwB/6Ss4h7tsV6FmupU7Q0qBtSAGOV
2Wbg7czA6ZfziRPDt09nZlvRo6/NdW2LVGc7CLMluPQGNwWUQiwzwZ6/GRkzl3NFPCrKDV5FfdvI
+cGTZKPeLayL4NyQRYo6MGx/dI6PUVKNXONpJMTsr0ZkjhpYrUqHxao7AWMCjnJvCqAVjXhL6kn9
3IBVFeivSTCd5Na3fDvwSgiYp9mdAXJEA37XXz7P/buwZ+oUDehOhNDp6ZH6ne4lUPQ1Udad/Ozw
XzSb+/sqYTmFPTm2wI0/McKC8iSKkleDs6GCecpOnZGB5Dj2U0LMx9N1fYuoeI3ld3crUyaivn+G
1OU7oUFC6p+Ea7uzs7xm/5agNRT4FmpksoGHaklPHJZCHf4XMSxxkjv+SYKLkZB1KPbCJyl/erb/
z21xEQGUJrPPQmGh6h0Lr8EEAEkLMw6gu5GB9Yhkn3vF/gejBVmPsiaVRg5A8g6h28z4yQhvS5me
1ROl47nzHuRVtEU9E2+/5cz6Z7r+YKE2aLaWpU3+mBMpF6j5FH9KGb11XWRv9xG0UA+TGIAmailg
l/NrwSg0NJ0yKBlplDnxsr/ua8h1ohTYKmj5qdzOc/QbS6D1/V4jGXde42LWctCSjHXFedqgXDs4
+WCpmN2WOiRO566mD540c1lU/TC62FRVge/BCCPBbY0ppYXDeKj9eIra58QecqlGaee+EAY+3C+B
3R4mHA7DEQyQZfScEha1GrHBfgHf8kgUm2NyuC5+O0QOAADeZBIuPNJu13/tPnz4gZeses1E3T27
zYhxcaYw7XScRPgztER9fuJ+henBqvlFPyQLYbPfvqAh/kzD0CjkPKkV1ivWE1ks+g1LYqpmRCGP
SWE5bWVEmyoRco0PinhE8dUgfvLTrKurWTHh3ct9Tt/NCvhVQ/1niOxlJPSeQYkgEUwV04h1Rc+u
2KXAHuBQ7ohxzR/ab4aeYf2hMj4VfEhSA+JV0JlXjK1XR10YObLv9sFX7hYBuR3FEoOUSSlwIlNS
V7CHOBkEXDcHsUQbKM4vWPlhAS8sKQNSxEX99zjLgyZiHqC4ddvYzGQ4FX9WmYmcSka0v5Lk89LK
3ehyAXAeBx2hGVlIy65Ntf2QLw81K64O4PJa51O24AeYug/wxxXfM521CeVSdE5cWdJ/013vkPmI
zfav3hMlQkvq5mLPxvTkYGeOdTOdPW3J6E76oFvWM6m27MCMR077Ig1B19/9gWsdMHVE3zlPuKuv
bHfyzz6sJhJCCkMCYGlKBrQG2af+7wINVGNVXlQw4osAlN/X3VX2GUFF11u++mQxmGB7p3eWMsAl
7C6ANoMZG903p2lIoyrYm6e7nJDoxk+qE7EIBIu9F1mBwfz8u91TS++2a6lAzFykkAnIQNeSYKct
llRGrLbuq2KtMaohdPkTfTK8UGaddeKuvxinyKsVjNZDOA==
`pragma protect end_protected
