// Amazon FPGA Hardware Development Kit
//
// Copyright 2016 Amazon.com, Inc. or its affiliates. All Rights Reserved.
//
// Licensed under the Amazon Software License (the "License"). You may not use
// this file except in compliance with the License. A copy of the License is
// located at
//
//    http://aws.amazon.com/asl/
//
// or in the "license" file accompanying this file. This file is distributed on
// an "AS IS" BASIS, WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, express or
// implied. See the License for the specific language governing permissions and
// limitations under the License.

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
nbx3WAsRsvDRfQdUL+R9iqbm2mepZqVfZssaR+hrHDY8fkYtVdXzKYrZ4vy6t9siS1LOTIKyqRB6
7AD0T4nyy6P1a+VphWkN98yySBszewEMwUUcLlc9/EJ0D+KuF/PEXFI9cDtSkgRRyFN4sK9V8KtY
A/YzFUGpJE1Kwvs3e1cC4w0IDv2mYk8ddAeMwakYCF0StMmlud8XGkp36mIm6h2hfrkwJrU0tJ36
qkSCQU92Q9O0VZI+W9hLpmOLoruPPEk38XLjGDvuBibwF6JCz0lLlkNfzMFFdHWdt2InVVd+vrSZ
9qtyz9REGp0wKASyJPQdsLpqfNymhDC7DfXHnQ==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
jSMIU0iIiep8JyIeN+H7fUlzl/Y7IVJLxZcIglvHeOPs9pymix0i8jiz3KUGUKAeBuCMkyz69Dda
6BnNQqt2nNqxOyIsDdDy4dLzGSJjq2cyXBF/+LqqRSByTe5tjIIwYAaNfGwTFAK8xNqOT+MOmv5K
jRmTzw0XMa4GdxHhwHE=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
LJb5rMxTVzCAG/CSmlyCcqfL8fC9zOsU9nXGRkJkM0JglL/7KK6kTLYm+mn5xnpej3YYDH0QmjcZ
fbp0HEeXbUcSrHCIPzOoqzR+O+TVVZbgLlHp4X1UE5+8h96f0ukRL/P3mxMd09YcSov9kOcY6hTI
V2KdAR/VG4u20Fs507c=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 38336)
`pragma protect data_block
u5AShdbi62xWfhhkJ07JbaynRuDhJWffGFR7mZqC8ApZ/jhCKIF3aD/jO79FMeDoG1+qkEqeGUws
ADoAvtNpDiznBERLutvLkJDeU4t2CER7booGd7Pvq23xvLAb5Byt/B5S2iGnoM3gBylhcLZrM1kn
/fmV7K3G1PJ/Gm6S4aBDuXbLyKhwPyUv3aWthBAQhpmcQsqxxEEBiz1X3qw1NfnN74mFy34mfgDh
al18BKEbCw2WNcDUJStOivvA8JTZoCdkJcViyvUggp5gurlAeY7XOMBZqQwYkqShgFl/kkjP13hP
XBJEZ4eaVM/nnJNUUmnB4snejE2stzi3mCAGlVYYVtnMAZ42K40tZw2ySmbpXyySHQleVUQyeHhm
ssdYnb1Nbpg+E1qtBDC95Y+BmBAJYO3MguSm7eUv/rV7ZP1rvxSA+MgPzSil3maBgbKG71Z35/9i
s70pKodxv7Kxh6wnJZhCye9wPRh64Bhuz8QfCqPUThCNtD+HwYrVoPDDPLQaUeN6LX+NJqqtdtMv
4ELVbhMzFx6/aWlhtgvp3NBXD7L8+wuCirOgGI0Z66hsNrBBkREVXTMEC+RR5NuPKx8jNoXBCdKa
8GgswcpSu+VW7nyU1fUcQRWzWvxGiVpE+h0f0ssnivPyHKbcAVg/neem/rm6EVV/cJttv+LpQsAv
DwyUYUxLo0IYi0lzEaSlDNjAjDum/01eG33ysStTm9wx+i6tGMBJEKHmORqbSsSeRlDQ/mqT5mKX
oD10L19AzJl5iJdQZm2dzwel9H8AOpbQVNPVVYcs8i/6RMTwv5siR9TVuKEq2eA9XQPh4RdorheP
W8P37LmExD2Wa7qzjF7IB1d+4IQ7z0w0btTYhOlYJ8/HOzyiO9MKy07Dbo7Tz0y7iK2yF7dG5bHG
HreRndN6IUoWYq8fxBro+qkPYH7nQVBbSsLgKCUV+grmx9oiOVovgE8KBtim9UZ3uZLmudED4DqQ
6Rs4+PW4C7E6PKeGzQkV5wIm+tU+EX46KixGKcS4F4y0b/L5j3YQGTfX9e8RjUXQiA58FP6Zn1JZ
2rI68vDe+Uk8V8nx8eE3zvNbqpblX0pHPE1scXC8CXZQ8N3Kc+V1+KUyD65G0BE6ZWXF9Yia8NkH
aVYBfNiJP/q9R/2O6wV+ZdAHWrFFs4tGuzs1c3hhXSjrYgfEFMMbDT1x3zSyd3oy0n/h7aVGd4vk
7Jc+oW1eeFjJJBvPl5rlk4eqttV5XFSKOocxYszGaWrKE5ZHYInysbOL1rNr0YxDorfqb5ux53X0
9wTYVuOdnlv/gCiaUCXVMj69QK7yYGvJ/BaCQA0x2uLa4Z7bK5OdRziMYiZKJ41dM3FPJ8F5JmBI
Ej3a5it2j3Wgv7U/qCP0zNQoNi1ttOt4bvRG1wrnwzlXMwFUSPtJohJ9k2RoqmFXPXbUnFKuuDAZ
uwMHOlWgnF24WJtb+DHqVkPx5eOC4bfJekzJbu6E+TZHI66ST153erP8aF32GoDBMNlclKTWdueB
jK39f8wBvNnec7CzAmNmAOEL8MU67q1DkUfjhQBjm1vj60/e6OV8TbqzQfe61jYs3uxRUbYJyL4S
nbpMidBgqzzJ84gDun0kk/uH0yQ2Q6cZiRlYsUTF6lUGPC7qEypIuhQYuOZYGdDhdnGg1C1c3QV4
JqwWhji2aoDFXsFPmUXsNOIM8JmTaT449VuHKew6ibD6Q2R1Gp7eINjsvqCzscFLGN8c7sgoyUAs
FqKxDgUEbtvDVQur29IievZe/MJbiUJUuP7nISpqQ1qqeuWoQo+HIqjTrE2g31JpnmIbvvyaVMzO
8vjPwD1qjgn1oK572lRV7FBskOpZWqaCcc0QsJB3BXvA1r951wKV+dDyDzphtLfkme1T9glAEiel
amaWGiFqr3Zx5s4YY2FsgZxG2KETdUp7MYN5/H86We+zhdAdzFdLnbmniYSDAFMdQSZ0nMbqdmjs
9G3b0NU7wAyZAjyh9w6++VFp2AKPilm984THOBW4RB5DvwCOpuGVh6jsGHS4Mrlk2Hcv7NfdUVdT
UraekvHU39XGDXfLXM0nKqK+NfxaDaUmzJl9fUA9i8j5hfNqxgpc/FGs4B+seahvq8f7v8aKUCR1
l3HktMJfyCJSeXPsF6M5AnHjc/JGSGpSEMmEVlK12yJ5n2xyPEIgDbN5hEpSv+fgTZk5nDT7tWBN
yKcW6lF+XBii+jmrr6YS2Nt1heixX4tv3oZHQyEuYX7ikPs9nDcP8dWSARfCqD/n58J3mYj6q3wp
C9pH2fWAT6Xd3EcDcv+2hrtfunVqzZm2cSHbCeDtBcBHsd1BV3ogTGL0CPabTkZDua8cZqnh0H5l
DH69CgkQ1mh9KrARUkV39oClhXiqbBoESkiUrX/98oNVh0V4VgpTaKpIEM9uc+VayPGYvjUAW2Mz
dGVb4bAY8KXA2Fn+iOejfbOemPWlMFEjhjlzm4cbD2wpvb7kOfaDZdkm8j/ZuD22RKDfCw7HDs+e
eyWHppqn2gBwK7E0uzlEcevor4MRjoIipTzlqJ1xkArmGbqFEUQ8rhPLYJ919+tSAWocfpE4bH1p
UAuVPPNFrM4l/opL1EAbA3wo6iSWQo1DJcuAOsI57Ne5bnkS29Gfrhm10acVbtepk9aHrFMC0PGr
p6h2yTg0pFIU7CmRtTD4QGF4W8CO0cDHb29A+jweQiyCVEV+GNdPuU3Y7ysFT1sEag120Yg6W9tb
yw++oxBvbAj8u82l0yfcaJYE7FloqXe305NWD1Yy0zgR7FBReSQCTtL8oleZJJWMLAYKXwkZoD0D
/pOXWFw+mIb16brgIv2B39wJ+wPW5asjDnVuHruyIYwv9bI9/DDlXN1aTr/dc103G1awAgTrPAFX
Jc8Kjdm8H4yfqU7TVL01ZlUVQgnpAe1vBVvJMG/E5qytO7UBU51e0QHwqntddhZlfoqyzJvyWeAO
uFqKo519Cby3Yyt9SdEQemUnU5VvFaoq6lqZhpE/lDjhjWPW7qpwV0+PBHXmS6kPK6KEdetgV8bQ
SWbFvkb/jrNwWVhNlHSBFQZtZLx/dZbMAWLrqWbDvr/wAF4WQfQkuVv9UK9KQNCapbb92HtTC0+d
5eKSW5iCOkQZOyV2ajnF90BRZEawdh0HzSwhxue12hIjJGNWg21XmMYBVWgkPoukSrWEd18Sk7zX
7zsYcqmVQR268eYF0+E/gm06h+nUwAEnQQX2NejIE0zj/eZzqDOq4DCGN85b8ZR3CA13JU+ZJCAI
Qp3yKn9vd7R1JykglyJ888lAgVdJ6BrwSfvU08nXyu+d4fXLAbbmVXLcJC4qmYMIVh1kJ5oCfoyM
X57AFcSflm9hAgkzIkCkmDUwYlguQkFXC8B/cc0VoRLEEVLAOBQbop0XXwSciDaAXbcgA/KfALzQ
7LaYzybxd1b94gen3YXlZ0UHzRRzNfDPrtEw7zHc3zNXh/7YLE1d+2aqUSActsuhTinz2qIx6vip
5wv3XluFU5eEfY8QrqWPpYuSXSGsW/KfsIIRIDStg7TPJyL6uQRSXG4bvV6oPoEY3hGXLsrqpwjt
RVM043jns7LE9iPR9/pODA8qA1UBBuwVFDIt57RgvREuYbu3kBniGu3Wte4zwxurreTFkwSy/iUx
Taww/CghACEtXDbr+IM1GcqSF/+QS+Ld0YQQOzhB0A2xC6Xl4UiMDV3+ZO88tFnxeH7xSElS2ohu
ql29jO3uSDX1oqKutMiF/X4PQmEM4fKKjWqIhF/+4teGvE74sqPP/UDN7ILGY8WQVJSky4+YLK1x
I45sq+HtR5Pn1+teixwagP802d/zWm879lJm4nICivBBxrAZkG7vLJkRtqI3l28mgwZwBR3ot+cX
SZ6mK64/JHzZw2TVshMLf8SrEpFeCGYxtpgoedNDEa7iwhCTcRq1Fd1GIPdy9uXy780Uz7f4VITo
Wah2sVEJQvOYFe17YHDg5zTR1xij2cUuo0eJI1n+DAHDkz1Di4fk8F7JCJ7PlCnqu6vY8ZQaHhz2
Uj6BsB3hjihTZ41ap5UyNOG8t8UeKwYV3wYFivv9qkcreNQ4GiPWN1uIb7HfVjLAR8cu9r8ccgg7
hRDLZiKkMhewlFNjhs1CmAWFpY27fk+BvytgZG8ZEXbLdxzOgIrk+YcLrnDPT/jDMVAwB1dW343v
ml/9sM1OKn4u3oloDATpaBy0RWz1vC9keZTwcpRxzpigIc3v0B2NGc7FMaFuLxkL+/MVjBSEwQEG
WFO8y28mJRDBhFcnisf20DmOJ/lmzmVYxpL3asa3KDWVse9AwEc0F8KQ25jT7OdTvF8jz9wzqbGR
pObdfCfDwbAi2st+HUtDV50CxgTHR9pzjvB4mKj4gUbsKuOrlb74++g90uCSN9OsNdCS9haNXVxe
cA/jcupuDcpiv57Gve31aZ0gsX3qeKdrGN2MK1qfdZNsvgrMoybNBYqB2IIssgLnbHS3RLuTmMjE
6nj/PlwX+VqHiJRrMEXVWY/Y/VqBoIEymZpQv0ZV1RNSn+Oc7oTK2gbqorZP+IYtH3xmK8eifzgi
kLYUcjijP4e/7Of9dMPIlURRzZMh/eNPvv+bMY6gtEfrin5IyIEOOrkPE/3TIYyzGr5tpir9Y8bf
YI85kjSsl7MtfX49Joes4TbaTfpBlFgTfuRWhpwbSFqfBI0pEYtKUWrhazuvDTFQT3agfXteYUXG
XtqzW17TMNpYyhgcedVckf1oeV5LqYZ9KNhYVBaRAwo5unpYMu7rQmh5dU3odPlaxE3GTEXl/4/u
TL7NkUu59U3UIQxeyvIs1UdE9WMGSVEZyCEtid4xk7reGDq4dCHxXY6QAvOFP+c8dEh87T7ofA0e
mMILAylASRaEPKr396tpLn3FS8i5Ui7cAJeFSFY1OXpoEe8Eq/JEDPDhM6WdDrHR1Dg5Lbotq1By
XaKfLRFKdaMK0PwWohC0EnF0Y7qdw/6x4h4gU8Tmlzj/cqzj24Ia2wNSVitF9LDjmGDelFY/E3Bh
JYEqNUIarht/YmKCYyf9PyDx/LmSgsyTN2NQ3oc+nnHRkliavURxNdpfiN1OKXsGC5ABcAD1sgwy
tvMvGFcjcKKKczf5iBYwIf5dpXfyx1bGRmuNY+t7zTNT0ht3kZQkXd7WvWOYNcUT8VcyoJ9jrU48
//YU/ERt4ADRnz1+z9dmd4aT/B7yTn+yPhLUNbWXP3WUlo/Ys4CiF9vI1Z1qmvt0PmDQX7qnUpcM
PA7U26sLV2THik0OdLoWLIAjtDDe/qBC/FGC4maGP/NQiNj+OoFmK5GpWetShMkXG6kY0nQ1ny5J
06QTY/Y9QH30iAoKXRQEl/pvPPo4rMH/viH8Xi75NV97zoGKrciCYfc8cl5nkHeVCeV9kjW+8fAQ
4YEJUkxfliYWmJASH9OekzUjWAH1QwDW56+D9M4RJXD01rM9potvUqegLGkOFJLm0d0X7ndXqtsL
Uh3KQtS/rI3yHBn0DjhUoXbpbjsuA32atw72zqN1D0WDigeIE1tiqnUiTOSXXlBCR38gMZN4WQqx
iCqYbCCtvYrxyEvzSM1Yo90ee9eYVjh3as2iyVMLaBGel5bOptDadITrdSpFdTIUXpmsRQdbI9/n
5lTBb+pvxMqWHVJfsUzABpIJE7RHeyn/uypL2tH8HfE07OBInFZvpbvAvfV1N+HD9P3A66wcFKGg
PUun5qECn1yzEMLiDb6uIyjMzxpDNLKwjEACHbmp/UUUuoOsqtwrWr1bZipjti/YsSVcdJM3JvU9
lrw4eeDnC/7aIxWawRDn6fLlJo2eX8uSV+iTZ9iyd3Bt2jCVDXnmLuDDuRT6zyGfgGur374x1DZn
wn2VwZqgroWVSgF4xRdJd63T3EOcp3UWTef0lDgEMGxI6T5YTSH+KsROCPFN72IVuUiPItrgQCCF
84hehRlpEH8lA8OTtnuOQQ+A8kIOX1tTdx2WFX156FfLBHlgmaQUhiElesuDg4mtYwcx3HkYGK/t
nbyMMEX44fdYA4rkkGSwaXqPzPnDiD9CIBNplLVxC1nQ+wTv5TBmsZ6wOVAhtadX2Zbdr6GJfud6
BOUHt3tgeCNnA9ZcXOYMhQ8AAHaki0aBKZiP02OQ+MnijKnK6m5J+pIkPyq7R4Cvq7ceMlCe4A0W
0kRqgxTyjZ3p8kTH5BcMArGCh/Ebn5Y6T53qD2ypnWxAO1NjkQK7pLiq3aTytIZOQErVxn4aPy0l
pF+6Oc0BjpgVn7GLAcWoueuXVYv8E4RdBTveqplVdf4urzvSLwoUsb7cxzN1fYLT1bf49t30mqDW
jXPbj0iEDjZzXNKXQP6Nq9g7AWfbT4wrykmok+pZSgJTBaA+3q2iWGBAsdJxPr15sRWf6edHjwiO
9Eu3Tucyoz5xt4+RJsBAhWxkhRQ7OLu6NHZibH6Hqmmf1xQEkpKdO+5GqxAfhfKX1T41JMcimD+D
vZXUgLY0jEXi6Xvw7/2dX+cHqRCgkNxgmCvPXjM6IAY0tE0h5Cd4i+SniJrdT0iKrI73OnDiSe90
KNLjGvZlWwHll2qpFOESA0sNFPdvzPeOnW61lMQ3a5JRKvkES+qQclKcjOmCa9h2emkq3avHqLtz
nUY2JmM2h5zAGe7QqEJtw1LLTLEgQbgiDqotZkmu7xeoJsF5XS9I0mlNJ6B75RJw/Jm9GU/fcKH2
90ClpmUGbB1nGzyPrNGeyxKYpR7zHJBit3FYCTF5Y8G4zE6BR4ktsWEloXR0M0ZrYsMGlm4COQbK
Xae0TTIKYdLpTlRgMitBF1/TSiBBdYIXoo3wjejyP+AZQU2g0hgItfOMEI5//etOVgs5PQj/JSA7
51jnd83ZgJ+7C/TY0uA3pLdi/936DyKSGETMUqk3J1u68THoKlvojyChBxCG7PU96qz7Kgl3y82B
2Aqn1RNkyv49Tnt3zSy8X9db57+VwPNdkqpQyCk6YG+UKqLlnidoUnt0VbyKkCgGQKIJm3aBHrUh
Wh0bI/twGq+waXLTz3LORX9+y4zUOOq71cy7oU1gG8C/fAurVGwhSAq1YRFh1+rXNANnwrUTO2Ab
oQ/ztlYhWRu1WWMkFP0bp516+tqeBMYEqg845OPhgkyFQKPPbVJU21gUYK4fnOxS7wPk80K+jIDg
EWEyRpZis+7yjlCDaN3QALA1graA24UD/JCUp5ypiAwhSdk66OahWkmNSn8aVerfLdL/r+CmwSL+
bxSxUAJQy0R5EMtwEtzr0kUq5oQ76NwV7LXFJS4aRppLD74FvM7rjg/tKiK1i1GhPHqvpf8MMb3F
Pl9M2UIdLJelrbrp46KlvgxLhfWa8pG6G4TJO++WGkwIOmhHeMGWs+z/m4FPKVjgiBGXonZZphGR
21MVPmM3IgGkHVaWCHGlqaAgGfmB75VBzqeEedUyA86occF1vuhaB2JtSfM6OoJWeIzvpLC2gdDB
S0ZOiCqp8GF0I7mqfueDVTB3/w3gSDUZukkYRO+fMrdL6rvOlP0W7iqvVzq0cssAGs0oXjXXBJcA
UPxh9vE88+zGmAsuVbxO+W2Jy+lUOckc7+9PYhlbeYGzQFb1zwpex1wpIMsQkJeSr7nu+S46dQ8n
5bKWIZqMTIuukzSoTZsEimm2KSvM1JKbaflH/IHAMEzGYsKKIs4rt3HPWtaGJH9+q5QRP3D2jQbQ
/uE/G4AjJZXNrzWRVDuXc5LWlINPEEr22CSlBzUNTALAI/6ifb27XcP2/eipc7RN9FrP+laLMPMy
7HSrHgUQ/jddOhBill0E8ggSWRhJQvEL4zLA9t3BI0zDRDxXrTUrARDEhkSsXhdKM/5p2SbbpRSK
Ja0o5d9RwsC2ykyIlKx5mDRadskbHaoMfjNasB+jopqNhUw5RKDaNcSzN0CYgXEdiFRBbUUXKbWD
h/wL5KdpcnuGUpPdmxqDrms+QAHdSptsbJgreNU2atHFWJTvshy3TCEPgDcrN/0bjIy1h4302cjY
d0Z3HpzWpo7blKoRjywLfUuMqT3HSMeTK7akEmuOALlRYoCyHOgP3kB5MsIAabm2zv3ATmvohi2u
iyaRrDpTp4BSvJ73vAO8+N1xTI75hvQU6+LNrB0R2TTs5/YYMovZwiJkEqwjSJa7xLH6wi8CCb1c
7orgjryolR1X/IIcI0RyF/g1im1ngBmJMoMa/4LVlFRwFoA87rSvgcP/auop+KzE4cyo4IuiYY6c
Jlj+JERo6EBFyemyl8iQ+1FAs8TWs9gqGNj1bW8LgsScNu9wHwdBGqsvEdIVfNOgRJh5m14twTEX
0qflv81DpUuuTKFhrWtUj53Yh1DSTVXfywzE7ILMG7V6yA+xrYSkyZSkpWfvT/33IdPAxnbEVVmU
kjqYI4L3y5qRz6OwAmVmr0Jz0WpvQjfcn+FByuPXYidXrV9BbyROqrDT/5RW3QoB76di2LGTx305
hYBED4x5kMCywfpUkboeqp2QDBBP48RzHTcSq7Wolg27CNjZA0HS5/E8yE42srxbGFlDa/6iCPRu
d+ghUd40ymNZT5y1OCtsVU3/HM090HJyRVRqFM5UiE4EkkRnZ/C3FhJuwZt8aG1xPusCYHQEHVad
IVwMGLBaZ2nZTOi71En9H6KtRZbkStg1LhAcRvInkosJXwh60C+ufrvKNFp+jeo0Ck/CXJLyhPyS
JGMJk0qKc6LENLZw5OD3zEcFIjKz0zEc7Hm1qGw+hEBaB8Tk0IzOIXf/9mEtlxk+Dxrn3TJQGQYC
+hRaY+dC8kLc8MUVWaPTZgikbn0s2EMtkZ0qJXlMtWCciejYvlLo+aPJxWx1ECWsatuFxyLOCqle
qTq214BXhABaYQ2X7XYZZnj2ZKaAUnex4N2DeePEDxaq68LOCBdLEy+2lMfcLCw8Ulp1vFQXnuEx
B9KaQru0dfpgYcZxArSbKDqu8rQMlHCSlgEWzLSRkvCWQqxI9jrb0zsdTqXkpuIW6flzzBu+WSUr
xjWB4hqzAzQCHemmyaclyI8YBKJjNcccF+uNJuoX/Bqwo9RmiegqPFbydvlxAXY9omAkR5kQ9qd+
fVt2VfYTHy38G0Helmgx8grHoDAaaDWfZRG1zP/MXvRFXIxIHFrrAHyYgFMeqLkAwOgeTPGmzxHu
ndxuC51Q01qj8Y12b41PCZAI76pO5LvTpD5u4r+QumBSpUV2i/5lTSfrN3w0j0busEH4uSERDnQ9
WLClZyfG3J/dMVf6YV/1w+CsU30FCAS6ORCzuQNlryf/nyKOYyPvaIQPoJcjrRhlB1TrGq2Q5F7H
vsX87WfxaJEcNyGbGkY2Zgea+3kDavo2bM8lmoDK2SSnImyTvuMpPuXn84WXexfe0RgWxdBP8JCH
a6ayPaez8RGP2AvPrDM7knTzhUzGDfdq3Heoa8c8rb7PJeAikX4QNpYgGpNPCsN310xMFAeOSs7R
LpcSL+nrzTnPwOXawvg/ylvKehOd3FTTIwrtLaAkuki8ul3tLb5vJXMi2JTH+48WTNvL+gd8ZURA
PZJr75PfDL/C91MoKVgyqKtY2Eob2Kr/V+In35OImTq7yQIoq7xtBno+lVnwuN6cdA/83UdY4O2t
nkTciOwL8CrNnYZLN8E4/7LTFCos7OhWNI8hlhaw1uIwZ5qJqGYw6FXK43SKTwwzbf8YvKNg3RIX
ws5vbVObeGDTUOO/sUHX/gYi3ukcRxtIZ/vK7eObyJ6zWkHwjolcLu4CvUSO2RSue0G7foitR3pd
utRAXjyQp1xaO4+vLUFsvnvItkco2bwlDZL3lFnIbt/b7qk1Tt20Zer3dOLH2Li0S3TjUl1rdiju
2KAnWrimKhT79gnJOE9FofeiwFOlqo3oa1URtvMbDJcAn+WQK2Zq9xgrEYqzZQoA4PSz5xKCTI6G
76sAwgsGXdgcMr1X6MKvWidtdgxDTxblynPfLsJ5uspl/3vTQ1Qi3ehdIzdvdwnYg6KLXoihyCFp
LroWvd4EjShiHUqsTcUpSmy+X/uR/U6U84Jnk5OlW3MMjsAuIUM+rs/ZYCggLPCs+Tx6EDGFCqF0
UV62tAIsk8oRQppckqm5VeOWD++yi6l7emh+LSj+XRqrQ+KOd3zfBfPMawbYi8Zyl2bi02q0Eh2K
akj4EAxIZ6uQ25XOmbCTi1Na4D4SaFRPhADWjXXYamobOmHspiggqeovgpf7nF7FB/DZ9jmY1b7b
UyomrOzqC+zn0bCaAQKjyk/CA7Ge0gcwhrhzMDr/pnJJDsoNxfcZik2R5V9kgrS++FHkJbtaiEPu
b8XTOEUXdSbACd6jT5yB0z14r0AR9TVDoQ104eKixb/zvyC29JU2LdM9EAVTRPGYV+J66unPYFwv
wKJ3OlFSaWGA6Bd11VyyA8fxqj8/iKd2SzvdpIjt5QvW5W4EPav9QeR0Pvbr2hKY/XpVCZDLDSjE
1ck9VCTEDXajuw7sduoimncgqv7FUtaSc8RaTjP3fqVqpNfoyTyaBLXSSzHrVzuuTwi9Wt7TbmK3
VkUR2ZcAvsh7huraokdD/QPuAEGHP2N8cAGmi8s6t4vVLPCFLsaHwdPQZk4gLwwWptj8mUAIUa/b
qph8U7KnlkC8Ez3O8iXVTyKesNQB6gnF9RC93IFileHvIZksowJLlI6g1jNVy0bghF1lkrHrVSYx
9mJcuRuuFcTjFZStqwZKbNcEEXGD9WcGYjd35tC9FqCLim8TrLZhPT5T9asV0Uf3Athbp+Zz63EF
CHAJr8WrXTGVW1n5GyBGi6JsAEk/vYhmEtAT1RqeFthUVvjzqQoPXwIanmehfMn3IHmHYgGedxSZ
FBgIPQwi85XJbpaRsdA+62CN2IWWQahOMxL4CkcE6qKUxXDZNyPdMGlC2vvS7U0tw+3nJsamxdcE
dqC4UrTMGw+6sWAcXBsOG14sX0/SqF547TCT/xFHeC1Dkqul7QO1S9tOcD50zXf8sjPFH0lkPoki
ccAAXlBntDdqu3zk9VJZZdxsL/Pd3wwQgiITbwdut/nnGdGToq1xoZlUkXauFFdMoIIGItsZjw5e
qx11ul5NQSprRfIhsMi2i7mWTyxsX9kou4ElCUDJAkM15utmpUpV0+ltc11j7z0/JXFKJDvIeyMC
H2BwrGDkiuYMgwERtdRbOKbOuL2AvHs3YzJSLrwdBL6eE9LwStLI+58UjB6kRWAt3omUW52CqVc4
SigjLv1V1vaQELwQG0moYvIcxvwurXjh0u3F3tRaWnePN/Zy/T/ptHhHk93+ptSF0lyHfJGPhO+t
2pATc12wweF2xYOJXeFBGyej6go3St+Ks+0TANmV+lWniY44Uiw1qWte/Jsl9i9JSWMU+NhBIUds
3rmknhO62hcKri3edl9P1Zk4Oo20vdeVGoQ44WRFoQyxPXb6kXEqipobGGFsYQE7N+2wNb8cXhGg
1kcp633u7DZaMtjukHJ8fo1n68PO+h9pQads9/GwxiNOVccYWojYpa4SoXy6Vf6OfJpN/FgsaN/W
mKxGEBzcoraGExpaMSXbcHXUJJZ0TuMsujxTZtvREQs2j/iKpANle/cJTlXNCzQu7V8l0iqFoz+b
D/B/FvTJxIb58ZgzEXGSCzkqkF52ixs2fPn8NfmTDFcl/8fIrfS2YL0QlyAo+JeLlfxVaZ51mxd3
N5+wLGV5PgPH6x6uq9wwvFo/TFwYNnaCKyhnmcXRISS/YH+UvLwRuDwAnfK88e19ketj0aFpO7Jp
/GLILFdHO4FeB8fK0RaFl/fNXMpnDQDerUdGXfq4YPuKU+YzGn6omFsyDOvVcRKRTINbWHmgqr82
GM38VYIHNbcrEfhWl+ut2qBOipZf8rJn1pgia0wq4kmaZ0pH/DuMOQ0n14re6ezHEfnLXEGhzu2R
TkNQmyA3hEiR1k5pMfWQrJlkTtps8N+oADiRSutZ1oN2ljD2R+eiEAvJ3AH+1yifhNuzU1f6UZvO
cazauAMoGuInI1wwFQTEGZohUNBEJekfqM2I9KWufVtY5+36M0UFSqQxfhRKTnTouzdNUOo8hq5w
SePv47tdl6nR459m0CxtqXLzWi9H/FLMZ0v71hicqdYpDR4HtVy2kO5V+UYkJ8t2GYfoeAqmk6Y2
Ljs1Sx2lCC1GeIWPADW2zdLPysxuq5XTE3Cv7xB8OF/tfLGNEy1PaWHNzu1dACuiOp7spACwqY9P
1vt6a6tdu+BaeiZk2ndB7fDjmaYUbkhqb0bB+dRr5d7/Eh0DXxzsi5a5yn7kI6+023mUGxFIPdPe
AffV3nxfEDIYNxBT2eAF+ujp+IcyhEr/v1wGP0rKV4Lx/xp1CX4AXxITUAsHozaaIP+11XPhZaJy
VJhjxFccANcQ+8Yv4d3owJFfbNJ48BS81HO5zvcE1PImCARoq8w96g/K4jmBp7IlcZc0lKwyO73N
WBfxu/emyh7WsF4BNtJXh8z37GKMoXvRvaMeMOernBb/RhmnG1gx5m+Y/s+mCN6SXC+GZQuIILvc
MpNNIJ2Didbg6f6HYct84H1+xwzd1bho26aEBpmdhKd0Z3z/k5nq2H/M54lkYu4iefI1ZVUmq6nF
ClxOBBYzr6rrhLheAkCyCNLgev36GhjAb0/LuaDeV9T+j7AGYGCg6+X5iMSOn1twP5t+oPtvnhcE
oilaiPHAMyzBmtROrA9mW63Inm8BvrPFekVagX8/w1hT1bv/DOMAK9KAXiluEmDVq/ZzAYr5n967
DxcPoZXl5iUYZZ4mjecGUjnFtASet7hvfuLr2La3gwaG1ab/b32cLrzFmNtxFYNriJwd44NshPMG
Q658M/LYCxGalDwn+rKzstTYG2duke+sqtqlaiKuclR/rKYpc9iCBfwS2IriEiRat6YDePIqQoeA
1gIaXLvnUH6/8/RiYc8INUV+WzK/8Lgpyp39aLZbT+7KcB0ha7ghGVx6+GF95NXzF0sCMbz5CkMn
SWfvYR/WLWlgDtQrcjM4vpZfab6fe0q2uZom1egrrywi9iyCWUkkEF5bPsk/ja+WVcb368nVpb1Y
xPFOfkS94lIW1JR3n4fAMs1C4T1ZdnCPjqdbXyMcEkKlZ/vQR61ZKndqttrtLP2jRlK7No27/vXF
9Dv94ZbJuP5gmRyJs7BqxMTDKKAJ/4E/a6G+npefI1zD7sBQ9T8d9fbT3rTFCl1GYwU9qQvvzTws
ZS54e4k1AVSzS3PphXynkCOiwmmqoFzdtuPu0w8PDCbamhi0tkCeG98+HXmxT406p40/e1hqvcSM
iFb2Xyeg2Xs0A+w4hVEbg8BvCFYnlQzCy1Pid8KDeCBlMoCZZsc+hjcIhBnHPw1uf3UeAkITXmWm
DXHZFrkNlqrrOWIrxGacJLshty3BIHgOkVoLCtQcMKg7C0x+tABHUET/cWAbZG6Ec8UO6bjb1c1S
Wd9vJq2oYjpoBUnVsiKjNq8avNSsGVs9K7DP8wv2I0zP58LT34QMHSZfBborduqWblKcNAM2RIFk
xL7ZSbybhbAmsWKkkSFItXAMW9rKzeB2sRW/Rcly4bZ046zne0ePTnYLtVlLWFnTxi/1JCPaHxqN
P11ua0PKmJx4oXcUz15aChZzKX7CM5idyeaCi0F8HL4mBXtopFPWEh8OC+hwgZX1Cty0Kpe7tBpV
rHxCTAnM4nhOUV+vBFTXsfu5HbraVtQKOdjkUPWy47bgsrmA9ghsmrIeiEM3/lvY66nqUacoVxQt
1RWAUqujxItfjCe4rqSSbC4sTYzVXT2lyU+q7lsMAWd6+Onj7tVKbfrGE28nBi3+AkiA1loP9V5V
/wILKeQjpQ9XukYP/8t4wj1HIVTtuGKWdBqeBcnQgh98c+HiUYDugXYFU4+9+xMPprMvz/m9Cen8
00Bs7cHGls4GBSDawZvBfIaska0lT2vJipfWwQB7mNOzygV7mhxzBAZYe8aZgcGwmvIXsaj/ZlB5
FvOCJYMW9HFHnN6Fc1aUx4unT4lsfrDaaca/Uk8o074sZCEvlIXjKiUZYNvR7KaxTpso5Ucc4gx1
wR535o3lV29yUeEoGEyQnQ9XVZCobQ82lpC54Sm+NQcg4OxTQYqY1GntMoJPCAj4BX8Z3dfL6sA9
0Au52X4SSCCrc8o/ZBnjqyOBZhE2wwOuvIRzm97USwaWAv6nGNJQofJYRDFdn+02XZSGxb31PkVp
MW06GBqFv6kUtH/DJllqb2Yz4Bo3zfHgpRddHHm24p1OQ5sqXAgSFiHJ98jmzDaAncNeYGbd6Iwc
bvtycXJbLyphT1F9m5SRPt5cb9mFyo4jwIVZ5yzWlb1uaFcLcQX6a96yJk51k1JVQGEA0+V21aIC
rgdL1mHVrHBIosqJh+vM1drXwit0tbU0xw15Q3bB8ePOwYs/s2fFGH2Kx9TH7jxbK04AZkXglppf
i1RrnGzScRWi0KTdCwePHkKe0adQV1nYIlyqJ0D4teNpdLNxufdnn3WsLG2XD+zk87IUWCvvfSwc
kXl3OoHGWKlxhUvlx4XcBZYj0IGy8GUlA0AdpbROBLEXMAs3ZdxEvTD7DfAphUsAF7XFCUsgP9aP
9HXvz3SFFSb3oAbq7dSWe/EG7WGqEzvK02MHz2/R20YZ/p/1hp3piloM5B0Vepu2B29YRTWfIj7v
XDUfX09aQYuFhi+fMs90e1jcd/xoK1E7bF+ygv0odCXSqIuGKU4Fi7LihcIqL/AK/S8MtS3MyE/2
Ur+2lNzMXIz9Zj5D+zRKCNPvCHfzWFTK3h3otkQ0w3FpsaM+mIv4f38bL326wfQWQR894zoa7ZK4
BdgZQBCNWXxH8cuPoy72G4xuN1xqLctUqDwxIYdaJPjqKOL2UuYkjg8HThstpbZjVsINvN7t7HhX
B2iEcA2lLeSNVD8bhyYXGFSq78GiGoUmn4Ek3IesmC4XEFDU+3ReBA6Xzn3ECbLVqBtxOaCsyvgF
/I8nPNRz+qZhSRIx6yw2H6cFsVwBZEvumk9EUK/x+XRYTPzoD1Hg+hijVcR4nO1IqbjOFWxe+Z2B
oNQNlRhvxJOvgzUP3Tr6nczP4uWe9uvR01B4b9R8RP2enx3hOf8m5TxQbhFZzuHXOxvS5yhWahZU
CQzyMckj7vMRmrL4anUXeNv18CALrldp7TEcmF3vx6iw/MydP6FZkaYhxgb/G6wT/UEM1x+Vk8cC
vhe+ymVKjfsTXaPr30ORSdC+C2JZCWsPart99tgBzBa+6P+6Cb6wlpEEDoj9SnGcXlXOTT+OQOy1
pMAr8KD9B0CT3Og/smg1mlMZKS7UwvWXYj0WC1psmyFk+BSvH9HLfWHgDTR2CL+wvpuxPSljUTfY
SD7OythBj2WrtTrS5FtEBlJ/rXMtSyMJ6j4Zim/+9egUY95PQ/fKQs0EoaFM8EDBnUjygG9U5Zy+
6SXxruI6OIgRkQTSjPPElPik+yLRchVO++WxgqhkqmN4g8AFrQJKH82eMnITudMkBLKBRAGyZS45
xNPyV9SmA969YCCy/dRGpD9Un9HCaoiwCpG/3Jdxxu2imLB9m23xWa8s10rh1LCzXl69DOcIw+nA
iBi/ySI5V1ejCvvXjALJusZyuDJXEK3s6oGVoAh68i+BwXXAk818zl2RhkLEkwdhWdgRWSOxrtpY
0jupaKE4IOLNZWus9xxi7skuD8+ISM/aUwWhDDU00FMTfzhuoy20rMWqZ447tGlVbSAKyQKNn7UI
MtXUjJ74joUTZJToA2TLPMLdhZlvNdvowmOpeT3CzoAKZ3MXInqArF2HZbSA2hx1ggc5tTAGzpmX
CSYqB/qPbx7tYY4JrABFYVPgzCFF6tEvzM9GP5LnWB3Jh7euY4J9sAooYkVxpA+EYr7UqhKYmVHS
+9u+FIjVdd//JcR8CS9jlm3vT0n1Jcw4+zt+9pzRfSRK4RSeTvrgeaGa16Khm+qso+GrIK8UxFmB
VRqYhpUhlWnqpaCCeHdn7hU4E3wynvPd616yXdDC0qO0KoljJJCyTazf5Vogjuz1X+6CgVpxvjZo
FCFv3fRlsicv9T9mmRSeW2fu/nkRAWVJk2B4nKV/zp0h3UGdublhmlISWgJa+Eyq1kGNiid7/NOw
CSY6CnwPBZU24oBZDVaED/dKPbEdtXjhRcB24Ju5agCEuZzd+R1YyRmMHvWXsbK360HOw9jZhhpD
XlJu4OtMeTyrE+tobe0x6H45HRalHGdp0ifgNDeEYIMe5wmtdSdAzsCQS5EgxmIR8UOpF7AqQ8lP
Ur4ZP1EKULg4TRFxrFpKqn5iFns/35Z5kNuERFTPof3Ian/hUS+PhQbcFzJTzjynmOnrpLNkKYEP
G2X7rDnf+osVvmQWiHHrbHm1GSse2Hn62lLwc1XBRTycyTnO1eGN/98ifrV8hdty/UfMQqAs2oQ+
tp3+kKc4hkH5+M/sRblyShhHerRvmYSRYHcIBwVm8w07OM2n8nNwTz/U5ldWNWMpAvJvMvVxkOwP
WlWDzPg0QYpAQDVRdknnHqp+CjdhrcKSsnjCKG39eAVPA3UP/QZPoFGqXbOpCru10cUNxqoETuYa
BqvNEsTwp9PWKPSAI5zNyFlZgy6th3qJ1zEsb1QWb3rD0qUud0F8128qX8iOTTLwArTcWx3ZxlNT
JfC/xYymQbNys+VmS3tTXtQZZYG7NBSu6v5aBug/XVOEnfvYD5NU2F0XqKSHSB3+AQj39k7uK1+z
b3cYqfSdVnkLJ9maO/fRYgx0kP8uRVQSyVujnHBXJRacfcn+S/ZYnOmAU36CyKV9ourJ0EOIT0Sp
iuRzesxHwyMpqCGBy8tFu2uoMEhmMy3co9EhJSXgFQ8OJfik3v/NRkH5BHJPCiFBAmhhupc+wvxs
a1NaXd+JrmLdE4eE7RXXXbZt0lYhTKSdsmH/MHPI1FuR1NITGJCA+0McvprtZbUfiR6hQ6kQFAGV
zvkW8hpdlhyeBNz05vTjrZgIM2SdN+6Gk7nFWTj/JRTVGbpVDvlnUnU6zveSVe07TnPl4ZiRq3Tw
j7rOUHYIdaKiZYL+22ZDWKmUpsHoWhY5pL6E9Bz6+/m4BgVv7WG1yLGTwGM8M6xWgdaDa2AdY+4W
UG5CrxKFr5ls11JwBdF9kcWoRreU4ONqizSj2ong0YMcrDM75IwGwxneKtTARTwwg0QY1c9wWPtl
A+ZtP7s10kmUNopIhUncv4tAo/vXnuix6dmfoSiu1BFO5lV01HzA3/f5FgTu9jopniHaz/oRrAnB
U3WUqJ1KkGbPCPqa+qY7VHinWsWtsTSy1dr3j8fFK+O9nea2CqfGvYZ/S9iHRjtEncDw6bdFLqWp
QlaXdM1y2iQGq+PfxtYRGUC5EdF1FFJ3fYNEqk2ulhklfp+XNFKCgfo2CaLx2zKfDTXb92VHunS5
34M3htCIV0PMSh8Dob5T6NzqTaFK8hQ5vlNoy0M5OdKMGOuZW7GCkJAyIv1veRMcqozCZbJMbdv3
l4iXFl9ckTcYqradItzNjSXgHE1NLQhhl/ij9BWUwmgLrwFOelGfAPvbc/NgBNFlPtqhkrISkm2/
YVOTTi6fINeOQw6exqSGYIi2vBfw/rv3fER2qYWRcgDSwNm4EzyN6pVHWOAyFb8pR3LA4LcKUAxp
yjencXD7OiPspVa5NCrui7G8UrQH1CFobJ3fEy/MUSN+o6k/XQOAlQk7aNUjfDalfZa0DARj5rbh
SVScj95uVw1TJcdP8RC3h9ymJAsNOFGUrxv4lrGQQRyiZwa6nHyfkNCqeSvyR9tuU+RRG8lyNSz0
OUEsWCm3RcCzGrcWshqH0NspJP99t9BoYTP9QHYlrvxoLI3D0jnhTweIeWfNbJBeg2qLgHuycR49
Pkm0l/gu/knt2aRZeLfn3Et/ZG410zg2S+ZLguc3Rf9VsSC2K5Yy8HLE/YkIb20KNuS/BIaoC7Q0
9u08SDvXgZIItyLqtccVFr2lnLrXETH6FMQSYUFaAvh4DBafcLrZ2cDfuiZeCyKip3IlQfINxOf8
LgZ/1FJCUDzGTScFdL+AZfuHZSLKzimqFQqIoUGLIRhNCW407cYy4ltlIv37BO3kmveUkGSSkQD+
UnzRxZxol4IReriIET+G1FEkdlmN7c0zhVa49N4BagmaqshNR7Sb7u0s7mQwFpTlK7lgeFF7MMNS
zsIEkJ3qYFg04VWvkR7e+IYgR3kl9REes9nbV16iUtDNTi20CGBFAChpruasJQ5sXWi9BbH46rHa
qBveNCAjZAy3lwB0une1Jyet5oq9s0W5wNRVICRYalscFFG6ulq/u087jnT8kdr1dxyGaQdtgv3S
jXwh4sR8PGHiypse++2KRVCc6JihwFWmar56VRoGK/LmM2B/o/W/bq5jJ1hMP06bBOeBlBJkkWNE
ck3wdbO3gIy5SHcz8kvFqqfqKuUTdKCAdpslhAF46XF+R0gIf/0qCkACwFasMl9v6qRrJAYy8hWH
0aRPcw7bEDq7JM9luOF1+IVF5BfeODEPoBeH7McP2jGylAOdUQypX/nf1YqceR30TlmuKdreKHxv
MxxXkfcmXlfwg+p0LFvbAjnUUNSzkrk4kA6N5oappNgfCOjHOllGUKRRJlQbSUIyYIqIpDvuMA3P
BSqjtDDt8t2OxnpddHKBP0P6U61nLcyyOgXBCsV3xFYsWxQKbyktBuFOpXydzpEceabKk/9bdNH0
R6Qz/6O14FMLvkRk0B2Y1mOfmQSQpxuyY0Q1Xg4IbZgnvfA/plCmVCHZzPAUdziSuOpnJUQXIycA
usmJgWUE5uFFnjARO4max/2hw5iyZsNyvuSv/8eVfxF8IRUpLF+hmZu+HZgusfDPzaFSDbylvbk2
y12qagwE7UNvil6l7qgrWR6T+wMv29MnAnL5UpeiakJ4ezva9l3GW96ZsgHJX1c2PLWOnjLIGE/3
84PvH5KfZDOLD+qKLYUxUCV4BXAVCHSPC3ftF1E/dpNT+KSlYsWCAcEnH/J1mfhkxBEkM+IT4CX2
ufWaFmIGBZdHfBTnEXUNQlxRLDD/z7s5JcOOP3Tx+bi6NGHMWFOVobEK9GBnPEoe0tVKGKxAv4aW
0tMGRKU0O36/KnqSyrKbvO9ua2JQ8Zo0Hur51bt9Sahpqtiv0Pr13pJxek7hFimMlauFoO1WvMUQ
gWks0vd6ELNU7Js6bTWBUFKLA1wVIw/QvhcnM1+9WhgQdxSDtcmTVcdlclGoIxvpv8LQyI132Blo
y1K4pSESFgBF3MJYpLgOkwdGHsOBbPFEhEFNmRdrFwIH10z+pDv/zgS7nApYK5mzr0CQejB5uNl2
nk7xy2wtXsMflR2Yuy5mPaIqy7VaBPBoWBr/bvlY8CPW9mLfVVFyPNEVi3j9dJoUqzTVccOMh+i5
2lOQm4Vj+4rqJQJ2b1/rjN0snEfJZH3hvpgmZoUXIE/Zl2NJirw8AccObf3apgrAWJBKFFm26JMP
Xgq5NSe/XpZlmJaAYeLq3GgUYHe5NMFSe9rt6BGFqCnkN66pyNnwfjpaRlGVlLVwAuyK1/Dl3gQu
Z5xg1/r18YpTydGwnD7ZxFjNayyBalEvAg5utZfeLxCjjNfDKMPN2wtiqORsBgsGVkZC+hmjURLA
JEqd2F3rjWDykt0Om0TH1v6lDafWzObKPkDpKclt56O9/UlEB9MKxfKJfFsO1RWY5NHT36/F1IIk
YikvJ3nbMd8p4tDeqPqL9JA96ewt+/nEPhz4fPt0+XaMoIbJzkl2k+8PUmK+SqwW2kz41lVnLt+F
VNtz36/Zll5FVoDMAtIyyxPXa0w2sCB2Yml9wI2QEVOnUCMuv/RksIaZc7/DczZWK/zFqU5+4n6Q
7pZacXy0ax5RyfS+cEJcINMtilHgu9qc8puXkygEtBCk2Rnw3AFCPfKevnmeb42GRnGJISHHLOEl
8RfHQjoaJUe52wQ7f0YXpuooC1nUR2iis89elUApH+EylNWNXkayClqaIkIudYBn1+AwtS2mvmRO
ycjEpYeVFVj8E5LFxzKaN2h/Dfcbhga+vvZzcYZyODKlDShU287ppRVQZQ1Bv93apslPGGCXQehj
WLaHQb1IACGmmdQRbMyILl1PNnooB6WS3BrUe10Vh6CoRETN/jBiATjnzmkItTEWcemt2hNpGqmA
8xKlNSqiyXNTAsAZQwvTgZ1V8d0NslSbkKGDXu77xrgKiaN7OEF92D7ZGA+U3WEHX78dtHRuO8b6
bilKgdrL/4JgykGGGSIjpdLfB2IEO8rwdQJawlDZUeXyuA+XgwuDP5gTOGwk1H80CfBzjP0WICsj
a4kyjfr0DqCHhjpqrLjZu6ZwYFLyZcgqnbewda7/Gcbnj+FS6MMeGOlIDUIiVgII+4VM1KT6ETQE
0X6ApXfCZxMVyrKZDFw7aw4VKQj9CF/X5qwXLrf+mYy6+ai7cEyOk6OvYKG4aw5TfmMAEXKcpZUv
E2THq27gmyI7VDNlGlsoE8m7SjTPY04qQr5vG7IP3UHFBmh0VUYAvZ2YoT8ZEFB5qAYw4Dquysti
0cydDNTIGlHAmPBCo2cMUeYWmajslcZiIpsx2RPIGWMxj0fGvVnM0UhAvCY9LSlUdGgaZxttVpLS
qstAsHvD9ZNrCd2rU/S8ONiTwrw7E8Usbe4GObvRj+R1uE6GqyPB56fiSDTUVA1AhNhLif1yW8wo
+HaxibT8DJnb7vZIigdTJswplSSyM3yRb7dMg9+uDPaduTta42WjsnxRVVZwLdoS3XX78SChjdiY
u/L9581/4f1m48sdYo3eiR+lLhGDYRQBh71W8eTwUFjppN/iQzMkTrO9/xsEp1Xoqb2UNbamv356
AJdInGY3lIYmgPSCAQABPHibQO/s4knaIRCPfthenPn/raCT779oXRMjM1y9x9Vp6e6uvlepkpQB
GqNlKlKQlVN8wrFMj2fhCtEBtIgVJ1mAiHSMk6rFykgbz4kjatmVbKgL7w5eLGBSbHsrNYaZfuJy
SKRAQv0fcoBQaOBCY7O4Xx+K1JXiDbo6FUtqs9JRFseAfHev/o93liF80HIG5hwfUnRpgh088Pnz
ir4qqTEHNZr21ISb6NzpBIlGWoBwddp2CfRi1WTlH281YkXYl7Vba2IGwJq0eFBYKHM2JEsSVFoq
NGWtz2UqVIUXV7Nf5092LQQ3YdYEcO3lmkYy4JKAOftj5KrZrXECIbLojdBpwUsQ/f1WpXHZO7Xr
ggAGVbhZPI9robTYyb4OqDBxumOw7zh6HNQ3Gljvf0/Znf1fPGTjhCxPrVbXHSCmEq5GATq83DHd
TqWfCzbQWOaUQJIx4hDvbaDpIw0Udo1MMmSzo4KDJfePDSmIPMVDcLM1Io7isyNsa6YVW066uGBV
KoY8nnbZcstxGpwhv1tEYihKdClAzvZUmaC+t8149oZFrV6sMYtoOvFYUTQIh4UOP/nbS+aY8clt
M0/KnqZ8Va+MzMMKY5oT1Qavm96k/ey3FPQMaFSD4CjYzqeOjAm6eqeDd1CiCfLU0ON67Ex2mzHx
4Ev+Zo5l4hxGTUAaQQdclbf6HpNojnBHaLBgHumqkSSd/XDNFX1eZzgD8ZQh/9jIBs7V/bLtfDYR
F+a3QauCL0n+J12QZSMfMSIZRxozxbgnwp9YkNw3JvDXJ3UvvzLZe5TAf/1nDhUEBJP6JFvp5/7P
0oHIWmgrwiCld4tl5SqcQpZnWYA2lLGOS18QXbXegOA7bMGFVKmDLXT96jYZobwmyBwU9a1c3u39
Y8idz6plp7Hf1r89KkcdCGK/QoOVUk5hR4VjUW4M+Vh68GhihAIgu55uYzXEt5CZGUE/IXFDP5uY
/CPmj+o+8B4njN7265AJOvGa/YliIGcGZjpzuoOnKwdLxHit5gYcEaVldh66Bvk+1RSOSb6SSFjZ
/MQ3JZk+m6tePotoXs3skHzN0+lchyhEvU1XlhIezsxBayeYG20rKg2E7oFYHoKsETYrZNOEDzsm
dGcv79DrSeGtQpZz6LzCrq0v0Y1/gYa9RRPaExpNhtrAFPniNtH5HC7iQB4+6HmvHNenM/sLBY7b
93gXY3HN/fk4KiipUqCPP/Exa84vKgH0dPnHZQ9SSkQplK5yGkzi74BUD7IBvZF78+Nd46ZgeUKw
PLckUAdrCR43GjC4CoBdY8Ozf2hz/a/sVxp7eqInrnQH268aVBPQLDvNyn3nThu869+hYao5drKl
34oJzBOkZq1Sur3ihupkOGbNwLkSsUyGiltVil59iTBycur5Yh37QJ0dP50MRv/bDcNsNVsksOHn
lCH4fLxPMDcZbaXm7nRdW3MMzS768okXRMJs8uLCwWnNmu4TipK8UvhtZOKMURjY6Vi94A8X0neu
ybMlIxJnd4vyhE+G5xZOInqBy7wjChimG0tB3142/li7e5LmXUkUxz0mA6+eYvUffPqOLy3tB1OD
1kBRQE1TW+CchG042pjp/O2sVf9EYDZvVNCx1UdD5maNE4qXw0pY/d2oXzCiQ2IgBqzxU7iFuVy/
UBVPFHCmpF29ANg2L0jVs2tkAPk1ai5uInedCNcbmERM+iG7zcZJ3uqvKieOfK1OK8YCPr3N/hep
xyr+UIa/rdBYppKBgt90EaFimwNukYSuzVuhPqtp0Ez3eu/uI6LclwrLouXdZo8pDDKCHwPgwX8I
dOaWmvzgBl6kFlvXsB+PXDTD+pwv7YZd977vI8qhsnKujkGYMuGKYVanylFpkvNUOrNQKHQg864o
DVsCg23PUxXYSaaC0dbLndNbgwSicG+guh4fisgWgJvkPlWkGY1j3AbL+JkPGqAB5kM0W1v+nER5
xDgiKSxwU9/q7ojQGoHroz1g+Rc3sJ3kXyomqNMuZ5mB9bwFLJTKJDN+iRo1wkCa/AhCrKLVSlYc
KhtmAbDZBkAxoYAodmqlrA3EATugW7jZrKmOrO85GftfuuZD2ftGBgX1OpsUwXM0qVG052EdfnqI
D8tAHcKin2IntgjhPtYJmHXVWeY1mdUEQfelRrtXGgMSY8T9MbmY8rOQQljgP1Pk4dXMe1f6u2dy
CKqEesJ6U/xtzJ2eOtxtWW+I4fWkPv9kYgvnncXLfjwwHquW4hXa8GvCvNvQtnwFPCteQWjSYej1
/Xxs2i/q4qNCVtGn2FVClLn0WCGW2WMgz0tpdXN+qf1FMSOCOuazCr5hXcDBHkEBcye2DIWOaf9c
+dgsPtFkcyclcD+UKRGjZHONWfm9ctlADVEMU1Ok7HfK0jCvNeahUR7A0A3/TdWmMql0P+aN9gNW
GTT04j6/0iH6siep2XvCVBMANPjH0ec5lR1I1yC8VmSMwf5EjdFXrRm9LhnMdelsCXsnpPnrFKJr
NsfTLz2YUuXPHNr6b9teuuTqhSoPgAcXmJPjWprB5EA6sR52IviHWEplL/Dm0CJ20XVHva5qtjNL
HkamQMXSdYmmQXc44gsBKPuTVscdHIz0ePilltVpJqP30Pklcnr417nL6FP6Ubof9NGXhbBo9sBR
F5aqHpigV7Jfmx6usNNmDxOCZV9ZYdarEG8+/RF5NQxFox7S+GLEQL4//RQmgM839gR7ndUY/VJJ
FdFuuIGUgCrqTRRQ/mjgc8DWaeODMBN9MZFBZjBJUR++HoXcy4R11SevJcBdrwtp/GePcL5E+yjl
6ILKd1OGY7aBP4t4m7ImLwkLlxsSnfMi8gTGE4A6iPO5rYBLMvJm0AKRV/9XzJomGXHbgg1pHf6i
TWoTwTl7aVMRQOvKeZCWhrM96EgaVUPg8il4bT0pM060/0Oop2NUfVFo0AgJp4q+IrsSYl54L+Rj
2LLZcmXVHXC0Zvo8HY92jArtskgI0YYtMHc0o5AMw9ic6HcVYapuSdb27L0xuLi1Zi9toB4e+D1I
3pHVb1QIwnBPK+PX7OaBRPBS3hgbmNYxOf+bs2Muwj/25th3vdZwtrOskW5q59AnRVT7Dii5N2Bp
RnS1ew0+0xlwPCiFzttqumzCtLkkei6su2r7c1+LTvNGW+8pdDlvCpD7u3utsBiqVjtDGRVpqZJg
/eIrL4+oM1j3A8ceh4KTRaX/uK9fTpNJTC72xiqRWU59mF1i6FWMPwIKk3lZZw/303+XRKZj9Y7F
uwhC/C6nRfJ8NTM9ktKEP6RfAMgQQXTPYSD0DNZfeyZ2sulVsv9AN2V2JmVcXLuthu1+Dkb/jgXu
3z/i4MoG9plwSz8Poqj6pCJnYEwCOvriZUZ1IHICdjbDXwvApxUfRl7Xu8gpPujFujWSe8bwJUW3
PSFMsZgdqWFI5i2mnewHGg1W0bBk8ZGRv8sEDsbnP9gt5IhI0DuBgYOBDNyI99f7WNYkumOvHL2G
kHqRm5mMm/5+Gu3yfp25CsRyvfOSAPBBOtsQboIIBnXOHoFxiuCISGcKC1Q4fSF7sUg6EuWf+8iq
FFDLnu+nB1YpGtFBsNChLgTweuWPoJcgYhTMtf9Ao7kJTODBqtyFB9DE8/nsKp7TJ38oI0p+SZuJ
f2wEpKfQ0sWMW+5vZa8DMAhMLFn02y9waLGqOlmwoYPUbZPNH7c7Tdz3n/xD63grrj1c9Kfm3uz9
AUxqZdQ7vhJjObu7uhCM6ZnQfcqWevGFcucujPDzgkHXX1FbjoYP9PlLfZkhhvoYSvVzXUtihYrl
3m9ASsZyc1d4LBICpwYsU2GX2UBb1MDkD62Y5Ms8w3GXsA7mUb2xeYK5qTg1hG5kmHU5AggOC7v5
OKi1X4Ss/de/sFIPld01AUHZ1YYRk0TCDW+qQN7jPii2lr/KXVL02XQBHYyPb1BzvW8RWZB7qFVq
IhGtrV+5pWMeRQwkrgvCwN4+ybKtG3QNFfiKg2nUTIlceyrYpaL9WnLDEAdLOTZn0odw2EKImuKb
QSal5TAUfW5W2uTLtZ5RXfUJPsNPQqJsPjlj44DHMGFcEeIEhSGblPhuWrk76+ny/QK6QK7FkHtP
2GZ3qtm5V1Rh4VqCDhJccmdeU80l9j9SJbrxrhkyq7bgXUrbuXUhfTLa6As281QsBrAHJIDskuMM
19zQ1CcZKqrs96Ec8oRUPAuLRY1+6W5ZI3PgGnWyT1kLGtx6fVOTX/aQwEVo6jqt8xtm+xPESurt
eO1SHOq3tJ2c0eRozKnFpbbpVfs9CRBZCRfM5mEVPkWXUSQ28oQBNjVzyJe/pw+7wGXovEa6J6gt
f1ZtGUEIK0prPzmupRjZMzRNnpc91C067COGetK6tjDaqe+bZ5kmkaRDtewH+mTzpM2K7JoniZgb
oEuvAFIz/crAYEpT6nc1/jI1qOLu6y9f6zgZcmeQ57ZuZZud4iT5DLLqWpbbBLWlO7o9YxvSaaFk
/rF5ALVz/k3J/DU5FAqKse/ldyaSQViuop3Jrzbz2UBDQu2j4pyAM2L5McPmXZl1MfDyLASAFodN
vX8pFK/ga4uAV1usGyNSUZk7Uhq505gMurh5R48/3Jm/5UOnr4SJt+9H/wqVSjk5ptllXkljdPQR
ccKvpRDY3y+OfnzC5q726HfgE3z1z67CUF/mD035SRJFmzIDvLxxYg3Amt83efXtTZiueNJyxC8q
kjVqP3KgaoviHJ9YfN7PedIhOQdhBgFRPQ1W/GiBHFbJd7lzpqg58O/nlau8uUkiTK2WLF8NQce4
WOdZCE+I17OpJSsuMu9pU5rSa5e2Q5JsTfWmavpzSsLQQY/HbpTjhKV3eBNCaK7ccuHfH5Q9yk9H
fz9+suN7Mek3QviQSayGPawaVOy6aqNnyMGH/48yJlwmJy8FBIZFHaNoqgYiY8ns2/66WA3CpQZh
ZOf3Mi3vhIFp/YGevVtE9Zr91h+scBk9x+ywsdjmAdHTdE9mlSl7oPQTuIlsoSqCm8wrgyIwFz7z
0EUEHP6t9HFTyAKhWK8MC5ekCmsA9FVfSrx8lT9rWo3atlu5/uLfkXR3jkespNXQ+oq4l2m4tXjz
WII3hH+EveHTLpDazweVj0Umd/r6MZCNyZiyepfrsv09e868d7sh233zAGg3d/XmirPviYDuRoOF
FUbMiDdvfnfI448hyuTHtrejcaVfbpRJopMT51jgbUmreD6iAPMGV71P/TJzMOiuc3/CftL2R35n
GADewMzgVqwVzOJG+UX40QSNw6F13VDmYUDrYdabBm68HQwBPvl4qLytOT8t+xesvCg27yrjeIY7
rvRG8ftabC1xsqcwg4cdjzyC7zmKMZAbaderMlLAmA1bm0KyMzGdBalkzoOLE66SJIEvgVaPNPA+
EOXai48p+W+OGeQUzbRXeOC4MOn1BBSUM2hZzbpOPRwzEIOBGS/jrpdkdhjr/kf/uFRdaQasG9B5
Qyrt1/e8wg4dF24EhX2f5rraKTFSHp7niJxAoCDdJR8J7v1T0riQvjBHs/StDcBZ9PrWjxE6bYw4
1Gawraw7tkVNXuKdbpD+pi1jraTBj8u9QMAMyQJSr9Bh+xY4YbtKZYRBa1+RG7k4jiAvmU3sCVbx
tT1nHKBmnbrv6OeiPrieUGwns4r3tIe60cIvqzi2um6vq+pBAEBlgY2EHwhN5/oKBg8gYeo4Cq4N
nWEN1Xv7TTPVmny0PZFrxnTTRz/38w4cnoVDBEv7Rw/SVx1u/uTssbBIDiGpXYBA+Fir1o8YL85F
OfZJvquZo8b9yHZE3P0aoBPInKxWT1KGoO7nyWTd2BUWj6BxO+b7gJ5SKz1JW+Ynowyu0M4Xj0mK
IuLd4DdTpO6daI0QWDbRYVHLU3ozdOYlnjAMhbZq2Fmp+3A+A4L4sHv/Ttnskt4JksJzd3bvxcFm
c8pfmE4pD5rWX8F8XvTB/AsObjZsW1F9Q907EXyJx2Z3upQSmQe6fTMAIDH07pUWz56dJrfl5klx
k97xbtNxYcuN2hL3SMmH4/grkg19uF1HWqgVA8GnUjlsJc3kxoPk8hjTOtJq96og9d+cf9ufHV9t
Pck5jaxxZf4EM5Q0n3B9k59vqqeHzYC1RaBqVvRM3G64T8jlzBTAJFJstTp7AEF17tu/TYhx2C2q
lwcdmC+0A8QeZu3tT/SsYj2G83boJqd4JYmGiCbzojjTw5izpM5lkLzuV37UHxDuLIRxXnlpU0Q1
iqaxo51E5fO4xyUeGsekjCE4QbsVNpAuuX1CCJ/7uULMdBzJjn5S3anD/KJgiH2q4LTkDUP1+iQn
6y0tsxz5w5nA0SJ1/JoEWA+llLtA5Cw7jYa886A9FAFQdcpzM0XNXCu8G9bPIAdaXEoJNdiZGAsj
HBlrf0qYl7muNJe3FoqCSfp/jIG/J2X+RNJaM1xkR3uL6yTLm6xoEqTj0ue9HYRs4/hIjzPv/+Gz
TxGMI2Pc1sOnmzGKMYCXekLd2dXhiqeJX+m9jsTc5NFU/T0uj/UsGyx8m1KK9esobSjBMJEqjC82
ewVt8r7i52EbXesLFQIKHhpXK3e2fFRWbZOY/RGy7aPOvaDqvb/Z+E74o5VRzKR1zF3eg7CsD4Zc
HWOc7ah1a8YEbXaTP1pKEQrCyQk/vrgEY6FT035rPUcITAM/jpGpkd+EDqnA6IRv8Ij48kIx2WMY
WFnYlTsXQWSzqK6CE+B2witIjnR6K1q4zX+b7D6svkUXWUeNd3/eQHn/HNOY5ixBUYfNU7rxMdhv
LQkWQ8iNwu+c27ktPfwyshQ5xBbOkTqsyU2LmgQ0MjZLW4trvZ9lDmRfK2CFi1tZlNCvOr8sWjTw
o8fdbslQ7lEJyresmenAB1XjQIZjJoiwTRNQ/uri+LlzQnRkrjIHYutROAHEGwdZ+HVcEaHhT7xB
vXh6jIEJh1TnmtIFaptSn1ExFxX8TM5xV+8PZVqX1P70ORoY0g6rXFywJnopoqjqXpvYPjU+I+V3
1s7kzHVx/9bkimSrBKV2f1/now8o8gEI/ZfyXBaF4br/cuVfLpWAxCyKIynr6GVHjgVEWRm1XqPA
zXWkdiys8CIgiRE8pHlUE292SONdLz6fCsr2KXc+SNMHIt82zqyaazzsfms+XPOy9MqqFnRDLJtw
sofOqZbvD/zjUZaKrUJskxDeJ1mRQZHVGODgA22BakrJLTXfhHxjSfZ7IueeQjAINIJ6CebhDMKD
f45HQL/IlXe+hA+IYqsJHJiTm8nQHspBIq/Ko888gJe2ILVU1PHderrnFAxkGYvT6O9mfhUwg7n9
qnHyy7CLWuq6MQRsNMQxPh1rWnLiuqXZNwbEMwbfqVogUrvECwMKGIfzmuyy2sdf3vkPfT1dq3X7
Psh8p6Mqs+JMTE0lt+84PCW88Nnp9QQ9QB1tDgdTL26fAsFk/FS2fhrkmsPYEicpn6I8jhJPmSe4
LfVm5ZothuZYdnVj4Acbvfs8ejYuzuZGqcjHnflWln3G262C+WtyOCK2GLfYC/45Q3YEVV66QZFx
0Q1po5JNYbXpV7xQR+P7xkrDsQjbDm8mN9nNRQwR+oWOP5iuZiL5SI0kTnqof14xikxGbFSeJfIM
N1Pkk7G7zj5VJ7etxM50i3+YyzGd+2bo2DX4T9YXw5SyUnP2Nmj/l7r0oSETX2n/MCEbSHFKT/8J
FD8omwCfa69aUj8VQD3vPCUH0lhMxCf0R+XlO/ujfmaSmSx1kUr0K38sGvKPJCkDv2mW5Mse8Ymd
HUHcGZO7ySgh5x7tfdztSIzVL3hxDsX/WoEOPoLdAvD4FTvQ0tvj/mmO3IzAtkjarL1F2/jctqxh
V/3L9cqxC813Yp636slHWvIdsRxJeXtAxbl6vavIoOVxp71yIUUuKnb/hkkXOZvqHsKF/ZwKKw8C
DJO/lt5Nico3owu9NxbEr3zCDES1fixKbBfKpH2iCzh9UKBgqrUprSuo4mqwKGgAvClovp9K9eaE
myOZXNVro8OrOk7zs/ZDPURTI+4CzQUMEy2zcSyxFJWnu4TF5YdgwK6vLjmlcePiJGeUhl+rGpAc
6CmqmPz5nn6skqrhL78IE+muJ9I+3XnuQV7KTPIak4PFEIm0iuxK/4huOTv9RABeNFt1pB/awJAx
JYQ0YIeHz/PKkp4xEHQ2oGBd6Vd9QVQHkLBE3kEkzIW/zTmT1AzkjxuojG+8eh5LU9zsc/RISCLd
VIt0Zwfo9+ZWAaNFaYbIlLuI/gZT31avcOjpDm/1JzaFfsO+LsJX8fmMUUo9SVsdpmWnvgBiSwhX
DnIVkL7ExiI+d1aPr0n0F23AQMsuMR0FND54ZhXToOxMZigZxmP8/3ub60dYwd59wkv1VrYPZ0lv
kZZehKlwjZ9kKvVqLHdLHUNegF8IsFoaq2+cN7yc4KUE96l6IPRglKUXxBUoJ18GMwnKS2pXvzYb
iFt+uoJxDH6OefLBRxDKf0nyPX5gu32xL+35E/5+l7r7IBDkbWBn2JgV6F9UBa3QH+q5mykmKSc5
/dcrLg7lnFDyL8FBgne7NIcFNYIyZkPiMWs6J1rgyatbxUJXjs2kEL41b7XlItu0R++J7A7OWpdX
ihmtnlj1QszPRjnkA/pxlCk670Vrg7Ps+bftjz1MJvhjytv9S3Zk0h1UgY1SDXJcD7aMznCOJV3O
CAIH8TBDrgzMUPrLNgz+Pr3zw2u+fRZeNmhf0/4ZZQ8FbpGw6qs6vtimFV1Xt22SBEvPAaJOS++l
lw48z/qAj6qggWfmtdJ7Yc+i/L2Ho1r1YDal+o3owPZpYePhG4MTUEOh07uNgst9bzxz2ldqZdcX
P8JFNAS3wx13ke2a4xPCiCjxfnOdYEOFIz1SjPsdF/1vFdIkQ+0AMo5/8TUsLXf36HthqnEJGlGc
5/KvBd8V6KSRkQj89ftbJ9rOhP8cLH6CQkBX4C/W/k9ufh6pnq4APDPZj/3O64tS8+Bvh5JftAWv
Foqm+axuVODjTHoERfbgKomxLnylYGeaVdCReGNWMtjq+xn2I7oL+mnI4yuoH0A471cLGiRbzagH
kyPMrYQ3eOmJmMjQtJUnqaSIGRQpw/mpjIITwqss14hwgEfyiEFpKCtpB1pGrX3yjPQ3AnQ5nexa
gAftxrCDuRcX5pkKg86aHVitydtLi61UFMGwu7srNjJFry4Dblbz2VdcSiYcnmxPG2kbC95FmdI2
yWELy3Rmbx0n4v92gfs5sAdDsfL09C6+P1qp8pTeLmFa6yoyzW1dkOhJ9VbiBGjVic1hSx9EVb6K
rRnxmPgBeUCHmzQs3hZ7G7Scs69VLq5bQ9KNG44JLj4YuiQoLItLp8QRuHurjk+QHGPzi+HaTW1V
99mv4mM0LdYnlQMx4bT04jwRwo3QxFdpYHcBmPZ12ksMnZSprASZCjR89qA5q3O1tH21Q1cz2/Qz
8wfIKa3kbsMUBxpRcREmFHj4dj8WSiUeMKA40blr/odbgouvYU9LQDrLIFQwYPHuG/FYc5Ujnbzj
6r3Ba54tPuzHrUbVfBPW3p8dJho42g2D2M4gpyWIn5hXPy6XMWlSR+7dkwikCMpvyEyEcqntnCA9
XA9u4eyWYxhiCnWvMO3jrXDRCrjRBjLTJtlM9lsmn+n7BAgHwZwBPmPffPBbA2zhpNb7iVScRXOu
5YYAqkaXCaRc3fbj0l8r8ELNUXeU6KJj4CbUggLd/NhrJFZleGzlk28pdYnkVGflMqQMkLnw42Cy
PrbMbQsKx40gJPl7uTnEw/slGDcYXSBEyLu9MlL3URw2tlWKFkjLjudPVOQnNKjtCKA7UzbrFeKQ
T7UU7ql1MIr9c1erTqljh1eB+RS4ZSLaBQKLeyVNDYp/KcGe3crRam6BkcAlD4bzg2ZJoQdMREic
HlPRA7t1iSK6JDAjj8lHBXrHprTAQIDy+GTTYuEP3zj/zyO9+pif7ftlbPVhKmRrtb67Qlv+LEPO
YLKT77FSy2qVg+Dyj6+oTDw2t6K8TQah0qLBLsfYCdwxOMhVAbARsSCGZYDOx5fFgm4DLBnTz6bz
UthIV60jt9p2kTRQGK4jfxUXBxWiFKF50Uy2S6zc0xWeecaxfL+fx7+6ZqW3eohaSbeU8qPIjDx/
UgWeLihPwoT79FSISsHpECtBsp+MmxY76k6lTuk/8XhaP+UtryDPpvZo8Nb2YHMCDQZKQbGV8T6X
ywUUwcYk2qUKYDmg0csqEstSdfofazF1nPrqE2qMlv3SZJl/u06wrzCHdWNPW7bg8v77+lXlRitz
S5fIjtItsEWyOptyepBzQi3GwJcJTnaFaKUqlhEL8tzE1sWrCyDnHap4pGVSubHp3/9HvjZtX7Hl
PaNT5t51O4i5hm4UwQ1gZC4WHLJ6p1Y5oPZMVoxWw7MN8nSqHJcmXyR8Gt9OQIeRx/HAuQmR1HfU
0uTtH1Dr6hnOFSq5xuWiUtlz69m672iQoWZU3tSEpVLws2ZT3wUXp/kiI+7MVpEEOoDQKOCbfaiG
a5DgaEOMts+fPZma6Ey56ZWSwhW9xybTH8Az4ORWJ4ZGIraHf82nBreqvdOk89odGnlWuGaeByrX
Q9y3hqVjvi0MpstsBO1TiqZvsOjj64YRCZlUZGgrBKkQw5Zb627OwD/8cJ4dgLIs4DyUu645rBQ2
ORX98Ax2gRAe6uQPlEXv6i0u1KaMGoycLPx7kEKtfR8PEQR5NkvhTKeuytTbL6yTbtzKi7ZMOPPT
D5SEAsR4+VaX2IQS+KRTxk8C7s9+8fHsLG3MDzZe6RSecD6fszVzqI+17wP+rAEfuBRDFvDbPN+c
tTbUjyGJE9ZwNklxvruhxKMAuBw5ugQ+vPivj1WjlDq1GEWfsgYReU4ofW5GZ9/0IqqJ2Y8xv4gT
a4LYHHtytOsmPvs6AderXhRc0HgsQl8e0qKdS3HTGDgm6p9aYF90FlLJIdlSRn76Pe5Y95h0xPdy
5t7THRzJDDP0yly/KOamGWRaj0djXxhusGzBm4rnuPkfU4QYKjc590KaTV0M4bA8I8kREU1qKgVx
BZ31IVwEW6AeMzST1Q1KoWt7OMrlcRP8oDDGjgmb3Lr2wubnPx/CsdFOaCCwJtIMqq2CoSYgL6V/
HNkFL9JQOp3jPZxzm83g8af5xcm46i/KgHxYfK/WteN0YZRBTGLuoDbdYr9sSXMR1WcoTwrcPnQn
IsdeTWGjyfsBrSNZBuGRUObg9ob4BxGSwzd2bIe6I1yBsssUR5vYBLaq5k1D80tlYaVI5Orn/zgT
8r2dUoqSENWuMqHWEQ24sMckPGlAQXRChPO8jYK+w3qrzPFH5aNltB0fCBZHWwpOlVJe/varU9cb
uM/Lpsden829J6Bjom082fp+Kz6gnVm8MZjePDrM4IUgmLdQSO18yOoWuwFd4QX5K5m+BXgCHxpV
VZzq0ovLW+x02MljYSkjWLLCql9FqnFDOsn44EF3AgJ7Pm6Kzqj/AdBzfKuRPxxMR9XqZb0GL9t8
nnYwvBCRHA40o/N6KHs4L+M1Yy35p4BF2qu8OQqGmu9T9jE+VprBTIJgYKw1NGQsZyyLTsC0f2k5
ZGLu9E/iOUbeIiNqLH0hJ+eSLSym5av8vNk+equKyQZ5pL5B2OOLcsEInxTn/4ROl50ONH+wHZAc
CL/juIFXFYOVTs+4Hik05gzCDQdoD0WYKdMMm0aiUbzTl8Xk+xDc0mT6kT2WX+Im4bZY1Llp26Ab
NDRHoNqFlkAhuK6c/bCBEHIYEfgVRPy5OxN2Z/+fJT/Yb0KWyH0zxWXG5+hAijn/QakwUvVDl1ye
WvRupI8dnK9xQaCDcrYu8zHgNYv2hXXDZ3HXp1iarYrLUv2ccFamdmCviIE1S9cEHbaajNV5EMN4
Gf2R9RnB/9OetpY92wl8kw4NuyLnQRiWpkNe1UEOaNXI4/pv7Q1UEwdYG4HfEKqlDY+U70jl/2Qj
DX+F53cuR94j0S7e0WoUxjN9lbG0GaE3ZucxyPRNcw19HLh5HKGlxQJ3BrhKblSbe/oD/hb636cA
ZL27qDo9tZARVoC3bEDDRbeBIjZg+tbET/INfinBMI93CkO6lZ/fwY/DnGpnOnw0OZ33i6nYupaP
1vJ4yQCV/jBXyFC2K9BPVQujWBd7ri+aj27/phSCCjSGDWTq9etxeRV5dU2LhjbI38YzX1AA3058
fDk2WcclGNbm9aDGyzNunn9d5r7hiYeIDCQYMw6DowiIsY3Ee3pqlpMptVWnzkJf2+VkuNLkTx0/
MZrnV8nGynkvTcV6IglVEpYPu/CS8Kc69UNz/Xb18an9x0styAJ+6hEG/9HlPtuQgpDDMfZG7Ljn
I/BwQejOP+PMK/+kl306TMPDGaMTrNTaOIKitocbqIkcXzVMHMro9FxCoqo7BX0YNUKt5trPaano
AQWwlRapEY4q6s5c/zOuy/akUPsKNDckLVNOBjjlBMGllprrSsQfImy+sfW2ly71kYfg8Ie+TcHL
99f0vv0okhFnSC4inBJc6BnWjVQYfmu8PnWiMsEhriqoAYQXEHO42k9VhjoMZfmnarvHLUlYUdc0
Zi5/MTHXlzzHvzVgmZ8udyyXNTHJm7HUxBO3Nqi49dUZ3sE0dXUTjwDgk9uhwJdJoAfAGLWUTimI
AYC0Xq1viSOFCnwpLBinJc5DdQiHKrTB+1GG8ItgntN6WnRZFqTYL2nSO4P9FAbexavmz19vNHW6
Bv3xP3S5gmto9rT9YFVzGn2y4o8hza9YZDeA58QuYR/aAc9WKcdP5t9ZYuKZhtVDf6Ey8lrcOUub
K1DsVIQefy7U6PIDaPjoc/XlnS0SthwXX45juoFOl+1+0rGQrvXR1GOr0n5vpDaFJ0/mW0CU7r+L
KAAvWjlT7uMWU/G+ayz4OArgRiDk1LvWTJgb6YTUpDhq0x80zo854/WvjvVpQuELbL11+/ychlfR
x83Bt2YgGDJyXTmowotfIEr3uGla8en4ouuQpatZjS8C0q5QA+TDBwc2jD4RyO6TsMhMirFg9raQ
txlPsGdnZwa6U99DNSXn1cNe/OWXjX4kv2APmhLK6OZz0arYOoifSg0lxNFHk3ZfBLKK18bhparD
IujLiXMZiplmEgBRdXfUkJu0nQ5yVzettLhBu7sZIOirhvvzGMZq2H4772epVCDFInRaHb9nup1Q
cLEH4HtgLP9aej0iO5rdSPbZJKuIZD+vIlqC+xYhCnfC8BwZOiqGaFRzFHKfAAYm9RVb/liWmpws
vRK9/+AJEwrY9dKy1ef4FSekJV1V5nW6Tr/AwquSD4cXy+NXGrAkMB/bq+MhSCgtXqVLanmFFeUG
3tBJbXbByXLS30rsE3aIUeJeClSE0WMBf3HiSRoklnukKZFBB8nAs7hZJqS8TsPCgXnuKdDLQDUJ
6dQwPCIyESrdjJM3mRwjVL2iCIc7VTs66Gg+NfVni09Gk4GZKMVVHRNY5XRZKqRTTxU5N02vr+/h
/W64RkuHEjCAXQNN5LzvQ30rsQTx1hWpEM9VC+FsnpqmtkkEvupLo8He99R7hDcQwJhSCjLS4YcZ
bwHcUUA6fi9INhxEj3+6j6RMDXDtufqK85OWNI/dSwccfE8sQHFChrZzQ9YpytuF1wL1HwSHc1NZ
PN6dw57U+E6YTjTkDQa3fncDmwS88OeWCcNwhrbl3YWUD8GI2Zea6ddrtWzIMlCXFy7FR4YS0zV7
CclbTqcBuRDW7W84ZI7wOdahOxQ7RlHg6HgPelSFarVVRlZJM9dBAPQCQrvO5wBc5u/dZx0iF1Az
vbmHC6CG+WQx5SR7/G8MGFFbaJKRKoPgOmt2xGoZ/N5qdpJNXrgD2oiA+UMIQ9kT0r6QX3RutzPZ
NCI0drJ0y9m8RD9INcQozprF5w2HKAwz1cqg67vUPwwd3XJVjKQ/zs+FE8PvgoIeSbUGCy85u3up
qIH69TSFVvt30M1MGYRO9CG/aBxvDphQZGV2Y9cspQu9x1pta1T/p51mzeK2s+xhztLvQAZQkVwK
Ri4Fz81qn2OtRDyenRG0+w5vyJ/uvfaogIh6TBTJ1Ofg9qHzQNu2nzWzGxK2O19mNZtLgaw/7iJ+
yzHvunMkuOj1a6f7nXrXApEzAKpU6fTgjU5AbVpw4SXm4SVetlkC/dQiESI4u9qJqLjYXRxuTPK1
4bIb1lOgxDNmbfm7dnoRI0JZDf3+3ci7EucCu0CdVaue6OPC99FvFCkpsf6n4lab7K3KBAnzPYXg
H2D6by0dTvl4SGQ1zv+71XZIgojRS0f1bnoeetSiIE9u8naHhHB4tfxFNcDXrenLAMGC71IKo97s
8UiK3hBV4xyhri74M1DOAcfQJxd2ToEY53k3ET4oKybux43e0GM3jiWvQKYNSyLvUhD2XixUZhJG
HyP6H0e1+nDJJg4wKAAYy/5xcSmfPwlu3EXRxixt8mhvv7yZCoIFt1C4mV88K1ZQaYYjWn0oanwg
87PY4AzBjPUH7isB1Cw4oUm3rO9OZeF9wHX6/vxr6YNOo7c60eoOzIwFWYThPmuQg7ESPkdNXfNF
0YzYL1R/+8hG75AgmJSxxm0wLKzbEk6fY7zUuBDOEdsr45orhU9vU2WXpXvzFiCFnIoIjT3NHKpv
Lfw5tGSB/hipZkVix2zFBFxoxK2cXLlPNUl5bw6nbi3uorlYhqpfIJiFzDG4hdfu7fTdH3SBcn2F
zE9eLCLoaQGv+RJr9/GX5yd61yyXS8Iqk9oiEcLx5ZXN2qM7CrSN3hQAB/taBUJ7gulPFt+vGUTN
g0GuLyz3fzT686eG56meLjznl78VcDx0YDvu2RK8duE6l6/CsVRqUv4MXmiyPfzPoBu2HybErZPm
nMpd/sxDlQnjwLFlM+KLpAV9X3xac1CuhCY4bFEagZ71q6Jey8u1mikmriGTraHhh796j5PV9eV0
Gd77KDR3F5HsdUKUJ4t2teS00Ssc4kJ+KGpKQQ/i4Epq70AFoGJbtjIsRweOFrPtXiYEqCK4PhNR
MwJWpP7oAra13e9p9A1CsdC4y5z4d7RRJhuhBoK6Gr652CozwljyBJ3yrkjbRMu/n6AlL33DXhJn
nzoZWX6/GNMSsOnB1+BRtjZI4REEScWyG/ic7vowQ/QkXHISBPbV9wZxE4WAgeIpk+yOMlrZW/uM
V5/MMdbqLpvNiV0/hgiY+DOcpUlrvGZdlAgb6ySF7CD6Hm6ePyy7crUNTfXh+/lBfYkkE19lWuZ+
d03lWuOooU6NhpAOMfZjURhVswv1VitZ6+Zd0bMCNm433ahH9TtgervcXNGKPVSqPo483YhTNgh4
2JdtHhzwW2+aifeIPrCSEpvEn8qVmdb5QPRMOTztPkmrEfNcqmHkqO/1trFetjQlcGyeaTZM2t2h
I59E/FDVMu++W2y4Q61ja51wVaHOWlnWfU0nXVqpZZkZMaBDNKtcCgXxID+MnMD1FVFhjFjvuaoL
cBz1bwc3+OD/4sY29aPoPeipRsu1CNwihErkUanqCXRcnLywwDAN+bY7U6aKCDvPb2pR/iR9meRg
oUvEYOgaAHz9baXM+Tyq9CowfBgLEKczgoHMjEG0d9REnuoBRNN2WZrnO4LuWmrsyvLe4Ly4zUdw
uuEYWxKTICTxITckvK5f7Dt/wQxFSr6d6LDlE0DgL940d3JTR6uMDqWQeFWtGpIVwfvDoONcjVl+
wUce9Ae1B7lPPxNbD8FjrNLpF3QX4cDTemZbLqUT6qGqKvfsWj+kwIAbVqq66x4eoKD5NcGKTfd/
n8DK8UmfrOEIUZq6UtGvnPCCTSKL7hiiNCTA6S25yzdANAOzMt4Pq/rHrLls/3ZmdKXB+PTyZblx
pyR3bdP0KfpyUYiuR9geJ01rDRTYhpXqaCPClHbTBwpZZuqrnTo7Frwu4vm9F0OPVWCh93UW8Z54
3RX/IaIewdaUvpS5PgpNzsF3vw/9zYag6Ay56ZtGBTLcv3o/fp/Rs/VTs8PnYMBz1DMYgLYx+GKL
5K1gXVMH4OjpYf/CRwTP/ynk1eDmYPdACFdsgirFLZ73hAVlth+Vw4YuWPfWsOQw1u7co/KX9+y5
0eJoG12VKKGCZYjC26C2PNjPXEfSdoc3X/zx8kf2lAM6883yQ9MsGsinxLa65yhmhtqzoZNwCRco
GyxQDTqfRBcRf8SJhQm4IKusEJP1BHC5/HywIq5q/hr+Wn59Ra9W5D4vRZGh5JcpS2r4Z8wgs+cB
Mg5V+5Ps8mzHANs9yhk4O02feP8icOtHRUPMYN47pLNgbYXJUQcpkDbVHB2l3IXcO6pnFZAN5NmK
s7wky/rXrXo9BelCJvX/QK3/ZHDUzA+HVsn85uF17h1jyxAz1au8xMC07d22hN++r+jWqLiHu1jt
N2KPn3pFYD4YYaCgrIQmYsXS5kk2lyB2V7X9N+8qRPrIp2DxGRB3EI74FEIVVO+HR8y4+FclFvd6
bXucYwiYqFmCqDx6RyOb+0389TH8tsnnuG2pYRnvwTWGBuBJTQ5z+fwL/Xqdops0tJ+OXjuQbU/E
HXQ30SAcEf4P2cqxZLoyVhi+B5rvhP704qWPGCf0RfdpgJaHspjzAZXS+X27QR2jON+MYbliKxkS
YiXqearGdw0fFjiZGtX0b09rt8svgKySwtg7aqlHeg93WWzQuEgxrRgosWObyQiBIYxw+7BecdlY
h0tQqGK3HgkdMNkgm6nIhmiXzEc36/BwrUt+a8/PLIWBcNlfmnqsRJVN8OCI1KzOaZETVd5xTrcU
sIAy7cZxGmOBOltxI6pHUjrTHMaJobleFCCCI2KAQLpE5YEQSEbPHXCmM4r4/6bhyWB86fSgx6wL
3upxpb/JthnZNeuPDMyjfE5mFDvP/D/C0dqqj0hfUeMg14ZuFVHbyPccQIDO5Ux3R4mtfRqFACo8
zRXcyvwQ2T125UA0/LIieOWh5mMtYZdyqLIHQdF+WU7SAZ23nowfcvsm/VgY8t7EDxBNLZQWlype
QkRAqupNDnzClHrjiDin3YKGeCrQwup6yNqg7/fBnmMj4ajz8Nt9YODd2Fn+cKErFTNsHjj7xfTJ
qUOitexqexN+1zLi1UXFI3pldk7mNyB2y3FbtyVj/eVbf53ChhyAqDskb7KWZGOxlATASVA6PkZr
9uhZHVzm18bGBMoVdWDqQN2SunFnLjFxKX51Q95wyOqFNH4weVBAGnVT4UJs+AJHPPsT3+KLWJH5
5omk8bWQXO378ZV2wQ5pjpN4erWr9J1wOU4vNfh3ITq/ozXQdoFJPDYDWR9H1Bcy7nemIBhtynVA
ITNzOpWbGItXPBbCaPYTVP1S/vPpaRj0hZmXzuIdREIAs81lAEjMXyt1MAXTMqGsHiyP/GfPfOOh
yNkaT66slBiRIV/9JGL2cRL6XnQg5PTZGXD0hakPjgA8zVRPGc1PTRNq2Vla3Jl/Y7XEj9jhDKXv
/FT0Sy5oi4zJ5nzOF7q7Wyj+cHzu7KvP2VoFarP1XaQdXrcaVmIaJ57Lc0XoCnxR059PLjIWtEEx
paWLO5fd4dVm3nW49qZkgY7dTjO9eJbhJ2EJ37si/VBBwVUCvi2rTux2EC9OU1tnkvFHNPSE4LX1
33cqIDx+3A3DwEg+e6KGldk2Y6x8bf365HeaUMIxkUDMu2binW+Go1iCIQWPSBke3gcEm7AxWzF+
yLVTKd0/tIkeREYI4m3CyU0meVhkwgqaH4c6Ism0kGI3MmX/IdkPtTvKBFB7XcrGt90X5X4qVXZO
3uC/jpbeZGO2XCi7jGdixfMkrrp9L6YqY8JqDlm/tm/iof7JO3GODC26JtHAoNoLVLG2iq3cxDQ1
BacDumuR8XwskZLgqZ9Gy5mazp6/WIcRa9d8MvazhtIJ29ckTtK7zJTXLy830yv+NVsQ+zLvzSqM
h+dqBz+6udq62Fs4J3weXCwPTcktv7918vsMy8TzSjuslTCpPD+PJODqndHcmpNuJ9QuaSxw3Ffj
tc6KS0KGuIJpDHtM4C+toZT+E5XancZEL2wEdzQyLbrsfX5NMVWCeyvyZGn5OjN1Y2VJwmzgwTpW
wP+cX38aZgOIClrvFWfc5l8yxpWdyIoIMw1qUU4VYUJMIAcZ81+5CoignCIS4X+v00y6pMFMABUd
gmWuLynUcRfjbYP5L6incepNIkwvC55VMqs8IAEHMfS2+mmMABqAYCUbf1GpK2iX8nXuHYTE8qv/
9OIzugdE9vay1n67Bet77V2wmrvn6YovSjZFO7TA1z0wI/t2WiK1LSykgwNWGFDXZIQbbT9IxwQE
HsyejIZLu9Irw7sAoku5upSBloGpteX/5Rmfqu+w7sbSmYRvS8M3oEcbFv9z/n6Mey8JS8EDWDtx
JOl1KmS27dzx81oIeHFhyMsplt9iF0CHcWQrU1gGJf/cJ97r7txlf0YmTxjTpRjxvlypJCkyiTzJ
pCTO17qi/hPyHIk/ZW5ZG0LL0xcrRzq95PVfQbFk5tG5feM2+DUWc/IozdSs+eSUSTMiLGooHfjl
+qGMKPZHTSCi0d3GcUksUL4L3XpDGiKqlMpbF4IY+Zhu5W3WREQn/Sa5d+EHrV7YjUjR/MBBuRBv
ili4VYxU2Ce4kfP+8zFOj9D0ayU31zRDHpLOTInS6k4fvKwuYu96CrBsYOL6ElfuY9+m06hRRsFb
L5eNlRjsmqmi2okEXh5BZtvlS+r4oYgeUtgt7LZOOr4UaQSIROABhpdc5AVWmvC4LugYLqc1nnXm
dJG7+IT6odPiv/2IakH965cYOSScJ4cxhSJyNv052VHeqj0Pc+xBSRUz2JsET0v73eBF6OOVzodz
o+4DxZGYqJLLuYP9cR5YqpiGfTTUc1itFl7xvBW5B4DiOlW15rVd/NsXOlwwCQppLFqq2L5u0TvN
m72SghuGivNqspMQNYbgwyB0zFLdecJv6+JvhUspExPh5UV7ANVMlNa+l3TOSQObpvD11Z+JHlYP
Mj5YpRWytIEJyzyxRSdzkW596TwN7tvEecOXYI/L5f39lXn51KJ2SOo1IZlF+jmN8/S3STtW/CeR
+49PmHg1SQigExui1SREgwz+ToodXM0ov+cMsv1//7DckRp6/eWIGbTPsPC/bhItxPeNMDhdsh32
5JgxHnT4PATtsx7vDAU2gksiNgQfs5NFt5YVAyOn1ARZEXLC0N6ADyNTvZqQpOVcNk0/NTdHJMiC
PuV1oGbsEXSyC3X56PDZ+tF0ML0/WTLLIiFLfzWnnsnsA/0GwM/DpkMK8gDrk/6bpgjRthHzQYDY
EHByMoErwYlxt9mFwbsBJSJAQuN3Q5SdO3CLAgbd0R0uzvBVZXv0cLC5jcDrd/e5B0wA74E0k/jJ
SzX3+9T3r2A2YJNDjm3plpvAfWsRwVjkz/IZRgWfX8rbOi4Agct7DrL2PwDkNZAnKEVHjzFanY5O
RkN9Yxjr7FObkm3HUFrhpY8tLk8YmYYjzaci6CgvdswQ0mAjwxTdtuNwGZowvVK6Snv2brqtO39M
ldgnMJWmACqLkgKXXWgusJ+Iz1mBW7oLtDjLI4y5Hyccr1nWPPZCcBdvTJGHB43FTW7pFZN3JcKN
i8GrUP0mHVP57c3xm/5a7vPh/dzLpAmjk53zmr6AFZXROcIyNNrHy03NQC9lBfWUYigbMH1wl+74
DfK/TuoEn5r9n2wnWY6FpFk84eUzdBKSmXQRqISQCffyoktYNrstVdyJnUtFFWhfEr+9prnpMow4
5uMxYl034n2+awgbz7qULBeaWfZIgrcHN6orxEO0b89cdl433BITjyLOi6+aQ4hmVLWbAWvXlKZF
VdsCopmonsUxriF0WN3lso7J92+BYX4wbw71ptLwILKiq15rorQ3GcNo0TVrrO2Y5G7juFqdYALW
Mo2KyxOPKTimYVxt74Lznxb5mwTt4JLBXsRqW6o5R93V25HO011mIIgjrRnOqFD/L2M1QkadMojf
Zq/Mofwym4vZTRI1aewfAMullvc6nOLdbvQ9lwVnaAG0IbNCiagNcIzx3Dfvh83UASTHr+EwXGDV
vZ5bO13XeAcX/MgF0BHjSiLuuRSHpoZIwtKU0e2Cyfid1ca/jVsTeB3Yke/jvy0s7O/74FDTOJ1n
GbQirJKNbMgdvK8xA47AaanVrD4TVJvjqWoxj07GrhBSXU8JOeonsi/OdTbLTp3SqShRuDVLvnHk
gsNFMxkawiY0PllQl2rmU1aKithtgmJPC//EkjuocnDq4YysfannWaGhQ5kLIj77fBnTsxqFjKa5
VjAWX8UoOHxlhYavcxDNWvJXYs+9Y5PQUFIT3RUEoJLUCpvxWoYxeSZEBvw2Cyn7UvT89cDC/IYR
7i96TK5rP28kv5J4kLncoluMbJxAFes8ZK3/qz2rysuj5AUSfXKlMlzkjdEPy+d4XJSs7qZJG+2g
4Wpu/vvKuHHykBXCBrtNLEnO264SjVfSjsqhzrECRmHRPVzwWjksk6ikuipF9EkHYEYyUyOBSS0p
hbgj+nyl5sj8YEIVj67vpP4xmJKvxjwjuHtHiraEVf2jvPGsO2nI84Sl/NseYL6tP9dxNs3WTmiJ
GywKMOIxc04NVbWzoY7jS3FEbO5vGjI9+fyWdQmwwOyfx7KDTdFlOayaCjMwHndCUPHUQIEyLjy1
zwQBHCbLsuWx36+uHBGkKr+xi+eUMJ7MetVPZ9P70tqTW8P2Ta/sMYoHiE45MHVLqAU+BZDN4rq4
aeIae5wlDaGorkvZphzeAGatej5qeIsrAuyGp09lc0xCSj5dmXIo+6qLVr2TFgxsVuwcpJTg6jA7
T9pLShcuGzNrvIGEsnnlJe5ZOxSv2dgC6Pyrf1U5Bo9gRKXvFbV+pRhZF0MRoqWTge5eDQI1Y7Rn
9AX4FET5qeCbMbRH11QYFMqWNfVQ3nri2aSl427Q8nFB0ou55vBdWAzT69D/DDbbskwlhhEYFKAo
sAUpQrXmmmw3SHKkHKkBN2V4X6TrEbC4QMoWROBGoJLCrRtlVw+Kg1mCeXRVWSVGmNRXWV0zuMIm
TMF8LbWrcPXZQkTbM6uopLIcPg+HSkO/6Z/Bo7bV1peeSHtZ5A2KSpidWSeYoPjUnZoDW4quu3L9
+erDmIoL2tPDsjB5+2/WzeUl3U/RTlLlZtyZAfRbyhf8tFNhpqhzqt/9L6B4l1o3WS2my7nEgbAe
wQhAoKKS6Scm8TLZ/YFrPRJSHLjqJqAmh89bF8OrDjcVTYhPQMWiQ42SyJvEInspiVC7UiXzlwch
iqm6YGihz7fdg1Gnh+ijld4XHTfk5kzo/Vfaawpykm4vopqrAE+VQnF4yr4dF+sfHp32aYNfR1Ak
sKrijauw337KJzQTZ1rjew1VVz64UIp1ngQYJpqqt21rQvjQLpg7ekilJ0UuDLGMdgm3wmQ3vxv3
NmnCVNeKGefitBAvYKn33lp65WFqd01TGq485ZlntfPqkfaIVQCiHWOPrRUGSHW6oJeUM59Z/+vG
FmT9r7Q7VWL116dIDwl7sS1RtK7Gcq9fr7ZKhtbCPVcBA1O9ALWoH5R2E+kw7RxpVB0e92m6T23A
3IhB8e0wWY2qMTtxgBom2/wZ4B3Rx4GWJfiS2HHnVWOpoe/87zWNHvgDNugnNrgzdgASlntJNTtS
ooz4B3Xp3kJFOOswgTWbaYUki1eJ3FfdaWzBwSeleYXLqYEEBusQlxzvXjyPMkih1m2nRhwbjMwk
Ecn97LbEX1lj2/Aqq5RlvjSNWg9TCDxRQdiYVkJutbckiOgS5u/DEZHm/bEFTdHZHZNUxJq6DoCy
quz31s5h4+pnk1ZYrxHH5KkfwFEV+lGJP5eG+mGYN3bFgWIHw9II9C+2NWkwUuw8TzN2tv3693o8
QYntNU21hmYPZdcXw/ToEosOMxdhPXu11jp5CXuBkNaQBgM3ktd8OSv2LLOv6gjT1SBPx/nR90up
C7aJ14T5bp6gKU2fR5jCOrEj/GAJ2IJ+2lkX6DvxXCbYSllA4icIYxAGEJo5nj5XJ2uM/Fpa9aYT
VyaoqPR7pj9EFqMIvaFcLaTeTiLrdXY0BMK8wECIofLq67z9z0X592CgP/VKR//hPUfY+fEjlb8b
fBgr4jz2fhSOE6iuk2iszh7OZRtOe/KvqPy5UUCV9HGMHavMuZFc/IZKSoYVNV5g1/U1mXxGH0m4
ZnlMlYUYH7jTFbql5tZi8nMgqCrBdCf7jpwXYkFWZe0xS+z3dyhMJyCdqOJKCR5FQuWkaGyevn7D
yV9W1ibAJEc2HPdMIkELVOTNbY50jvTStfSALWpyh9GELXD+/oAgH9yNf7Jtaw4M6r8lnNpMYBZI
IV4/cr/I/CWRsHBhXfMqVMVb0pVK5QIqc50mW7yo6xERJJLMa6Rfmlquy9kuiKDgPeP84s/slWbw
k41TwqYjV21Y9NQcoozRz/f/2MdicA9vTOfLWQumIVt0IP3f4Hr+1JvkRyNBdsO8hm9tiVYUPIoa
1qIye3xwKLfIvQeT3buxMiiYvMvY4iJ4lfM1/J1UgW34AVvKQW5fLUSrMsYVn/SeTzvjrtmg74pG
52beZZYnQWbeW5JNUXP1hWsR2rq7/A7RjcZ1FaTE0SuoQeeVHs2cMSCzkzCz1J5fZILP3ZMym3zY
4ajWZJS5WwUNT06nJpHxulggcHBie6EG/RpmmU+j7rNW1cuJKcWyUJUXo70myZgugKTHGGlXOOfs
OXQeU3Z/9JzEb9ufmk8C0Cin2bjnw9g1liHHNNLJYOPMfaFOk+dx3vrVPDe4cZgJ+91qFFeMK74D
pB52jGnXHgcIszJtvjRvvW2UhRQd3DX3H84zmCadCaMKEjW/92ghi1uhR+i5FeEyYfystKTENfNO
Bnf2JbC4u5HLgvvqMKpxVwrzlqILMu6iqHNIqI5XNNsVkWg/OEZkSlwJkcXsJ8boUrZyipZncAbX
8p4EcyULtAsr+JXfmbTqtdIQU5Yof2oOdqEFP+qz0999TFGv4A9yZhPCd8vxf3DJriCxOljI2yrv
062MkGoFo/fsgRXKS2uY0LKokHseRT6JXbaWmL6xVH40/kRdzxaByG2V01AdinfwCmWQo2lVXkBg
B4fu9AJl/DaP7gXbUWignMqxoO6oWlr/PUozh33mNt5L8GrQ8OB5otpgaqw8blzh9qWaA0rq6poV
Ut2HexNAL1i3q580REEPlMc79GfrhElwU/Ldhu7g7m6jXa73KTqG2qLawUNWI82mefARR6Q/NySd
3JhhJ+vA2cA+38C7D5g8EyRQnyjPiJ/5vJOW4HE1ZUkB74j2nVOxkWxyR+520yzEhJ2Ajavse/bv
lcdrDq5VGlRAXQbgz0H2FRSxMc9WrL1WuJpDDXQI98Et3b3azqwIMAAQukvFFKsnmdq0wtbktyl8
jpjNTs1hIU3bjLYCpzDo04cV9CGeDbw4hsv7n8dhQQGIXJlYqCCMAlt7CKYVH8bEgMS3IUj9xQJG
VSvlfQIwJfgivamz65T+nUCAqpxicJZvvRJEucpw93tvdKDLs4VLwr3oi0U1BkyqjSxtoIyFhJ7G
tknBOafjFWIKAvMZcvdCrvfjRvisCqqbNQ2QlyLdunKKfoL36ZY1TRWz7GAbc1nEy/w2RBLrfb36
HSinLsPLKB2bFbbfcls77H89hkq/asyvXwbwY2sx+tqXhKPpV9JOkUt8GEgeyhyz8UqO7AlUA1pJ
FcRkJxJYdtYHdcJZ8r7LtNYFRrXfl5IYfW70y31+vbbzypaFfnLkzW7IR1KjC9aVpLkXC0s3l59K
rOjiL4FU61Kxv+t6pYBn8gT8oJvKi8EvXWDyIQqUyyn+5pulZpUOwXjNbuXAr4X0kpkFkflR/7mo
NnuafMZrq2aHThu20qc0e2+RUpWiBzPzF9+8VUhhaPJroc2hBB3uf+6XrRjJq9i/5Nd+IH4WNbIc
su4irgo+0TpA7X1cDWrh70OcNLHk5sFGFKBvTsIwrgGaMWQhXRN/GuocFIvjvt0dn4Ce/OSbyuLx
ao7zMor88Oh1JedvUfjy92pCQasJA8DoxvrUOpn1H0bgE46e/ErKTbBaXn/UnOr+4Bv+mVdMUxqm
ue2FAd5YPpSLVTO/GggRk3MBI1nwBFt1H0n5j9IOVCQDSH21ByjobWSkkspb9RblURCCdg23gHEs
zalQncc8K+0CRn3QOibkpPyD7FotmExA0QrF9M/GDXME7dZifaOljtuJlTJ5pziMKcU3JkCPQG8b
hvyEFk9dTmllAtX/6o1cPF01Go9xZy+mavJZlRQ+3Ly9r93HuY8aDeTtbZdmlbaySLC1gsTweZ5Q
olQ0l4AfDM38YATHEtfTWrzS+FwcRpCsPWMdUWW8vWtAzUk/9dtGr0ktvfp62GuRf6WGYQj9/5Gl
AZHiJvTdgkRXTxQf+7gjxwyJLsux/1K8aQQLbbD+uQUgcwZg7zHxqlnb/T+Jw6eAe6nOMMUSwzCv
nsMgiZy5UbgWnMVI41P5Ec/i4zhF6bGpNTXkQYw2pbomDW56ApDR+uZyi2ZD5AbRmHXPlyO5m7dk
PZCK5t7qRm438m0SyWYKYJlyD+P3R38oFeBxgcRQqPi0KGx4OdIohF7hvshl8iHNx71pS5FFdrwK
BvKjyWWjbYH9kHj/ocL70CbnW3SX4qLxOQ1aKIxbiU1tWoyI5pRfc/bDqaTd9GcNP/m0cHzfzKIo
FWRBVXf3sFwzzYBp8qUcpupphw2DImVRbuGB3xCnD+fopOrWU0QFmI5It8zGdnvk2Hw47726GDld
zvH9MCCFluL1YqSFxEIaRtOApbsZFw3R0iTySjahQNMbiTutf4bcyM7K0C5GUSyt6kKrN4YYayBf
t4TxBvm68AyWaD5Bf/A5s9jmZ0txhOX2pwwxurpYj3LbQHtWFodNnjIKu/Tg7JPIoGDE/v78IRs6
IC+Cus4qhDjAmahjkJuOTvUUkGUoC1d8gsbObJdcVSbyG1ftoqIQA2i2xfYkE88zNXJCpyqwPu6L
2oyZ+RFT9lrJVEQDmEW3L5FCZXmJ6JO+oPUhvHdmGZxSCGYSDS96RzgPhaedwN/29NdhfaAdJuUk
4CE/yMSCvQdNk3Ya2HIvMQSghIWLsB7KA1qBAZ1Np75ZCZK5TInCuMkdsV2enlKc3V5ZpVz8DBVY
d8WdhG+9HOgSbtkrvNGd4c7f5ObEnI9qePHQbL3iHSSLhb+4yV0+F5TNKRbX9ZP6LfxayHpOWwBQ
+5vaGouKe73b70Ps8Li930AjVp7uJYoXm8JguR+STdEs7DzCGa2jNCnr+xrf/uMr10/Dj/xrXrMq
NzUjvX0adZfL/KTEQC+BHP+Wft1tG+jTl4MStGCSfRvBxQwszIhaK5GblO62DCk/PdtfDRnuqn1/
wgZge4NBqFWjaJM7JNzAXy+c/lbAcK4c1lQRIJX0d6G7am1ltT5Csr5+A3wvbFFnJLM9AqT2YrYH
NLakYv+GJ600qu1hcQzXBim9Bedw4Nwtsc7hxyotNLnXOkCgwyCh+LRyqTbMi+rgaRYffcXPKj/y
cVV2YPSQy6pH9Udl8exklf/FCUo0wmbGssI5sl0c1NWoGHjO3+G/ic6jvtSuD67HMNigOo8K3l0w
jMS8Bw6Ix1PTuK/fDx+n9Gf1hAfKjpRcDbcteERGalSP/CalVj/uheVbKrpXbOsZl/J34XH//Ycb
VOu3Y9305GmPjO3nbTSMfcvnCa4cPxARk/fRNdLhC2LpTzFOp3NWcujo5PcphSl6V9L9NN2ydpBI
dtCGQ2XHN+JOnDPeXKoGOPBavyU/OSrizHXVf0EuQDohgyFVetAsHSSpydIOpyZb33rgMyjzxQLY
Vk66LFAXI3roE6ZQMmRZu2+7d/eE1hFe9BbCa6bnYT6N64zbicMHFwGPuxqM4Nv8fR80upJGlONG
e8L9EomgwiFvi3ucNXWV1lIq6g3fBect/daY8620R6SbsJAb9rlNaMbSr6mBCWjknaeam/0C4xRR
XlxcflGkqu8lwJ1gqDJpCzJq3hSppgtUInNQT6N4RveEtSfQGLg5yxVHtotWb9p05JiNCXuaAgKL
Hm04m6yEEsI8f6UvoOYlaCP+Pt+s/Sjb2/9dI/lRaVBuX6aIcJfMqaGrpSi3eRtDwM9XLiHEtWng
zhmEENzIpEHHAHxu0He7HnXgvvoNSAHqXt+Dfz4nkeFpxnQbAf53vhf3sckRQe17qRY34WzmvtBD
u/1RLNboxz8jIkQEZZpXDEVJt0J8NiA17h2I5phtACxVaiRSUBn61mgwIlkD4kNYrKmzlgzExHki
DbN7fLMabDx+zqhjrb5W+BzjKrTrjf113f6YmlpJVVnDf5w2TIaJtVlLabRawf6cP51l3M8BALZW
jLwOwJsSNwbAl4YjMeuUTvKSNYyRfIls0mKPhBsREMsLsy/6IFsNAGxEQGtW3KpLWs72ql+UlCRd
5QDT3SCPSgEp6NALg+T5BAH2NcdVU/nTSJ72uOp2IcuO4jim14olgZjGBerUpNjYiSZSECj8xk9e
vSMCJkVqvVT/grEtW19E4I1kQPXx0aO55ITsp6ye0Epqaw14/mxlME0JVIFRR6Jxz252AEdeGGHn
yoSpdxuR69oXzntKn9XkS9JZhy0OkhqSzxqHBWvBAeuZ4z2Dw8RXQhSquiv0GE0Wq2VqOSgXEdRK
AqHLINaz0TfEYgwUd1EPbJN+LH0UlgjU5Wujj0rfmW3HsHL6g7PyjDlPCNU9tP+J1A3Qlts4tguW
krQvWSdVKYnweTsipjAU2Z7gyf1pdKBOhPFJwCrz8PKlRrq2Vje0NWgcjjghg5h0Fpt/ouRx1Yht
K4Bo3L+odZqHZMkJzeVzM2/s+WjvRklt8keAfHn9gRf1L0kwFuQj+dTenQ9ji8EgCtjNENB9P6f6
zpJc7GVh0wAKWEDYyNDUz+HEBJXbC6KPf1Ent6F0kDuE1dDo1dk12TFG9Ay6nRwpakTwJI/sKFiT
Dlzn/mNeVE4VfB49vb8PZ/uCqj4qxbETebbeg/xjizpkTRwsxEOSBLF7R7GnH8pc9Deg3/az3wrr
vUOjiuxFtbMm/ELur5IY2BNd3Jp5t6EjiLXBJOlwaFVK1lKP2BGbs45xWSlo2jr3JtoiIhRO8HBe
GPM7mbyOwu0IFMNkzMP/GLtKrSreOmmRQ05UwgMQDl1tSP7l9Tnu13QAUQdTCRQqwO3nuudJUVlO
h8NhzV6ewwrZpRgb3FfNz08zBLVOzn2twpcyFn1LqIsKNISRCB6xR+gy5F5veyEdvQ0e3BcqIPmv
vmRDNOiIaswN47B9Pspbk8BA470yR9Pp2x1b+d3gG7uqOc7qHqIs784uS3FpA3TFGZjXSvTBno/U
Jk9LeHNfV3YtOo11XL5RiEhCnN9dBkjRkqF98Jttk7UVpcA0oAJ+6DA7ghC4ylvh+M4QxRVGI+Ma
1jg9BRtA50yuwUnCaJ7ImsaaKOmaZTabd8FRyu1WxAjUjDo+sTjdPa9yrbFcQvy/w9LKB+s70kIc
opySkUsWEfPOwWAjM9OyNBEzmsnLpBLyo5mgpn0s2L+IfCMwK6IkkTdcrRp4Q0Rbj8usBuLvp6IL
1hEPFunNdcI1Ps3nVQ3K6UB7eV+T8uOFfeCLel/vi/Ckucg2EPaDUoUVGKWHMTivA33jbmsR9cC9
3V8DMLjCrthfKxdr24K9iRfvVCAuU3eruXDZOl3pQ0r6DxbPJeb5BOxAL/wTsTB5bSXIY8m4LmyG
ih26jYD5gvBUBgSooBNzxGV52xLidxetdrEORHuU7wrnTsCFPSlaWn8tYOmpGLJsLG58qbtn+TIf
uQW9wYz93EnxSYnaxUSEGuLd7bnFfUQ1HD7VygO/4oSP2TOjd9z9TVTDmnQ8fjl6db6Mo3Lsscx8
HQ3g6hOPdQcN+NrgVXjkBxZvPYxcYZFP0lg9jxy6+eHnl4ipuwReGwcObOh26VpL86UataSrTeb5
qDjgwLammYbAK1Zq4qdLYLYB5ejXVrj3m7EWKS2oCi2nhQeawbZqKjsKtk8CFU+5IY1uh0LS1qmX
Px/goEhlc7YD7MblixgCbSXi5jAQJwWawMU1bOJD4sti9Ezq+mn8UMhvi07zIehbzTMbkVg5a9TK
GhCrjOOlqDbnIk9A1pYOgVUqd1PSLVxGG9sNpZ+xaWPvibxeUau4qc2i5TOP8Rve07g46NoZABZ0
giSDzLKHAbR/rp9bPYeh7JkYPEPM6i37nIQuP2xP3Df9GLQiSxxGNuPWjtkf9yPYZDJkGuPGErPv
ORYIHLvZnWJkj+5laINun6ElUj0pscVI7XK49j89ZvySGcxyXz4TfWLKV1OtGB8t8KDEJLGz6XQc
D/+2Pw+mQKEKxK1J6TDryOf/qCyL/nznE31LHop8/ML+ptArW3oijQTa+pLiKRDdrSV11d9ZdXws
BSdxllGctgNRoRryLGrA8ydydPiptpAOY7/P9ML5fzzZu8ufenQLqR6BO8hT/3UXYYV4AmfaZ4w2
MLdiUFFQn15csFOTaO9PzKhBTu0VYtYIhmuTEkQ//CWNWmP3Bs1LVAHx3BIjpMJOJ9hjnICTFSV6
pdW+mJKKK7KxAe8oRbI1svv9ESAS+E4D/+2efOWKcEhWhdjf09ubuBdwqsP1tpppXVxqwMVu96Rf
aSbsfDhRRGvw0muImESKdBBD8BORfqGYqRezpaBGhaBLGSqA7IxFzfvIkiRC23YZB4gRf5PLtqrp
ocgji/w/QDyRSioCkIHq610s+52JXbU9FcfKlfBacwxVIK+7pW5o/B41/lpnN7LmP4RDmjzQfAlf
JOvAQsIUZb6pXjl4pA6Rqbr9EhZU4tIZwO+/k22A+W9m7zhkPs09G2TOT7j6ejIN+4rYBW0t6STA
LwnYVbtlBNJc6Sj12Sk/MR50SOWTPqGZOdklKqzZidSia79luyhp8JxA2OS2WkqLPthLBpvaBzGW
t8LI5k/xptLEfwxbtF5+a54A1iNCH8fj4H2RSOx3CC/o15oSxegeBarzlhb/cQ7VGkRI10DmTnNR
6aPLhSLrd3eQPH9XPidMEDcfJJSu+4DfRJOrvOw4IJVmBrItIatSWSXl5x4osRKszV0hBbpmR6C7
osZHPaj32nHj+hMs3irhWgTiiOotNp8eLQUnfINMgNcwrPlUH+/CN9h8++PdlGcKNKomKH+VExd/
A5iKXq9pk+Q4w2T4JfC8rF3r5ht0QcsMVWU4k2pKtuZjRua6FHb1R2Vuj7StkRRAx+ni67jOQtyk
G+4tG6QJTKTfkWRYa7uCAk0t7bKCSGI2yvFdyXgp7iarWe9aKixwjSeH+nRSrrvmYiLrGQgXuDSq
1HuOO0Y12LdQa8k5/ZSjaSUGtIaYsX9vPPgadM3jP9ybcLyUBT/9kYAcNpFBD9fhHz3b8XRC+Ned
5kXXkiAJpka5m98uqB+3eW4D22eJC3rdNJMRHV9FNdCxrwwzx1gzqGFv+1/F3GAq1Pt/1mODxNVb
cuJFnOfqaweXC4Y7whBj3CDfWJI4tBC+I1jv1nxjmWlBD0EmqWPp7b+9RaKYYCftaoq9wh8Db1Fm
DRtfvm3gJyPEg2ow+vo+bbt9Ss1pWay/wcm4gojcDfBbWFSLGHlEpHjjtflSB4b2/gtHDbV5Zi+r
RvrJKicermvkaGr3+5DzMm5JzlZB8xRifKOffplY6m0QcW0jX24v1XcMFun+psUu/wxjhG9lAWeu
mOm7gjhZ8tBV8re4cqQvCS09tgCMaqT4V/uh6RRyD96Ca/8Vr5NlV/S7V3frXVVTI3wYhAYMXdAZ
mkxJG0qdt0gKIuU+VeFXmT8GOUQXJI8j/lIVcygA3djmftxljppCQkmr+BNTiUyJpNvYwxV4t9/9
J+7c6nZ6fhT3qcvdDPo2ySIYhTesqxGS1XWWF+0gKNyRook9HFM9rD2bmdYW1WxHVg2d3HJVbitK
rem89tRc6EfNU/lsPxSEEfoNpdz5/wHfeaPXAxx83jqdJlKhmEpGcOEVr0+dHMYavFIriTOrBdeb
B01dWqOiKA1KNb6mCq32lhCyihIQ78hVjzVt5i1945UKNXsdFfH1zZzMKfsExQK+1AP4r2yAVHfn
eAnHqaqRrQOzhKOhzfBxlWy9Pw78zPHLcm1eN0JTYFhOZkgQQfoaUhrdgTQkGdwBE+MXunf2/JzQ
me25CUHAquHdJzcuxfquiiCbmRElym9dsQlhZqLyNz5cPi3OBUB9U9vr7yF6eXAAARnrxs7s6d4u
u/Zv52Xz5g5bJFrJkskAabK1qE8Sxp8E8fTLoBYt8qGdRqXTS7SqT5KoGq8RnC2hqlMoyDBUe/m0
xDFB1k8FTefxvB5Ixw1gk+vqqW3lXX+bvsG+mzx4BlUQPQI3VCT+F53BFoJ9Ko4Zy90KuLgfMCtK
mMurRlUIq/mSf7eEEA0FBJPEbC/Jo8IwX8kuBCnqkJY=
`pragma protect end_protected
