// =============================================================================
// Copyright 2016 Amazon.com, Inc. or its affiliates.
// All Rights Reserved Worldwide.
// Amazon Confidential information
// Restricted NDA Material
// =============================================================================

module top #(
                     parameter NUM_DDR = 4,
                     parameter NUM_HMC = 4,
                     parameter NUM_PCIE = 1,
                     parameter NUM_GTY = 4,
                     parameter NUM_I2C = 2,
                     parameter NUM_POWER = 4
                  )

   (

   //-------------------------------   
   // Free running 125MHz clock   
   //-------------------------------   
   input               CLK_125MHZ_P,
   input               CLK_125MHZ_N,

`ifdef SYS_MGT
   inout               SYSMON_SCL,
   inout               SYSMON_SDA,
`endif

    
   //------------------------
   // PCI Express
   //------------------------
`ifndef VU190
   output [15 : 0]     P3E_TXC_P,
   output [15 : 0]     P3E_TXC_N,
   input [15 : 0]      P3E_RXC_P,
   input [15 : 0]      P3E_RXC_N,
`else
   output [7 : 0]      P3E_TXC_P,
   output [7 : 0]      P3E_TXC_N,
   input [7 : 0]       P3E_RXC_P,
   input [7 : 0]       P3E_RXC_N,
`endif // !`ifdef VU190
    
   input               CLK_100M_PCIE0_DP,
   input               CLK_100M_PCIE0_DN,
    //input              CLK_100M_PCIE1_DP,
    //input              CLK_100M_PCIE1_DN,
   input               RST_FPGA_LS_N
                       
`ifndef NO_CL_DDR
    ,
   //----------------------
   // DDR
   //----------------------
// ------------------- DDR4 x72 RDIMM 2100 Interface A ----------------------------------
   input               CLK_300M_DIMM0_DP,
   input               CLK_300M_DIMM0_DN,
   output              M_A_ACT_N,
   output [16:0]       M_A_MA,
   output [1:0]        M_A_BA,
   output [1:0]        M_A_BG,
   output [0:0]        M_A_CKE,
   output [0:0]        M_A_ODT,
   output [0:0]        M_A_CS_N,
   output [0:0]        M_A_CLK_DN,
   output [0:0]        M_A_CLK_DP,
   output              RST_DIMM_A_N,
   output              M_A_PAR,
   inout [63:0]        M_A_DQ,
   inout [7:0]         M_A_ECC,
   inout [17:0]        M_A_DQS_DP,
   inout [17:0]        M_A_DQS_DN,

// ------------------- DDR4 x72 RDIMM 2100 Interface B ----------------------------------
   input               CLK_300M_DIMM1_DP,
   input               CLK_300M_DIMM1_DN,
   output              M_B_ACT_N,
   output [16:0]       M_B_MA,
   output [1:0]        M_B_BA,
   output [1:0]        M_B_BG,
   output [0:0]        M_B_CKE,
   output [0:0]        M_B_ODT,
   output [0:0]        M_B_CS_N,
   output [0:0]        M_B_CLK_DN,
   output [0:0]        M_B_CLK_DP,
   output              RST_DIMM_B_N,
   output              M_B_PAR,
   inout [63:0]        M_B_DQ,
   inout [7:0]         M_B_ECC,
   inout [17:0]        M_B_DQS_DP,
   inout [17:0]        M_B_DQS_DN
`endif

   ,
// ------------------- DDR4 x72 RDIMM 2100 Interface C ----------------------------------
   input               CLK_300M_DIMM2_DP,
   input               CLK_300M_DIMM2_DN,
   output              M_C_ACT_N,
   output [16:0]       M_C_MA,
   output [1:0]        M_C_BA,
   output [1:0]        M_C_BG,
   output [0:0]        M_C_CKE,
   output [0:0]        M_C_ODT,
   output [0:0]        M_C_CS_N,
   output [0:0]        M_C_CLK_DN,
   output [0:0]        M_C_CLK_DP,
   output              RST_DIMM_C_N,
   output              M_C_PAR,
   inout [63:0]        M_C_DQ,
   inout [7:0]         M_C_ECC,
   inout [17:0]        M_C_DQS_DP,
   inout [17:0]        M_C_DQS_DN

`ifndef NO_CL_DDR

   ,
// ------------------- DDR4 x72 RDIMM 2100 Interface D ----------------------------------
   input               CLK_300M_DIMM3_DP,
   input               CLK_300M_DIMM3_DN,
   output              M_D_ACT_N,
   output [16:0]       M_D_MA,
   output [1:0]        M_D_BA,
   output [1:0]        M_D_BG,
   output [0:0]        M_D_CKE,
   output [0:0]        M_D_ODT,
   output [0:0]        M_D_CS_N,
   output [0:0]        M_D_CLK_DN,
   output [0:0]        M_D_CLK_DP,
   output              RST_DIMM_D_N,
   output              M_D_PAR,
   inout [63:0]        M_D_DQ,
   inout [7:0]         M_D_ECC,
   inout [17:0]        M_D_DQS_DP,
   inout [17:0]        M_D_DQS_DN

  `ifndef VU190
   ,
   output   sh_RST_DIMM_A_N,
   output   sh_RST_DIMM_B_N,
   output   sh_RST_DIMM_D_N
  `endif
    
`endif //  `ifndef NO_CL_DDR
    
                       
    //-------------------------------   
    // HMC
    //-------------------------------   
    
`ifdef HMC_PRESENT
   ,
   input               dev01_refclk_p ,
   input               dev01_refclk_n ,
   input               dev23_refclk_p ,
   input               dev23_refclk_n ,
                               
   /* HMC0 interface */ 
   output wire         hmc0_dev_p_rst_n ,
   input wire          hmc0_rxps ,
   output wire         hmc0_txps ,
   output wire [7 : 0] hmc0_txp ,
   output wire [7 : 0] hmc0_txn ,
   input wire [7 : 0]  hmc0_rxp ,
   input wire [7 : 0]  hmc0_rxn ,

   /* HMC1 interface */ 
   output wire         hmc1_dev_p_rst_n ,
   input wire          hmc1_rxps ,
   output wire         hmc1_txps ,
   output wire [7 : 0] hmc1_txp ,
   output wire [7 : 0] hmc1_txn ,
   input wire [7 : 0]  hmc1_rxp ,
   input wire [7 : 0]  hmc1_rxn ,

   /* HMC2 interface */ 
   output wire         hmc2_dev_p_rst_n ,
   input wire          hmc2_rxps ,
   output wire         hmc2_txps ,
   output wire [7 : 0] hmc2_txp ,
   output wire [7 : 0] hmc2_txn ,
   input wire [7 : 0]  hmc2_rxp ,
   input wire [7 : 0]  hmc2_rxn ,

   /* HMC3 interface */ 
   output wire         hmc3_dev_p_rst_n ,
   input wire          hmc3_rxps ,
   output wire         hmc3_txps ,
   output wire [7 : 0] hmc3_txp ,
   output wire [7 : 0] hmc3_txn ,
   input wire [7 : 0]  hmc3_rxp ,
   input wire [7 : 0]  hmc3_rxn
                       
`endif //  `ifdef HMC_PRESENT
                       
//-------------------------------
// GTY
//-------------------------------

`ifdef AURORA
   ,
// ------------------- QSP28  Interface F -----------------------------------------
   input               CLK_QSFP28_P3_P,
   input               CLK_QSFP28_P3_N,
   input [3:0]         QSFP28_3_RXP,
   input [3:0]         QSFP28_3_RXN,
   output [3:0]        QSFP28_3_TXP,
   output [3:0]        QSFP28_3_TXN,
// ------------------- QSP28  Interface G -----------------------------------------
   input               CLK_QSFP28_P2_P,
   input               CLK_QSFP28_P2_N,
   input [3:0]         QSFP28_2_RXP,
   input [3:0]         QSFP28_2_RXN,
   output [3:0]        QSFP28_2_TXP,
   output [3:0]        QSFP28_2_TXN,
// ------------------- QSP28  Interface H -----------------------------------------
   input               CLK_QSFP28_P1_P,
   input               CLK_QSFP28_P1_N,
   input [3:0]         QSFP28_1_RXP,
   input [3:0]         QSFP28_1_RXN,
   output [3:0]        QSFP28_1_TXP,
   output [3:0]        QSFP28_1_TXN,
// ------------------- QSP28  Interface I -----------------------------------------
   input               CLK_QSFP28_P0_P,
   input               CLK_QSFP28_P0_N,
   input [3:0]         QSFP28_0_RXP,
   input [3:0]         QSFP28_0_RXN,
   output [3:0]        QSFP28_0_TXP,
   output [3:0]        QSFP28_0_TXN
                       
`endif //  `ifdef AURORA
                       
`ifdef I2C_SPI
    ,
   inout               I2C_FPGA_QSFP28_R_SCL, //FIXME need to hook up I2C
   inout               I2C_FPGA_QSFP28_R_SDA,
   inout               I2C_FPGA_MEM_R_SCL,
   inout               I2C_FPGA_MEM_R_SDA,
   input               SPI_UCTRL_SCK,
   output              SPI_UCTRL_MISO,
   input               SPI_UCTRL_MOSI,
   input               SPI_UCTRL_CS_N,
   output              FPGA_UCTRL_GPIO0
                       
`endif //  `ifdef I2C_SPI
    

   );


`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
rfn+6xSOaWpgyul8VIbRDVm0zc0GOvDPpzaRHhXKosUzcBaROc57c90iiYvpe96FJa/CTbs7psFK
DwRnsXwh+7C6uY81GOTvtJqEsWIYxqTBnLNEvdPbu1mQzpyYINtq4zwAbsW/FhKT/aMjugWVZNy+
M3zeKeJ4KbFD18oJcNCPT5FbTTS1rzvExU5JGau+hEfq3/pCpxj8/s6XbTqICTB5ljfd13pq5pM4
C5DARm/uQxCGgZhfI3rwE40k7KutyZ769raJ+OcbPq7mgmrGfQTp1x94Zthc69ABoVa8e2HsFvWa
Wjp9hxuX0eKNbQmKyrx5veTp8Q4dvjUorvItrw==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
b3H7oqTKVDjPBqbdGpgpelJfGe1FQ93TP026KYtA/c63lwiDYFnsMcqMtdyoWU7Y+8Moq8n+3JFC
KzR7O+srcL0zGlcxtcA7eSSFfXodI+iioy9x9ZoO2aFcQ4tlgYrYopih/qzk9sFzjphxLd/e1clk
mcIMq3g1HFWzAg2FSE8=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
c9/kHRTRfHf6TPpGg1hp0xq3X7OCH/zlTHfxm/0mrHJBka3KdxguE+NJpF7KVoO8GYHsHZPgsheJ
8FpyD8HvNUxGt/eTWMQ6CP7tagXTfKF3TtvDdD8hWma9f48FyRQqV+0wlF7CRi64vo6Ei+6leqfZ
Delay6m3fRclFNIew00=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 39152)
`pragma protect data_block
XlnkcYP572+jHyrDmZf54QeI8IyohDtf2Ch2bFRfjPMdzrtt5tm4pMfRTyT4Py7wDaKmIgCbvmTy
p7abJgNxVkKd6LQwpZiYGor5YVmbbc5V+yU5fZYl1BgELJoHFFgrEIZ77NCEJPc3hXSL0VkA+K/k
gQwEXNwQTuLb04XfZZEjDFzGcDaaq5duW/Oukv1wBCNdqpmiO9qd9BSM2WbJRvt8xFgu/SleW9MX
ktx66ImBHJfAlOr4a4xBADZzzaoqTaa1+0rAkO02WLFen+NafLhH2lmpHpF2FdHGycd9JVQJyg6v
59H62Hq5+4ab6IFNI5rOep4X21OfWnn+9hB14gMvgjIemEkFvDzH2/OpFJknxBdIMV/XXZM22umC
yO46RovoY4m1Gph04JcZv62rnXWiDCcfvy2V/1dlEz1KDfbRH0C6KdUP/cT+rG+Wzv21yuhMovdT
upW/AHL33DcZRKxUJ/+Qu4HDq5IimM9bIq+ZW/nPTAWKL4y1Mop9Sg8rDK7ZYQgHHr9H42uTQY9M
6ZkI9s3370zolJfb8A1xoKlLAvEJyv4QBoaXQ23aLw6EpcZ5pr39V7lyMg3q5BJrqjP7zBN7QmXC
Uwl5IaXEuAAzSTxyh+pp3juBTq7r5IX0AqAQPgl4pQS0gN7MA69csNLzXfeOsKYZW8H5GVSHvvQe
pJrN+4OrRG7l7IHT8dK8OQHEwiBEIv5l/Qi27OABxsF5NhM5kkijrYwuRcs3ZSGYdox2M5dJrZS9
zeC3aaRPqkYCS7CsKNKWklMu+n6vz0NV0WA5hDf/5SJUmGc0D7GxE8Dv1zRCvlYGK23gXt7pD881
PSgBnn9a2o6DROTgrcRQHsGgxZQeh4It2jk4A38b/VTUDOOxT50Y0s+PDtTZXJ1+/nTe1lVcna2C
5S4p5iVnuVOMJLu06YCzEHztJ8s6FFUb6EqfuTHg6Z0YGRlisyeq4ngpPSsoZ9GMgsUbuCW8LZYE
BvW6HnSWxsuk/ecmkT41cn+fbOWpOzkB2BpxFA5wLxzZ9PpNfAPc9Wk3nPbDpwQqsbjfHUlp86Ju
n174/m49TaTsEUpIaNI/03oF2QAvM9sRa2jAAKDwndGNuV+HLlHnd7pb1ol3mRpsAnRGJZ/I6c9r
ENmWc78zmkEgsbNRXPWyy9FykIKrRN4zd26br0NYaAYnLpN4Lo5+yipmT1Jha0L8SywEc6aSipmf
AnnzO/n27BWCGYHXMDgzO20Sy3aePyusUipVp0bopbat3E8KFYh6fAoxgMjnqFN3jIo45mUfUMPv
TGU2UPtmr8l76hIWw4uxYh4mPcTGbHsmENnjCJXd2lMtJfYA7zt/4DCspEXETY11l1Cj8tbamanr
9eYPU9SNy8rTBzx0ms2QExPhi+F5gmKqAPY3BINLnrIbyFQp2/5f1MWEXaIWrXVX9mGp5QgV50rz
MqDMkDZxzTXW5KluAaOJ4Lf6SNUEncS+ea+7Y14FB50vfmjfTFNAXOoLY5HYNKfl6vfDvmb5Ml6r
z2cE4cszWZQ/rF4KyD5VpX21wcadwZBkxbGCKoexAcQuHYttxYEYb+jo49gnf0jif4igiPLp3BR/
HLF/S9Kr3JBlL30s+jzscxfTh0z4BrOdAa+vY7OIChdnv+Spfoy8pE++rL4vzK7BHJXN6vuMLQjX
wHOmoweH9YbGcrhI7JevdU5EdXEgf1BKl5EQCmpDLN2E29w0KhHdfDus3zy+QHQZlj89DAs2nmwI
kwD9lx9rGv/XZA3/WSdtSMru8iSFvjjIsHhA4A7MhCtqn02TI2AwuiKfc2jqsiJax0FKxPU2mVYS
l/UGZxmj8X8dHbtlrGGda6tAScvHJLA3jC2RWBTPNBAM2AKcRgkSlOIUrQmbG93u81vP98h/rcOj
+s9i3xeOyU0J4mY9t/teiamzD9rWjskGsuRcJTT+LW/xhCgVcHSM2I3g0oQGsTHYlv8aTCkigtaW
3Dphd/ia66ltbtArneKcdwum6GT4nKuEUPwm7Y+jzuUD7pRXnHTcOOvtHagr5AH6y2ocl0GSZcZ5
21lXZt+4QBc9e4TANpPx9WSQOcy13K3z3qU8D+rmTVs5PUiKTD3ebA9K/EQPe1z2WgGBEV5yCT5g
tvKO76DtYxstlUC+vItxOPkOiahW9J7FrzoupTAlu9i+akkEbum3AL+mqDx+ezY8DS3QmqORXzrb
AQn23Rn4OMotG/GT6IcQMKLv8EtTzRLTReNmbwjrDM6KNIny9hCf1SkFUx01sigGn3jAgHmM1m+G
qb4fKVZJx56ALJ+jc44JH4UkJffQXd11KSR4Vf4+JqVzZAT+IfJjcixzej4+KDherimeP0vHcy8x
N7f03IM0OFV6OP2GZxMecSOypNeNeZpoJBc2uTpnc75xDr0hhGG8lLVlWb7TW89z2j404QPaUndd
9r+dhI9XsPDx13zNKYf3RL8jDEN8sv62hMIdyhYzW3W10DIkjlHBEg/lR7LVWnbIMQj+2VIf7Tau
qRIRWEZsGyqx+94BkhmF6J1eijaR/sBKMmvolmj8XHH0S4/W137ctldOyCxY2wEd5tle3ExqzsAD
NHO0Dj765mFX3uRO2pmses1HyWlumMrF1RHENxyejkXk2pJM16Ny0vEE6iSM2su3RPjlJ04GOlja
H4PxqNaqfKwJdxuGIaOXKz098E9F5NeQSmp3Nw5c9X+7raLvWr3jnO7iixu/I/NtEsnxxjowuFWC
V+grTJxsPaSBHVR1EyMnjUyTQeYl5CCYrB5q5Buog59wFgWiLNvC28Wn0ba49minnmQT9qVlRxGi
2Ps87+c7JAk5QpArA48yjKhFjhdZeoMQ/pj4RHgjRSUpEa5G/xL1jqtU7d8fmIguHbbsgNjN62EV
g7PIboYb9Ymf3VY+U3ydhisVMSvY+YedR4+avmvIpK+z7TzbpGzpNf3pdkmWRGBZ/8Yv/5r0bJXJ
z7Iirh/avSpF7zWKVGlvdyVMiHXY5VphdL6IcbfEigwRyNoKr6WVYYGS+EqS35F/CL9gE+ebApCt
wP2/AFOO/JTDa/kV/0FSezTovqDTiI5j12gEMAsS0WKY83RJy+ipBCq+C7EOuC9z5hS5F1Pgr6mi
Blu0RNY+pBZ5Ih5Vf7YPknbspYvTJZ1Dm6hjdGFk/6QD7eNNRP0jHCrb0zTam96Az+aEvE8bTToG
6P6oQEkS+yPLdP9/+YP4RKqlUU8i0ec5WdhdiR8mAcNnDZt179DDjs+PWEhV/ZbmA5C9OZJRkFRh
Jk5MNedxwSi+DYa5xic47Fpc9Dqur8puJt54xGjoh77O9J4l7jTYL5s6BOfGFQjlIMqTEjLZAxjA
H41QLoTMsD0XYZYxOW4qK73te0nly+kZdWCZSZpbh+68YNdNxKLwIte9hvKYcsG43W/25RzRdJpE
N0ydbJPLr6wNdJF86o8F2alHgIlNPqmo2fJLyLKoESFDw60RSw6nbp7jpk4mprisCSfVTwIOB+3y
CK++F3ildYdQ6eUT8sxKud6ShsUjX0tv7Tm+0S3P9GekGWL/frnqyj7Ge0rOU0cCV1EP2RrN7Poi
lfUdMNG722+sIIqRWJvMlly9/yhV37ukZBFK6GFb+UVqk43BMLJHRaW8059U+9y4HsL64QE4lho4
kKmCj9FqWqugBCoUFQxXDfmYIEzzLG8+yrBz+pYzUzlnlsbrLYUj7bgQ4zxGmfSUw4JL3qkKMCXN
1WRANaegudm7kaHNY6cyUHkmDEefMExVrdfPny/HNYBTeOQgLtXwJg/TpjuP7Oix1C3U7BC3CnxP
ykxcyrQo2cFxWABypZIWDa+IrWbqyJppDf+yU6WYFJ8GSa4Vr8z8ZSdIg7Szw/fkn8HMfKOw/+NZ
LXk14vmwQb5drpaEoPqdJ3VZoAr3C+TIXKUgAX3QJTLZEKLhyy13y6/LToKt+KXCwp5nM7FORGBa
FJ1k1ogDVPRtr5N3rTRfKbhl9K3pwfSS4xFrgpO6JMNlMQXSozSNXaW80NgnkrHy0i35m1P5fsXo
FOCWQdpt5JqAPi1XwX0SrDEzka2QIE1o/aZROWOR7x5fO/SIXXvIyPRvVDnk6U/Jh7VgRVdHP3hz
JIK2wNPV01R4Egxir1NN+ta9pwUB1Xxi6HI8karnVtwDk44omODVn0r1E0XG4HnnVqdIVyvQASo/
KIMPbjmqey6XT+fgggOQcufFxg9V+GVSEilU5vjZnrq7mkCqb9UuDcalem9HnMzQiIVUa5Q/ilu0
TSNWrB9lL9GBst8JD/9shQrZb0qRRH1yI67GY4du5LcNK09HCbImt3H7ncbKuONiXRyL2LU2MC7f
+ebaFH7b9qbkSbk7pO4AIjPrwepcUJS2K9IqK9FH7AtLQi+5cqJR2B1yG0u5pKDXkaCJNwV2BzLJ
9LJ5tiH5hj6ZvQUEaVV/kngkUERUQNCCWxrZHaR3GkJv6SLPEqZu+AP8rdqBrdTa7IHIv2PSTTYx
20EVnjR5U7BOIlUJ6pQ2nrEzyMQttl431fSXANbHg+vR+BHE3XD0MHAMgMwEnfXmw3eqzTJ+zIcg
XjJ92iROVgNQEIU0L6Wxvkv0yg3Duipzn7yjbqhjDVYgDAoRStHjMEJOY5pq8u2nRcguI1WvTYSD
iYF9Ny3m+KKLcD2iPO2dD2YhNo1ykmGgovkl5/z02JxLq134m7ESPV8Yq3uJCOIxlbnyX1RwSqyI
vT42WGEQj3fHS8CTYxKFyphxlFzoLrJUjFt1dn9fdnqgUhoan5m6ysec9HqEhn/uTsFrHgwmHZvE
oV4ZfcuYFsAKYjWjfrDfM2JDpVEYXSjRvPDwbUThVklGKsUMsiXZ2lsnZCPCy1IlA1X63+wyoxKo
XQHXxfLtWvD/8XPYLJ6uabPcympjsTVtsOIlv7+WO6+dZOwN6vX36QyJisOjqQHMq+QY/oeVdPK+
QEm1v9GUZ0oOybtZtIlaHdWhtTde6n3izYv4yIzBl4YT/VTs7Qsi/RP2XR4b986QRP5nwwrzSW/y
BTvFhS/Jtjb4czYy9N7FEEplJNCe2vLzkcJ96OmC86m1StlZ1trdodZCtonCMdMH4sKl2Z4Vr9a1
v2UP2BwSvs9ItD2q5Pv3DGS8ND5dVo9StX7Cc9poXtS8vzo2csAHQCRtk1vsW0yb/8R2qWw6bggL
Lrn1mMTbeSxv53Le3y7UGB+6XjynAyUMKWTO+tjzIJEv6put4ldojmBYkSVNq0r1vB+lo2YsyYfe
DqhXeY9+zedrhldTxvxuFqe6yFLfrwhsIpli9remcfOUfMf79HsLIVL5kDyfma5hh/mpSeXZGbae
Y/0iQv7CEgDrgZGF/7bX5oGlOS0cG1RVMcv9HkFKZitwlOhTZiGYSmk5qBCruku1aeZqU9YFusp/
DqiIQjsTnG6uk9/vw5JosmVgqZDwFjxrijCw2+FooUa+r+vbtQ3BiKeXgTPxcwCQ2g0r5J+FJW9i
HnuSFFCnk3Nc2LApmljcutFFnnFQTu8DmFbiDLENzBOj3g+eBKqXol81VA6GdMZTFMQAzJHG4ES0
eKyoC8PY/vIBmsjdVVdyGY2MugZ8UWJFcfeyQaw1oeo+N/VQMapvGTQaC0keU+HJ1whCW39aYDHZ
2+tEKldMfLYE0Gj9/TUUf2pjYIGpP6S/Ab8tmWsqF7rXUoWTfbx51mfmFvLL+yvp/j+2UOPx8XJF
Sm6VJjpU8VWqwirwZf8hV47mcdH1RP+i6mSk+w5uAwHRiTGoSeN8qMgCiSjQRtfFXELruktypA4Y
0DM0YJjD0WIZJEu0gSAa3bGihgsfr0kB1Ff2UgMt9vmVEdDE+XXve7XDdCbpr2vwtniz8947XWc0
b7LplPE7/Eg9Dt/tnkNLGifGegT6espQqV2fjg+smoHRYDK3MXFI1kQAPvDaAasUiaNE3c7S6Yql
nZKRfq7b+2Ky9w0oOPygwwMwiSkohNhaSd088OYyBAWHyNAMCo5qO7qeJZ86c6Dkxkj+VIa/XBYI
wF/OiSykMgMNMBuF0BWTaZZ1sUyl+3TaGp6t2x4JDyNR1xLX8OoaVoXtiyCkIX1SeuiIxfOR7nOK
MBGgNiskfiuNlogy5IzWSpKC1wa1aW/22Agp5NkJSb4J4pFVuio6A87b35YH9uCWobuU8dic3juz
2Lcfr1W7CJarV417f1B/4qPePO3bgp1hOl8gdOJQf6faFlnvGA5Wz26u/JMHwX6U7bl3G55fS7zy
CEFzFZ0OY5pWas0/h9WiA+OJe6HUVnk5RRCtQXvCz66UbUkAOKmlEiKMqBkRYUdAVmcrzslzR7OC
gPcrfQKqd84MGjRX5IbOfqyb3kD5DveY1OsvfWM1QUDZs6x76IBtcY9qaWryO3FPeXtpRx5C5TL9
b0AFEwEmDHwiUKUfU+Frdk5/9AjMHs+nyBdRiNoR6E8LA54vD/nQIfcc5QBcUgkIgQ5lZm8GtE8w
dn4SIAnJowJSZs91YfU/N1BnxigRNV1L7uYdm2eFQpO4RMQ7YqQwciCYqXaRvy79ayO7+EEdLzWo
ElggwJlpuYEByW7Y6as1jiRe1XjgdX2Jtk222KBkDlynRgE3t5kGMDMchIZb4NX5kXQKMHyWaa+7
TGGw6C0FqgJZ1NRkDMjb+nHwPlBlJfm7AFdoWCxBtH9JCvRuWH4TBIIBekO0LfQvLj+v9d5TWKdH
6NLAAdASuTlM5c2Y5lZ5LQ+s8WKCy74P7bY+qDnlwgHMLxwIFXB8PfCF1F0MYXTHUeySMuY+BwSh
obGovR9iI2BOGet0wal2xKEju/nH5hEkR8CFo6kc+qWfLKuW021hq8iFZAFTujX2e+Sa3JtaIBT6
nUQHprxCDSiD6lLrF73X7q9QJgURzkJq6kK4xiqeyg2dczHbsgEPu9GsE6XRN+3UAX/EGzS9fEHv
FEbsYzeNqITaG69cGcByhLNvHOuUFvOrOnlnYAL2qd3dYvnA2k/rOvVf81Dsz84fpM13OQgrvkgm
Ja1nX/iGKVeK0laZWCyRRQJsqqVNJf74gDrB6iC+PyPMD5jZXviv2gHF5r5Wd8UoyzFnKUwkYmXC
w8uVYujzE9A/fFWyOOE790UVsJY0372SQgkH5hs10OmQAlrDLdLhigPkn9VZbaRRESZ82CpX0VXd
gxVR3CGczeOIqVZQtq/3zNCMLDMnT6kocbdk79iX8cMDRcamAyjs3texYztFN9P6kkCLwOgOm0p2
OSIwMEhDVDvEnKy4y2OiDeg72lCaemPjoz5KndFmdfvqfybin8u3P+Lzs+jAUfkGETPgmeWH0t/F
clJel2ManS6a7pWQcswqgSgwfLwcZsuxftBrtC3ZiPbClICWOV9Y3ssRnapHSrjJNj0kFL4NLNuv
He7VTijYyW6a4ZG1pr6NWknbEN1mRC7c2xngV6N67nvg/UTiGIlQOl0l5Fp5lTZYiMpnb8jMiM47
eLh8OPiKidz5FN9lBooKiejJ0v49/g3AwwwgaC4a0ddEM4TUFXH7d00Uc+JlqJkz07PSDD3s8sF9
j/QpYUCY/IkVL/mG2Mh1FnS79tH4Mqxmc46hQRsgM13f+zrV9XNxdsTE1lhfc7ykdyFlg7I8O1H1
y/KSMhSV+zLTk8Clj9WQu1VnmeDJMNRbPSDYvtX88ZTc7QSd7JRoSMgLuzXQayZwx5abd2Lq1iSR
DR4rVUNwMZsy+xBwdhXsssuJoz9kg7LDQJM56rYN2sv987Vqc9ZVEBwksKhFTtw3Hh/auiRoKHE5
H9Tja3fEQyh6BuB+NVkyF96/xcq4YZLG5BFlQqkZjiIL68UiKZBKopNCz1zeokfUlRhWPtZnzz0W
7d7WoISJyEZZiHyExF7c+ms+Q+306F1DX4WAutGql7w64FmSnnuTXXY2KOxp7MCtVwO4ZF8Oc3Al
300K8HRWpxKE8dsguPzc5pP943uZnVkSD4Fhbd4KVHc5BbzErAN559hlNC17KO5EPCk7GHI9sAVH
cS4N7lbonmXVRrGLUhg/md7Wt2WnSHTc647cP0zumDjLhF44KAdEeBVECFxGLwD19ei5Pl5snNOU
CjGRHcMVEzTzDOzDwyFcl43vlN/r+sLftE8C8IYgdA2potOxmfH6YRt6KUMu+C9JEEloV7QFfpKC
7X5k2X6bldwKH8TEYHNlMFOiyGLCot+QErG16pUgFb7pLQy5ytpAKyyJfeugk+89mDqnWB9xl+hD
rkH2iU8WlOC3UneWVfXUlugFZ5t+Eo+Pc7QvR+htye6J2uB+x3UrnaSOQosT2Edcn8Ox6fpTXmX2
4jYYar1Pv8M/TyZ+5zkyqnaMJLUmZOLO/gepPoMxQIv9rO4MAOM0wYRlI1EhhKVtUrT2zAU62vGh
Ds/OGUl8RQ7A5o54ydH2k7BMY7vUpYwJYcT60LzsGbbATujb2z8S5tgIF+2nHcXL3aTE7QXvKNej
z1EHJHwrg4vt5puGkKFaLzFkgCJByaca/lSdyP4KJFXJReuN0YdMJASd49n89qWSih2CJITCBSkV
5oVyBzF2hjnM3OzPczRRb6XYp/4FYPa6wn7p7MQF6KrB1/rSPd7ixH079IdrGzCU+9KwfB9ILPn+
Lj5WuRgMX0u8Ah1IZ4nHik+qVN/DSz+qVsA+SHk+NU0PUpBQrFrRvltF+AhcHSg/rSRSl9QdMnnU
p+F6cBsn51yN7ks4P/hEAqkGTVWzpIgumCh6yAqQnds6W5LIeTal9fiqI9V6k/r52vx6LTNlVK9v
AoVxofj8cE4M4HLwL8VMqkwTnTJ6zPbLf7Eju9e97QcEFfKZQHLILmuWYDdYJFmh33JrVXg36PDn
qgNT/AcAGL+L193l8+Ovb1EE32s1IDWlTtvq3PLQ5o6/4aAOGkJo5c2MzW34kldhnvHJMum2O4E1
cZ6I15OHFgdhVqSvOFLMe2BzYqG2y9tmTrm+mLM7MSuEWNUa4huw16zpnUXG/PFCJgVFFSat+VCf
bJC+kHJ4FyFiVVdBi8SJH+KFhyveZivfZPxEJ75e8DSg/z966ox95xHjYeQ+2c71pX43/bj3yGAi
pM+b8HK/bPIC/PZMJFhVouUZZc46bQ1LmIZsfUk5mPMbr0wM84ghQ+T4pnWuxhP5IAYr1Vm1QHsM
u+LZq8Y7Eluc8nzARPu+XSmeZjJ5X4Eg5ihUMuYnY93Uyiu6lvoBAxDXrNZ5JpGD1meWAkpa23ll
KAJ0xdnkL8k4lXf51tL+nL9yUhZiTONLfmI3ZJRh/tPw7mXWJaK5Q68cAvMDCU+9VJm5pLDZthLk
g1xxIzLrYd34B5vnYBI18/ZAGr35EoAcW4+TCVIM1my1q81S384YbyzEELNDSMovf8JZwej/mgUa
hb1fwX0jPVh/6PFIROUWFWiKDVyQRFm6dOWcjS1UyaRl6ev8Y16SpGtpSQ+Pl/CA3HK79tuKR3se
5NBD9+LACcV8hwovsMP2BUEoBbnouXTKXKrvnrkslb90IRXkWf9hCrk/7GCsR3feOGX0ZfPOp/Of
1ffvFr0XQUBBnromcgzV6OoXG0GLWoj40Ze2UkUP0gCAPHlHduA1OYeYverEgiHdRiy3okKMLk0q
9FHypQClLLd2wKbB0sdVZLsZRpRPCPmq0kojYxHnEW9sqTpV+Bm5Km25PUY2KSzud7Ib/yKxMFj3
iXEqk7tEi8XOOYLzj5I9BrW9nePSyqhty6rJSy1QYXdLAiB42t80ByOgR+h8enutJSSIZB39qO5W
OeWjyz7z0hbCrlFs6PvwIODZQS1sxA7ZQ3B7MFOOJAk6egVDlrCD7hjmR6GOaeu44SlpWddCzUFR
YbqExBVLvL+06ApHWMVkxFKcb6TZGheGUw2Gh9vG2R1DssBSPvHIxY6vkTEYsyz2AdWJu3F2WYqd
Mv578FmF/8sxFaB6M5PVsbquJtq11zd2dNujpjv+IBTOyE01i/oIZMdWQFxC8DG6uuE2OoZTFa5W
T5M9lIIeBu6T/77vx0uH+4uK0susfjz1FXAtdpckpWnPqXhyWBFN9QT2thUlIWbLA3EUR94Ka0s0
ctW4d7CAvJq97IYaNBIBoN8YzJbRO/PLZoLCBfE+vd50845+Ut0/sBZnzrIIumK71rMyR0wS27jp
GDUVh7LuARv1F327h1PRbY2roClqLp6bz7TXEQ7mGGWsdIJpgCapWWLMnoeDsfjO82X6xlRrwwiR
XX4iNTgna3l8QtUc8IeHv2eMuI7LhvhjViLmH/sOyLrLN2fVKaR9Ge9VLzYv7/xafjmVC9afW+fY
hqYqtZRP8DZXyuyDYBXqbdnPLiy5rctcmv6eR+COXJTvFHeY13wacI52Oy4ngQb6hJ1+RPmQKzrd
/SW2wIQMqPoxtiElFgTdcYD1Y6qk1SwIn2bU+8Zgn9weDdYiXCf1dyAeeoshas+IFNpxqMXv3s8N
m+OZx6hUiM+fH5F4BcD2kktvDRTVv0N7mBMAqPfYuynNbVa2FlfPpRblfIlGXznssven/YymMAh9
+kLtJRUbHAlPZBqR0uIHmlokeR+N7i6vawX9tb2Cz69rKD2jAJ2IVfQYcm54xJfSVpXsTvkUgg/C
p+YIquC3UbLJM4UoJmrEIcFf1gRgQIg8JzgPkQh6mqx89kowYC0KXerrWSMTocc9V+LzzuyWnc0K
2bkHs7qH6Yv0QXwXmatBzCVDFvLttUUsV4lOlKNiqSlQglQRcFX6DOtPYrmQjze7gCfEx2kUu6mK
XryS9yF0ul1hQ9Swjus0IMaN7t+Ex24JZo/gQiIHt7W/jZXX8wYXspgjFrHJ4sMMiLvUbqOAqi8k
EMPNcQodX/e1ViKNqto8BlwqM2vqhptar5hi6PSdujlEKnmwPFTvseJWCjkwHxmhBhvPgIZf5O2b
sAi3BvKsv2n/R4ad8Ib3w9YpLBQtyWuZ8i8o9KeLhn7LiD/DNkoTbdXLMhN+JoS9osnp72+yAa2d
Djzs+iQeUDIqXeT+0DSnNu2QGfi4yRp8ldWqMLzZeU427rBxIqVsYtDXD6TgwAn9NLVdw7x/grFf
+e+3fBrJlVfrUJNMlrxrM3y5ifd2dHqGIHKzkcQF17+OkxwornbgyS33gXlCKlWByBkQ0axSlf7d
LxX2EMpmqZWJnzal9U3C9PUiqmXPAvq3zkSsJxKBDeBo2bdL+d203Pyiu+Kig6JIVyloCEssS3CI
X2MI4ayxMHDIngGEtoQw7Staqa5+gYfpno6QoX5mGy7ZjLCslLcZDv67nlpjxTSPsGkR1YavUEOW
p7Q/2n+rCtpAiSgNJVb9IzUTVb9ykFjDMAafaUjPZOjnJj1OG/Xu5xXQ3x5jq2L3d+V0GmpyyJme
XCC+TkNiEF0h7oI5SVlAqb4crT7DFbH6CFWXyoRUILj71q/++zVOncNg8ipbtaJ9cnQo3T70HQrc
TWUmvqWzt6cRtia9xFNNI7/4ZqfsOmf3+5N+VRb/VGa0GZk8JOP6pWw4oFJ0BxBFqqGhlZg/5uhe
zpflyzpOGA1Eg/9wVfab2dbPDRCLh8Mq9zYrsLVBwLvWPVPf+TwxpLrZnfMocf4y52/7gQjfmmrG
FhVQhOmB1kAf7pabA4QMlFXZo6YZyuMFQl1BApVg9SEdKQ/yhVY6GrXCa7+aYhl5ZZFXyivrsHsV
gzV41WyAbbnGnHxTcpxvquwjwOyahbQ9WXXgOwjMcUg/X2Wj5BjD8P6JFcENU2okemLhRp0gHKSR
2dKgPNHvH+dpH7d/fuuHGnQYbogiBQETj7QrmK7bTn9f8FhhIhxbtdj8KPVf+BF2cLSCBz1LVq4v
NzJOUilVofaUcHf246Y6RLVsdq+rFv+OLNuqesV1khJds/GI5Bx/t4R9PIlUU3xYviCm/broTtpr
vrVbzf6Xj45OjjkGeoMSV9NQjF56M0nIydSBEdyf43nBKe3ep+xR08vfnrNVYUwx5qF9Yxagn6vi
p9y2uVBbQTE8nUKuxRtlUpLRIuEJA/zGXQ8OogzRZEywFL2Onpge0/Hc8Ar+BVYoYY3g4wLKwgb7
3GvR25eq+mS8Z38JhyhTSWEBKsD1dzf0bNDkYCbOOiFDSqRmgCt20vrDjtf0v+fN+o21DdXiUok5
AnHc5ebfV7ssEer8BaNlHze7HY/M4/vQyJpHAkmXnrCR0FbVFXHTxVphpZIbiTami8NHzW0lqTv8
KkbWP+GKcsNc7AOmXljIOQlEKZJqQVJJLXWR45ZHA/ahEMddD7bfpxQGe8osZ8y1rpTruQi62eZj
pZYB6uC4zeFht1wj7sPfkqFACPQ0TZB5za4Q5/zMZEjQPJQldxV1OC159DkZetJ7Klh+3985lxQj
vU54REWBO/Xu0+UTq5nFyjd1b/NTjCome/OQ9fH/1YX9z7VuK45XsN4YuAsTGJTM+ZRSgpJiQvgx
HHmR1CxW1zASw2dwj1o698CGd0UpNnV3KYotf6Y2kMyqIQ04V+Y0WFaLtjI5ANNf9O2zNtL69U0C
iSNpis5uV98YqgVgswR+znMrWyUOChX2dYUNRbFPWKBaD1Gq/4DWIbDKIQ3c71RyPLRoQ+748Qw8
QarDGtzey+/CE89s5MLaEA2WXiwlXgZn99YRLYxEVGRykcyAXx0KKHlZAuNaEIDktCZEiCWf0Lk5
N9JTXfF8oinrNwbqpb6XSn3rzT3tFfNcbdWHLw80Df3IUJ7GqP2ZB9EVFyAUPWY1oau8nzYoR422
68LG677NWPXKsoWdVyaAng3STVmrLP0W1+aW4q/xmajqTEKzE0f9Hcn1Om/t86QYqHmt8ikCw1l2
DyoUhsocvcziZVIh21ojSR6D16c8auRbc2scxXk804aRMIHbLSh5SN+Ls9mU5lY33XXN4fuCmOpl
doTFqrUqMK69hqatV/CASihZOkkei76nwPj7hBmasMzkH8k0vodbAYUWA8VBeRX8JSk3R0PpOXrq
fMd2MluKJ/PujdRkNhebkRVCBcKmjJvKyZXFkSImpMlOAL4XW5jE+x80yejQXkE1z/sFX8y+TeCF
LFWxVnPMA65qIeqNirwVZSCqNiagp9OF+VE5UErQ7Ejb64eFeZSUP8jrdExBV0qTfz+YVJ/tXcQB
a2dwS0zN9Dnsgisgj0cY4cTceo1PQ1qrDFrlFa9hM1kie/uJgihz+z9p3gmtE4I3u4ex3DS9Vnp0
xc0hPxmfeVOlDa/lKk8syznQwdUw05c7lMh8Aa6/TXXdjW5gcdbnyXVwvbz7U/calov3ZoRWXyIk
2e+1CAnU389jpUsSDQihsIPqPIfgMJ4EBweARa0L8bPD0qRrkMPKO4k5vSGNviYYVX1Glb4psDd6
dUEP5KM4OrRrqJvRUHo/h90vVA5b+QvRGaweju5VrjaUeo8+hC+GR/IocMzQhChZy6q+YgxNdgab
k1Doybhcr/HSJqmTZQpUK+zyRLp5eSvTq+QsGgQ8RyqtPucIPsCcxfZiXNsofyLiiYsYF4RwmdPL
U+/FpjbdPEVQ5Dp69M8XDV1VSAJEqdOi2WDc6SrklcnNx21IfFzJ/D9qnc4zvdbceP6I+y2Kv/55
ghTJBFKV+aUgStZy/N5qkq8ZkJ/8ftp5OuxSvjUDeo1PjqBmZZHHgwwBmBPo/y6FuImnxz1JaV4W
gYdmQ+Xiuv0Kpz/6+Wqkp0XaPnDFlUknB5yc8Nl3/Z2gkG0a+85J5E9sENUdbN/GcpeKu3TtZGrV
Tqh4GztMnXm+h3X/ynXTpCx8JDvjCRUa/I48fuvMb+eboOGNlnU8HlW7Ihvr+0regjvO6awbAVYr
UdQLqKPTLFBdmf3ZR8aHABkxrNZxfJ+z+2YwevKBHzdsFcLCumUg+TzSKud5Tte6bPRuBYwsHdIx
/3fotfiaiocWuXtOhL7L8mkRwlNZWWPmsY/oc1Rtm9x4w0oAqmFRqJGxULV1njSjf+kp2yY+n9bN
QQoY33J1ipw8brO2VbEW6QMRYzxzpaaow4LvcQGps7H87ntpBjTIT7D8a8M5+NB+wDe8f+aAFH7L
0PAyILjmHg6OeMgjkLMSEzRkVMcpXI15XI9see/xKrTDtlRck0mvKE1upDKs8U/7WpYMS397LxVN
pZKmnCIxKXhDkprTXbJ9pxPj3rbYIDBWlDanOrGqw/z7Tq6LdK6wvbcMA6yOd0PrTEZ3sH/VSCpK
Lxb0soKgrz5dTJMziYctYWlW62tFoOd9wssg7YXeMV/qXj0RPSme6gIxVgKDXvgVpEA0FAKSNsaf
xiyaHLqAfKQ9LYRcUd9n0bZHLK7HiS8DtjCvJR73ShSIEj/FyJZiJvzS/8lJD4mCm6WmJ/Fdtx2G
VYMklXTxZfBhZXfE5PVUW4Oq5k8T35JwNgOH4pEPKG3HliW15em7pL25cxUnu9KRAdKDDuLPLt1I
IHk3UCFW2OV1O14n3WZW+zjpmx2UhT7GYEzLkanepdso/WZpccLSRAyF/5y8MJLjCOm0WooT58g+
XTtnkgoZKb8ZiyQnb9630HNgnLrvBFKlJZKwm5CyCwpAKFiKkfMSZHK0ONIK9L/JEBIjrzYxvPIY
MiSxVe3jXp2urC/atUjj4cjhlG+qUKTgyUzui6QPLGDFGwiFoJ4Dh9zrsoNZSV2POodoaWvhVH1i
e4wmvjaE8uC5F3dzVQxz1qfniWzlwQrk8dLrVhtD8/eVXVg3GVbfQPOaS2mzqyv9tsx7zu+zdb1i
CJ4YrtMSfGo1WoFwxxIflYi6XRhjlsMP+7BiVBluX4ThC69rbJsug5udz1/bA3x/GlA2SPlj1+vY
8IkFQ0NBmRBwZat6DZHHcxo061PjYCpKIGjbNaxPi7SU8wMs/xZ8XKNdeccxJXHmOf1op+UQD+pP
qPoywdraaTyZwXkfW1KRMCaH1vQhn53/KCTore7r5VhXQ6JrATz3yIpVUGVvQhv4mND2bmzdVMVG
v2YdK5t1+Ue+gBOqVqxAtRPAE3PEC10gb/0AVT/T7WqKw7zLouYnsy6BUfyG1ptHZSkgyWpzoX5k
mTGYtj72vlNF1m9yeka+OU29osV89BJpEz5NZfwKQlGNv4ZVSq80MNZxhKFGT67O4vSeijT/wTY0
zMu4nbRv4t+vK8HFhNPZFvGUKBz6Iw6/OW1GV2B/V8LTlGzLtQaHCMLQK+xHx+DYbKS3fRGgDuhy
j7mdBbC6LP999FKYUjtz7+gKOz1hq9SLyiJ7VlMkpne42C0iUG+1IPTcWoPvY14YQ38n42jGQSQn
G3s8cW7i7cxxsXeX+1XQETxurq0lLek/HQ6Q0LOlxXrM2fn8YeGmjmpuiMC27Xkypdmup9shwNh2
RNd2niNXep/R/v/TSZ7aW+L9HI7oWOQz4m3ChvF+MLwDBu6yZUQrZ38YbG3yaNKk5Nwu1B0VOKcH
lA+xqw9uREOnAIVfqwAT40kpg571FJgHIvwFyZZkBHRwZI5slDm6LYz1q8IKeSjJQ32/qLk4Nc2Z
4xaD3x6MRh4SATGrtbLhE8Ry/oUBb8nFaFX5YVeRW+pEpUsFOnWeAUyn9t7IJayb+f0ZEcm4iYvg
0sq4ZJpDi1MMT/IxdQGUiqWkcdSEWt6O2Ue/oe+yom2kjdGWCzndD2MZBxmHx/ykepqrzu7VtLDt
FSyxYLMlSUQPYjN0iDofDdEqJByjNfMwKVivLrlr08/etTPaZtni2ypfSU6pGpSVkAcxevYdWVCf
T8BSCbXXw1CNcaKwx/M2Xb6HFlh5qFQ4qxvJGIEJCW/vExaXskwsTCR8pUGn6HbaEiG0gZMnxIqK
7spyOUWJkqcF5/gsyHTlHQFPEQA24P83rXSYB5TD6URATLGeQ3sbGDPiWEyqiMQA55JRxIVv5JZE
wySKMrus88Z2JP6LfZxoOnvTCKZ+pV6745lOgV1a2DhAgrfUtjvA06zC51xar5HXo1d/jwxlvUuB
cpLci+owimtHqMKq9sdQdPtvtg1ymSQqG7FNlcBeLCxYl4CRPSJQFeouWMWWClIGyT1uQMFAtWy/
FVx4WxHT9mPyQkvifAEnyh+aVJ7jwp+5PO2HMGSOkySQ+j2pICy+uujhFnsPtblC2hv/QNNU0/++
x3E+njbWrbeqHjYrByt8oZfIMBJBibRNTen9P6Bp6tUNMRlt+DvnwEGrx/C5BIDAmBmVZzNhTfQw
7lHCgr27U4402A2bDyDj+jFIXT8wJqHgRaJSeWWxzw+gOeryspnL85R4vti4ByNz599AG3uti1vI
a0ydaU6Pv2B5VMpeyY4r+iH82/0Xy8/OBO1godbHk5NJz0a7ky+yrY6xUnLg17sga7wiUKtAd8ab
9yuIvnr7oSLk20/UYeTXJ+Zq69rLKf289jz4X1o5D/gXabuCLRlET9OBSPEGcMnJuoP4XU2+YJmo
NXDsKeEGjlPqiJf6YH9gSAXhT+LQkz7+IM+vwHH/XR5I8UIDNEQjNJAkDojKiZIPtxbtazQkJIi0
9tsB/S8dHAyRZ8A3UihM5YsDL51NvMsoGc5F13JTfkoz0J1TjzdKvMKFW8RfeJIivOI2333DdplG
JzDOj9bKR5FOK2uwHzNEWEF/6IPIz8gr4+EoonEizs1bQiFBps+hBGUs60i1zTdrKGu5ckEYl/t6
PGZz1xouLVUY5pfgceFDsqfL1b9qOfuZuNJcL5jwUGRHM1hVuxsNc1XktJUMtd7PEEG3eRL6cgeq
toZNRicLVuKI8yA07IXP6x/g+uvkh4BACN7DWmf8xsSshzn9L9BpLO7LechzBuCkYRt5E076hxjU
xdd1uQxRrXhSpGw4GBR+FYLBmMq7qOV2/LT7mHNwWXHXA5Ed0cWAS2omgR9NQje8gwUT/uS00BZp
qx+JN6bakYKqPN/RdsNZTEA7WvXm7+U1Yw8dwAn5+ChFPe3fHGcz/qsTTy2Lal26FzvRFySW3i/C
C+Ziv3k9BB2pX66CNzMVwKwVY36rim8d/TNMRjnQaZ2NTkLyDotd1P3Dbs0bhHPg57rkBHXKVgXl
d79BPu9S3u0mJ8mT65S4PSvwhsmsbS+MjdxGxp7GcaMT5PhWLiXq9/38fU1vXw+fO+YPyJMVkmCF
Brc4GREf95YlvNjCDDGgE9g0XHWXFQONg7eYZlsm2O92BEge53Smw1oR1v1atsqTAFkCsh7tytk3
shC2Q8y81zH7SCv9MfxzaREpaayz7sQ8iVn7+X7QIhHCSeRWcBEpvO93YWx1bR7DvQkQxmk/W5Pd
jkZwXKe6Yya1CupuVmWKxyPz0QfKP2c/vZPAf/XnVgNHJGLEJMywpYyEQN+a0brZCC/AVIaV6FsQ
P/0HRzgDlooJ3eJsbQQWNl2MB3Fq4rjLd82jQHd7ZrVlFiAgsSMogBp2T59WW/qQwY3zVICEcsfr
2YlCc5wmRsGB8b/eEbIz1lHsTRz+x6TxB2pw8GBP2zoonKmzHaV4U5y1tYxzts2OVJD0wtxJiXJv
tEga9SpBKhTdDfxEsdW6J46PUMrBx0CU7pI/HixIx9g8tvLc36JmtQjcgmu2LAGP0KuEAoCYkAJz
EqzuESzbidQ7oGm9LCgDEGZhz/qtqdFPruRrPsO8bt/O/xr74NQX2DyjjuQaGUHyCx2NKdLGgBLt
sIkXNQYlptxKSOwydkOt+WaBb6QCxS5dUxWG+C2phFybjVk/63l4eALmkgfh9dsXoaF48puOxB6u
4PSPqErRCSRqrdin/apSK3PFSRdSog2xJyttBfye7FvRVy6n32MINZraetuzd8OYO01U2Iv/Y0ZH
3ofHuc+53NT34ur7V+SBAWhBAFtRo7/Ek7P6shSdgcn+g3Tp+a1p8qBAgg7MoMN0uCWwkouwowE0
uDvq5WFYQPRrcOw9IB0LSpJ6NpD4uKW91MzmM2g8+9z0GGO5yjKBFlqT2NSA/04yZyUFk79dftIA
sUGxOGy8KeLCITa4AhSUfZ+B6Md62nXsWo+XJIMBHiFH7z6qnrxUZvUsLOpO7TuNAsHSzAWAFs+V
iBxPguUu1Fkrhy8KpvxbUbeXMnlZLETPOEPMQinW2be+NPpeR9Klxr1MARS6Ej1/R+gssrbS/Hnl
v4Z7V/X9LQtP8etBLwzfjEUkliCmnXNZj5RCziHL96baPUXoOUvXxpme9m/LgT/mGa3V+KwNCy2M
cBitwFkla/qeaJ2mFju75VqRLcv/AN83pBT/Ei1rY/58yZ5dzCEcrg9s8tveBEWSCLmP+5KYkgjb
NMNRpGlz2apQ8QFIIVRXc5WYl0ECVhval6hQFVLxVgokRLvqNAJNdCOyZyFZKj2HB87k6Tsa9ZUq
HKDg/pMWeWrQ6ybFdFzj3XW8394lkkB09JSvNV+WZepFWgCXjPvxNHkd7kyCUkFnvoEMX+DT0idW
Www/z29aB/ZAClIw8P1pjNq9PIJ8+4Y7S1rzF5fBeU8W8JkIxeZYF+Dr1EvJ4Fv2F2XIWOgyJ6Zq
OlK/si7Wh0gg9TVDtkBXBb/TatdpidE4SwF+Hrb+gn6cnJZT7V84mdluiZ2WBgn1iMV2GrRJ6hrD
a2UjUDi5KIBH6WHEY9ym3Jtack7g+pyyq1LwnqmAw/hFhqTvt1IFgm8i9MojpoOFsEVo7WDw9dzw
7toM9vSZYsBf2K+8Sgp0ELOV+s0Ohf/FHvcuPaRTjTsj2yjigoQcifyCyqLwlym82yFF4I/lRM2k
EUmguhYjRHaOfpfdws91svas80XupyM2oyvF4pZU4c+Atw2Eg0DLfxyMEm5Bbn0APRvxQfn5Dtpi
qtnRNVarVINCXy+QTc3curaEq0acw0O36d6IEjoJTt/UodsDSdYjlmkkzYfk9goE1zorzgPWXOLh
C5CiBfVWunTHT3srAh3NFGEtSNplQ2j6MeXg0ww7Gfn1QOCKTa7mavaN4tmm46Hv+D9ba/LbWJTr
w0TKJUqn++xoPSMAMR9Xin1Lt8SEpxJX85WHSIYAnLFehJo393+VAZNMLWfSjEr5oIiaYdvuI44Y
GIJj6L+mKH1tLifxkZLT/SEQ+8CTTINYPHXFdkHuz89OmQo9aBrcv23MfwJFseBiwA4wviLQO4ch
AJiPWkZfl+2yHjw6+BObD2vJt4skyhg1zNyeKFKZyJXyrZ+Gfm4HWOZWhk7A6K6JHkwmToEK9gYg
VOpVXDxOP4GBSPY0rvyreF7Dw/rWL29fY8dmGZ+XtQUsJhL5sGcZXrXzNrXwms1Kk/KPNBrKAi66
a5MPVVcf3OEpggzsESUtTTuMN8NbLte1nLGRZyiRd7bGRax7OjLGMqxIekqHBD1+VmIkk3s+Ga3Q
jJbFazHssJIXz8EsJeZA/ytphk3lKF0vcGFeTROsf6jq6ldghHo15ZTnGZ4wipa6/XSrQCQj90LZ
iZjpg0TBS3+hSVIJwIdw39CJXwxIm1j1MaK8LMdzx5nOQVgbRS8lY11JnKI63xWpto0vKDZTqJpM
EB9C3SH128uvE6QM0oZjUxVTlGLq1Y/H3vvBC/FZY+eKHXKHUp2nxSmabGXz6MGr+rQyWpnHOJAW
+lHK009KHjssZQGrj/3sofL3v7gZ2aq52TyCaqNQBkEF98lq68csN0rLnlEp+NvrdRhOWUmBA/wS
3wt+m+jrdbw1ifO7izBJOjwowFkWD7yjXWWEzQbTID5ilqwmmE3vMp4eMcJ/tiQAIE8ZlI4PzKe3
tbTrxtcD+2WVojoZJ57mWGCbQlO16idHvogF5G895RTcuHeRNjhIPOF2cqIGIkGaKS3jXQZLVXsp
17XZWTKla6VcnkOBVQkH1IROyeawZQuX3IQbHXZvwV9Ah9kl+JZEPz6R0KXqYd0N2dl7bulmziwF
IKw293s3WOfrvqw/QgpHJGPXhbnooByj5I30vf/5qJLBihnlFPvYjQF/POE//jFJmhqfy/d1ZRFN
U2KKqH4ldMEXqbbYZH2HL5UqanAxz52spdidAPgIVz94UTN62XKF4bKCbE2aBJt404T1rjHEYUe/
or3iNLPbCbTvmL7e+oazpsC2zB9R8Wb2F5MwaL6q74xi8GJcnLl43BYEBKvpL8P445AmYIIkquVP
qZuJ62P0CC/D3nJV/9y3usuZLJoHJewD4LinUgrQls7tze38IMRudBui8Zr8YAzK3mYxv8LYEaxE
dV49YT6dNwWc7d8x5i6NaPOAKBwqSbdv/9poUW3y5jfvK30+Shv3sOpU89KXo9vMPrZ/+ugf9Ctn
vC4A9DbzzD1k8kMu/35h8blZmr84NSIqaNODobmOBaayVj/+VdSsfSZJoX/pKvcaWpoKCmtzBbJm
mV9ZDaRUectdHpzmC4mEByuDJNBBLlYhiX6t0A62sU07FFTYcUUhZmXlu4XyVGPpkB8pZHQIUC0o
Zd9MMAbrIxEjT72i36JRePmF9VkRUkUrbDd4A+Gw99I5h0c2kpPOpzj2CFKy9UZ20N4C5597PYft
Arjlys4RnSYcm4LpOAGbstrlmnTM5XCy6O7Iiti7DYSnX6QhClzQCMw4SB+EkXcmSxvYMmVbeG9n
ho/kxadmctREaXNKu8C/Bj6nEFb5yQLAmwgSRTH+nZzuC/0Oze1KJdxa+Wam0hx3h+Lm0FKZF/Nm
PVXbOmACUb3QBzywpBYmjJnH5X5L7cqzS5LjS31MQnYdVvkJ68utrnbO0cTNT+EXO3LBXEzHwjoj
SFJ2Y7Ylh6BiSq7ETRi+hqbwFreKPRa7fxwz6LjZQtQUEYr2OM3qic18s5j4QcbeV/0XUg643lOe
ZFNKNYwv67PgN+6Ojgm1sVha5baK1X/0cC/VLsOPsNDynkiALc2E+p0f1a/gcp7QB1a7+/+UO+Bh
+a+MK0GWQUMKGZapT8ZjxMU7z9xBe7H6tWSlp317xy6sYTfl1FyxXuJ/Q52bB/9Gs3hyO4Gs2EqP
VGRYgcYs7FMWBtkcu5q0QtRBzOefS5eZ0dSCNxJvZHByYrMR+lPm7Pw7GzQCw6th50AUk+jx5tZE
orIn60kAunrSwo5go+LyYd+FFod6hFqSprWKojUsu/ZIqizR1p4i0KzbiaEqt5kssiJ0xARyvpEk
sNZJ7blJiTEnD0Tff4KHUiD9vUHbdag0nL0EBIr1qXzbsyOklPZ2l7/yA9in+lNAE/TNpmAMa2DW
qEkAuJa3ew+gDPMtNIR2UW+4/bZev5r5khbGvPqpI38GjgXQDacujW2Oznh2q25ovdyCy776R99n
ARZWs5KhcRyxrjlhzX/Qc7sUxG0yMdFW+NBC6Nx2thG6hDhVi5XEhyiZugSBGlY6tYX08xnC5Jx+
nEa1u9sRslO42uKbQ3/bOHnB0Mj1NTzHRVfYun40DffLgmbRvniWaPJzkUi9tniOa7qWcp3V/qdW
gPvAoTFMmKQOIkCYSgWnpH2G/ZUHliKV+Y0Y9nBK1ZlcNrTxQQo5yne6McGZJuCg1NC78ukd9Lyz
dPuDI5ZnyZoSiD4wN59HT6UhIFJvhXLJT9nCAxGTBmPPtSbcwuljhosDiHFp5ATxGV2uvL1t7uqY
8lYWqHcHCGJfzPzGSJFcvnz839W11N2F6UU7WZpS0gm3Mm+OruqrIBlTTIFlRBXmHfbyfQBOcgnI
lUhqKcG97vaiBhBTA3hMSmZWKGBUMrgS2BQmJkx0E/poIby8Tvaw4r6EZ3ZtswGNr4nAIw2CRjI6
uwtBSSnwwfQmfHHA40Lr4O43iIfs8kGQLW+mH0i0w5KnauFG1jCc3FWekLcbNk6kOr3czZCPDJwM
QilJ89gENk18BRHg3/Qumi68+eaEz3VcIzH0XRjSgIHVXHZ0i8WbQBn+EYH11SVy3gUWZW5yA2pm
o7yXH9HI6nZ/JHRS9lREpBLAuU8JwZvRPPvzk3GJSO6OX+9OJlboC3Jb8As/zpUD4rIwOYdZDWdj
qWVd26K9VkvmEsd4R+6JmZMyo+Y5hu/9gSxp/YCwXczNp7COCYl+vwjVPiHWygyHX3+sDDOZmvec
9KpwSK2Wj3P5vwIb5Batb7KhJ0bjOtcD7CKr865Bhpv5Kjf8xGpE/AG14tJMVrhBczPJUJKlLuz6
1TegnwrHya8RCZATt1ql0u8emyn09rBO/pVMxOW+CxufRw8BMO8o2GhhF3QeCViZ5jVHdZZPLw2T
YBgWRJGnZBrLF6B959kqwWtTYLXwTYPmwJ7AwD+AitCs3tvGRVMdP1GOdHiVjRl3/R5U2QUf3J2H
8fMjdDxfMugObDoeUDUB3h2oLwOngo7MOkkYM2ib1W/2QflPpuqlMcWluaW8orm7jDNQG4MtxGI2
LT2pi1rump6rj3kYvHBSmcyZqRJjsXygqrno8UF1rNUYoVaVhbRdm2U6dJsey6YWdgtVEaugkS4u
Ms9WgUjE+jLdUgzN0Qn0FQBMbDw5bI5c2LjPX+9O98hj9FF5aLgRWCd5NskTp2a7xCatXSF0ww8B
ZFDpxPuoERPWW61DNiAojfecwJDrMH38HMjB2fv+7DclcptFdyrfHshuQ2i2fnLBQ3D1POUdN1l0
RGBoWHKAGVPgjdOnGfJwvBVV7wxOiMv5hZgIT9Dyg85Kbw4ZAwiRE9cnbONJTYIoOKM54VLov96j
bc9lUyQlmyIXTXGJYZX3Cv+ECqYTrxmUC9rcPAD4zAsMivuB8kQSGForWwmnCjO/gR+XTsRk7ree
YDN9gL0vJkra5Wx++0mF3zj0dqK6ZfR3+xCNiKitLJclT3i02dANdMy23WnmXPYufszmjGA4f8bt
Htcv3glyrc0/+0taKr5AjqejwGwgvlB80t3vX7Ps/yBzhyyDBXWS2JApH0PF3i08iNqxJvcbVb44
j7Vh6TKwD22OIgLbWYlKsd/Rnb+AncbMCFj+GscLlpQs6d1YE2lDYS6EpR2lsaXkWVLhsQLAz05a
hcF2krd2Gt4QCtNYxD9t7vjyp0O3ik9JrqZ4KEiq71fOFz0ocf910aAKFYG34mWmHoLxLDpXdNGK
xhGk8K5EC4lYlAZd9/eWTVTbZYImJsvNI3YJ1y3Xxg33bmB+FS0pvLfBssWEHGqkc1m+boz9y/26
ZB5JYbcstNvYHF48krQ+dD5RtMPgehkdIfs3j03JIWGo8TGFCAtzcSk3vLntgd7HPYvtGvlHyY0K
Gymn4lc9k7HzDW1AbZs3cKo3fYh/O19tNSO75AwxUYKxU02EgjnNfpFNDU5ii88zYnY+DznpSxKu
PKlB3pVZHMGhTnjgorK1MawnqlwueVMeywHc5DJgwcCuaCOZzsnF4sAm42nIWsYf/xZHD/qPPQcE
dYqPndaFIjeTdITSu8US2uzRTPdpK45NyDhheIB+uv7HmheRTTZf5CEcI0LhLkT0qbVunucleb51
Sreh2i+ic5YUwM+pi1mnCoTgzHjb926XRlXdbSVsEhfpK//sxgQBN6f4MDSr+q39c0lF/jRjjBVW
ju7a/CAbSI0BJTMd0W6s0ZqePK0AcxAOTDvsCoVG0m5gZpkye4R9lklkIkGchoirbZBp4teERyNt
oVVjtkn0PrpmpHi5kq1AC8PEQTlFdRvt+/hpqg4fRGRtEzCbP+hJEqUxzE2WjyTfjDqsg1mCMEFz
9z1M6SnS+izXRGmmi6foWEeenWGmsGtie95zr6wdqozSC751Eb8JBtDu2CncldEDK/q6LD0edjw3
9bOYlfX1Epvu4G8NSVyZcDW9DQ9PwuXKRrgCavuxeORR290kRXll5G7TmfSp4LtE4Xi8lu5woiKK
VOQD7ik8D3ULdgiAW+dsW3YS3DmMRpqIYi8oCCh6TbNbrqhCkat7b8Btm3kia7bFDj3ghDGVELXC
jhof0aUI8R00mLN+YZM/zSGVKJ9JoQrpF5g9P2IrfiRhI3Ai3RlHqjJ8i5lKyUkNaAeIHoVuank9
pKRbBYkZ3f16+1DrWrpemJ/Y9F/1T7k3EBZXbk6R0GUfYutx5jSAV18L3jNH23XG4Wrb33K9D2+Z
23Bei1F9mhhz9HY3qI/JWirzwT6Jg8MGEes1wrCIay0eE/NpIq9wpqiBbOJcjeNM0nWkHlkkRRFb
Pmo85VOqLxYeUzqjCmQVHlqpDR4sI/eLVvElBvc486FDacBodjMpzLM7460pxOEk/bCHQw3rx4Uk
Wl4NB0d2KPUJXirdbAUTs/MPRQ7ITZdrYLmlDg24I2kLfkA6uwtB+/t5B7CiufSLeHKVz6WBYcIt
AgtV0vpnIjunSbY0QUxQFujNILmoYqnkgOIjmpE+UEfKajhni22cAZUDJLfwAIvZxx0gbnRNYYrl
AHyApLzvjzXL6kfEd8XVsGMLmBXiE/HJrcANL4dp0Z1wdFpkdh/NZ/aw8YhHFO1bcXY7mcgLg8Mf
nRWghkva4tnoxvTABym0hGfMBu0/khsYaT2olbvhZxIXHfdLS6nxHvsWTdzWPUzy1pEg9qgySKAm
bkQQ5FS99r12KJ5qDOLxFsyw9KRTccDlH+vAtmowmvsxgJ09T2jq+BKoNrOt83iWzdR/5GgNvS8U
UwdIwGzJuJ34FVw4j8Xbg6FRnoGb8tNdKBklrY/+gIeLPpTLtpX0TFkRKzhCpE5l84Ek+TBIQ/MT
3zECFqBilwIiBqbg0HCm1jYYQw6/wl9bihCIWWSNNkJTDtU+y22gcP/7TMIGTB+pH1Dhy6btFaEW
kVU0znnta4IsuJHamxIxasFul/tsIkMGuHZ95D2F3mhbYKUXBp27/fG7LH0MvaLxg9RVWMg5nEuG
WlKPgAaADxamFMieAO2UeR8iXacHFDwzohWBFU/DjZA2ChkTpUqP2/diQx132cBoCKS2XlqENWAl
YgHNdPEjkVO2MxUQIpiduq+TmnP+HVC6BOlTPGag+8i+98EpsUXqPqOj0CoH5myePx8pjNukkIRn
cfjBMDCS61g12OLi2NJ87eo2md72Gw0Eujt9cr6drOcxU15gZb1N19haJF+3QtXoy5ccD/o0uFo8
XxVOcw8DjLKAOUyGRKuWD6ItvqDuBbgNiAl5ia4iYdO3ggUhZYF2Q0aKF71Wdr4Sekea4jbRF5hH
Ec5qR9Oqkxw3ADMrG0UJ+B0IhY15xTswaDY4P1ZlfwNxe2q0sPL/rclPXI8VyWzz/ceZfxsrmnbT
aimIBJTYEgnPMwk//ii/pIkd6+l5mHNy2IgcK00JKhNk499ld4TPdjX2GsIvCgMHEV/sQsCsZEnv
7pCO+Xp9nq9wycRrXEndLS58UK7KVmNmFJMpyWMtiXSNdQ+3m1OpwSR82g7w+qo9DfcJZrvInyIY
qhdXFhQZsQR8UZgub484nMmrv1ITBS+WYq+3WqpP8n5x4ISrSQeK+QPa2x6n42Nod5hnNxnFmFgc
DPSuxkmL5BXQPrDJV1+/PembGIomjj2Q/gkTIVrmbhpdFDSzryKp05ULgJUAUdtAJt6Mu5vCTXRz
T5oqJtQwjDtigFKyDQx1Mz7SX78LH681UHi6xVAf6eEsDqzI+wugAMBgJy7ZeeYZGZXrN1o6eLCB
JLZEaMgOeEE3dEi4PcNkgaKQX38nH/7M3n9MtPSOwoKAo+xsBAZP1Vy5379jG8U3HYPUvjwYAs2C
sEVrEePlS9eLoPc8zajT7pPUhcreG2iWPAQlPyQpmrfkCDNmP7ulNHRCk42K2Vy57rfpevITenbt
22KC40Mz9c053AW4ij4lc/N7ZwA9je2mLe8g86ncUssQhaDTxR90q35bnfTUJBeHsn3NSlsCXtEG
eko+aVhc2VCube+ldYe4cX6rLXOohzvmsQsXteAhbqWk5K7/EEBPp5oORzc5CFb+/eZ7ZZW1a3xD
YqyVyL9ftKQ8oMwtHMYFRMVbbPB9b6bj5vsGauEUsvKVGPNZjMpgv52k9hv5lLMFCGxSqjk/ybn/
e5ORI0vz7rtmCZLaPlPAolTgs7rj+xGUn8s1MU55f7uwj7Oh5toWh2teGQiIbbt5CqNz+PuU8Osm
HJgqpPeV78b1p6D5uBnIHaHf0gJeMELUQKE0ABkrZLgp0ULuK7TPz0taKdCKPg9UVxF/yT3KnR8M
OIniyzcNLZG3Be09LuhtvFG7K92S2tFw3pmRFQXaX5MCh9ePQ+bVYna1cV2/kJ2x8ow+FT2ea6/V
hvupeUfgKaXgKws7y6n/rTKLMQnxFD7NApVIbgHw78ZosOMb3lq/SDsFxtY3C+gm2BDYYN/o2qw4
z57vuHAoG+2fTrWiO+dEt5eMsboSM4t88R6DpGNvvjlHC/i7ut/onqiHTQ6dS19gwjiieNFepKSb
BXkuhw638psfU1dYQ6DyFzxxO/pMQsf0W+wZ0Cz1JhrRzmjW/A9NO31PyqDKhE27l9zxdKNkxvmq
czHkN8OCMBzo+ZnIxH8dBWXjg0uqlILXPV5shj4g3f8QXp1uNRw5lKYabvQTZ3Z7jwB3nbNPsk/y
WKam0lbrfpQu8tRQpCXe4NflVa77Q4eqyHr6eBeep4eAeuc8nBHnVeJbmWkpz9+H9XunvTd6Y94o
/eLh0YdzooYHuO/EH5yE6bS03HhqkYrW3xIWZmgMWl1PZMrQTvzO7aeJ6EP8opc50OOVP0gwax6I
zHfMcVPcWDreMVP3fdYe7lkzCKpHupHKvKVJRl1JuDi5ruTy5NOClzXcRXG4rwuMWmGUOg4ECDwb
+mP3VXOJolv5NKDFrsKx1H2JgCyPKNt7sfru9Xf/Yb1NpX30qXwp5rAwXZK0Q9dfJQcW6APk5QgL
poQI8Xiti/GrsSz+IhYevak+yQ5WyP3mYXM74oO3DfraN5lOgikdkvZpKdWJzMsZhecIrbpc4JR2
5krlwDTGjwvLOX1ZMa+rjIkhbLvG9EhnOp0nRpdFkovnntUIXb3t5AV0cR5VIM8e9KSQ2q3fg8Ii
9mT+yCD00UTiLwoFvr305qKGkluH99r8PxMwS9QAoJun9RvB6w2nO2IwPblGu1JOJ+9aYgeYM7eD
S2ivEMdPi1oiTlGORyDRkV+YMjUE4kcM1jwlZvReWGrQeIBABcAyTsGmG6WvBl+7Xp3rWXG3RqjG
Qn1GNWG2UZ6xBgGOuX0s17+PpKzucEwo3P4O7YfiINnRFrSdQrmqoa15p8wRJFdRwGJAbikclSBZ
NonmflXPPqp/wpr17+vdFMxe9xIv9M9vkwLH7s5QHgC05mmHt8YOWiyZ7oPxr/pWY1zYnJ8GxqUo
HLgR8bFCJcfsl0IxBItW6NxQM9YQLfg1nhMDGH2Fmvjf+cGGEyATPAtZu4Gdlb7lxX5CVaXB9xT8
sS5H71aUiiDcEFYyBPsAQ2TV8vzK2uLf9CvU90Fl/s8IEgVldZrGV1PSdEFC4uF+lkdpDtcahbvl
Pdo+VdgHYUTfvxBQdKt2O8A6ivwmnt9Dh2CO45qS+Ry+yLEHPGqIJ2PfEZ1HbU0WFTy8taC/kBhQ
h8URW0BN+AQ+O5ZGXUd+IiL5t4ZTiCllZbVSWeSKJUVZHliU2hf4TLPIqtAtOtm3iJcgxH2+sScu
gQztPuNm7eQLd+Kzv8Ej86+Z8Z//SLqd7Xx9abOVD06PsoHbrsP6sGzIWMuVMmqbVZMAD2opq9UL
Fp8zaIE+MZDzm4wy6VcMYge8SZSMUrrox8m7qrZ5n9R9uE6Rg5z1NW7A0KTMEDHYP42u3QXLCnSF
NKXGfvbwAt4xGiUWv7OwzEKC8Nw5XqN5Z0jTkjIlhCKLs8jePSSwila9wrQl3TqBEbSci16R+pYx
uk1GU8yUqOwNZ1ehUqT0gRJAIjuf2GMaPNcFSwDWEp5bEWtBvgm4+CVspJaXD/EKfKGsfcqcNq/a
NdYimcKoy+GS8OKaOQkQboIbNWUNALciYM/lM4mQoa40kSWRwPIftUT6000+/M8vLlOzkcrk8A16
AF1kedj9H/UJhcoWzPRJtICuK4ItBV3kB5CQ6aFkUzmh96DOujSYyipY9K41K6jp4ewv5s9qVD0N
uvj6KqqfP0j7xXh8Hs0IOzaANpg1IsgnEbZ3kQ3TTZbSfO3S+elYMLnMHLKCSAL3C/C1RYhLkHke
9ACn0SsZoMa6u56r4NeEwbD4DmMQnQfNGBZsEgpht75FE2mIasprFsQcada1xbaB+8pUIX8gmSDl
pANyKMWiHsbnHdwJYXtGTz0q6nUfQDmrdjErdpjSWok+VY+a/4tHFygxB2PZbajcAxxseZLmh7mM
M/pnuYzZXHWZrXLKRVZY89o5H+LU+oPUphF90dnBAfXNr5N4Rd9JR5dFMQ0SaW69PVBlcV+7RKcP
YlCd4PYL0T26XwHiUguT6l3qi2F4aRZiFlyzFxNo5yMyClo9iPxyQbKUaTicYvawNiChUtvnWQms
lAmKyJfDmf0GQE9TMhzKnB3MuB8DFpeHYvOX2IjwEKJKb0C6/VyCiP5opjaVyWo7viAYHUXgg1uT
0IdibPcmF28DOj8E5TVyxTIYDCulvK9LQ1gVWLmTdaMG/CqQOIsq71Ds0YPg/Po/WhMONSUPIUPU
WAgng1z2ppYeJX6FhGuyRHxmwqgnT9rb7XwyVd3Sc7cek/ZjhVTPaYxEZfdYEWIJ57j8ertNTi2A
2ff5tVN02z9aihHcp1R7o+9dVfpHFsWarzja0TfZXBNe8JiiGkXyfvLC5HrNnud5d3NeMh41SIg4
AcWG0a2ixFqJRTa3gJipL3reAlKQid7uKk/JQqatgxYCV9WflbZ+9E+O8W00pHFcrAgxJTEuz2QL
s3Q9o1kLgjlKWU1lWo8xLl6oW4X3xmWu5hxG0e5we3wpgXhWnYwPLEbQyPMcDfMUiQBNJwKoqQzH
9iq5pC0xp/jfSm+gco4mF5hC0fPvVRyvI9BfFClSCDlEbwHekbOQ7Xnd7kuwMNeoWYqplvhcdxlB
n8UjOXTHsLrpzsSVaupTP5vJbqooGXIkgCNvT7TUj2aIJHfLVYqohFClgatlYa7vG+WAkLIfnXFS
9P2TSGgBq++UQm0hdXZTFwIV0PVYb49zTuRk+20txiFz9H0lCczG5Gqj7Z8LL68r/4Yf5H4j237d
FORI9Qb67hrCrmY97kLsfaolf4luijczMworocP6EAohRm6qVa8y9K5Yk/7MlHdcozoJ5xX5nOLa
h5NmcCfwVbqGa5YfCxIABNzjI3ON3R4LDFcYSZv2C8HJ6LQs942Dh7TlA4TvHdbv83UqRNL9LM8p
VUM7w3xbkMsbsyrPYsSSOL+kcaW67thFWSTKuP29aOUEMskh6ym5RM3r3o8SpOFCPyjfWtE92Yii
EcM846zAMeh2JTxmfBrhRbsKwj4/soXi7b6/ZxmgGRDh0wXEn/bxcS8tX4BXN4m37+ACNxpEWar0
dK28OO4LjZjt+dXeAXkgVTPojp0TNG4fjwdL0P6b0rfSF04n10Cz5JxP7XqmQaLQXRDAHvJYG2p+
jaRxCN4YNaUdh+ZK88bVMNPwHOznZoaliCUmLsAjhAX65BwXKl16AvxPc8GnHdXdqT0LRhm3S64S
3aSsxuV0fnbABH4ZII+7nw2OaAG0KMzwAwW5FwX6sXGII8F6pomC0vTbHDXl9Txt1yIFPWZ/SUzU
fyxyD8QPU8acYDzhypi983cA22hoL96F+bftIWSdBvoQN4szev8n9pWZa5EW7WwW5v0XesbKy7SA
0kEo4xj0643mOH2CbPtGN8voylA5+KFAXhYQ05slck8AP2rXHs8ZCM0qBtPstrdAawZ3Ebtos1bd
VwmhmksxyQ6LITHTmq2uYDPjIK7i7yLl4TOi4m5ls3vFhNj8zEm4RuN0LskgG5MELWCHFRioTbC8
2IbPoeVeI58LMHd1WR3jeDwSVE8ApVNvY3Jco7kIkVWZzEUkf2HApO2UREubtYCmDt2Nz2lmKy69
U863Z3TDe0mFiKL07mMuZhfCxHLvTug9MGiqPvFa/z+Rk7MkKRTymmzFtsQ0j5JCf6sCdrsdk0nW
KUDFuywqzJUrtcwjc37Oh+BuZoAfzJt3Y5kDO7KEfq0tYYVP4W5oPVqogwhJetOrCzNBLHvM9AVN
tPS79Q0RWiC6I4Bb067ggU32VT2xzqnATdpT5AmHBck60PKJOTQ8ZkrhJDyl/5YrhAz1jMAB5TTR
0Fclq7SroVflTZpbRA7T4wb/ZZbSEPcLu7dC2r8KQsisBMkLhHA3oQr46ESW+l9OuDKIdLjiEjbM
DCK7tFa2dc0uoAblAYEuV6fVTnw6JvifLGUEHAaARJaacqSI7dNFjlruoWrSJ3cTTzYo/IK8Zo8L
RRQPZJghsAdRr8dgIoMN+A/g5LAJJm+rAN/ss8Vq5rMMOE4u1tz+XbfBFTEjJzFbTvfdgkYX6ZGO
iqqlwtCuOvnh9ulW0uRYukZHAofUMrZfv+DnVnYcm7gwpNeRbtDkJjV4LWonBXxhQUplN5avf+j1
cfXDwR6EavAnRzYruk1BHMBxTKKk1B6frh6vLuvy6nnEbY/t6tFkJ/Gep5X5t61Z2smESXQX8mdb
lBYVkIANQMTfZ6Wy94Sv+v50eVGcvf+nt9C3Ck9QiW0yncqRQx/PxKOIG2Egk3UrqUjOMy+TZWFE
l4U4rdA9TK+D+0MqXb4VtHlyCWhih7Xmq+aooEaD8SKSfoc7ulnvtm3iE+NqDWavN1tStm2tCvLZ
OgM0AUyDPB5AbB7Cgpw4MUx0UAyE3lC+uSNyst0pPGHhX80Npw4RGPYbMepz3HBZBUNbZdiHmRHy
JzO2wdyLmG0QHskjEkT2Gtb0d1CkPCql6+uRLBZ4FhuYhRl0JCcTx+zhsLa7E4p7pspFLUjavK5v
d3OMYn97dgfCMjwdgrPEKLs7vY+nUSlNF37oYzlpjkfPkZ4XU35UbL2HKlQDwt+N9Yfs8KoOW08R
Q2ivj/5IDJMqxY87wH9SCGKlNy5dRx2LaBrF0w4dXCjQIpkVoTj8EmM1mswVeScDbRe/PMEd+HG/
Xl57aGLLrnlPURg7FLqUkUPCMtID4PNXBBR8NYTPfkGwWrI6acYrd+flCLsvyZmSyL6TAYB5bfTw
OctEpI7sE0Jpx8OA+XOtZwNF6ZZnZiRf5XfeqdICT5N4rx/ErTV/32jB4Obnjzn/XczGpk+/YyMM
86ePWEKet6DoF/1St4z6xYaC8A4XstBUub+p8pEMFVtRD9qioxflwXH54g57hnmE6hmO0usqOTPM
KibeKdacZ1rusTN5dp7DCJcQLsm9VFnLFo51e4Ou5xMbhmwlSGmVm5K1mEXegc5bq9zPF6pS78de
7Am+wq9NCaq3q4xqJKNzXMRk2mpij04ze5TVTNP567RQjjDBvBQ32YG9wVxQoANy+iCfqSC1tI5f
cFuKPowY+x6mH1uY8XYOBhDpuih0D3wddiXQaNPBIxLs7VkOV2BwxPuXHhHeZLKZR+ISwm7rsBpJ
bSVN3GsHohMpxkZT5rE8AocxoNVSH7ijRbniGY/R77oiGFjyBm7SwPY5HcNoItdEN7UQK3JZuQ7L
Skz5us1mxJP05DmcANxOD0RP6rOn22pYDihlufMgfFV5mOgvUXonsqR/OGDbPH7laGbCW89zZ7kX
uWxSiFFuPkfPG60fSramiel9wuffeYfrjdnY0yvncjyfhlX8N+lzIyApEDcAY/BMlMC5bKD7J5ay
fZxWAPsJhp0kNxsPoaxkd/elI7B9oymd8syafPcZsFzNfdDBE8u6FXGjDtHhcbS6AhswiYZDC4T7
TDxnZlZVSxTRBG/rO2CYdZDCXxjiDhQXEy1H+diCcdOqM7KGrUgsb6lGXyw2VcjANWloo0b+JCM/
aYycTck1UhwQH44+w7iMPQW09Lp+bCzWAI75Xuqhm40BgwISiVfGCmLe+lkdirnvLvGcBOwDTFHs
/hsRfEOJEBEcejCWEqlFZJAt6q/gGs788RO+I4mZPpSJ84wVd2Kks+lFkF9jqTN8CMKSUX7iYos2
goqd4cnjKtRf+sC0K4R/NbFaC//RsrT0UxB9Riramem949dvCMzzIKPkJkjfPJCS0O0QTw394meP
89L/a5HLOG4eqkQyNYpnHBgZf9CKrq8+qw4Grh/ojWnOAhEexvvFeIwKhVsTYEVtrayrO5WqrG6X
AH7sg0gCeVQ1bybcFDIU6YBbMB4+fcZD089PLXdg+gRQG7LS/HDx/VqA+IiaCdOsUrkk681ud4Y3
4DDP4KiKyVKtD8xTJeE1GetlZShWMpjtkmv91W7mHFPEJyc3v9kHWCrGE3OxezyWGgVr/yjCTUpm
t2YXu0SVmp18C6GMleeYqaT+YJ5hQUxio4s+XyPVtNQ6RE5++Z53dAse2LfXouAlARjxI2rQbSVr
o4mWeBxYj59SBnCkAQoAZkWLM0zP9FG1XIRxViyOnTxyEpVjIDuAPjIjhVIdh4xYCXGN9wR5/cBZ
78rf//VvAjfzn++3+mV0thdJ2TawMeS3RZMHZQOdomXts6QSb+dR2t2hAVTvaGFF0yJ1SIq3PcoZ
s1IgUbBkJjaWMwKSY0qp27BIvIDdlCK9G86dDcnoo/QF5PnjJAbm5YCxvHFldt4AGRdzDt0iMX2G
UydFc13Qe7+AbTXuNeqWjSWOPzcVs4xpY0lhVtvAjgO9Tr1YRreCMp2fPbs94HQJ5Z6t2y1C//kp
g6HVEtdtYJROFscjWSSeYRzLivawf+reVMK8nwBij7UrFHq1hu7aljTsS3ZNhf9TZ4RHRSgi4HIp
ZgKjhZpRCEQc/995/Hwd5S8hYUK2ay0spDM7o6OEytZOW8Ka5DERby4eajig8Q3jgI3V4JMPTNvu
VGgelG83t2CNMpBG/9gBuffj/evsSMg9vBw2l6ZZQI6n/15O6OrN5xRWW4CWKQsmXns23sKF6Gsj
X1AuxnIjiiqA1kdQ/b69MsHE9/QRAefd9wDqiNl8WV81oQ10/9rt6XcVt+qg0gaLNO9vS5mde7v+
pcSeMWEYdwWc7sQ/yMA2YZOkmjtGWp2SjedwyqpikelIw78661EkjNCq5TIlgPvHnLp5CuDj587+
82EQeAb9ccuKcGh98GNLx5BHYRzXiwjsoPk6N2a5I0oCRoW5RILq8kb/sEtXfW0bLM1twlQ6C5/k
UCicb98ASPVAM9HvJRB2owUh45kUlnFBWZ1hgWv7BijniDAotMOb8d2CJa+LPGBUUt+9LjCY+OnZ
f0POUyni6sQ0+gHlBVgmaxME7PoQx7+auN7joKBTpKFwPjykXRTorcwTUGesV9lLUAJ3/JfS+5v8
Pl4VrYz1b/zhtrTkYb9qgU84qoAc4E9/XZXNSjX31BWSf+m+Ob7K+Gy+d7/1zb8+6vFYN6DxCs88
tVoUzyz7TcY3uHWNDU8NfDLiCqVnCe5u1ZMSagLqiyLr1o6bX+d2JKtPydIS+Q+FYDQ1oXovvJJ8
kEDM0XZkqDvDBGJ/+PLbug/8sybYkSk8EHDWrZngNl3mQPTB+J9f9avm8OzunHLrZOMkXtX6VWep
T9jAVLY3dUYcg6Jyy76EMSb2Cp2bKLnnGOzyvxYzbtAPN4n/V/QryIiXcqHV2/vKG2wD0pSHYPkv
0qjt67vZ+4aRWv+rCqk3XFYV6t2lHz0oqm2NPXkRG5b9h7snNde1gt/blxfpeCcORpy4znfQW9/T
F7sHLiOokNbRkOimfty2xIVgQOUM6rkcF6PnW6kn2V6YThEaBxHW+TZPRxysWqzIZ3xhvpjEhsQp
s9YoHF4U7fLq8XSaX/7xjbQquWXFyuvYV4vZaABupPkfqmW1AKGRdmuKTT+KrSS3j4s6wD2doHgy
Fbq7v53ZpzmHDWZFawmf2wKH4/e6Sl641Gn4608g9a15HeYkL0hu9MEEKRsS3EuDDxw4TiDCLaW+
AYkIc+p3yVTnfvLd9aNIP+0luq3jZZHCP5+9uw+Qnawb+dvmzlDh/1gtM52qqc5DCzQlEdEE3/zA
4XPqeXEschYDrZf0509nE7LqlJADYB+qi4jYbliQ0M7NUQSVA0Bvg9o01980dMw30OF8gHFU5dEa
zuF7cFz+JWb18pB9wlH/F/F7/K37ZFu1Yl6o+5Vs1Oog9jZRz5UpkmZmNJbwoPDUi4cg1yLYvh/g
SHA/D/dmWbMLsK1WyBI5M52OqA5QOoDuZGpxpxui7xReHq3yFqeTRxDESTS2BQJj2UValLOStPIX
zaBJOFNk7jynJXkFz85zTWuONh5AY4zbKykz7SrFp/xV3XboZhspkLXuXUhP/IqrupVkkWcTyKKW
Rjmhg7IHdog+86G6AIxWfSAD1o2Wm/wWKAjd2H/mDl94J8ghJkSBJXUjkaQwegIAJ1RHXD15BYbp
/k+mfP3iw/OvX0+6uNddDBSf+pItfX2e06K5M7dhCTcbyMB6pdJMP+xT0hvlp5G9+sU+gfRTYAXZ
g4TNuzacJMCeMWN8XyNzD9sJi8onA4oUgccD9vOEw+pYJ5wK+QrIDmOl0Mofhob1sMY57LJqJ2Lu
qXf81iOnWEU2hV5n/XMZe9/OU6dX4GHchizlON1Dp3jzE8o+aqtnxyCiBW0j9gfP1svjQYYofzKz
sM/ORYiIkWpbz9+dihUkS1Zn4dWNDT9ZgPHDZuHyKQwEoSGtBZKo1V8c6xHe9vUxMU2xDs7zDwy+
Mosfc4GdDdoO/32WvuS5MbeR5ugCa0zFqflYkqlFcIZ0ndLNINx/XeWSTayubPTCSmW984D9DjRK
Anb2ft82XowtmtnBzP2YrLVO47sZdCjf2dprZEol8vNeDyqDDp3RwWjC0H1gcQIz7L8Sih8OWLZy
jnOWtuPLMxYOJfNVwLLLNTG0/JHVboXfv4FMNcJejPiDocd7/Obt4qzxdMePSgGKb48dLU/fxeJU
9gq0VZ+hHWREAgka93CvmzO4HkN/48BwYhAFp5LTN+dkGJXBP6NlbaoBDliefeSCzS2aj66Kg9TC
rGJ9cuTjiri+O0jTLr+aJTm96lxgwPO5itcXe1I50wjCQlNmV/l6hQuVG2yG8LT4oA/h9QpeMqv4
aSiJAvPEk3/KQ3fDi2KvNbNjZH/BsYTzHilvV+YhLQlH11lRgsk1CcCebaP5y3uvV5pLDbxhge1d
PdsTtOIxVwbyTEh/1vEi41gbeUaJXFpzl143nNLueAY2eYikkLNwu2iQ4vxlgQthMqQ5jrCS25uA
JN/jen319CemaIht5uowQqrFx4FrOD/abZgCdphahtmINuf8X7hgZtiAxyZlC9QwbUgduqUINLgA
LmLaMarLuYQxwsjL1OapI32PcKUpe+WtXhJ1FdI5N2GbVuxYl7nPkc746y50IlOc2YIXcW0mafPk
tp6gFfHmeKR1Le8S0OxLFxhVixA9NSgiOP9A9L+k3q7wBMCp8CoSRZx6NQiwzLZcRwyeN2tZSMyN
4tAXo54BnEcU9L5CmncKB1KfxHiokmUlFv1AHzTIZ1mswLpfVeQOYY9fJLwaHm2domeh1roIZbiy
jMvr58CeyzFb1sGO04T1JNzasuEvsjR1c9M+D2NZ6JYSW4rE24mR6OEKXZH1yvsr/HywQh0BQ5eq
LylKW6ek+jyMTg0pExEh38hdmz1F/k6TCNAudwd6NjyzoErjzHoFmZOnZjX54625ify/zFbLRSHQ
N1P0B2/8d5vcK7B44lzF6KpkN/q35X7EhqVENsJaImzGAKPfPWLmNK7cFFv4H74P4mLYT9Oy6Cwz
NypNWYMOqUotT021dG7KdiOa1OzeYW3ungMppbm/oyNX6Qn4nZZ+FgWN/F23uaU2cqQJQWFpg9fh
6nxV9zXWv0NQrq4ElzJtQ0KvnX2c29M9YodWE+BTq1nSkEwkL5VotlOP821xR5/+ue01nAejj1FS
xd1v9gD1ZMwiZoorVX3VhEgVOFOS0A00CvTmDpTrb34otqLYa6MAQIQnWk8T0SO4kVoFiqqGDVtK
aAtVVPbSf4ifc3I6vAS7+lgVq1HfaVvWAM089ZPtNkXg8QNypxcu5HiQttHKfWG3q7WzQCSHiysH
apsOtlH83+3iwyohtBBMLtD236yTiSgcSah7aflw85S1QzUO/q1FAuofDU78V+vxqDMfWGSIBvMh
UoqbMqUyJ/m+ZomQFRe79wyUJJoT8gzbNd6Rvb3YKXZ/m2JqCUGgE+N78hwJ0jS8FRRyAjeQa8GR
+ZKFP9HDYe/GxH+dLYXR7dhWnLFRYrOH1rfipXYtwhUXGRJXk2wzA/EvZdL+vim0CyGUjMcYQBjg
CsrWTxLoW02FYX9m0SyXNkyvVNEqlGBH/leM58+G7VcA4mZw/YuAPAgbST7EDE/kqxaU5IcqKtvM
+H86yD6ND4gli2ryfkPaV3Srg3dhfhsiKCY2HnG9lqIq065uvu2onbQsORQMYMqXckCIXwV4WBFz
Ur4k/6GxSyG/T4sLlFdHxIKrasZdvgR6UoJuWnk3uDUrahTBVrWB8iIk8EKSOSp60aRJaU1vsETT
G1k2bwE/Mpgtrziyz3dHDzObDE3ExI7R/bE9L5pvOweK5+KcCTenFpLFjC3Hk9mqYwVHRQDjmTfP
RfJ8jZP55p1bYyEYBI4Rj16sldTcq5laxCfhBxESzyqU5s84OKExzpavPmpDEktFSFNEiNsazS6W
b8MfKsuaA80OKcjv2yt2ZZCytXL7m0UvP+F2HrioULuxdSrkhfMhpbfjF2tOq/YVjG2lNR1zKYk/
q5fWk0XJ6O2pbMyhj2+5wNUctJoQg+xTRV+r3Vyu8gF2oM2O+X5f5bKh+iM8/hUyAjxfzWiDA5e7
C296XmasPixC3ApwBu1VcYJdUs5FqP6+q3f28IWWcVWwGX9bgK42ISDC/C63wJS363SbJznooJKY
dRYvn7LEyuWupuuaABIXx/u+/AdZ+sg4n4w+LW1UBeDjzo7IRy8z5wDXTo511Ly7I/6SV6phThTS
e4PDyz0MT+niBVeR5ne0SJB24wMzhcZlYulbZO+zOnV9dtCfUaOYAOo94t149DTRiakELpZa07la
XnZMD8M0xLOxYXUdO8IfizC7I9hl6x31GisTxGkfuH1/7jQ3O1KxA+sLOxOWlhEnFkZS3whoWsnL
f+ix2eHznKC2cgNJqc7r/6fD9xbt6Lp7x5nekHrZpI3Fb/sQHPSZxKDui3FJOpKWS6nK8DSsX4eF
cq1hbejUG4RYO8e4YLzpXPmjX7TyC2BzNeLHVvHKNKvReH3ilmNFe5z3AxBUf+dYaXhvIwJV6PrV
GiLaSyH8i6Y/wf5rf+ARveenW/dIGDUHj1yRa8ZQTZaaIwkNIVV5sEe/zerGPR0jgyvKreKvSKuE
d3ssYWoModRLZksF3eHeQ3TgubJCGj6FvSV3jkzo0lgvW3G1NSPp2iyHawUCZCHQ6nRTEZ217D6L
lGDGuRf9BTwZNWDjE6Xtrp6G1FLYiasvQBEWtC9A0B8+tE/LmA5rm4z9IOLyo5yMEfJIOVjTVKyW
NkX9LW0lMZTbTrix52lQO8Gk+k2j+Hsj9Rsx++MqVq1J+mW5XcUrKlIufMaxLPAYZcFyoy3UqXyp
p/arzhzYod28lhsoYd24ac8TfuKsrHibZuR7n5tU5Bs75dPxP0m/UbpbkhnSfA/0/o1b9xrpch5o
UuojtY/nRpd4yPqfP21fvRDWm6yZVN1+ysTUGmJmoE5CctpYpboWCK6KQI0zIM+R1PKQqAzYelw5
vzS8oj1ohHvid8mmZFCeQt0xHlZAxVw07DfuVN8xSjPET9fTIz46yfDFo9m+FG09o9f+vZ+b99u4
1o/XN5B+TvgGA0yjjd/y1t2c+cMq2aMRFks3eC5fiTxJ+Ild+XeXYvdTInVCgl5L3iA5BhH768YD
ZyvuxNZshj1TBvsBFsnTu9fGCrxJ0niBP4osiRYCevdiERamwZFAV/1bWwbuWgWUhFhQVLUuFDVR
L7qeWruboDBlxMksOhJ/xGeR/5dKN8MU5EC+WCAqLgBjakyLZK1EHJ4wHcFhDQ/lEznHGwmmRJjK
SFL84Lqkv40bbljSHKSfwdUm8uRiDsnB1T8eEog/7ZSeHYM7yV/daPvJrVPZX+NYe4J01UUaA3cm
2yuuFiSp4ln2gToajn3/nDIuO65Kjo6OVeTTUVgIinSEtyVLmZRJyKedHvSOe430JEUJfQHKp7KJ
LXxAefPzJp0jnLGpzL0sIaw9xnMXPcdsIgMxmyBq2eS9GtYDEYYzSTC8IdlsC9P6NclwKSInerd/
o9fa0B6e8d0y7trDhKoe6yZHJD0wfEE59Nc7UsfgHQFK9odrjWWq2Vw1uB3m5qekjWMOI72x7eNX
IemA7Bfu/wopLPHUSWaiAAkwBeX1Mf7VmHjlYKIeFX28TE1q9pjHWcxbQW9KnnQ89ZnqOvS6DWee
qQyNBvwy83me4OBRmzOLt7b30uILpT2SJnTmJBPNlnMSWjm8S7qHF7t3rjgmp6cQXp/Jl37/ojbW
fClTeWSXFdxIzCgquAsP4D6V5JMUQzB/GzVibOG8ppUfy3A4qMe+4G/TsrYIvCAFWruOthIKb+jf
MGq4vStCXSGCaRp9LzhWA3EByLp7Hj75xWzZBhLH1mUIqmLdWmlNDFVR8Fyx/L9cRzq06TI+n95O
QX/iVIO6inXFAQ0GnLZY0ZTW8kDrcRtK22wdg8HWaNS+pHfyXnQ090Ey3TDttsxGr+yVSeExcYW7
bkawWd8G6DYFEyXV3w6viJH60srevGgO/NsVr2PiXpirrCILokNjzOGSmKECO0fv1H+uQI1szMTh
dcfLuCstFvfKD9Eh0IZCZsPjQ2Z8QH9Wx4oK3cOg6O2AM0HMzZST1EbETKaS9yLDWQooXHZv/kUO
OM+CWxEYADhOkurXBiTaw26HGXdyeYG8A79Lx/vCuNmwegVDqH1suY0ue3W4I7iLE2HwXxU4tT7L
KJ3Wq5hTcbuk9BUT4T3CKuC1CiKGjgVP8qlhxzOWJhRskTmKAoQBTEikU6GrVQ9aBylCzJ/qehyl
YXJEKMkav5FW2viqx7bVqIWkJmiZsuJc3E8Bx/DruIbE35kygaz1e77EjGBzjR8NhoNcfFN9OqLi
TBCiLLGHTKOfzLWLW1x2SfG6NvhxMboW0yLCIReXn2jroo6bFdXSKo739jv++crP5QFV1DlyrBet
PQgb9ZQ7XQVQwULnlf4h6a5nR33srVhiq8oqAOMFGj9I/rWILM4oprfuasnfw7X615sFq95N13do
uu/ai0DSpl9PoUfQWIvUSCIW1lCvJ3+4lTgq7KRPgOBN4HTLZraqVh/CI+Tpm/8iPS7H+FEqkUP+
XqrqR9RgJPQW8TfZqCddm19+JBZMNcJa8dn4JiYOSDtB/NGjpsTfWXzKl3J/fR9/7Q78noWhVJix
jBOQCCjH6R3XN7S1Pp3gIhbHDRF8X9Nf2Bt/g99LfI/a/uTkk87G5yJqjZSEeTN8NX4TQvYsTl0t
98sT1bOnBTIW+63EfXTJ/Xi/rnu7rIDQsHLhy9f+zHAMpWP+PWp2TS67plOPKo/znF6ZYXPDc0dp
gMrGpkMjcgCoVqDXWZBxWcWrDK15JK0c5SYWJVc9ZUO+RUqFgKDPguBS3GhFdJI5LlppcF78JMqW
Zyo9nGEeh7DeeDrC4n+ep0vGjGMGZUSH9tN42FksvNCNOp/BZv2Nb6T7rpjIvPdL9usLsHXPIiCz
txN6zrMk/HCfenxmCrSDa1UdP5uG8oK0wbJBLT9KxGegcfrYZat4NLYxfqatTNmLcBrdhKMj/ry2
keXmqRyoHqKmQopsIa8haC/ypzyJjf9r12b6WR3B2dSFXETcaGGh9lqGChT6ztXa8qmIWr1CKrZB
PnPc+unl6ovIJMLmn5MfZKkOhVd73aI3ZsuJpQw/D0RBxZRQtsiLL7OlqpX9xEh1DuaYQyfsao3W
quFzoIln3LOf5UM0eadSzqVOAF4gFBtQJtD+YrnEcmu+4Bc1NCSGgFOZAVa+/U9YjvFaT9TvsQY5
6VATKu4Tvbmp9txBdzEJtaKUA5oE8/iD1UoOjdRuZSEpmNDWJxW5ofHq6qQ8aTw8UHKKCAewFCib
mFpLDy6lh4N+rl0aGkBX32TEaNvciDXr2/DZPox5iNgY3WIlb+ZH4mVT5RlvW2nEWMlpW72Zks/3
L5Z1yNn8sJ+HJKsALRLewDpIaRcED/rHWz9nDPO1BJ9FErOV4Blo57uC3pATcNGygZXuwbjCEUHO
NQHkbICODNPanFtDthYrtJHUv0TldyRfse98AmWoPxI0bReUtM70dj3LzHMhLtJRimqWcVVkjAs4
73UEIzJOM0F7hor9tSaNkHoqr3jScBBmWBfK14Qde4uzPPQACWW3iwiln4ljQ6W2zpXh11K1i8t4
VTN9PuFjS4Dh+PbeMryZyFyRWLcL/JwXwuA17qidunNjXQpiRuFX7DskBgVVpqCFwJEu1+l5yWCs
KidquaR9rX4+2gCHz9Me3CzYrUjp0E9jQRwGpQjYrnK9j3Uo2tNPgr6bdmsPEJdiCOv/cfQ5BAYB
N9VXZahy5B0st28ebbdE55KEBeal6qsSGfNxQUsGNkjKp6IHRnMTSSWbr2Ga7dKndls4+sja2J8c
vA8WnUlYCaqMSBHlgigebhgEipQ4p1WlWuKtMv9rumjfrDa/MtZa3bV0dQGl6ODN0h1x83pCCtOC
WIbFO15Xd4lwmK0nF9zPPtfSnZQNhflcDHzXVZND0bTyUIZlPk6tNJLHIr+JPoY2WmGUA8an6/ks
keLOSCVyjrfzC+HF4AEtce/KwrtD5AJEoDiRVMFSHbMYfJu/sri9WUUmSDm/zTpKQO3rB98gDmrc
i+UfW2NzC9JwWAA92lPTdANgEzMDuenzOIAdLv+7TgKEyTIFo3+PwgSl3VmUi2V8si1epHIHkGCP
HCt+NvaG2ZO1Qm2WSg3G/V1BLYQau2q6Meq41r5ZHme/OgvnmVdwoGfvOXoyCax/jYo9+ETSJelu
9PKWdmfkp+/I0rGoneeCU4M5qAY5NUDjxtQHnIpTV4P5TeL+5UfgUYMl9IYtDUIrnAxNPFbpdd99
vf6nnmfuvdDBi8pbzkbUsx643xUdh0CVHrNX3dCzXvdkXJ44773pifSAVY3a1UVDk6qpklV4P6C4
60/KGHZZ3ZraRtrzd1szOgYKN94vqe1gDseOxT3vFd7smVHhGeBvG9o0TLUae2oamqk2fND+/bXO
B9S3teXBSe4u4+tD4ivjrBeDEMOSveoZhhF6YCw36bMynhq6jszuA6wtjoui3OnqhWS2BhY+d29o
sccnEqlOY9LcXPVHJHlSYP9iCo+kq2JhSKwzd8gld7N32kzQPzF8f+DI+hoimYDWUmnTQgwwNOQY
90wUNEEgXgN3MwX+bAX6fhM5iFYxwnz6XmPy0/U5mepderUyS2JvyjNjgHsdHMBr/3uVutdDrTI3
Z3WgaJaGfCWsnACTMVaDKlzYtC3XfIhUqtjNaYvnJw9PpGBN9BG7oDarLP90c82y9/Ii45JuGMU3
WQN1rnuNsnkjIZPIwmorvjCg/I96lwqftxs9A16is0HwemYUQJoMGeeK1DWOscsr9/eFRe5tOJbA
NXD6zGfPHL2cvhAQPshp1JYe3qaTohicn8kAbexBwnkgjwwgogXlvlPCL+aWaCVtEHUtGzabym4s
0maLQNiL9qFWgKKl+Rx+P+UwYY7okUzHY96pwjrNtg6t3PfWiC+xwyw2DYwaTjnGMbYQkekPrf2b
xZ0N7XVQyKoZ1VBUyYDioCbnp5y0LQWrzs8Rw8WtKCZWujdOOqOeL5r3JNsoCTaX3VGWbkcEbnLl
gebbvArCT8FtXKu1gZOIvkuLnMDA66QqpHjZZB95bs3nnNSv9vAAXiV8CNFKpf7BbmFPakLlNpK3
mJv/Lu8jlsE5eQWpN8cjJTkYqMdKE39gxI99jwlbwGZrxKlwMDPwIsMgrAi1Ma6xm49WLt/t5NmC
8tDWMvi0uUbwxWrnBQBLfbUfZ1f/nbdDzlFnd+fXsz9n+U7mimsJHrmuSeobP/l8OdO4kwk5MCgc
s+sHKGOfJ2rFvgsO5yO1ZrRG0e1BcXJ0+LbViOhurbIPTLFjHD2mZGXFpgm5DSlqGEeGyPGsDg4x
ntExnU6nSw3VQyweKpinpRvA+INYnOOobAPGjgTMRyj4oJIj0YLO5kVJaa1YXcgMzunw+DP5pA8i
bmunpma3WTybOeiwhF6f26qyOUionhUwCHfG/5PzHhVaCUNanSrPRnJoxQd+tRfKVknXl/Wu6ybC
cRPAc8IBQ/N+XJTkMKwvx+CcKxA2SbAcTwTjwSAi+dZ+JzIs5VonVd36n7UDqsOfbraVYeKACk5M
gkgKfeQpa4A0unFddqgTbnDNY8nja9vSWkoI5jS2W5ufDUie99IMYImCuPZtI7dVyrnZUb/D0O6j
HLg2QcpgTFXh1aPWLE1nTdowPfNz9RZB5RKufsU38X5cRN0wuddzoa8Ljn/s/L4vGxpWXQUoEc0h
C3rvjdfSo9yKw1vVPL5bQUJQ/AR56BMo6qIzeh31vUVdkssQPRFMBrpLiWAKBsFfW1fSCkhLrNAE
/sEufuZrgnxZA4Af7LzzADP1U83/jMsVMXhAsMbbH+otFc4xrWJ3HcTN0rP4Q3YYt9i/Y0PUdctn
iabTclF5kNUjh08SXrvVlT4G++A6O5Wy+MsmpEoWTYPqldNyZH8qQEFO7ZT+D96z3zDGsP9NbXkX
yW6rquNCLg70TVZy0uK058TFSfvR0PZ6dh+g1KXmZg6xu0i6V9bCeQBNMESwpuFicFZRubQ7pEA7
nAMwN634O5ViyfMwALnjHj/mtmFfiL61XDVEArQlOJEstu2dwe833fzrrZu8D4IMplOOk/BPU+Tp
wivHw81KN06AgyiK7i0iA+WEfHzuJdyrac1Mp4x6hVh3mPQfHm5aSuwDRwyX+m+lFIJsnKa5puab
POTt5/tzYVHAqDu5QLe00T4XOrop0zTvFFeTB/yoXLrnDzo8HJTglkEwWw2KP1dG6r+eJZa9q4oi
oGa+Aw52fnrotT2Sa/jmV7AkKKu/JgebZal/jR1R+ylI78/RVe7tgQmBrbGGSpZQG3O2IPC2UeMl
86RiyvKJy/QrGdGfddCqjNOhOH5tj0tgRQb+YX7LkisRdr0eiuNw1AhLxMgt+6JxldEm9f22KBG2
ig/ZwcFmMiPvHClpRHOet+GAS+xfSx5m9Ruh8EtQfwveKXrFh8qYaXO4ZHQ1U/VUzc+ZhMrZXrTp
bj/21NPJYW8ya+YRciPRfiW0QkQJuDhbm/6B2HyjBEJULgDpTs2UTYaCST+VXjGSDPtJDKqvegYp
gXbggdueUYrkL36uNwBuuQCkvBI+G8NU8umasAJdmyKj4b7AidOJ5O76Zs4ehtBzt0SUrwKC4Ahf
Sw0yBrLoVSNecbuTY9UnHhbkYfjjsZbNVJL3MEXOH+M/eTqpB73bXURJVkp3eqt+E5XdoRJMy447
5YpYxqXDeGQYhSkAcy5vPS+0Y0vziQu+zIv6QaAq5aW0vPKBqKG6QJea4uf/xzII3u9W1zZ/bLrv
CFHhVqb5eEKZDoNx6Hm/Qgef6a9SZW5jltWTr8EO9MyyRChamYdZ8B61XfPvtYshXq7zHRddZTpC
g+BHzdQRcTycjMfrM0Gv1AEV7KyCMhaYIQjOED8SvS6JXyFSFH3JaEHEVSu7a9RarEPFoXrzeieD
Bn7xeATGASAaiaXiE2EWlXV7c3EPBZCsRN52rPIKsAfmwP7Vn/zlo1x340/RlzmBRK/m4P9MVhdf
TnQIHr69Eu4bpqaqr5nrBONrxeIGtwvXRIDQ/AlYDQZ4g/KLVpfJvkWdQN1ECkZCiq9H1LPI2R83
8SL2UYGkAFvR1wsJTaub/dGBoXFGTFajBuYRk4MA5LFIjlcjGF44pem99Ap7H0/PhDGKkb4lt3fS
MkJkTdIekoIRhoAv346lWkTyesHkjY/yxqYHLlKfVsZSaYoiSSWikWKz+CVmQa4la7viD+mlRxsx
orUfMwLgt0PNGyQndrH83OAVaL9BXlufKXuA0rzvqPy1l5ftlQUP2EgT7S5CxftN+79tMFt1wZUM
wpGaz5upJzo3DPqsw6/DhOTEFnfVvXcK0pmvnI9mbzg1zdy6h7zuhSFyZAwPHkwxq4aKLgEjIsS8
r/Ik3POnGSlQUxYmKg4XgFEDQvV1x4PEHNESZWBQ6d2awn8c9aOE9UQimpwS9apkyC6Kv4Q3c6Ac
5lQzQKEckunDsICkDg3aLC/qViLwKPz0MVCORqMEUMhwaFqY1tMoC5RIodoS9r5OSi/euA7P5VhQ
wRqWWuzflBGLqiC7xFW/2ImChacOFYDbp6E2jhG/wGCsMryZxH0VG+2LVxSXe1j9VQ+FbO0yp9kY
5LVrqeLisHMqaCQhEXQVU4EzUgI1Jgb0v8M7SPjD64p61SYSXaKZ/SDZZbj/zb+2yW7tKL09sbn/
FRcbSnth+i6KdG+IP7kEPujba19ER/gpREhBKxG33iTj4qlMhPXFtsSj3qiA6kBbMwzcHurBUsbd
xGO1ImOo4XVj9BDMCvK3KxsJNaIqQN/bsAAVJIfoanbB9tqdPZoqQ5v2gDWI/y29DbQhARpN3zsx
MxQUyh3taYVVwjaNl1LnQd3uL5FdrNk5W3/0kQLgU9VfkkCFeq9g5Ap/cgn2CoiUULjxzAd4P3Vv
kpQSBOw4QNpMCWrKwLrBDHjpxDN/F94q7WrUi3ugox0Mzt38So9TJawSglEELGqTRNd3ksFqo8Po
G40qytjYkaJknZkc8E8CzgAHUtfmu4ndx9luEASzcsJaO09Q6fqi+lpU+bHdVNHoUmhC5huMAu1G
Dpg504bKa5cDiUIkguMv78xst/Rus8HL7SyUGFY8zhA8HIZ6jQyOYxdIQBYSvJ6e7EbVIzr/lGWo
Arc3R6sUq8CEezh4csSrpIX4gZ27Qvndb6ASyy2M8JLToCyn/dBHPm3xSIqZe8h0qdf+ae31r2sn
AVg9xC7bSperAbE8nsy085lo7NrEBodC88HaJ69luuXV3PIcoa/zaEHxIWJs8dC2t7kXbmCQ3bFl
A5oIfDHqan1PWISWmQrZ+XbUeR/nXe2jBYVpUkj3jd9yVIwmtCsnpJZHrNazhQh5gyY3FQPagKh+
EHJDtZ46Wza9uHDXsAyeVmaHTKCPMbdkcaNH4gPwJgYFQcYVPZ11xtFpXxycyd6XL1I8uoxHoZge
VZSCUy6biVxNowb2KrBE2HveCVru1rPNTNu9bpn2etkswAlGRQYFkXAc4A4UvocdcRILftQRVhc1
qeDEWc80txeI3/XHLqi3KromygUQPOR7B0b0gH+D6DSipcsX8DXBJjs/k9v7PnYfzHAF7MgsxcGR
KKUM9WSUX62HWPFmoEsHVE0iaV3vfThIpfDX4ltQmNt1l4I3Q9oHZE3xrkzlXxn3WkUK9UctP6Rz
M8axzsZ/quSoi2mlQs9KpvNOAKvaLylJG1Hd9aDvlc02mY6jDMvlEN/XUk630uHeOvO+WgTBkkpx
BIQN1VgG0MUHLOt73/EuvBPk4UP2WvJcUACANW4MnNWRb2lQvkLwU5VzBz4viRHj4YxeyW7NbshR
EPK3D67ml4eH1BgZ+JE7WiXmvLAgkxF26g0E+jgcatF4ppmSsq2sx+xl7D1Tw8DaW42Pk4uVzJeY
OEu/1S65kyc4gkcC3nEwrALRd51zH0/j9clwiUi99tDQPrFxN0NZl9Ulq24uhaH8HVOGUEXHS+eW
30k1msr3hXimT/BC+4bQnXfAc2CT3EH5JSgTfyx0lNT25MAAviSz4J0M/QlP1oJ5C0X5tLO4a/Oi
Ad/bM3JO5My9vHOrfhMqjRJ5IEOcKervjK9N22Xkw/TE2tAqg14M6pBdhjJT0mpLoxGkz3jWYIYb
XbpUmtcbxC2c7T99ZFwxmwwXI2RGZJy5KI7197jPcHJTSj2kmFWR9rFQhF6oWNKz88yN4OG5bOxY
lSbYQl5/9bao0k5gOocaoWim7UsEMREbsNAcD1QxTqaGrP+RTpAfaDPoTevNd7T46E1rFidR6baj
R5jv7ySG2CKQp/MF1wV8IiYVMZV3STIjjM+ovdMs0us5bv54j9/W2yq6chVwjjMaAyP4h+722lit
Sb2r2twB5TbYavpB8RY6zNlMyZJla13brYJk5pGWGFwsPhAgsPQF+f+ehLjiKxHMzjvn6rJGYfqI
76t59VaDRZPbACit5fk7gBoT3t4GSLJpe/Fo/8su9RUKRAArVxFEc62PHyimW1XvmqfLUoCCcehu
xbxRmY5yD+cNW72zNzfRyhPXioXSPpMbkS3wiOttP4Io48m9FRhXzjqcYcMpf930XBbQsig2Kt8F
d33GT6OF6zxM2+aVK5pZ4q4wtZcNr6dAdpqCuFVoJV6KU9Ar3Ly/qBFsSL00nLI4HhblOnkg9WVw
j4+S866JODoUhogR3vMVMnNgspgoRKbSfXB9zlNWPf6vCvUfy4UZaAWJVroUTjK/KdiRU25uvv83
K2UF74zP6heZGY69LUDwTClkISMY8QckunkfP38NLsd4nfMMZKqp8Y5ZoMiyh9B8txYzniqInOso
AMdyvfnVwuTc8aQIsyxpglmsihUhrv2uC3AibcvxvC0zbhtx5qeV8iwNyCv1oTejklQZWUX2ToAR
qUszkUOOAUtIEV1w/uytw4RgTtw0vq62DxIcpYi08Umewoq4cGQAEHxz14tCP5W2q7ocuKqyb4MN
wCaeKY0tcxAtgpJqASuR6v0+Zt3wXLAYuEIZ8SmkknHOw8mqwOk75i1v/X632tZc1JDzxWZKFGhh
75wyqWwCzvKGNm5/9/O1vkUqb5dHOozQnvBXON6o5Nu0KRE6VTrMxrAngZr0Rg8PCloonW72Qn1n
kbqfy0Jk/0bMnU0AbwV/qIc6hpvzMNQgGbBd7eK04DkGdjahEIv7WB2AcS16v8N9GmSVwjA/hiH5
TyD0EK2rhxP8W+/ahKofCNzzfu6GCZnkHCN2s2GZM8ocH5v9MmGLdzXUDzfrJYfHyBaM70UQIYGT
MXqylaC2Vxm/k3QcKmUf3Fh+b0jZajVUlXxWor03MPUwpu3VxJ5+AhWU2XvKDYODPpfYHfRhMe1K
hmqoREeH4Yp7I/q9yZxEymV1kwMbqO6NyvhAnvvNXupJp1guzYMKRGhHT9sn497TBZ8NIMuDDTS3
MDWPjUb7vChCI130N0DuLVM+bOHUdI4grEKxd0sXejUMFcjduG/JOPzFxFzD+MyHqFMRVrzwLNeq
obWJdhdX1Qrb1+323+yMpjyHZ6KMX55M2ucwd4e4A90ED8pV8py38t+rXpr4aKldv8DwbyBBov7e
aNMe71AQ+/SRLzq5dfhfPKJE1IoKqTSjDH9rDkHWMnOl5T2H5Nm4s59yJfw97LFbqxduS3crSXxu
QYpd2/4BBBlp4CEMmqD7tEYczt+O86mlwGaCSxWZBzJqCN7ZKj1OJfk2DTTKAlRYHhU/e8V+DEds
gUFA9R1MAnD8XvjSMjuMEcIMYeHQbC+Lng7nIGO0jQJi0CZvUwsGVkMRaKsRJcXuzhfq0NeB8gI0
+M3hqe5WrZEFtFpagc/G8HBcdjYcFQZCkhlY/GOB67w1d8XpYiHfkKLfH/IDuRbhV4tMRQm4Nx6C
UawiN0NTRT0znzjKQiYlRYE/skBnhUVq/xvQhX3X0cUfVhXfa/+EVsO4Yofd9a61a/syqCunQIwM
AoTwJgojtbXPrD6FYPpjbX+fAhU8fhRGzuunTDT4lsz/vj1JKMAB+4T+jmh9iAmnZiSTol0eTSql
tCpSvZwuWqRgmfrzDFlmCFkPgCInwfH/NkWjL++7ZiB/4Nhf7XzIRDIgxrpIieuVZ9m1CwZXDXya
4h6Fdl24yCbK8WqZO0KuFaOUsfucgK+bTir4R4IPa4sAEbnYwllNKkwZGZ0DsIeKdkKA8YjNzU1X
plYGo3jptbwGy3s3tn+fPPJvwmwAM1FLA9lzWnnyloT77FncM+doRFWc8imwhE1jt6MTBv3vy+5y
cSdD67wcH1N5eHFD+QHwkbGJmY1yOUkounVga3VBsbpEE0JPCsQ2skUeOwRh5OCIHahncnekMKiL
8HTZh7/NE2vl78UbbtiyCaUToO7cuvTxasa0F0GCrqGpZioCO+CW2Jr0GsFX+eoKcUvfGzwXq0PX
gxXvZywhj8mBue50AmC37KWgfaCQWX4Dd3hIqypDn/t+y4B6hMtPoSSK2B5SbQQG08rhAbdpnguo
2rqwG4I7rTtOb5TV+qkO9Brmn5ZW8BKOhYAbYPegC4ePLjGAwCXxCPqQpB6S6otpCO/5ZIs4zfOg
HsNrWLbQAKcOAPxr94mgu1OcxEmCtXE70oaKleqXifdQGQ4/4+jzUU5xLk9YNm1ZP1lsbn+IIG0z
w97UIxZ7jwRiYaPntBIc3lHFzT11ulUWE6VH5W0zZAYySF6YMb3lCMrFVcPx2313QrnbOAM3i0Rv
tZiXVOfudQhR7hlFso1m+a0IYJkJ4BKXpxRBwgn3n9Y2PB3NYX2nShPKWtxEOZziQRlGjGPDup8R
Sud1kW3W5ebDD9RCngoIjJnbfOgBEdPtBQVCPstsfnwhF7mr3iGkDMOfp6Sr1eeA6UsJIsCi2my8
C+pojP6blQzBphh0VIOiQfXLZXl/9cevtWmzjvKe2y7luR8nihdaQKQwG+P2ukqLg2dcw9XZuUTB
piinpBVdzN0mnNGDQVgG0NjzCn0D7OKwHblgWUGhEBq/KheSCufbwZOD0ENH7TqzFn1NGB54LMlZ
ncWTuRLn2pGWPp8a2OMYjy3Qk11YkjmdwfPrtXBkR4bFO71/VuRQzeK1edhe/mOzMMJAw6zODLj5
zZoplgk/6ARe4qXu/uQxAM6KPONuXU1QyRL4zMJPXJD6XRnfOn2RUXgLxW6ALmYrZS2Bc0jhzzug
8HZXa+UrPwK1/cgBt8dv9zD2jKA4RBMVOlr+mzy3BvMdi2wWhKyPbXNrZ6jj/+i8d0NcZ3xc7pmQ
DX2r0tTjWIRdvfZYF97AnKX6Wfy4w72tGuIx/qNojxZm9Fxe6MHZ6N/mCH3U+BMTcr4HBSWmbh3z
bPRGN8uo/xOiyPyVR3MWkcDNpFFxeFRpA20+5Nz5Mnu0HGkidSmYi0ntpCCtZDVbpE/ag/lKbk7y
Zt0/GnXvYr3gUYgIclUAgY3X5mYqArWXH3fuuZQPgK2KnvCGjSJyvxeB4shQRONu91P5EY0hNDiH
CL6dmKya/iV28ma7+G2RMStD3lhbns4Ye1HCbE1M2OfMRlMvH6earJ2vhcKlD/C0zD49pafecyxe
RNQr3tvIyswRAF4PqMIYEtr6x+F6xNbNqbtrI6RrtL4/7HScyjoll+VFpWEt51fR1Rv5Y3M5xf82
uUGhiTYELWe7U/3mG3Da58zSv0m3HDjDDhsiY/VHw9aUDuRnsP/bmoqhbPG2xutdhJh8Y6TwuDQl
40+ZxMLRgnOX3Y7UW1J6RcuzPTR9EBOFtKWrDLV97paPMIdDY4ozh5nt+K1grwRlEO3WRh61mFfB
U6T7wRGTodwdD36vtmUhpzeePSgoJWf2GHv7MTQeohtSGXjquPA/u6aEKCxXmj7cEJnD2RgqfVyE
Uh8GMlnkyQQumllYU0jzQCsYDXDIujb32ZKI98eru0uZAQIBhXHnrh7VV57TQYvjmUzrtLJfS2Pa
4+G/aScvnOkCe5OYb8bFIX34raCbtYLkgoBqiJ0RN1mntEiddgHvVQYgLS/kvSfdA0u/ZNB6nenE
1Fp3Teu+pj1B7FwYC0E7s+5CZU3yOaz1Svyi4XF9pMlixJEw54C8dlD06MOs+qWWSMUX7QQUMSou
vrrzDNqkujArC8L41SayVR2MMKLyDDwgeVgHpNfZWr2V2DJmdhwyPELo3nH4xFmkPCA0hasSq48a
wFFd0391z2RvXaexb8gC9+GCuUB19X7ZjluJngSYYqO2xbtatkPfnnn4mDk67Ipa9Hjjcyjl/Mu7
REUSJc4rDfgTA40jV1h69Tc8cESkb9CyoklwTKFXq9zpep26kdF7Q7ZyTO9Gylpak89vuwn2GRHZ
WktE6B6cbnS6/PkegyII8hhyeFrVjAub9eiHscCAIPmvBDljQ0GMaEXeTD3BRVmwCmueszakUDA5
2cdVJJ9wUoPpXLo028jU0ZTIFBtNYHJhuLHdpDbqrfpHSO6DwvWXn4Tt6ixfrLvsrt+8QkzFS/NP
yEmZw7VtnbZRuSq7rHBhDGcmXNh0IoObRFq8OzBxI/qT088Yw8f5VxMDVXyXl58ysMyYEN9MEIyH
NVv7xD8qERYnuGSgHAuOzv1AsE33GEWc4OJtBwgLaFfyr348oUhGMw/HKmm8RftdnBpAYj8QNrRV
X36fhOHwLG/yD0WXihPQBXNr2E9OMAx7E3rc8qLPauiNW08ioxAQfzCf2Mj6+0FABMavnYN3Ka0G
Zs+ftiYOmviloWb90BM4PgFbVJAp9qu83kSYPs7NDboKMiWntMb56xbqaTreh7IJj/ld0nbtoaRF
wBuQc0WQVc62rQzvuVZtP9j87NhSX0BT3kJhGuP0J1JY97O+gCtmaOIVRGe/6d8ldofeaNyel4cz
ntnJj5Qrdeb6eSnL0iqg/5+IcjxJ3KTeNfIkC4H/3/SJxRBiix2gCNJvkWh4ZbZqKYjOeeLhMb4P
x7gj+613aISfBhLo4OX47qqSDzflk9rcHaqIJ2feQRPBGZTOYkGvDcx86G434OMqUo2g7DYCGx60
VevsRegl9eRpAipP/iskbjoezAgy1/EbRp2OOBGUqyYbv5Bou7xl7YlrhJ224/PCgA+eqiyTi4M3
7vCfIUjC2ucw91x44tRjho64hEDep0UdTn/blJLcKNWgO1JqQ3gV733ZVoeXDWAtKGlD1yG7S421
weLuPsp7dTEpomgZvnkTNtWnKiMZx7ocPb2osFvMxclA++CFvwgPGqX7KWFbnJ6uz71VCAaz3z85
cgGx8hYw23UJTXFouCDXzv0Ru99zskiMz4UTo+CI43imp9uA8mvMsVRlRnwuJOWB0LJ1rADthYom
qRrnb30bVfFUBsy7Jfsx2VDz+dfB7O5JQf/G8JCtv5umyZ3VgBj2XnX1apwNeYW91o7LBuWP4cqi
IKDoNwn8TXM1gwXLJiWkdAEllbzrFgTbtL7SQSAbVrfVgNqHeuOv8D/71XmSkm0pU4W7Qi6Bmk72
Ixb9gdy1Jc/JTpVnTHvmxQbFdN0rtJkgHOXOc19+drduCRK+Ckl/zQVLy3XQ6rV4ofgnx4XKXkcV
Ktwt/xEfeIm2MnkDUkJ8Jz4fvVWpqh4wg9UhI/AlzjLXrGmNrM5jGHWIobn9PyyXPEOJQtkkhzXy
wEJJndhxv0sBdUWIxi5H3vYwRrLaAAjXZu3d+A9Zfco8Pnqic3GX2GKvGhvDCYDcZWkKpwqRU6EY
wH1XpMsXWazbht8hzEsH8j6QibmnaJHxFPihxHgT7cWM+QmBDqXA5HrH5ERTW35/1no5G+8ELW8t
8n7Nqjrr9TftHSZhpqZTqzv8AQ8nfTNmIOsJD0pAsMKc31jas/cYfBKfh2CpPGugQe39WYQz9bIJ
1lbiEPvxnyKd1eR+5Xr9bXpZCU3jhnIwRVX77q0YHffyu42kmOmrROUr9VY+bTrROKXH7U/x2raj
YCeJrtZOsXKlK7+l/Ug1TRgZZ83BulW40KJWTQ9ivlO2QwDWh3LDTylz/HlDAgxB1RrXpTwdokO0
DQRtVXaxk28rDUev1FfzlSeeWPZ/PgnvML8FvIQM4FPfhZraft5Hib3YackAGnfoLXg1ecLp3Avu
rVZRvPUFuXRhXJz2TIEZITzcuBc42KWB/u7o1NGLDx/nY7aRUYkin+VLkEv59izNXKs0tLrU53bE
0ijMxogMHVkW1Fkd17C/nUkRcDqBxbXS29TBZFUgmP2jxf6Vr/Km4qtfJ3HV1nFXPStuVN0hFv7s
OoK4ow6SNrmvBUdmybKJslGcvKvIYwePvQnn0K9HxjGOF5PS9DNmo+JDkMKhyQbsj/SKhTG2q+rG
/EY4MkQCMWvoQr6dIw+Cxgq3qbU0MFGlYXyhfgUb6+j6XFhq/m/raxbTxhLV0hZ9D+lsR4MLUgvw
/d40ociWx1gNtjuu/YX6n6I4VKo9OEwxSAbsyUQUrlR86CEsGdrdtUOoMHbA/EtRmTk24mKufh7O
Qr7Akmye0atu9Z/3OE5vb/ZnM8/KwMHTTx5sM7iWwOdkHcFvLrVyDdpSaUSKCnIFZ1Lb51Oi+uTP
/IfJd+pKYM6DY90fPWuTTCpZNkrs3I8a1tqcF/AAXW6LmVBbWxXvJLKZBmiz8JtiRPLFW0h3584Y
rxUnMNXDd49g/blOIV4VxKEYJ/OvTTg2dQkSuY4sOJwy6sAhQ0kF1jVLXoeOOsnWv2w=
`pragma protect end_protected


endmodule


   
