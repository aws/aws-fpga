`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
bQK0SIEcdisfSwb3PhfMRoedAPSuEP8kLN+Z/JolLWRiZvRW8u4CK2rUaRpgzEAFkhHqNsin8hts
DKffVru6GJnKdjbVfKOhZM7qgl3d9oXnRDt6LlHaKvW9BPI/McZRxhet0JNB6HvgtBzeIQrTubuq
xYUp/cV37TX+ijVstLYpOVfTWXyTt/5XeQ2y2Y3xZYDPyPTlwJxby1Sp/o70/U0dC+E9MIZ133hk
1IVqR5TtmXLq7SrCo7oYjLf5y3LaIC4xfeFp8z1RxF3074IQRFbFwSyDl2C2RDaf0Yf0+fuaZgKy
HPPeLdw//cWutGA3s4OScBlQWinzWlJEYD0juA==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
WV0s6w3y9TeM3zSkCUcLwrWy81se0feGcu4DuMqbzvCitQyS0IuUXyQBE6B6FKHLUaL76HVwSWI3
oKmUmIPpM1TUaFszJIUJmM3+iVmxisCpB+X9/pO5qOfc47t5wDToRAOc+H2yKhVdlKK4UUQbxPAy
SqB2ioNIlo2ZWXIEvHk=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
mg/SRB8yKEr13rZQwgzxDIjVKVX5DtRLWlhLoHD7TEq/ASVYglJ7rE1BBJE0AIJNmGyTTiodQtkT
alz4xVSVUaSbrQ0dExDqNN7Gj2lc9KPEEwPHQKGOaCPNn+tXekQYjCSeWLEaHe5PEt0SMXmtrYNM
WAm0VwSFEtFZ7q/otA0=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6880)
`pragma protect data_block
gE2At3f+KkhV8eM6k26zkPrukY8cV8J3QQzaceBYLyfjxtlPwkEw2zFGzBCQ3H0Z0NlyHEZ4j9hK
KhS9/7E9i9TYDdfYr8ctfiO9noKXrysIXFvPW6cwB5caCDocWL/bVu0QVrV1TSySGOTSFJEcUwxO
8P4FnUag48uLB8UQKOHToBK5asDWzhnT0Fy5ngLBS/t7/Il2yBvBRihnTJy6tIStNBbHsFQ8mAiZ
fPfRPuOhqss2ObVViY820nBPI5WAiQValpHWIurMWHAkBwS5V//tlIVbSKSGZN9KXh3+YyBe8Yo0
/fCq/33EHMnJ3M4hz+6o+4ovL3PaZQMBUuF2y/PVTpeKVGi2yQTWEsuahmNQZGsIhdyIHLMhqkxx
AY/kFUvk00a+Z8lVfj0+MUDUw4QbdAahRlGrZ4MCIYt8WruKEVWndJ558J9DgUmWlEiElOATRTjs
kn/hbrnlbHxn+XfeX7fhLCVsfcOvLbH/gfAFzA68P8ba2OsCXS43PwYGaX8GPGyMvQ+lgFav8ifd
fdVCkQVzlNmnp3XF2iXGQS2gOfFyIpOIZl+3aPYtgQtYAztspnIPwXCLoMp/oaFEh3EZxjO+Dy49
wRIRdfsPhN4BeRjMlkcB82M9wvug5goOhuSvSTy6BQg/HMotlDYQWXT+iSGUZyXYg4ozSrpUUwPB
vtcufTlDWq4PAW6WLK2Y6vrjEWyckONcUEzHcQo9wfl3PQ8/4rqkqZUpI19FTjCaZdCbeAj4dPyG
y+556kieKHz39YzcFaQ8Gp5B2ONUU+XuXR3/D8vHQNVr2YYtQIraObQEJ/jjJASqOlimdIETWBGk
bRYmcEwpA/gl1CqquJn+plzk7UjsD/AD6R3AEc2oxZnFa+689EiB9OPzJnshoCY0YTJlnYJMernC
7onoN6qBbjUno87YuBQ/Ncw9KM3wo4KzwvDyTRieSTDAWgGi5sw6GjUuGajE4tsLQLwSmQnEtE6q
ywqqcdcEnXoHsSlI9J4dkzV/olgSLf/tdYhdKbR7lacEEDY9figuuzteAn/8jq4NZfJfZ8iICUN4
e0a00Yu0ig3b/pUT0baDgPiJA8URcf/3THuOc6ROhcF/NTzJN8KKed7CgLySKNARo/X7hgVKhe5Y
1A0kYhUgUVl3HiGmgmkXfSI2JzKg/PuMR9H7Qo2muUsFMx24O6ggVHd75HCj0WJt6XMRmHMlkKFS
TLsbG7X3NkraOp648Oi5GxQ4qLNClApBgrrwRxOWc7kg/xiwdVHEZRMUtOdhFh7vvXPHZa5lgqMV
5zdkonc8aQVwYG0lM5FrhMywpOjsC0suQoYKr0Xu9+GHWdYX0ur5aLhHlh/M9nfXTmSqmjf1mQKq
WLu8wGAsEJLWfSRb/VCQCbgYttlxnm50ivxhUw0RhoLrPfpCG8zrTiE0jMeI+Up9kwIv8kwsme68
JguvXLSsiIPEmHSnuVsMsLTJkkmZtV684DAkqbSEQbKf8wQIC9spbdLnL5IfxWHkIv7YuSrKJ1N/
WdIcDmBZzUDsez9bv8fe2rp6QkAi/UAzuDShqSbGRAybCmzy/td3UOTZtmu2FCchYaWRhrHNdz/B
tBYYdKneEeqJQ1zsV75HmEet4NcwgZjmdexgj4AhLtPjFuokG0dwU4lVuXkUrKcDHoqmyhlTti1J
tCwbicehoxM7sBNPkiz6+ee4Cqt6Sg+VTmuoNZKCvwGZQ3cb70bSWT32KSx3k5ghcUR5OU7TF+0G
Y8/8YHoUdBYaSOPOIFw5WS9F7q148i32+hZbTyWRPZlmn9savvRNe6nhjuLLoCkWQ6bpwX18EbHG
CZezLshjYBU2721uIVCk2+5JRQMFocTeqQnIxPuRykvfy9X96+sq/izFyfi0sbkwranzNc26pMDQ
ktjBbwxzGjsSahl5j8Ks+q77OO5q3mp3BeYi8BSoN4jo46dcvNxTgnDpRU+XptM0lYpgcd3m/VGd
j1SLrIwqbZ1TRMtTVOxm/iUne6qGP3KiUX/cz2R0Uc75o+HOtZJsPIWFFS0Bhw3oR7ddKy9pN3TE
taF5ahdwihp5AB2SxUp6t/ysLrMiWj3qUTdpZnXh5HRhqEfTCFtJIVfa0gDo5NY6geU8kOBvPYrN
p8svA/iLEG2Bq9SH85qiX72SUKRBPcvvAec5JOKikjyxnVWjipKPKG8ZKb+vk/WH/w2j2k22i2r2
7TQQypfUJkUyUpnassPgMtpqLEzl2N1oEt3BDRcOtuAVljNWh+9lyBOAg5HLxiiK+1CeCITa+Y72
iuMj3eZ0wtjkKwua7hKxgZCwddYVmXqh3hn9IoZGgcc8qWxeF9mHaJrpGXohxiycbrXiknK20KSA
+FME0lG+iwHODrOrPO+Ov/0PzBo204LN00csDf2nePdHrVydTwCSnyNBCTmfeIKAiaMJ77+xev09
WBqn2lTku0Kz6NDMjh8BONG6s7xDtQ2/4q8r4OjGqF/HRqQn+lqD7O4qz+B7FA2IC7Wzoiztj8Td
zFm7IDzupSo8ey8GgNAcLayiMR8fpaLpS4q8PM9Le8Qbxm9l8bGjdmx27mKUgkSi15a23Jhk/Xmx
CJk+K5rgwfBn8j0IQElZJXVnYve91FYE0MHKkEB8CJazctoNDmTz4GIz3bhyCsZhw3QH2JGlYBqr
4XTdV3L5K3N4595UPUyQKPOaqUZxbPjGQjeAHCsojJ56AqkKG7V6nbusBIZjRsfiHrrQQTyAy1f1
cq/kP8VYRRQ5opTc1rusQ7wsvumE7XLhSuqI/RZy1Eu7YwOx11bVmZK8tJD6V6CpaCrsmyZw/8F6
poqDvc6cJTK1+XuSsYBe9gzVqwrag0bXv0ssgWke1J+9LtPiJsZ2p0q5OICoSLFiohOTtcK9pmp7
akl80Zbc4jy0biEq5iyy6PWBqAzdOg6roKDeo64OUIgqwzrOZxm/OKiqYvYgHyXyUVvlAU6JMFEv
9PfJ4rB5epeB0KANFKLTes6vK9n+iSJ3ON4DlfxdSbrRuQ3ad3FC4XWbdIaaAXFnaJIyAW/0qd1a
7YDUe4MJ5l5GITrUwQtTmdEfWyo+HOEVX2hO3RQnK6uytT8xPMc52Nbt32uv5moO7vz5wENIDkhf
WoW7fcAw+wYTe12P7FlOAHnIexXac1BUPgga7Fbn+QoSSPCmWQ9G+oTQMFTXlyOwthp3mnyfaWBo
W/l7UXmQu7mPCT+fd3GZIF5sRA1nWw+NXV94ydi7eNyxMn2CcEO9FTNCbIVshsDkxwORZd6xFDBB
Pxx8hzqhRnsHxqNoGTyTMcGgAzzj8lv8bgLC0hwrBA0hRHLX0rRp3Fxg1HaSYivx2K93FINb/RHw
SClU3iO6jWwQD77VIdthudm4P34jwnvslKsRVhHsGdKcSbq9aKvKOH9BQFx+JLhxst8fXjfh6eNE
pdO1g7dLEGirQER9NleMG9FdqNDUKDaeZaC5BOlrAWG/Ju679b0h4bbuyP0VWR0aEllFHLv1omK1
13f/IG5YKBIJiNeC5lzzDHF+AHydSDaEqtgC17CmS4i5dNNwSVKVAwbaEMi3VUKc/pni+6tf9fnd
ItqAchk2ErmF2ECe75wOCl5vz8KVDAEGJQxw5Xs1FJbTJATGPVLH0yQFFIWuJhM48yKp9SKWQkth
Sbdsrz8fvcSYfcWmCHfwAJwccf0Lyp238yCLQFld2nLEYK300wBVN5OzQHbZwSySvYjH9J+XNGha
gHope8wVsTe8Meh60KjCOnwzVSrybMirA2qlUXpABhnnqDfkp3durmLjQ/8cGjH0MCLN72uGQo9F
J44Di5OHCasPWiDN0QrntSjHaMg7OSrPpDz2kxIOXvxKCi8NRC32VXv/qXAR8B9PqEi1l44qbaS2
/ZPTMt/LdBxgyvzzCNJWHO2+N0eKFUDKzhyIN58vCchfXHKmw6Dst3HzTKZ5TkIVcnGjqBWBq6cF
17cDJxLszOQORTp3/INjt+X12S+z4cU/qtD1i6D6MYp7fbxNP1zoC7A67CSqiSV3U+Ly7abHfxj5
1Q0bo7Musyil3ra7I35hefEpA/Y/50IAmrLLJwJkAb5QZjkwDc9QEkE/VwN6MCDwcYroMOSrOI5W
C0VOu1YhnIBIQf3JmO4z/cEsa5NiuiVjKWvlrRVZ+ZCnwtTW5Zgy7t167SeqfYUqWy5L9JTzGjmY
tPQTJpBvNCYZIH4iwi8EiZiXaOh+URmqmh2bg/hYhPm5PpHTzLrliNBWDHJodxrNxzid99xUtxhK
tY8DU4LOjuf6NO/t7w+oe7HO3sCdp+YuAyhEhhpSjhet1xHdRk4OzNodzyPCR0AqLrz5Tyi/9P2j
/Ux/z0rgh/7D7w4+/TcYe+GZ0XXBf29JsWRNp4zFzEdDDBZPlRpYfaYS7O9AtPfDhzGTfat2JB4t
sMP2tSTByIyms9a68SM7DqCUeLiifq8gZGQai4QoYjqvQyIdPHmc/Ii7mihg9xgCu+ZwqbePrWct
okWMnDoGB30WbuTtb9nVZXq6HPKqR46Ay5FENkGlIC33in0YOoICy2B0F4E4f2tHdVPGgFf2hqKT
8/3v4fx8pO0B0U9/delhtEQ2mPtQblGy+BCPzc8QKwW3sqiLOISBguHFucJHmho7R5QWH2icB8F7
T3JGwwL+2mKUPx8CCC/der3l1wSfGSEujE/RsMSvy2WmWi6irad0ZUxmGlW+9iZ1jFXy5czFYNul
q+qmzmquPT0leIA/nix74gPC0cWcwdXhDxqCLcCXXckkK8VlrwZF2Ziji6ErxR5gkFY43IlsPcHe
YnpruucImUS6zAEb0PsabD8F3AgeMEOfYkklP+/0Jz7HLiGpDnWZ6EnQe1MnEptrDv8ir3Suu35Z
TRU4jRis5lXOzvkVHkBENtYFdmCf4Kt5iHDBPxNo9hTQbLrSYU1QL121ZAJ0uo+oD1e9NfGWDtHT
hS4BLgomTMIwCGCjug1iMlVQkj18udGzOYcFczJJLGKbMAhIQarAIwcwGaFzn/Xs52XE+zpihOQQ
v0G5zBFJ+VBZ4/ayWarcFke+lVBMSZTmL7igQufVUfIVK3QcOqmhizQ7rWcpHgSoJsNuNJf096KR
jsLLwSmyy/HTKZGoTGXVkKudpXSUSFzS+aQoePoy82IpYdB/H914D8S12+VRyLSQF1438p+Y8Kv3
mL++2udlKFuITFOUc4O+1yZrrLjDuoA2KPl0U4EC/UmfiWV9YIQOnq06xOjGtMpc1fvPxr3IHsHA
50OZDUAwF24FycSKEf9806yohgjY0HY/8fgkVSPLMYgbBscJE1EVizqekgGRQkyHWD8gbpXlca0R
PRVM+liAa5MsOgdNG+UxnqQfihg+7jEYUFuoHMK7zadTOFggRwNX0OHhf8cSr3pWB0vVx7ry3cf2
BTnEovmrqzX4znXHq1nUAwMEU3yutp8cUojiUOPx2pYB5e/2et7lx5r1C0oyGZW3OkCMlysARfnl
YU9b6nELgmCrah7GpRYkCChVB0z14LQuMIMk7Chcm4uJYm5BV19ZSsdKiV18x9FHkLmobvu9kjvp
cGgkFpMaDBo4aTtSitBCtQavfBdt7GNflQVChOop3xntN5Nx+rjPLBvA3F9UGkyWyChBNypG/sMA
dlqRXbbJgrErCLdQDIJT8W5+UdcLicYx6Z+ucmHGKiS3YkoMY6KdhTDngEA9bGEVXzgJw/XPLcha
j3R9SgXZNztC/YYvAOpGEOcOTeZV3/6VFP99QHnoVNCP4h15WQ6wgAt/XKD5DnkulQ/kNoKu/YQ/
YEnLekRNb5zDzZsyObKL3Cy56+RikEJ0QFSO4OiZWbu8pglKl334fNjhUvei3QgAdbROKj+t9MUa
FPprOHvxYkqOlIEM0EhRcfIYhB73ihkBnzSyYdEv32oqrSNdytTZwltvm9IXKjC1IZRLdvBqdzak
ddhZKOufIEJ88pnYYqhbSDqMi1kRb1DQ2TnB02zlmevHpnxxWnQF3OnDV6V7k3ABp0PCmwTjNPXZ
bUSbwInelD72deoeyG44d1BJO5e83G+ooMJ2o/JO3aAb53kEjdRPpsGSUSXInDBQByBq8m9J7v9W
mYLn2L4RhmDa1mR7O9pqqwBhc0JgyOaJsN52Dth+XisbEObLv3mmfrqtYX9YY5T3COKljG1YHWCl
Zj211g3bPTDnv3R6lUF2gd7vg/+AmdHlN7VJvm1y7QlCOEO/ujw6H5XdSS2K7et9nVLeK7Z64fcP
5AI/ndEE8rmFNBSaI3b+WF2teoPsYLGzhdAskgLetpY2V4SzYXRUM903uVJtYcAwSRoCPTxrCyla
iUAUGz6JJRqda7hvvg1tjn8EiJogSxF6YyOEdfB/QXdo1HTPBJlsXa0nQypx1Csdl8eiGa0DkzVe
JTUHM4X9YD2FXGveSisEutKdgnnpEpWWTjStkt9Iz3rO9VoviTajczF6dnaid9h0fa9eIM6qxZ/i
m5GavXtznFTMPQVELQH8ixDt3zD/AnjF/JGKCk8yOslVJOWLkqaiwmeZyOy/YzC+kcoEw5n+zBUR
M5QBdHpQnYCF5BDdLg65KzHJkRNnIIQZilns4a3KQcG1ZwSQ+fLVuh76yWaMT51jtVRct+MPx0ON
dXeGVIETUd/e0pVoMnQzMVDm2GyBUmEZ/vnFGB+iU77mPA0mfsv8l+23+lDcuHIrk1aCoVOP3etK
nED/oFg5W6PIlS8hVHwc36I+kQ5+W2jullHXhIPcLaEctuzIWN/qHYur/MCNNQrANWxvW1yaioH9
6HenbfWqLSj9oMMawST1QZorg9Dx2T3VusPcHiXGe4xw6Y8EuN0KgImN/oQGFd58rqTYVrvZbWNO
ddmYhWlk0SsVkxEOaU5iVmfcyoDzLVFFreqWhnp+1/JXCUTlpbqAbUGLE8pXTidqfavqURmbhQvm
RjFynxv1yyX9jl9zZxh5hb9lS22gjOEMdzSBijgN8QvPeBgJBL8raUgY1oO0A9o7lwlfKtzROKD/
kTMFXwBQzN5xBNt+nvmBMmojgoCVIfNtT3u/ZIcybEv5UB75TWu4mFHqU2huatZfujW4hqfPG1Wb
aXlMSfG0+dWzAsfpxcheyHym9CNt98iGbHAKslTXEkYrvcZpBiEdo6ANYb0MW93xyO/hwuA2fVX9
4LwgClCcWpguHv7w/Mu96JIRjBRufti4XqhV0QvdIVHuOyVzIa77Ppu1GH2J6zydW927uA7InQOk
E/4FOxHMPBhqAINk0MQKbFAmIJjGgikOu6Hwe3NVN1sxYwa4Igs401omH14WeoYWdM6fhRXjYfi4
648L3WDAAIdzDADxdzoRDVR5orRMb1y5el0exhnvP0J3/Nb6/2uILt5jyoMMKaelPzKamxvg8X7k
94UIjiJFuGVyZ5FtNfG2Wt6XueZM+FybBgOcAcoZIZV5By1Gh8d45bEI/JSg71yan201n60/hWK1
fM5UkXG9qviPTRYCge8gDC22uhbkzO2fKEOGXdiy+OonWS+a8sLMHVGx8OmwGXwVw+aECvIn7t+w
TaZxQGTPjzcBIiU8RFEAAo/hd7e/XUE68dPT6RdnXBVWLdQ/emgBgpkh1BLy/U5UaoHWm1tWpQ0t
7L8kIpzXET6yjIHAmmKZ4X35rz8uW0j/ZbY8Ccii/Hn9aL3i8kizdnkTGfPR1my/C9DYNxjn/AVs
oDJxueRPH3CpQUgI+B4AatXYorao5SMVTvhbxgjoc4HZ6l5LGyBP97JrNSnThQOOpJSLtJaVrrjt
MNxdpP0XUyZdgRsP+gCPqtREwKDwbqhFuIMs4a13rVjTZZw0TYzVcVua8JKVRvE57UtemaGMpEmY
Ub/83Jk6k/T8Z7+IHws5mOT5zNpMu9wsSp0HhLLOLE6cQcuKZkNTVonRGlnPZuusnIXW1qzgp295
dfdnzQ0kbX+2DAElBzr6hFUuR7Wqcwo1WBCbTXI5kn8JwuhY8Tt8wIdeG29OArFEsN/x3uU2ORL0
hqN+ftHPrAKvb29edxbItC3jGtnL2L8tm47UODJErO28zfFfXo0e9+DNtmmWXLEne57wGFiN75Y+
0uw4Tl1KpM1V4JkFseYbZyq8O5NeNYGOwtYNK8QrVYQYHGFi6NqNrr67b1aQZUUVqFBkSh/s75cN
rK2I9OPQitcx89Lah6rXzZD7COnyQEOD7EJZ7tulOPSglROEttejqtxbjv/PSc4J3F/lRrfpA5n3
e7JID05JjEu3suWEkc5kf174RZj2qcC0vFFKCr2DDo+5AjYlBc69w13TkfNG+dCKvxuqIEMYvT8+
cDAaRMRNn76/Hz6eobrIPeM5tmh3yZb3T+fD3er3rc2Lmv1gmR8r8zbW5X1Hc91RBC4whVP+49UD
F12+MEumAHiqOhqbVLMoKJ8OQx0vz7x42Wl3TVyYg5gWWK5+15Id3RIlfo3q9KWekMN8nNxtjfHU
O5NeKnrczGEB3cYQ/8v/BFWJVWyP1hVl/x4Vd/NM2NHutGiZ4vjbM8DIcNU1WjXJw33pIAvlFGwy
LPrPzuZ9Ed6W0UXjcqzgiuymxST0cp4BKVnq1QuNYFsqj5pzGiPFQiV7JF/HilwxpcLG1jpJO3zx
74bzQMk4CecQeW5V3Rti/zHBXWQFDqMgaQ9B4coWX8biyxx5qObG+cIyDUjAVCcm8taL+0vIPExq
Su/sitY3QzDVG/mnCNc8+I/2B/TZ8D4/31e1VQkqnrhrKEKQDViXuykcoVXTtdFDMVaCGVU6nLPf
S+UzpWpejkKYIc4hbDcfsukHoqTCwWuAUCqwpN+pAb5+gn2wMbTpE+TwSMVsSxDls62oTXuqeoIA
BVXWurPYtv6F2XLShpEfg3GemyK2zKQRpsF/TUqc46ZTPPPyJ5SCCk7lLMm9VGHfjZ+SdoQwQpVd
7F3EZSnHYjcXBCIaqETbpk3cNf77HVbGlazpnWuBlIVm216UNf7gdMCOjAyGT04M4U4cyQWfAJaY
FaFTEDdnUtuE0Z4j/hn5phj+XVU6fy/vbuBX1OXWJ1jIejoSImyrJdOIfDjk4N4RqIo1SkcukD91
2RgOFX1pVn9LQFJWZONjiAGxhumeVvtFQmX4JrQUul72cfOkDCkmi8/SFWNg0Sb11eTnQFIWSzxK
PcNt4Ic4rBplnejQpFYPxPDDT9MintD5aXi4VuRrsZUHuStUmmKGTQ==
`pragma protect end_protected
