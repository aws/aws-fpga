`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
QhqE0waseJLdpTxAkWsuMtIgQNLnSj5Nk4TbUUXhKosdy/dgRonVYIVHpCWSB1ID4YbH+kfifsAz
P7Al2YmcrrOA66vlzdta6iQZw7u+BR+we4HHpu7vBaOiSKD90N6ASfXUtVwEFw2k9s665LWsyIuH
O0IqGMaq5Pg8DpXEhhM5C484yZVCp7RN2vHfpKMO4wRGQAYi09+Uk9FIaByjxu9StKdKV8RAQHhX
inl7opKa9VvRAg+KTZWMUfxpl4yQaxT4b/ga1BIR8jTiyF56UJPMur0gb1Mh/Zw3kU9KeeyeVbH6
4fxfSxUA3J9azLnfBYbrKncDMukrX30u/+mwPg==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
iput4jyIBKVHH3SMHYSWrcmPYC3lUxs832J+A/AeUuLogGkVBAeZxIsneAT8yYQbKEAUtb6UNZaz
/OYgc6bXEvFvNeB663M/QK0LK6rkbeanIc1iUw2WLkzwt0VFpItQ+b4XnHrcRRT7iLbDJESujwLn
9V7MDK6a2xDRJUeBPNU=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
ABEHsTTELOBx0o47eKlvdkpvOIaCnZRTbsdl3b2VfuDqjHcMy79zfdiBL61H0K+inDYvM1i8kiMV
t2tM0tAet2ugUG7vy0vlnc8XulbQ6MYflEviEO83ei2bsHJFoqmByX9InatoYMW7urp6IMgCnTE8
K2Bgi9WASz0YrxTwnvk=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4208)
`pragma protect data_block
vFyOjGMmSDDFFQPrDc4qLjH6pF/iWqdUMgB9kDJCjCHkmZ+zsX6A8vrbbooXT0ay83ZlQmeSRQOD
J0SY5+KbrO9uxPFdRQUbGazJy17sBjcBXQS+7H208rfhFP81XIoTH88blfZEh6EjG8sEvqHZwRCC
UPz4iuNm+0vF6oGtCyMhUM2Do3rl2DapApBH7vsaoOxG7sUDqXqTVssws9O9uzDdM3nVZsIy+4zp
VHz+33IzGI4U6SdN+oO/Pbr8IfJ4v+2iyQsr71jBeEiPMMibZzJpn+C08HXVcbsKSN1RClBsx4nb
Jm8YolF3PTPQ1dFVeEF3bhHW1ihw21uYhFMY40N34+yl4S5Y7bIXHOOFwkMjS31XbyL1OLt8Ls18
9ilYog4SQUr7cufStWwGwClAiPPSxhMSp3JfbvnDfWmr+tqwPDvv7lGLaHN047T+b/GVLA/U4i2X
bZOcbQj5EVEW9r9f4AbMiaWVC2iiIBWCTanRHkFOasF31uL+jtOZ42S7PTHesdlRgcaRgMU66QIL
f6P53+/uYEFbYfO5kXw41Xm8Sf+tL61Td+bD+ck+S6SF1ZqbjBRGQ3f6v/Sj5vmnmp7PWt3U7sqp
Qi/2eBsQ9bO8O8Cui0cMa60pKaib0gu6G8tjrKj9HurfHdvZROO5KaXFYSBGw3fG//4wyNOm4Jhl
FZCjyHsYHded0pAMz4FqjUMIN0Uh7YsDOlQy+P/4T+n+f6zBlNzoIZTpQf9v+63HC8XfmdYjv8yF
a4SGXXs5A2PH+xSUjkS8VhyO048MqbdohJtpQAoWimST4xKllc/yQs7iQ3b9IxVObazBxSszjxgA
bFPJN5hkf95pR7pp7yKMCCf++s3xUcgkOGpI7iPDr5mPZI3ghScocIHn6YE1v2T3ndI3ZIFkMRgN
Thwzxf7frBtsOuR2xD+iPBgEnqvbi8lHy1dbQfPAqSACjhl5S1TWCoqGN/292tz9x4HE+dtrFb3m
1soGfa828iMcxCy8uy3TE/h+7axYZNdbfpJoLWmj4F5oGBr6817OEbJZRSewpVKANeCvqvmr5aJL
jCPcQ1/lhIhvDmS9sd9gZY0u0KtPsmt4lyvxJSpg1soOgD9sfzuzx9Lso4qiyVFbNAZmAlmg46vR
FTekQruwej9vwK0b2nxKWP294COs/3CTmzhaeBpQLiUdVKRkhFyGQq3opFgF01hNrviE5HA4295Q
HGJ3XdoiazNRv40KStJ4LJE8/aBCgGIc8GTa+8s4KHpSeN7XmFIJDqC1u5fv4g01S5BqpZ1QPmnP
Qmfqxqn6YlsTUrJgxdxer7VcRibbcG0h0triTnK3hb6pPKmfj4rFY9pKLQ4frk4S/xLn7FIYlXLq
7ryreb/yD+D5/px4wW9ND18miLH8vn1Nne3SBMXw1DD1jGk/ssmCnaqMqTfvi9F+O5tnTTIc6zTp
bi8fI/v3qhjmhucg9RzLt78vJJ7DAZdJ+8AxCRT79pZLDB5+eL7TnYpBpDLz2HgyMszhJdVEgad7
vPhLyhSbMHRfVbWPJUazbup8zhJnKlKgbAG/ttm2TBOzpFPIpzh597LbKVlcoROYZ/k1UN5Frm0d
VD/dTSgGJDpyO0I+xfttYDs76MaRlBeSIRmt6B2eFiJg+MZPzD5L3SrPqx/UQQREBXkQr0yyw9u8
Bwiu8Tj1glSs0foJtP7rI4uCjp64BsA6dz2GgtgIZpSiX4lBXsFGiYRE75bZl3MNs91wXD9hecF2
GoXrP2OlpRx6Js5Xs5ZwA1n4sjW9xd2BT/I/ICutiatRmAtCd262zqe9g5731LI/uHdqGFdENN3/
eov+jaYp+WzPUKz1KSQOitGPm3o2neZeu4mVfxdKDPsiNuYUL9SsyS6V9O5QzKacsawM9gc3LO2r
3DS/DnjFXGBzE0A3mz2nFmnGy84CD2C1LuNrsj/On0wcPTL1H8xXLtLNp6PGrv15PRdPk1zfMWF4
T7nUblwYgEJHNLOPr9rNvInWmCEVfS9z9lmdPShx4IHQWyOB97lrIXazChUbgxFqIKhpCj0x0o7Q
hUIjHP4uAvRQzVN9PKT+IfoAWTnD8ZUctZxYWL/fagAvfQ6yNskihedm8OVnPH90SvocQdzHXDK/
pJMPatd7iNydQc4ZGK40r8TuNXK8o4CJMs3OhfCi+39yCaTG53NGS52NjmgysxsulUCq0F8Qezy+
w4VVhn6mXQnaswrXLcIqzoNF+14vk8yzlN0mab6cEHzutPR1KFK8NEdHDRpQ4oahqMdQeLVJuJNG
NJf1+TsScoVv/hdvdbckPe3m0og0qQlMTup2+WxYf/Ut2V68eTprL8pi47kSb9nDqza/Buzamd/O
hTtSN6vt3ecFkMdU/9dHE0dfCpoVvMmtDqsqvzGTQUiyogzyAF/40xFlO9uqZNAx7Uwk+9pcxxX+
IW4i4dlnGCr/ouaatcjSiI+Epb58g+iASDnSiTBLLNRZk3s5UDb5IrSSNApn2rR7nGIWu72vZ8TF
dMEXayI+kmgrNqRgVNOMYosCLJov5aGugX1mef7rqkXfquaciKXrW9PXhMTRec4jsnzEaqjChF0s
zqpO4gSbB4We1WkT7qw+1b5mc/3SJUny41h1bQRB76//gFFG9tR6XbE+w68upzuzXEORtaE4okRR
9mB+ryJqOWfiaTQMIGQ9LDFm2ru+Enk9gSse2UBGxiLdneNOsbCWv464iW2zqPdpH7yH5GYsktqo
7wX7WxpbJKAXl4D/rzFFfI78u21XiNJY7ezFIVESdJhIQtmJDixVLTqX5wYeFr3TGc1rNFmRacaZ
LQWlc8ixgh2zhcN7/h+Qjzb4sKiia/zQ/S88ijRZA+9bqphPJT87zsBPPYMP7mXzUXC6A/y4F7F2
UE9ljh4B4o8GEG8u9skQP1A/ux8tAUf1XBGjcnCqjy0MPZ2zrWteBByt6Xmoix5PE5oTNZNB0Xhy
KWbVZ+2roCcFKtTbUtWyt98TYinYVOAREEmD8frYQfIc06cvG5K76qmLzAjf8RpPDo/hjMoN7CBv
qpVx1M/p98fmdCmJiMlG6me2C7jyaBBakKmkM00eNEbLSXfHBzRI54u7r34OdwirhzMBpbAx4Fja
6aYfEf8JFKxvOLswayEmx6HkjPnp4g89iMUxhGHTUk+jM6fqgiPexix++sTyr/iSmjD3N8LZXae+
tT6zh1Npd0NtliGBUc6mW8bmP3HsxZVwIeRngN2jlpexDOcXL5BNZSlBMUnO8CpwCAerybdbXvY9
C7hGd/eQf6cuHJ003Mc2oQkdDfHpREvpUL2zBfS+qVPBRf/FqSGXhcXFL9zfVqBFmWcj86xdUiQK
iYBYJtSt2Y7NbeUGi+ujPtvPcM3EpIEDEUsm8hxxUpU+/8bogz+IKZHu6pWZUPNz7ow5SZiEkHPw
JeA2qi5X+JXK3PDgGT9VjbFJLBK9c/5CHjf75oxJm+xPyXaFBT+MwlYCys3pP5vVwZE7zJrFk6N+
Qna0J+FdZEAcUMNUZ5XwpUOH+PWHdQ3pu7JFey7jUATXBKl5+rDOd+cN7artbft6jQz5Y2TmQf3S
8MQbs0QhhOLq67TxXDjetH3mK0HjDS6KuGhKHl9GI/MaRq0dKhBCMIADhJPYIFn7X41/5K2wO3Dt
W6DHUdT56DQ+25DKk+QbX5Gd5CPw+FE1gwvgeFVrPMWYyBjn8j64aTBOwCXwm+s4gEeBtAKHFNfb
/+bf4YOGmlvjHj2plS7s7v9WHT3ixJocA3or0lpAlThm4lUFBJ8GPwf5WY8l4lqMXtXGhwvJMd0G
0nR3O5/nNKgWQdoypUmRgCeIxijGO2KzCrU0olI2GTN0bGhz5dTosqB2JfnGNSx3mxevIFMuHVO2
GO7ESjyUoztooUgqKYhsfzQzc8Nja/IIXMNmH/dkRSxhF2fIYpA4/QerjgoEA4JsMuAu7RKFRkyQ
7Nqz5wf3ABaOSIUNG7MDz2ioulauXc9LYETM4NsbDw0B6Pmkg2i9F66q2ercFVJ05XHJtw0iiFwt
imp9+H+f3hDBleY0tNtzd17hdq00m28yyMF0W6RvZD5RAAyFQrYKLzxGZmogrs/RVFZ5Glss59xH
l4AxIQXVbjBapRP+XzUCZrDxv59cUnFT3LYGnLdNQMi57zW+QPrayPdiYh40IgvaMtvjvzVZ2qY6
VkjsvVRBDT+mfTsuhtr5b6ffr0C1E4aGlEBez8xiQonS+yDKcnXc9P5eIWAHg7O7tpLM8G3Vno1G
K3ax38WnYloVQxqUR77pVp3XVHkVChIZ2mWFbc037HlRBq6leOO2PRzS3ouRfjSkXoDIBrQYdXUZ
JqTaKcf19sOcef7wEE7h5o9Wr2jTMFpsEndsPkOSOuvrFLDq+JDPwkEWGByawom0nytaTo325tNB
IyHlRU2JPIUSB8TJyS9S0/yGm77XNmHHxhdD4mjc/TWahqmg+bDiINlYVh1zsrfx/2IELo2VS1Fw
+qf9La000uQZqfe3p1hbui1I6UFAkmTVUilwTqPqFDZrIpIz/YZlVynw6kiuJS/dfmEOzmOg8X/+
IMEBrAeDo16vwy/3SJkWjBxSsLNuWAHOw85XZyhqjmaRgjfhZDN5Tc8IWBtoQ1acw/UM6pkACq/f
CMNChqn2f3HFEpCIpAnRsWS8Q1kfg4xXliCyc8C8GPxfoXjkWkQrWucXBLXyYPCpAM2j08zRxT2F
9UHgZCVnaHHzrCCFTxVp2FZr5AkmdDQKQJAok8ku7UJMIr7LwHQdS34+7k5sOO/P9Nv4vRxWTOyZ
/Fr8XrZrVgeZ4OUV8iwEoSowN5dVZUAYOpm5AyI+8+2gR0BuP47uRp8uAJc5ABFYIpIFMSuxhODz
9kN4CsenKQHvluJanRygzVbL3x3f7IdK85wOg4kagmEtRG0XHNMbpb0uejfMI2lBeSgP6c8mRJ0Z
cjLbIy8Zjvvmdva5G0BpON4QqFJSmCHMvwkOa8Jy7yBjPwr1c8AfikMDElQ2dwE4v2ZnY/9ZjPci
cuD20vnFmw+It1bUADSGHV5DvwMWU29Wv5GuTMRj6dlxkK2C36nM9XdMCgF72uPSkEQFwwcjCN5r
QQxH+TZQ+Qw0GpGTEOe7Lq754ZcGnCfIrWtI19gtI8h3EhEQXm6Ae9xG5DcQfUd/qL+1ZQPDRoHB
PMrMZPDCwUWbQL0W+oEpbO3WV2Gs21LNGQUT4WSe/1I5MB1+ph2b2qKBvoHEpODD0h2hoXk1VqDa
ZDnI4J6F27/S2lb4ssqUB5czQSyiPsuc/VjaDNSi9LQta1jqWjJRXmM5ht9cx+yVXLT5Uqce6v0V
PX0ABCp1dnPUHotOaqno2X2snhVFtsmsFQzO6At/3NB0q9Ege6DDk0AYFlkh3Ez4QrLLvcvFig4O
SkMrcnhUaRhqz6bqZVojrBiNB/kwrW2mWjCU1roR3UDYiol+u8MPl4tVM1SfwN10eSSlbrLoX+B7
gP5ZfblRZ07/TcjvmgevkfmTXstdrW/cLhAVg9IjOzSo150mAdnMk3+W2PG7gdKdgib8o/3f8Oln
0p1wcLJz4PTKwDJtByJJmgI7rouTBhDKfjft1RQE8EjPh57mTBtdk1XPMymw0WI=
`pragma protect end_protected
