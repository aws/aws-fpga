// =============================================================================         
// Copyright 2016 Amazon.com, Inc. or its affiliates.                                    
// All Rights Reserved Worldwide.
// Amazon Confidential information
// Restricted NDA Material    
// =============================================================================

// Value to return for PCIS access to unimplemented register address
`define UNIMPLEMENTED_REG_VALUE 32'hdeaddead

// CL Register Addresses
`define HELLO_WORLD_REG_ADDR    32'h0000_0500
`define VLED_REG_ADDR           32'h0000_0504

