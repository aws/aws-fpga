`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
EvXSzYKSLuX9ZUaLe7E9k92+cHyyiB7HahjHflYlNFuK5ShizEeVctVCgBrKHjfr9vZn1+3dmvmo
JRTub5gwp7GjdfnZIfKSjaR4qQ7swjOgl5JkSR0FhbZuKIIHVlenqGsuuefn+ZqmQftpR8qI4Tev
kWo+HGegffBja3PGYYEWpf7J1iQVRZwk/GeTym0vqQsdvdEJg3dxftCZQRtIXSs2siRRq0YuIiK1
p4ntTJ95bYpFQdURpfz8EriA7qesVCVcZG4vQECxXKECFD71ik3mN47VOJvFgqQ3HhoMdknHsrIi
EALCqzvXaGADS/mEaopLxlI/ZJxbgkV/v5S5TA==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
qP2S7B/+ZSUArnU8LcPegaRAKwil4cTZ4MQhowAk2dXSLG2wmH9uN1iLjFnUSiWbdrF42lsaAoZF
P472JK7GXx/LZ/4tgG4g3HJCUD6x7wluBdbX5FVHxvFW7svgChsEO21v58HOxOo9hANHh8jzUXuq
L2fyDauJPbJhSWok5mQ=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
XK+3R6UMy2sW6sfvvkGu4e5W0ztOJL/emtKjK600oekCBviabz9XFDLvYlu9n+COcv3TyTMtq0Ug
fW9ELoricJYEATbv3krYeFmwxxKTFIRjKzjtEHVpveO3Ba3w6SDqaNWpbqMWw6evbqQgOUJnGZAL
ucof0nWkOdHV6aSmEs0=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2864)
`pragma protect data_block
M9GLBetb53A3qZLSsSy9h32qafQvXyWbZYnU6rkuCmMmq5K6/HL4oSG7RAuoCHZpomiKu2bAf8rl
G5ZYjSahD7feil/jf5llnOEDrchxbZnbp1pSEYP9LAl4NmQW8btwMCgGIEubLWA5APCceKFzXA+5
xOkI/ggeXyLW7t5kC8GhyB+Xg7Ye2rAcFlLf0CXgRVv2JAUGaohDOFr76It6rEGgyd7Q04M4iAsC
aNToeWuxg0BMAifXY5DEIgA/Gobomh8U7mQ/VJpp9WyLVbDgBqHfdZrifrCRTnuxgjHRLE+g3Ln7
wjzxpoIQKoCh/OaHw9AUxGd0L5qL8PDGBTOXSijRNOVQwLpRPJ+Q/pVxRlH8+A8EY13KHgekG3yK
H4sZbSBcJhVKRX5d/VfB02tsx8tebdIsTY+SR9LdRwxswNlu+xuI0v2QGQGx1Qmie8Szk0Pf5b1H
PoBU1kYhIHRerP8WtOKr4bX4tItuAUTcP6DzeNNLcfafTULnsuqJboyRfw/YOqL5NFxDK0IMR+Fe
jK3K+fL0PfQDQbfSNsit26OMgKIvBUTLRodb3krKyG5oelxwmSJN0ziiDJqGxNnd/d9pv0EpqPPz
uehkjfEnISnoxcHMCIeBFZLSScvg4bIwA6yAo2ov0P4kwVH0BfuM+9dc+yrfXkRYHtHMwqaldwgX
wVoMTbQ/GDod8hoRATcIzhjn3zhO/M0Aus23ihCRNOdTdTO9T+VCcTAoKL0Av0GdFyfIzqMJ8haE
n4h4zVdp0gmgGVuMm/alhwwcZyxfLhHOAq1ueHNIM2Y4ciidMrACfBGQJ1Zz4banrKmMrxCojajR
1bjDbQFsPcLxJHCac1ZZsVxjtGeRzrmSDnxCbOgnRiHW4Oq4Ike0rPLEaQ+eNEB3sNc3a8VG3Mfo
f5+oI7vCZNE4hne+vnAbw5TC1Q8CmFdLTNP91kJKfS9PaIZHyZazcMXk2i0OCtFQbqZTXBPwA6o5
yRwVPAEWSWKGl/RUslaNDWllpjDyRjrs1Aznl9muHcgU9N32VodDAGxWFriUzdMzRm+GWNp0pP6h
EdWzdLgRMYW3TOKt9Z6Fe5kioxyMUOAmxZaM+2KadyYcgHK9Lkjsujukqh/kj6ugie3x3OXd0lsa
csQi32+k0YrwT+NNpGieZ7MNC41RYUizDBg9bHx2iQwZmot+WN7FDzwDF9PLb8tFdmuS4lF7mCmz
Vx2dw8ViOza/aDIJiV95yqO3lExGhwoyu0lRtAPQoIHIY5XMI4nq1qmkfVJiOKoKMvyf++7CPHsp
onHaOR/p5AtKFFM7tsdk72ahtdXt7wLw+f1IUbH5BTozySesvZpnlRSOm4bxEQD0TBIk1ymzjJqN
//i5ygJ9GcMLVTu4GuF1wG2An75chI2YlRGFv9KPAzTlcDzYkAQ1Ahf76qdkmkW8utkfSPTMNVhd
OUdDKumRCO9R/XtSWF50758DUONnP/NjKyQT0JxYZ1ytcL+s1Za5HGEEIgQfQivB9Ssp2lgPhPnY
zQGrhUcZTRH6SPR1bQ2B9kOI+y3t4VYiLmkNalaMCxzm717HPmjG/+3Vk4wYxPg5q/G3TlhaXDJ2
3KNw//LPJDZ/bkChxWab5xC6U1WRcHMZhkbEwgnOshpVL/t0Ss4GdaSsB5aDTrMPoOGqh0Z1x5hj
Y5dOKSJbcD42bEjPD11ObxZbpNd/upjKf8jP+SN0+CVaJj5b/qiIv/CABbauBz4K4SbLIr39qv1i
rD2NK5gu88hf8XyuzeBOl/MNpOIUQT/LAE/yOy8fCAv5dLUsByMyUYPaURaCEfZhoF74GJVbc2Jf
STwhIJZAB2bC7uZ8YM59Ohf+8C8yzwJ+aLNrwiBNpSV+Idmt0/IXjDjxgjStElN2xX/72UN2Hk4Y
ssvCCgd9Ur2A4gY+F2+wQAfnBq9dJT0E0MMFu7aEmPIBbxnJWiCLfMa0OHqZ79J48Hu8lPHIZ12L
J69OPYI3ZjSVEjKjnz0RRsxfWzz1gTfTiCVAevEXKScE8igI63wmE/gxWX2ixlX0zJ+I6glITf1f
gH3bxcibzVcNlA6pKZ6VUPoxvhT4lPSEnY28uUgC712Va6XfuvIuPFCp6DG+5bugeaIcv0o5LAPA
SMgoeYekNyYyHU4dZ1SpNof4jc5LrI1jD/qmuNRv9NNyfrMQ5sxxv9dVxzTiXol0BCDw9/Sp4jGA
dlELFHc2ldvUkc8sPKJ3WoJX+IWnSWxbK8gpSETHmDKbT8C+sNLtx7smXx4cNSdavP97jW4anDz4
AliuYW1gO1SQdMcZUeYh4bJlCyXr73CIeKaHGxQQpJSvGBqQ1plsy7iF0teiRESa2wG0wu9FZ3Zu
9P8XiEfD+MdAxLnAn+b4IyWwtRTZ6sAQ99V0T/ijbH9udFxhwbRO4NSo5JCjjZUXuomH/9hM+0LI
bhNHrIB2hpNXpCg5AkHkSw4KA8cDXOdVRVxGM70CPHgmk3H0GEErny3sGHedAy/izEM+ROStFEUU
8VmtPYVeGoCD935W7FPEL396cjiaTx//x8F3FlgelGubt/Ykf0+SFcsaJGVJWHh3reqV5JGQyw4w
HaMt5f9kXpw0DByag6PEYV/KkDT8xSmU+o/vPm9wU1zyTabAWCWjR0Zy6dx89HFlsiyA8q9MuWkm
+j6IXZgX7HWhy5l9G9SmEsWhowUWVaIC9f++XMplvXQYl4rNz/zGkRTPUqQlgrKudoFc5+YPf9i6
9ZBenz6YF1Ow4HxRdLQRGok1rpV04n1MxtHn2RMGoLYI2uhn3lUECL0L0trglc1v7D35nvsPLvSE
1/JHNEjPgRAbD5v3kzU4WU+8uq6kdww8jLKwkmvpdOuVLbmoklrQsJTZ6qqUFKjqE+84QCLS2/k9
/um4nY905Mt+3sCu8eaJvp1TZxOr9P9hrhTPu7bGPbSK2Dqp9aqb3z1x4bdJvibiBDtkqRjXq/AA
nqEex1QYfL97zt56T8FhPJDKvroKlSiaxMYLv89TKmX3J1++XasIWKKb/Gw1HSZMQO3DgpOaHr5R
JUPa2tP/ZGbe6XxVcU9xHCBNLDs5OOYwYbl/E/93AhYGiUuFFwj4yHUJAQlGUIHWLvrG7rpia/Vf
LJpfuyHFe4TG3bpDa983rQJRl1JEQ91rxpiEbUMdaQTJdRywx/uOI6zjB1ngjqojO67TpV1O1KQu
yZhu/6qMtzs+ggkTQQZDTtr/jKHNk0TnXrrUPN2MpNOUqmWO3LY+88xVRTqWDOQaBOxl5USxRCMq
WZXCkbnWPPptfo7KF3PIIFkSptF2VrGw11cy2tIpFvSpxjWbGFb7zfUFN/5fpi3m0Dlwt3diqS7d
4zdV8GqBrabe3jGINy1wg7LdEtjuYy6PGSfLCD4K370T6pl3dMOyExqFztNNF7Vkl2pXFFmal2Aw
BnPL/1SJsZzX2rOut+UFK4UiYZLPt377euEc5erQs2alMfjo8Pe/R8sbRqD8/8AhrzBrvvoLYweD
zPgaesltBSTlAH+bQ96Hh2OajNrW07Z4cxxe39feNYZiA4OZ8HCcf5VqnzWx5r7j68sVJ/Y8K9Fl
xrwwCZ0Xl3VF5jo1Eno9uoiWsRAePuiQ2ZhSH5Q5Z9SzdHNxFjjZgFGqMyVIPmuys98vfgzDpJ3P
KcjA/g3E5McHwNJV/tZrR9etECKaBVyPI6hn/xtjcb+TXf+RGS0f971UgkH9rGBnYE5HyZznMvtn
pYHyEnpyePUP0cLhLvZX2Nr02TifZ6FKPlVkWaQnx5nOSA7Rk0IFuomgybaqF3mQaqBnBmqtQ/st
2EdFR9UsuhrR3Zj0f9Q=
`pragma protect end_protected
