`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2016_05", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
tl1xVsb+rkY5WGoIgP7xU1TLRP0uWt+MM7ogS4WvX1mMhgD8rLgvEkFEELe1qmrGw+qJ2zM45QFd
R7h4Q3xK4gOg0bKrVVvf/owgZw0ZKgjkrJnj/dXOTBNEc9gAWIFEeMt/9gBXUNFsmS6i0gnj9Jvb
A+rq7FXW/PMh6NbDVk9ao5cUqcJOzmY+o1gdFQdbKR8qI/vbIdolGbM1KaHQ7sQzRKEbXLMlv/1h
WFI+WmpFhCnzjf0VGdjRKGTUPgfn6lEmy+5uxbGq2m1BNATkLMU3t2TusVIxsjGvYCkBSXRt2XWs
SZJEuC+Cx+bZI7+4+W3Tw912DVmlix1NQnE8Rw==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
SDOC+oRszem2AFEBUTK0oLany3V6TCo0rvt2tmRzfsKOSxVaVSrfcdAyYYUwqYRHfhmoJ2BXWmev
wolwT/FPtlfP4QXWMZWaVV4inqWLbUAwg3A6mT1+W7Wd+NYsM9hWdlBHwdeFQ7GYKoYSQVkDwNVK
pn2NTjrb6VgFLVwnGnI=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
LnbN7MZ1YmwYDP+TIDZPLRnYvHtMOI7IPCrTDcHQqh5OEymsFC84j4tzGoT8tUBkwhdtXkd+72mG
W6VtfxTKFiqhgxwxvbycsSqrCJOzU0Y91tkjWisW0EzH8LQv234nkrTZ++3KAOQEvjzdMfeh9KWw
0+fQIUyp5XUTyDYWJds=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5824)
`pragma protect data_block
GZ8eWzo/zilv8gQqiq8Ht6oayq36kfEc77VW/7sthZx6ODW2qIVj4W1eg6k8t5DwbfzjmT2fBPQl
cmHu3EKmvrlP3g9swvdXdZJKkMWbNY/4NgoYTQsaS30o2R78856j3i1Iukc4j8Z/iu5f7qXzQROk
IczIHqkz0WC5O/dABYXZj+uSP7W5XTZ1V70i3dPJ5d7KLacv512PQn4QtWC6iGr/qZjj1sD9FNFh
ct0n/xum6ao8FxkwzsJnfmv+0EelbxmLSraKbF3HS5SbNO4CgwKDuRdkNjwP8ert4FhDqBPE9T0b
5uxiqyl2qjxv0MNHfFlXaYsSXpHjJ0kJ1bpQge6pts813fUT+LmI2kgoF+lIASWAGWqjg2SKaaS1
hlmMVOqwHdHTsstkCdzqanLSn1esjAp7fPtdjXSTY7X5DmA39oZCDO+P37SKkwShqoro7jdlNAtT
ALf2gsNFvmGBqXirRobxMV8Xk6Tz1tun/RM0keyAipfKxaqySUk7QDpPlsjeB96esgDr07ytQ3yH
yiOjEH1nRQC+Anqank3fRG4H2qnt29nND1Z0dSBJulUoxYT2pgkRq7cH+Qyf4hAws6IkM6idyu4t
wPyx7/9P1xLvdFouWZpoz6hnpXY3AvHv0K0dn7qoSNIPhwiqyB1chcP7tsXMKEg5SpR6W4YR+xMb
i8F3jurWemg+hOLgkdb06FCLe1cME6Tdi4Wm4X8a1Z0LhGmsfFR/rw/0uXiOjXSLa1Ic0XxDFEP1
naW6KTI4cqHZX+t06WnmxdyxxX7GfkGEc5lEMnD3iawEVr/EhDwfv/mLQmLCLIR1KR4zSLB6yAGH
U/O+5bFE76WqpnUpNO/SnETuqwfYeUIbnWFTxqC2LoDiLb0XsBz8bVJfofvMzvHa4KvT8Cyyw8st
E788REGEpcFQ6N69udlr/oHVjuGVKVp6ngSwi0yhHQ34tCqgfjemopW7Cfb7A7wZSO3kWqxQS1Rg
HJcQXKMRb8GKmP8672NBgIKZTAnSCbzBAdeyhJ0W5ug41S4uaE9VCt1paTae801ThPjOsU2LFA47
C+Ek/m203AGHtQipgBSA5MQKMFAFWMz3Gv5c/IyFh8jk1KEGo83dVRxTSh2NoVpHcxfqjjZ6L3ut
9qchtLhAy+zVQ5q9g8QurZlP/YB5KAZt0bjgzDJgIzJqG5i8lg6C2IJPhbLkiVNh9SmxGDRt3sA9
NI31ySluIAcvP2B851vVA/rWqDbTTCEGbHjvvaIsj3EPgtzBCuJFjMYu2FyfVHrVUc63k3QVD2yQ
PreRTmG7trmDKIxWOI8sa7mEP/DNpIarXN5dsWfE/Pg2qZUACfK1x7zltpDoyqGd0d6e/es6DN9V
Brap7JRC7JKDhArdOhqnUFWexeYcgVHg/UUBEUDueQIA/OINIQO4FLvMPlNnkOfKGVhlxbEh4C72
sK5wih6GdSclfZoiTWzIMboNZpqhiuKTbw8AQ9SPZbhJ22rz40Mc+JUnIPqoOID2PbpvzHIWFmyR
9Eqq/zHFb1sRBn/smQCJ2wmT0SPZIxys5y0xxf3HtttAWKjHHDhNWChNroQrRN0YepQGgwh90T1u
/AaGPyBhbMmp/tknHRVrbxH6EVuqAoSIGlwV3BGjy7RAGq+ObjaIof3BXQWe61yCk2HSbQ8N33jR
NVkxwj6d796qNrpA6K5LCIHuBSiVM5JlqiJyW/I7FD5lpLvbYqrkuVkyDnEyViutiZ6szGCKP12A
GcJwduFe+SJnFJ3xvJYmSErLyvN4FUHqGy9CNF4LDgeZ2KnSTw/VkxqghtJbULJ5xBQPCzFWPhub
hueqM2ZK/dhQwwGNrRzA+C0nzdV+17atM9okzGsXet2JYK9b69cH/e0dHMZ3NLWKgYCguE9uLQEl
ZDcy83rk9yzJOpQltU9gHraNVoWJmaCE3/hog5H5RnpyoRptCkVI2j/TSyodG5vaLei5qYJr4Tvp
NJgrCvG0oR9WFHmKK3Y0N9mJYqr5yHiAWPjeukHraUbLx8h81nIz38WRN+I0JVRZMDlcs+j/Dt18
vy6Smm7Ckl4tHNBJcoJDTfNtte2V1Nvu1hmVWN2oTgRZWIwMAkwn3h1Ze5awmSMvtdXZYCpn/Xfv
yNtGLj7Y2DyMG4AlHPY89Va/jBgz6zQMOdwY2qrh7MCE3yeixmKEeWCgkQRnKZz5RlrNh+hUr9fO
X5vHKd+0gT90EV0Du6mIK/K+s8hsIFvpLK/fJ4EAoI0oJW9GEdROC31rUszr0za5Gllh9HdaMM2u
pDQCMzAKofDdeWBOTDIzHhjVSCfYr1vFd81y+la3g0TV3la9wnCgEjF5STQLtPp8d7NwGE0sCUsr
JLrZiOXX+O5p9PyE00cBTK9hWd+YaKmPwgVQxMfiWZSe14mrIoZ0SEuU3aiK2dcQ4h8XEA0CL5XB
M02odiAFupD6K8iblv+eYvGQeOwmy+w8cnO/O4NYMX/apiupJP8BQgfe086dhCESoDnOt47Bscw9
aegMciLAq5aPmvCGhMfwZmqJCq4A3cw2v2USFoeXneiuTkEX7//eCGaZGnVdpG5uR+1v1QCBIUJW
haE5MXarcPglRit/vbVYnfTbikZtx4tjKMotrRs2s1SurlvYBCYeAqC2qi6uwx1O51T5Hys1Uzvq
as3xK2sCUEooXzEZw6ja31+2v25BsX71RmYxzL8buylxcyGlSqqS7iKYf9Yj3Xi/USf1Q3lvxI1x
uVnmKJprDicI7BCulJ1PReF2Y2y7TNt4eewVI1VsNCA+OVR373jEXDZZnek8HMzkQBrerMUutEGk
w4lZ6lbfJRE+T/HLBpAyWTUfiXCoqr2G+fiT5eCIDKgHgn/NaxrbUz5lgpFf29Ik37au7UIoPZ/0
L2UC5Zy+ym9BmDlc83QEKC8gcWvgHvaXVypxRZ/+g1DUceYfEgO7UTsYQ7BZ85h5I/cJHQp3+4Hf
jsa9YWJqYOD+rCv6dVN0So1VojaWshxj8sXOtZ3/OIV0TTvyhwUuU48xsUYDCm7c9zysbUxHHkuI
3juUPjAuAoFk9UzMQcm6g/DWY88fmNSUGXrZcUnYJuhm4ALGZy4bzYlPQIKYvVQbw41txZKc45HM
tmjfvToJqRSY4abQlwhSL8zW8EE0CD5TOWMC8fqyNdXZ1bAZj0MnqEoYzaBfVPEoIdPYSxxplJg7
Qi/YhJwhGOoYev5CSVrccdJeIZxjhWe0NAxOXkFyS0Eiij2Up65IsCLGnb9cuLjQj0LLjwcX0ZjL
jEH7sS8G2TAwIOyYa6NKKMbGGKSzb7i/898pTH5FYQupRNqIVmkAm6E+rvFpp9YVdRzt5bIybH6w
ApnDbU1tpU8Nokg2oF8CSVmi30aBfp0E055FpeyWdnPkUE/YzwJXhP0NA9Xen2F2sAeiRdNJwIVC
7MI4BTA/qx+MEF603o4RBbk8mhEOq/FY8MSfC6Pmc1A2XPuO9o0KgYxkIvIH7c0E5L4lzxLOFngL
91laYWK9LqHkfHWTHo7FOmaraSYhidbcmLWfJdJt6Eqf/nXtAFhQg822mkbauuP/H9H31kcDcqzT
zb/4U5tVj7+GT+Vd5xSRtl1pZheAIQlKKXzFoNcpu8RwlRyvHEM05Xqxb2KYsQGGDpfc3qrTHShK
4m+830/42ZtlLxuGf4jneHAVpPqJ+gKxlElfn2oIl1ynvLSTark7nlCWVOcXBo/1CS2OJPpi2+zg
LAf0VmKMlCu8NEJTc/epwO6ZoASnk+xndGlMd3shG3e/T8OOqQ6bShNveodS5i6tfFaOPfpc+yKw
2fQDGC8fpEFw6LPMGrNDpP/yynJi+YN46yRdaks4hk4LSHF619ckeVsmG1fmJ/zuwGI/NslwBo8c
+J229L/i17MlXRIxIWtsmDWZvj+IQfiNHUs+wv6c7UX38wgV857o0iysMUdnOki47bu5ejXwS/dV
AtXYsIovmXdk29JUNO6maEmcwJLO+yyzml5CW+6UsoxW1JUKtxegV/WpgAo+caxXDyQXcuZ95RGq
PPxCErVTNlxv8ew9StOLlEn7Hn0Tlfn/3xfg4bFAy4X92DI06qfqKimR7kadBV87OFAFwamGtPCI
2hfR91uX+oMJHlQCw+VYP1sic0dm8Nw0FsxYbqONkz7Q7oFXAvvDKhHTL3PHopszyfc+xwdHJEko
n6TqVpi9md7KibgFXYYLs27ct61skqdH3XXYFH3mkDaCDCSYKDTmFXt9z6KJ2bZzPHGd88GK+imG
bf5MAy2G1L/YPr/TFmlDcjeQcdkGK3Ar9gqedcCZxrVD2AVpxOPww4Ew2sbqnC/IxMcDi2O/XxaR
PhlKP7dk8qoHlrwalz8EB3ma7wCPbNWyw6JNqlBltuL/Pz872+vHRH2yDScnoH20B4zLydZwxy//
eF/AEWV3lAI4p2aqghL8bztWmr08otXOHnw9+32iVLMWWpAquU0Fce213bCwzjce2ZlHGD6HHsPD
b/nBYBq76GxKoMMNFWoXO9xDqNGDLWUtBRm+KVpZ9/LKRGZUcaUZND70afn1NZMj8WCc3qRNGrvB
v1v+/ZevoZZJvWWsxuCSDWC23OfWK26F5qs1XO2zPkiQ4f0dJKrt0eazThtSsfJRFQhSIpxhzpGi
/AkmjQB16e1rBDzdQYwnMCauv3D4llpxVd75nX5C1X/dd13xvKNK7MeWlw6zoGYbN6tWj1fYlXiF
3pQz/IJzLPR+bTJNV1wDYOwMdObDPQWqjtsSbvSfH2ILpwiCzcq4xnWKksxvYak7ClAkLbiRhS8G
f50V9Kzc7NyYisZ33eMe3JuPsO4gISN8AujiLOnfnK2BVBN070Jlolz2iwBXwovCU1IzARbChY2i
7KsuIhMJAX7Q74bZArDOk7WYvf+noSsMbd3zPMtcYCoV81lh83woDlvzSeeRkCQDiM91aF6KJLL8
Sc5qCfRlE+4617jkSaM6GidcK+jdh5V65LVmEftudvSEolNxk6b1E9/0mhYU0Hvn2XIIWmeNvARm
xST7h+YnynyXCX2/M9agGVa0GKxRppkzLS6bfKUCGazJhK4HrTMeCy4iA7dnV0i3gXzUw8J8mMn+
eXlYcE4M64SYTDYbAmDCxrDlSAlY/QePEj3XdewaFjR8E9RAnoFAbHSW2G7sGlphRpQmMtBA2EBy
CF+GzZffNYUKxHccQRJRbbymB7qIuYKGiyqAaYHn+tDjbkxJdyZqX0rZ6qJJy3djPHO1ZD7mtKpv
e+zX8feLd229OfugWVz5g2oTBi6ZaqLBvOeaPsUU8xS+1DmKVcWGeVRH7EdEZVOYOK06cCJZ0Kvm
fxzmbJtxp+HP6uimsEUYypKyTICyCeDKQngDeGyaKZMWLJkxuv78K8kZMgw4Iu7ZbakBzvkT+0+B
1efnUNVTNE+dqD3AVjUOup7Do+dECxNuphoagZpwFO4r/QmmygTg28OvyIoI66D5F3dgGpYzGToA
6UiQP3cTUNncukpqQnKMC4TGAvTq8TeKcWlaTlnDfawwNiU1jlO2DNJYnsRf481ws/mQWwth8ks+
Kn/2QxqfzRkuqQ0t0q+QKqKqn9o5ht4jiUFSxwr5tE8tH9O36KVk2HPLLWDTBommxa8rLM0KsQm5
LxWW0s0BccGHzIOo+qNEg5wRWkSTA61B1E237dcANdtALR/Hl67MP3R98DbyW16+0YNXIQ+Wj1Jf
xi+67aW1ogCNOcHLit18YMrHyBsSf7tKwmfAFRqC5XkGzcyaqaxhdgPU8NPl5VyyTPmsswnaXWBx
UCQtXmL1dhL39qvr/fsxRg2E/OjMvNbzBwxp/O/zf/hJFbh6xKp6iJt/Q5E2OIyDe+YNa583LHgD
fJJkw++eJ9q1ulaRtv7fsm/IKaqHM8+QyiZQSyyZU6viz8CdHWznQSdzdfRUJchEyv3zLUhAUs8/
YL0cM9BmYFLGKq/MGTY5VPtqxADTFAcUCqOaoHyEGhxR5tm4NUaGoPt0nUZFR5wGcZVlfPpFUdkI
VtOampMxrfl540jIe4YmSSYpiYoldXr/usog+wH9mytMyPCTsUMUc9Pw4eMV/KLM015kv2zMP3Yr
+D+maS38j89AFcchu7XZF1R2YHQgpLqIMu0bxsBulwW52hwp05zs12RHMxlcvM8tsFQbwCaFOMX8
csYFA7S2s3InXUnRlDHG4VTthvqRcSCaOfQXIKg9HMA0sJsWKMpj0Tl+1tqYu83PybqYry4BW57B
HyDea37ptna0+n36EouVM7UStD9p78Y1Ae9X87XhGVp59JfMQQZSHwdioEtxUeHw1jwz0Gg82lmA
4bt0WIXzhGKodgjI9kQA+S+sSqutH4+UaIwi0qzSZ03TihLuxrOJR5k61wqqnhYURQteP4C6VCBq
FjVPt7QVJEEZWLUVB8SnAkxOOGvB8DAYm/EZL8wwzXGHYO2lcy1z7w/d9meH1wv8qTTu2b31LUCc
JFC0wlReoTMA88ZvO6XJ+hqpAnx3lVHwk8DjBtUixP6aZ4s4lPMyfKztYKAN+VbHss1aaR5Mcwhs
/aTGkDPFnoZlXT36U2UxCURJer0+tEnuoIUDLkIgtIOpiLrC9twx7zuD1y5L4wFIeLVge3y9k2Oh
5gzI6E3PdSSF4D0Uj6ePfcR6a3HnM9At5p/tYBTPt7PI37lTdUpRElXnTTIojXbMJHkUTXGTO+Va
v9c1dDj5FTJvma2bmNmkUG7wTDYFVDbE+wD6UCEKGQ65BUrJ23pLJu9Xk9TNOPtPYxCCMgPsafk2
bn9A0y9ZK3slNsukBX5yY8vqSeDBowmGd5vSNdaPKXx6hkvqqFr/O8MjolN+98ZEM9yO6sGeg44Q
14rQoyg6uzaIzPwedlBWX8Z5A3Tdnw10mI8ezLvpVYJT7UrlLfIc8PQvWxHjeI7IRjy9fM2okxSf
YTPow9RJKUQLcaSMPGSu6eMa6Zfz09I7W9L9zyJfkoLSKOnmqAgJAaVbve+nyj8HMFP4NnIgYf5F
AeaKsCMh2Bn/ySNCL3bKQP06wSpZ/4yv+FsKiYcF76ve3UrjuOQLA2CJAv0TVD8zhwdGMPMxuEfo
+M/DX1vEQH1fUyNFtyk6xCxHKPCOAmt5bU/KkwKyS/RN+EKUgIDeg9Jan5/hhETNihlvhDTQI2tC
w0ThQQjCDXrYjbCSr7TCJSSj8PWW2OypbcUKV+rIhziZWjmiQBc1MbrUpWorwdOcBMofYE0Xzh7T
V8rn3DwxrpcdUjhev3S0yI2OBCp4agYkKhjpNuNdrb/JrK4aERhDnpByWQTNM+Ik8tZBL8RSLa+1
/cV4k11dC+TA+fQYOBwGy+NvhjXrkxHvqAb/B3tWCh+x+7POR7AaLkX2KBbPLY/tprJL1lejhprG
QElnaxKskW3+zb35fK2ra5pBg8toB9QpFT8wbZZsXAJZ3gmdJa5uNbdww3qebUuRoGlITyUxvrde
NdD0RmqysT1AfVd4XNXRRUr90agO/evbr7r8zllzZaA/K5h5Gk4t1SQxS6ByRBgCF5uuexMdqljF
Uwnhlk6iuT0F9ZrZEINxdt2pxBCJi2W0bESpZyVdGdXt/ZCBEkeitrMvV+On7HIp+qLcxr6hl1Ca
t5ESJCUV5nIcVgGYcx+WsFPcoQ/1/dgj0lyv8jtaLlgg4vksbRkFiESysheqqZU+eJB6zJsD4BkW
w/lR66Z+nqQyiGpFhqOA5zC0DQdSl/ireL2L84tdW5Rvd86Elw2fwH68b93+XQT8/1ytdrUGJjWa
h1x1yL9DJ6MFJQ==
`pragma protect end_protected
