`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
kT1mLiaaYa+biez+hKMiiXj5YWPeVKgpyEwJvVyQACAItgJ2XSKs5g+gi02JBhwwGtUYHYHAQLw8
BukTy3AUYhXiVxYVqv8aH7QdIu49qwYmkPjFjzol72P42JuY43jozX/7aLzy+p689QQobVlwhrwE
NlNeMFTzLW6EKTt8BSCK31RkPzZ0qNOkA0ACkCMrmpybH8jl8Ac3wp1Rij3mlX3UevDKOK3r4lIz
1QSOpfXVYDg1lSNbQ/yBcNzld9E8DPWG3HxXQFyFv3hIb5a0o9Q9p8oBFfOFaA36q3/0p1kdKiRZ
D8BvpyYbJMdL5gOKkavdasn/fCa8RBV6g5lNdg==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
29J/+rOk0LLKX6hBGV7Ci/2kt+CZtq10UPl8yzg6nAXK4pW3cfQlPufI6q7q/f6QS+gk+ktkZJnC
FPqAu0J5AKS8LNF6qjAmrsuweyx+GxxMmH2zO0+1mGLRoTCYO7u9I6Q5H8fAXds92HREZlHOCiLS
G8uSxxoXCdnorVbqAN0=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
FYC98DdqhTRbPn4asyr0nK3uX+SaLamh2hDfG3we4meoRQBI3/vF0GWrEoNvT4IoorUhA6LtMF4B
XZdhkVs4rDAgboyKvJ1QLM7Os2znz5CXG6iCcR7rpSi1AtILSi9Oj8aGWnedgu2a3KTw/7GThXp8
uIzCbhcVhgaCn6YkyoU=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 704)
`pragma protect data_block
UmLH3/HK6WYYSIyIv56Gu88zENuDCiPW5g1pgDRfZR+BUOdtsiKzB2O7jeHWLiayjkW1pBunOSdG
7R+5Td4FjCNn84VY7PNGycXPSc+27HO52shgfYkNyKouuGCsBgyOBC8HpIeME3l0Ez6lrlT3Bnl3
5JSsp8ya6VwPAYVX0QxtFO0p8zttRbtiEfZnt/gUclFLMMv8oXUwCS1+U0SJu4C4DUiJ+yHKbVIB
r1rbRwkUyYdHvEf8RXsyygWOgngP1lwaXQradcBNAhr2GgucfxOmRqEdSv6RdJE5WE/4tToPrtzI
Y+HF0HjbzSAfYp5zZpFGZ8Axfi+q1B6BF+IiFvrE8g1dcC5Ba8ytGbYg2PIygvk7Q3AJX4bBuVJi
Hf0TvcnXnP13kZM5NBVH3LOmoca+Op2m1DVCAFu7eKGQtT2ooaE2KxNtKIra6+1sm68NuL4db04t
RdLa++uoQW33ZIsweYNU6g5s+u1mog41Ng9KvkfIj8qlY2At9R5PpMwegvArwMMf5eB8JRVfs7/l
nXvRsCEo/enjLBjHBuFOQOHbqbJGhD4VNKjOB9pPEF+sMXeeCXMVu+srvaGwy1OXriI3yLXZvFSd
IX4T5qxQ26vcilLqmbEPM7J/v/pxvga+XNdMIcIoLL7MNa33m/kWljEk62BPmWXSzXR8KWjrZxzX
5/Sz/degeYW92sF1v9OCwwFOp3Q8LkFAqPbBGpnqGci+ezDSta7pupxsawlrOLU7hCmoYPdpQgqY
W6kAv8qcDWeXLpc89HA/iBRA1fBVoIuogVawc1g1QdbG7jdmc4629m3tMYlZxOYkLU1SIaljbQj3
1EI5RmkvqPXCjb+AK3ZzIWQpzIW0sFPuel6GD9sqw8dwa5QOC3tzrrr52OlJs4ertQEkilVRB67k
4bEvMeO8bxj1Cgmxft5nnXY2YWk=
`pragma protect end_protected
