`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
JkhULQwAJyDWP4tjaGP/HqVbj8K4aUJSXBhBzsUCl+7MQ71WyfVpurd6JkzzLxJZEWPuUW6FXvun
Qh6Ke6Kw9hqRYn1gR1lrJAgogFSLwJVY+7WBMdW0OAqoMtLHQMYWvBlNub2+cvqGxhzc+3SrTPOq
/hvMB33T/4m5wUahF8e18wD3GrNM3WIC6h8teCwt1ff8rfasWFFzCKBfgZpEwGVh0cTdRZJkh4Bx
0Ci363v7aEYLM/pa7Qkv5lGmny1ucAQ1wMfwo1ypyYBcgIDfAMhBa8+SVILwDpAvavNFq3y2v/Aj
eKpxUKYbDk+SVcJnFG6IdsZChS6rhSmkZN/Ivg==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
3QN4qN6ji74NuGlJUScWNyyp/3/EQyUr9rVWd84jFCYlf6Dzv4DtuHn6HzZrnp2iF2Ra0e+tpjGA
7IozS4qnEeyDQWt5jJBSp/5+ORst+ZPA2YPtTlMjP9+QDSHiqDsjufSyTw43mWTG+tPg1u3b1Oy0
air28ylNBp7EI9d+OPA=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
VulqiLCnLlNzi/4+Q5h/u50nAaiY5nObim/D2MJzhvglzCZI5A5AzJxX3oIxat4KU+LXUcn2Ha8y
7EBSctkygj1RkuVDb7MxOzFIY/kIXSlQOVeGJHjqEkcq0IZbSmYEp7V2lyRPd821QyhUaCxQj1E3
miJ5wHydK2Cdyp9429o=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2864)
`pragma protect data_block
sWtnIZkqbQa8Af7IoVimOB3Fj3sn5cgdQqmVKthGAIrgy9Ho1MydB8L06VXi5feMg2RJGYUK092L
jWxpaG/5OOsvQBPbG2FXJXD4tqK7OKC/gIdYFBtYaq9h5UHxqeLziPr3/C+XFIEyym/nZgMEUgnK
Jq8gIOfwH78wUUyAbLRzMk9Rguh23sYXFqF/Pu3X5iwudDMLVcY2y+5y/U7wt8uC6rNXFw7WiD/k
DcOATK6Sj6a4GEwcYyzMV3PoqkVUv0kJAkpmGgJxkhXozZlpT2jxK+L3e0mib8E6MzqkrB+64v2O
gEf4Y2Yf0iHnRGPU0ZEzULAJdvGKSNmVqhNPaJqhaf4X5hAb7LdtN1Utjgjsg3Uf8lGFahy19b8u
1+Dt0Fm2lBhpUJAUrKtlBywPRM2MmDa2HNyTeNN4dhbcsb9DH+hckFNtAodaqrywFacELDbk91V8
SUq9x4yRfC8+zOAAOJ53bjjaH0hbBtjCGskOpkCkZR2gGWFqw+Hn3Ox9sOKBihVMnl81WvQNaVxM
SkjbawHLvdsbv54NEycP2Bogb4YnN/3gzFa55pE0+OKmXOMgaiCMP5QcpU4fxdiouuq7aV34fyBK
gKXdzhfLmxlw3hfrxb1lUg9cfHOETL7Xxrow7ycF7yYeqVMRV099TlrJm5YsfpqwgeiLQUBjDRHv
1V3nGbqyin/gSeb+GfCDYMpUW1gc8S2RDRjuAa3Ht4UnIbZHGPFZhC+uTmIUY8+wXK0HeJ/CBawt
6kEtj6zIwNvU5jT44i/DyCPwgsAvudRGAkILJev0/PA49HQicrC7jM2ebsS7natqlIbHpfEKsm9Y
s30evqCShUZaunOXZdzr6hd2BwXC1S5fsL2B3udr+pnL2TyzyWQs2hzWoa0mlI5ri3U5atT5mVKT
TEEoHhdMzpGEselSQv6htGtCYlh9jpEwqTaAn0gRCFBd4Kp5vZTfyWWVnNN78IMMnzXwC5mI56ob
VqPykzhVJeoUBpo4w143AefjVsTMQwWyLw2VrZ4eRW2Toh3wRzSwQpTipev4fm/a4WsMsJUErr6k
mgAbThcBSs7wkXbK2Sfb2p38Mx1pNGOGQB6w0CcFmlYFPqmN0JZOyX74/OAMSwhMZHCioEhNfBpY
YBkvgujJRhtek9kLB8wDqDuXAvWTX+7vLhKNEarCy6ZO/DiBjH/ZeZJ1dTeWe3uDMc1GZNoespop
B8l9FYAQXwgXzw36euE8y4PJ0bzCdudclCPFrWV0+qLh4olPGUbhP6mHoMkHGRztq18zcPELu6WN
Zvdt3DdlD43GF7zwtNaproyPItnDTww+TWBcZCmZxJM+MQXxVQ3PwnfYkUMYtq3oUvy+67XTMfCF
zmeCFe8qGAF3YL2JqwbHwpmMlWXWgOklDcM68XOFk7jULr9URuAdqpmP6Zs9dmRA8sPhfZpECf7N
co4KEiC1G8bcCCaCLPx4I81UyEI6VeFXEAUuWpdTJ0NY0SAiTXJWZWy5C1sTXkneuZ8d6XtGhV4P
N9aX0xboEkmqm8Nf7kKDXLmKSfRQaTm/lr0R/H6Hi7OgZL0Bb7ACHwETZMy3A5w9bsyp8DThOGuL
Pe6mKHXFasDoCKgnUOZpTokL7O5rSjJKnDYhQhtfvLaa6/dcb3w6c3+sXshbgTCjLUJuly9UdqHg
UXz3IFMjqruJnSH4sX3f5c/bf6HACTyVXV3PuEax0ou25wXJjMasvjXYIApiPcAkS0KNr9PY5c2Y
snDGNjCEfAL+eYXzdw/S8NoYH3u+yLIt7c4b91XHjsMg+81BIPU03IExOged+iaKn4zsvS9VtGtQ
+WURIspfx8HPd3X239TbErSmuBjGz1gnMD79XxdlDIpi3Whd1hzoXjlUfbCeDW1cb4zsphwwUuRU
Belr0Z8TbRYaDsk2k6zB17Xb9KSAdHC5TUdDtBHS+SdmuDVwN+o/asHZfp0MqHxicHwLtgOJdyOy
sVekr9Jd8v2fmGbeB0AzFGunEXuNOg+w8K8EAzG6sX698ob9oQEzIKvaRLgzgb+1XcyLqrwkRvV6
/nls2IqS6s0PqFUldiV7oqUfLJdS9xWkv+NNa9ZoR4uFOJ+5qtJ7b077gwVp6OFoDE8PNZAaCcxo
b341WTvH8AhQA0YtwTj2yWnQp5dpC/v9Df1rlgyl17FGhN5lg96qzqW+Yilh0IBg/gEG1n2PpwGV
qboZ+OytPb04vFGEPCRzKED+yOI1ydfcC3LWAP1BmZmDsEfTaAFlarX9xgbaYl/oE3g1X//2/cJI
hEwVmZpt12b2c/F4HhpmMSQzged0cxeHl64uHqdZRHu7pSYQZehG1h+wN7YJ+UJGBWVy9IR65kih
dHSAncb+VjXOMUK3SiTRZYmJewqNdGaKHT+KJ74v4S7Q582iFu31MWFaRUInoPwsOAiwIoMUZZyA
tMP6amBoN9U+fmnayLNCHUAwAeJ91XPMP9ml469cZcN7CXBR3hAl2t3mq59mnLxp1bQ5NnDStopf
ff1T6PjxqTJp2dTjnKoAOEBRa9n53r9IHubwci8Veo6CAE1t4PhZvywsj6slzRy2odj+8i1WZ2AH
YtPRZY1rQLS1qJAh7mRChOGLh/IX6abOmu+D3iKnwt6AxctZSV15MNtljWKlYTRROlHTcmpkBTQ8
4sW1afv6Avvf9pD/lo6DKVApFvCzrYlJxYB+mRzFMrqcgO7YK36yr/ZJzk02R3xVeZsVI9popDGj
1fGg1BNXymvfIRSRuRdr94a+RBzc0A+gqOlHkU5vQMlMDtdX/YjwNXzGca8AvpZTuRIMeisitn5g
R32/hY9U0h29WuFkVHYoLHJ8g7cxH5iLD+T4iASX85KKRxoxPomUtU22JZcYc8j0Nzy2I1f1c3zK
Prk6DlBOTr+U0Kz8N+RDFIGp8re8TrLMQWdqiROazaRnwwemNFIJFYc3giI4dvbPU//owlJUCGe/
WlflblrCNBt4aEDfzYPyI1tse+XZddZaVDKb/eg2qxPN6tsrOvUiEBfdcxZ7qtQuZgyHgYn1MigB
siYMgW0btCHTcJPqaVtLrfn2fwmRE4JTsGa2n3a71yZ9wF8TLtnDDTzsTvRyu7nRyfVMhRV5xaHE
VWvc5WAKVa59r3FrNIEcYSiJy3j9gVbEPUytTWlxt1XcEn6sPjxtuX7TIhXfp8HiubPBse3PrWoO
syzVGwGPSCqNjv5JU6/NxjHlTouToSkNlqGCxiih7MbsGtAhIjPFCg0xp0seQmWUaZOcXVErl8LR
kAA8KgqLT2E8o+gNNLMI0gXfBOEhHNq0dc0Nk6M0lQWNh+P3uPpbdnucSbDKf0R2IxwZQ0Cg5zmw
uRoIi8dZgBMyoVV87XV6sEz79LN1tdkOXmyVxGG0Sov1T9uTtQ68Uuyvc3TjXrW67+xhzhuzrsz7
5QArsvplcVcuZ1VXcHMArlMsD2MmbfYk+JDNbI2QdAeZbH9ChjVv51FKKhFQxvn93ks36I1Z1TDJ
cBFAti5oA4ITp5zU7KpF5sirO5+qX1wDRlSiEq3n8NDRt+DjhTRkoWhKGuOvs5Hbg0NkHVVndVjE
CBJyTNVEl24MMvEHkiqZAGkX5p/G9Sgel5sngEsKTOhC/tAVY267JtKy6Ux0+G0s7mdnRvrmTQib
7ERQFcSlBR7COibIyE0IKyIi5Kvz+cRRYVU+qWjiBWVL6SEmd+K8FVfqJVLuzYW13p+v+ytIc3Oc
ofWpdLEfLWcoyFCoxafGHErMAux7nFsWhDOkJAa3c8qFIX/PLXMeLkC2JQ+ofDdGgEQfXK3mTHTY
btNU7fe9s3T1pxl3OCg=
`pragma protect end_protected
