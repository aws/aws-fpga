`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
epMxLuG1uJpu+SIOqdfJPkO3Qhngu9wd9jnMw0iJQ7Rt9jY35f8p+MAAouLh2RbIVn2cUUhoNqiD
D2QgsZbd4Cp0jbDRu8vAvcYvv8MFBkOEXBuu7FaKJpOdPvVGS5nHyPT1B0rWwXEs5zJgckKZr0xl
bZzQE8j/eCC0UChehlRbB57nneKDSMVkcOFvtkPhs0F0zhAesH2ntHwnn3vDlvBgYNPCkMczqzCh
7gM0WeTgIKjkQFjuq2bZ1yfs+WJgCetR6u3Jy58k9Lp0+scqwzLPKQqBIws+GjhfxVbtL4gZvFrU
uTJJhSSMZcz1gyj6ACkucJBIZC9OPR4syjLXTA==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
0UBGELifSf1jckay6Wtn7tbr2knWdgcPCs5iVXQwkUxoaGjHDe4FLxk8csixUaAGMQV0w9J9VqNp
UA7VHHsQ+FuuX6mu5JN/hvjNINKYsdUDGx32+TSZ8CbEH1QaKPtiGwddtmEZ5axobXOcNYIFkEjG
l32bikZljvUlHm518Uo=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
FzUKbuUaS47yMFXsJ+abOrG9X1+z6+0tmGKiFj23kw//zVeTRalcHGyZ3XPRSDaprpQC8dwV2n4Q
z8xN90Kb6zw1PAlisxqlXX8Uj0FU2wgKdxaOKXrjeRCKKFc67+rebTHmn6Dp9PT8MTZ2ihye1487
cwery/FGXzqKDuJBf0Q=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2672)
`pragma protect data_block
7P4dDkaLGkyX+eoCAVSWrzXyj5BqNg3nQcT+FD8HoVdKf+UlV5Prye0YcbtheyW9jxT2oLLExqej
eeqhVNMHKcK7UTc+bJRZfBHYBUEEPROEMYv6lcRMdqjS1h5VoJgLGml6aft8FCwJSIuuQ8Bx9xmX
ap5s02nH4hhpkSU8JxYrLDF/sT9cwcHHkLHbsYDg+eEOIZ0+TZDt03Ko6MdVKF1eAd3BJ9QMOVsF
Ga/8n8ldP+u0aR+U0G5COOVsSrtBQTm2JOI55Gub9OQZ/pbtaOgN/+sPmpgznCI8d4gzu7/3Rzj7
Rj5eToiMd1zmCgP5ckyehpM+htnCCpND7PuUMVOD01yeIIGUMpcP5+NDe1Zp42aVC4Bir80xy663
a4oXdZVhKSDW2cJr57VqXTKVCkeIA7zjRosI06G0du5lMBKIAnPHyM5pMJDUiAFeDOyCS2dtd2Wd
7LwDpls09EkjxbGpRr2VbO4un61ZTchUnh8teNd75Plr44N60s+OY/bbwMJ0WR43ENGJbwToLhbN
8lSBqVtQoIzCiPBFRSqBqmJ/Z7AF1dvegs46p9M5BOYMuPUgPw1dCGdFJGGnpf3bYzFzQbcMQOa2
DGVJH5BsH9QEQb2s6yrjhIHMj1japB4XUWyPwnzEDUfUl9RrEp3XK4KAbbFM34vdPGuD7sfE9dCP
CfAjiIBUpO1zvjLVt7yRfeEPrYaAhvSIoMrchc4MqS0kY4sJkZzxeMf9N/EzsGKXwMkYoMnCx3dB
MKeTSgxWVG+zzIiF/TURB0QcSSBwqo6nAD4r+vgamovqdVNzf+YErQFOxsJ50uo69jUHrM2/OgIY
UZj1Opxjl4ydDl3aWcJ17rstSzerPDEgS0NgRA8WIQHLGH/Mh17bM4FNTZEV4e6DuNPaK/LruAcv
Nzz6ZcN0EOcazjdD5uV9Z6JEfnpr1fHiNzsgJajYEIWaQujVEs2oSZME94hUXq2A9tFlXhcMfSI6
cZn5GefA/pAr3eZmNTBdhVTno/Y6WsJGewnQH1PFhKmteMyC5e4jZfgOV2IAHxvVCgeB7P+qr+XG
2NSs1NVq7Ws+e7+bb3CBGWAPVniy2okrfaVnIGy+ZMgMFx8P6ts6LEIiHJw51PTCh1nWRYSkTBvx
2o5BL6Lm1bd3haXS8UWQYTyzhz1GTeB5RRiIrDcDhOETTNAVXEqOpOIrtVKb+We04iR0kerTrqmD
aQ7yszIVc/p+X20z+QASR7q26gR/AhHxgbvVPIZzhxEiXIqpaEyZIg4cAh1MdHwVTBcM5nOmyweK
y0hmPd3Zqx8DMGJDsDMxc3MDLdVnLIOUN2vUJM1mkd1Dd82JnPyBb7dgY1cmb3uT/+WU/dxh5OLT
ObqPleeaRjey1tzswDlYhBcOdco0TSqZIhyK7hITF/cg48LBbVDqI29jUNzukwHNM2WTIOCMrIqg
McdgpW7wZjEPMenfRKR12YDvMLbrlxUCAk9W/vHMUA/nFmlPG7JuDVeTDqlMd5YRfd9E+cXPj3Ga
O44qpRYTUC1D8D49tUlaopeZ3Z+ixdpnr3wy0DsIMOSqNeoa05CgnVWemuzoKd1+f9FUoLt8/NcT
iHkX3ePU3z5jt/uUMCGiG9tdq6yHD5vCe6+pfaHXHHh+PxIjol5coLd4TmuE7pylByhTJqFlRcAc
K7eVCwPqc0K9hbwWE6bg6W+ojqGJBXaMfZhxfkCvTdMy2wfTAnj1iXp3ASKLzMyS3gwUiJhmsIZP
AXN6u92uxJvPzV0MXfvG5TT/BoJIvkkNvQRIpeG1wKSd3BXsbGad1Yk0qVfL9yULJLtC//oV3F5f
q81UVMOXFO9Sm41vTcsEw8EHlLD6dAT5Tk938K3xS1szg3ZZf6zbuFIKII93aq4aJGVfLNOgmHXA
MKUIcKz6KduFbPBPyUdQt7O3OjiKFm2u7iObsZDiDnHs/DemaGyIYgMktTE7J14cKGBExmffenOU
36FnvYhDe8L++4g0ZrIa8Lo7o3f16OqHN26lS1A7cSaJh7hJguswJx/+T7Rg8UAXcGiOX6vHvpCm
ZBO47h+b5yJIKMN6T5ND+7pif2HKPVc1yrnKPoN79L4QZ6zRydWOFKHPMwylwgSpvvXquCfC1uD6
wDmKaieT0bRP2gmcQDYR7AB2Rxh7rXKBy76C3YFFTCnhnOgoT++4UV8YHe5XeAHqArli2y/A43Gs
IxQ7lUxk15u3UiZg8LAhnsmwyP93NEZgkMDsEMitiWkl9zZrtRa/GMmRAB4uGFHS0B40h4eCoY7r
RzMVYHeYtJAxekNfgWirzdvqETUNjij3ou7XHGV4qWCjMzM6rbiDk7wwedu6O9SZNvbMXGFD3efq
g6pb3M1lLwJqj5sSgl3BSFXFjiNZhmUXEJQuJECCz/JwgWUZrD3VcwQ6BUKPKNmq19fer/AoZtqn
jIetcNs2nMtynM0zafJ9OvrPqggO1B/9CMxJWNY/5aJ+a0Qrh0Qpotmv0jEn2HqFbqUAvKujOnJ8
4XBj7A5/ehVUPtWblux6cDaHvYEfpvnEmOLJ4Q7M7T3cdcp+EUOsDYzSLsLctEhPVVjcEP2g5eAz
nl84k0Clm5efJAPsJDfp8aWoEK4+qWjR3Oz4MuGOJ+mYTwBS3uMqs/3ggR/JohkKY403F9d4/tFQ
n3EwALSJv+/jqBCk7plwOjohj9yO0kia+pX3HBbVgSPhfmJnkmRKKeyIVvniMe1qpxhNZXa2SQB6
4k9xK5rS+tJ3HlcolQBDFvB/MfPzBvdT2e0F1556KZ+ikvVkJUNoBduQ4UHAS3c4gc2ZNl1iaGpD
qPWXgS2zH15PYS0pHAKuzAhr/IRO3m1OMDbX28SHXwsXhmtz0qrDrzODBx1U2V5Bgvn3ZQ+4fMq8
Z+OVezinNEcAAJwuaMNfaHrmbSQLm9/p3MIyBauC6enX7fxTeFODTKGnsWv1YSEZ7/LWq0X5CRbM
2UpY6Jx1hFqSsyMapxL2UYT/L66Qz+gX0RyrtFeGkFN37hJ0cD7cGbw6hvEwW/tQPJRgUmH+z4lI
Xny2HqEzTzjzuHFwXf2/EIm9w9qnxUby2mRAWtkFmW5eZLPKm4lOnKekfSnmRO83Q65n0quQdlQ2
wZaR2v27i9E9TD2VlU05VtMZoxO4hZdQc0Z3WVDizSdSt2v9Ii6tDxKJtuxoQq708NxEEIU1nCZF
lRk4yQG11Ws/3dLYfw4gmYlGyk82MuzqH11Pkgcw5FmWRdLWGrnYOWPfkuXhMwA0Mjd3QGBkeD4u
9YM7HjSGHW9T4TGwLyMq+lFSk58a0XQ0tEAzZnnzMXFV58vMgxDmPkYrHQyjfxQ9ITlMDeQ6hJRC
oIEWiMXKH7rnFPF1NEe/OQDqTR31UtqmQBoAoL4bc7+5gED4GkARTqkBMuPV1zp5/KCZ1QOP98j9
kdtihIEt9OE4nbhNpEGwV3YsYazNvXW1OF4dz5fghe/639D7x7IbIjzRWNhqRLzwMC26lJMKLDW5
0PVTvBrykCh/RNJXd538/Cel7VdELZQWxo2SAUO1OtYwOTmbQecmls+mKEQrvOnjRJE=
`pragma protect end_protected
