`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
MGNOQArww6NbqkmW3Az+ZSDFeuwokjBjCBxM47PR533SoeSDMAYJQkJC+0B5yRCZ+Ex++g+daE9n
NtNn3MfqzjvZfBQMUlTMDqOLqiyxLZyfenYGsz9pOYjuuteY0/BbEgkPPhSUKrqsQrRPNEkCSi5R
p4OxGxnA5GntCfqxGFtMiFfDjDDRfWVVveEpcY4acR02WjeeuEfKuaqYGKVjrRFp6i3TW00ZEb9F
oDIGnvNnywNm7dxT7pjD45QXJ0vfJT0clUj6CvOzN3Mhp6Mk4D7DZagshOdAQpcV/MBNToOT+tVa
e9HpMTY8ASE8Dd6Rq2lI4++Nit3l/NF5ZQzXbA==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
mNwtFtv+7iW3OIA1qgG42yU7XN4zGt7FzZBJ1J09RNQEODXPydP5I1KTpE+LGNf/Nxfo/WXA6IoS
7YjygSfnxr9byh6QhLg96l0SU9F7vpqXbWXkzjvBaqn+d8Oicq6vtin8grUf49wFusl3RTjUc1B/
SSI5bK2k+G8xIuxZyV0=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
CtStOiDbq0TlHUzSoEzQXKUhHQ4Yor61J6X+wH0UWmaxGEIH00VnC50XXyCO09FOCKls4mKpBVye
BzOkrepmNgZnRu373xR1tswZ2zBEKQuevYWWcy9i+42cCEnUYR4/JMef5zIPCGnlTGn/fiQU9ZWO
ejPE0QNjOaBTcg2kaig=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3024)
`pragma protect data_block
lXtICizulJ6NGBadrs00ghkww2U8oIDBXsLERFNPJsu9w/dqDxxR89kUsPOaL65qcFk/Q7lTF2PF
LU0hVVubuPu23wDszDbiplSUvWqd3xnMmXQTLOZLt+Nqv459oq++9R5LLN0V0mHB4a0XNitT5hXx
XEQNDIfe1/EVhR4Qxw7e6yxpXE7YNuNtIWNDwIlQO2ybe7OPOifV+X/9BTj0y53Hr70X5QSGqkx3
xWyrq5baDuFsj+7xto4eJFS+2u5TJF+Lgg1r6DUamBfM1fcpNZ8nA7+IP4xZ2JXyWq4BKMgqIMrL
tByhrDC20B95nt5sE2c+++jxtr1oCVIJ5q4uIN0tIrZFgYnRN0DaOrc4soFupOm6iVpP/tnCAdDa
XTZw/nKOl5C/lYdsSdciElmYoiCTrPPPvMapkwZdCCO4inM8UiHr6ToxeyGCPbXlaZH2oI6fTTun
hgJH0CGUaJi6Efn+5W4+YGbPDsYUoiVvUb9zEFHE4mmwH8XgMu5C1bzp/3i/4UMEzhILwKjucTlv
pLdvTcmQrzYKl8ifvEmLdRuDpZOHGC2IywEAmmbXXAMJMBU0sKXP8WCy0JSTFZwVPeAOQPhYrzOp
19ClxkfU/DPuW9y5/5F7SpPpK2CLpW3uijrpBfE0Ij5JwpJ2bfeIw9nwzJ/qdRWG+6HOd37XWXRm
v1TtrHGxHqC/NbG1L45V9gvp9eLAayQnqx3fK2f1FviSgvXQjRATEM8GzKHg6aF9VzX/fdkNJ/5F
yUTentACTQTgNpee6l12B5GZf8eIZca4SRJpeGAfXIyZZVmONgjjF7rngpjxPvZ9z1+sJwlbDZd+
OzohYsu6D7890JxmRbplGMzgHbgJZn98VipY8t/+yf4cWcLCAMMbkCiJaUk3PuwS1+rNMp5wieWd
3wGaFDJqt5BoEeZRaOLDbCPcC3iQKcTXwqHg1MD3ynDP2sIZFBmhwZfqefofStOjSzJ16qv+WoqM
FMMYY6xpvn7PCMoYEmQkN5OnNe/3PhYP1Gjdsyxm+x7V5PVD5Yn4iGcM4MLCCF8Cx2QClOcWxRFB
pnizJp9AgMDvQ3nG8e8LlRVwIS0FQGxMB2o8KR1xyLMQ4DmC4N6l9qao4V6hRw3VhXYoBcPIp9TM
jJ43PsC3VWL1tyOv5f1dpSh7SnF/Q9Rf7twf6GsbRG1MwK5nJ59Br4NFlw2nhki2kzM+oM/ne76e
+JP2OiSQr7PqnKQu15RevA4vycc5voupJTsLBOBgcAjWur8podzrSJEWLSyS/vDHkYLzXVVZyj6N
4HUJdQn1WcFYA6KlHzoVbuGjv1JwXsDPtJAlw3AlDDtbvv9fd182y/kPF0OQY34vIZkVASHTxRHu
u20dSp66iCkn01/BLdPGOT8B+7JENPeD56Vl7TVxLz1/5A6UNoxjjRr4UlR1r35ZMcF07rnlGvxd
N7xMdoBN93j8iez43n6b5z/ihU2YGgv32yT/BKlBwxGJX+oLNRbYTrlwsrtM2yTva5jLM4UwBT9d
QrTrcmrw7Yvd8p8Tz9hwinLfFVELU2/soANFotg52zK2mkPA/voiBuItWCx8uiVkU/Khjz8AY33Y
jjVuCuVlaw2JaV2bYLGcRDWHWbgqJsppBlE3qKOOS6aPWLCzhw1b0saVCeF3D2gYjbPWrVcQjiIL
WuO8ib3fFXUVkn2leG85pbaE1kd/T7U/Q1EWHf7CUpZwwnb8qw5wIYNmRH2UwW/vSyxYIzdPLzPc
B8ZrZMIeRUWYfwyjUBca7M/jccadsOpc0VXEDKMnCIiFSjaFsZpUWg8tTZzZfIhuUyGcyjd8oQQa
PvvPCWpexB0CZbKZa0jm7q87MouFIGfTpzVPJ6O1n2AVRo9ch0xjDaCdnGIHv/jnyZ0LDu7xgWny
1KvqMUv0esh/UhBogt/R4s9+N6A2c/P05r8aN4jUB/1sYiDOZlJm/RNIs6MYbKIenzsOMq09m+j3
rSy9esJi888bkn8fg8zHvIuqmOUF6321272/Xafl+FerPSfCTrl2gatI3cnV61cgfZoK07LJzAkF
Uqkfr6ANlabeBodT3YfiQJ6LyUSzTWc4tv4bj4sZzE/EIRSRJq0NQW77zowaQtQRDn1Ga3aO7tkS
mTVzyl5uTABx7YZsYxXe7vrOCmmLgJrL4rDzRVN1iNRoJDqJ3bJo2lanWhzfnRwDG+7JQ0M/rSsb
7q9gyVqNgEpKKfSZTnZMiqkro/k0PXfVvB9NI10syePG4zTJouG92+89z6XH/dvXDRZJehIn6qAJ
Cz8uZtsH38PwjCS/Nwh0UuuOhMJC+7n0SoioHihLETNTBGPo3x5SdFIz4KdwPK6+L5mlCLET2rWQ
PCRJmlhLc0l6Gy+1AnWomWr1cJvdUn+uJKL/RlkUPqsb/xuVmWh1XDzsu78XEXiTjcwOTZFgXarP
4yzW+88n8du8mtocNLMfAjPFySQk+Va2qClb/AiPbpkIZADCuEZ8GXt4sslb/qppojHXJ67uzRcW
mKee3iF7Pzv0wCMFjIPyPAP/KdFX7V9pRroCRbm8JmUpw2uEVy4FCGOd3ge29c8OpPKAHikufCVo
tXAqmQdqVjNQvH8N3mr/Z2OQHC5zWAqzcM1dtQe8B4YYN9q0njNaYT4B3QBegR8wO9tKueexRzCq
/B6db21OkIGAWwbqdQF9e7VuoB0/5XdBkH71gyvpVlb6Ip6gqXH1/Z6zMVByEUz3D0LSrTDf0P35
3ZcsCp/3Oqju7LUNtPt7a3OW+QnroHAoeJK2MFGOwKcEzggpXZ44zGCXzmuOj5i97ak7XMee6yNi
l2rrLBc6ZvZ1gy303ovK/m4zu3kfyf8jeJStLivEre+dP23YWrabiyUKpUGSmvkNCNvFssN3cjiA
xerKMmtq4MCr+u6GrrkdLDbZdBFXjWs3DtVZo/dAnv90k9W270XM2fNfsRqwY9R0G2kNdjlgtfD2
+rEBydf4ueBlqhAgkNsE+8r20IVL+lONqGJQ1wGbMv7WrIeQdcjuBOn0sfwW31iegX0fdkK4HErg
IVjkRi4VNEebcKCDBFuuEyGk/qGCNcHE5i2LbrabfKbtshptKhoE+Ugr6zKotxn0RHhHtgHBR+BA
Z4sJZkiWk7dlcug4a70aAR1bhqbxdFm7LbneadaMuOym3FJ1f95vpkS10oBPe6vNvgsAY0PwZ4Aj
rw7SKzJO2JYkknrnwK7PBBHvwXggfaklz8UEA1cxsSGOkHfitqSAX8r6FA6bOpyA06yPmCP7o4Au
V5IneLXojd+/n7HFM79dQo3n18vhZtm2u3t8SK/69GCQvIgUXdqaTpzAnaM8Sbc+kVPkELvyllYY
DHYqUPlDlHLw8ctNKhx9hYD6+3uGsS5M0+I7o+CwOyaTOE2T2vZ+TohF6JzcWgPgUgJLlyFWlT8a
ic+n7To4CzvPiN6q8eOD+v+h39ZQJaffU75BnAuzp9Vst/GOeD2bD9IJCdqYHLs81U9i4YZ2vPrY
17bV23/hK9rWXmLs+ZwEdhJyBxEX4FqZu/YV/MA83jsDJBh2f2c8NE386yKkh8aYsXIVcr69C6EI
WbeEdS7DlVBUDBk9PpjmmtRSB6WaCs+I09bfoe9ODFa2IIg9Hzd6S9WUyVeWd9sKZWUBOK07FtOn
KWMdLSTc7VL2ri5Zz89ChzFKzCY6yqCT/JWnRSHTyR2BnQxyUnjP7TUqS0yYDK4GDK8I9uM95j53
5R9Isx0meVGqfZmlPO6dBDFua+jYb7aBF0933+xPLxQA6lmY43lny4unVWv8qjAGRVcK8NbnMkqS
cUX2P1sokPkaWIY7HAqgxdWWu0m3mCYbwP1lXqkVp6aG1XO5IFW9tgGcuMwju349dURbUEYoOC5c
ZbE/qjddt1TxFFZWSXEWGN6cEEKJPedTHOnO8u1WpissKWbjlUs2F8xWRlM100SUoKpVfot0gsPA
JdOw6DbYQKqBOShrdTa/P8Rj85x8gUAHuToXpqGWbORZKIUjeVPBF1AEgSoswWeaCf5jTL8JoDUS
9gJN
`pragma protect end_protected
