`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
rEqUBqdNJwQ7a47zwrxfaS/3+QVITf9KOJeVQ4XaRIWXnJt9yO54clQMHR/tZUm/b3D3Um/k576l
gLW1D4bIL97kxcuQwcVdozFH2koq61lG88pmotKcBHRmVBx/FMskxGjf2va6uenG95785X06ncX3
y6zrspvZ8VXYHsx/lgpKLf6xQjm9T0iutyn4cvKIXYBGPWDDSpvgkMr2xKxfP/JtVxr0WHnjBPnM
UTnGDPg18QabVDHBkBcbWw+b9FqNEhONburu/bf377xUKqFBYK83FZ9Az2lThvfU9G2gzmpjmud7
PEyIooukXMxce7atrVMmwjOJxUgGkx7WqqwvkA==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
rBcWlPV4p7AZFGRP5H+SoMxPJ/OxajTLiwlaM3w85FXlLIIwglNxOn2zBsIQZY5QzAx19CxPJ4GQ
Yp474UWD+fXHMF4lZ3+2xZ2ZhCX5C52vYHt2TSVet3KK9vqUIQ97IESzdoZZ+ttD8G0xSIa8IM6+
CZw+XCv8htNKqk0jvVw=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
n7p6wKX+UXCUMGXFyssIFqtsX/hhA9lCePNYrznXYAQFCESiPxQgVM2NYavAsxeY5vFhFCrUrvHq
v/AzYOXvZG8XfM8PglD8Q5yzNeSUn2chi6eS91TpQzy9GzraPhqXuRfobwwaaywwMEMpkHxpJELA
KO7Y5T2/dB16cdvnGu8=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6880)
`pragma protect data_block
y0NuULivEGGOwnP78aYOLKikE3y6tXqHoq11jj1g8uo1PU3/wXz0vD0AaTiU1h3GLEdcPvqtuBdL
VufBJuG8rVRzPeRb4egIIcmQ3k3hI7WqUs8ibIxavTiHpyVhDt0vmCAbcVAw5p2snff/VKvlZjJA
94IdzqAu62rgMku+QyoMGK372hszE2EKTHLzWGigP750YuWRdFzNvu/fruCCDYFOgVjt4KPFy5Jw
c6x5VcL8bAU0OfgXGHLqQZvuK6Dli/z1sNZTEryIkZ65Gv0PI3N0O1xHPlKs/M/zd86RTDSdgCSP
wphQbIjr1sUwV29U5syOM7vummKA+ewbyhLSFemSVXi0fE9C4zwHTUrmUVuZw++G5jN6oRGsDcLH
01cAMv5ZvubSEa76DPbohBMakem/HJkS6N0ZBNdZAzEaH89ykh0GCVoNxYGequcPTwspEgTNNkow
8sw6kr/bFFjXmC0h9JUU9scVw4AJfCJpERue9jFvVT1hrkFisOuBIOrZu62fzbw6C1XI5Zh0j3dh
eAwmf/NVU589Js8D1Zq3EfNeoYz6HQ0OcyxujESJpARJTkOwe9BtInUg85ozYGDxfsiUi444XN03
NdmpYuc5jbOUdacfDkDEW5YicyEr1dCq4UaFzQ4dvfv7RGmduG71wT2UfZLjc0eiZ68niQht4fTF
OTuxzGNVuUgb5wFU25pvtaewIrtuaTsakXXpNf2bLfkDpqVnFlZuVuF7A5G+Gl3TgnioUMKPYG1b
JC6lD7KAzWXrW34KtmXPYR8bBLIZpoW3fwYDQAg8TLvRwpxBHc7r0ZP71dhv43SCxahS91XG8jY/
IIE3RJAhXGPigTosI4qAM47ue9PZ7ydvBtcy1JBtERFJmmnt9NsUmP0Dr9VKtHMIkWLihN8gFuNh
/vCMIvEfQdmuQTRIliT4HsPrjzsuInPJc3CwuHNhH3tnlvM/ZeucyrwEC6S+IJP+cSFs8d0xBuer
O7t8Rg1QoFmDcCMSe1tQK8+vPg8XJgdrBI0QEW6imwssvnqKgq3Y57o+Rxg6oNvIP4Df2JOAUssR
QJn+hSsvVEEuaQwhFYSUcXcQlIfDBKF1rOgpf+8NEl8ZXM4JuhkG0D1K2KE94A6GDmWJY/varHQh
FgsAtdJFChHF3hAVhH9v4Ez1QmAAwc1F4t1MyHJCBjN6+3UwtSEWda7IR+Pe73c/agmBa7Se9XGF
oRzGkthA8SZqNsqRyJkvZ8XV3cdmlDFDa9LKtbJskvhWiVhfa1FmMSoVwWFrW7Ofzx2DcM4AB5Rq
hF427e8fqlaxGSJ022KjDrwhXah9U4jwkN/X6bzhZVdmKW1CP/I8YlAFk09i90AfReIpbmXfu6v/
dS/+OnbATsGBkGUBg5RckiJi7q7sbL1fdkGt0qG+Xuy2FrCdoOQh9v4kgVvBXU5DpPxj8o6UdA/2
DEMlFkij/i7Gt+s8zfgswjgVRg5BRm2SeBuIx2UlW7l667S8yguRSpEghuIXKUaaw/2ifSlJGTm+
UBluFOAuSZ63hrsYaKq//pTepKCJekaGWCY0WjnzQEu++vJrohvDCjjcjhmRS91wURmC3dF40sAn
HyvAZZfdq8Q7IYdxdCWTNlbA5MjQqJHZeaytKNcMi5a3tHrtAhVZtn2YI172pdmOZ6MVGWXi0GiI
KN+raT8X+mR7GzdY8MIMR6/ikgb/Br1WBNzbqcEfQihu7SBrf5FHfDF0ZEOEApf526MwyZEIcWM/
rlwaRdOGbAOwsBCXic01/LcM6Rram0qAa6KZmCe1bi8VvAl1W+tM2zrlgvDSTfTrSQUbrlhxVrW+
bcfa0Z8gOgW5aCXbdwTiilcYdJhIWnw/wNY3AMi7l9G9bWCWFl1F9NpKHq+sJHVBTym7LJ5eJU77
JqafWAusqyoiYH+NfUY9ki5BX1WuOOcPFcogkwY13QQy5fRYxwjbSGcIf8vnkz+tJbEC06ZAyjmS
2L/UjyYarpVxPMWOMMWlr9+QEbnfhMqMQjKULmYSAG6PIaDo8eTO8uwDw79WkpXwf0WZRpc6S6jT
GC0XPAIo2925mJg922agTdqP0FFi4HzBAgS0zMFB7VoToO15hT916xbbLmf9wa8f+dISYw0UeHfm
9x3b/2v78rZlRrHDsji8Y6cZiT6vuNHVEdL6Gc9DVFIzCNI8EIevB4ZCprmBRpWx4M2PcmhCkiBG
sKM7/oJhR5beeYE+u6/Q6wBxF/dVmlojcI8jVNge8dX0Vp+MCOzqh/GzYd6id2Chz0Xl4z93Ud4g
8ZGwdO85VYGiZWTzAKBpU7bCa5a96CsK2IitxKhGrw7bw6Z2hPmlznnOhJsdo/5cVAiJtdkdzkfR
ZKkYFIer0X0NWok85rXbeOWLKS7jdc5t7/Ye/hHdijsi/WIMWS+fHjSlzgNohmHUokYZD8GoXsbf
WiywlYG9RH9dIH0mUytqTstGt6Oa2+t8oqttjuFAKCf08ikFHUkFNEUxR9pY/P67ibOooko8VjVP
fo3OSPl86chIkJKoVQajnV892/JhrHaL04KnoXrZT2WU9MKorsP3L+k7rigyGIvoM1v0Lk0EZBS8
y66Dc8BuoaHVO5jOBvNSYhCP8tKJ+fTfQi7jDWJtxnmdXYHALfEdoc+RrTppVei47Xltv53DC5yu
FPsbWN2ercxya6Z3DTXZwuap5C1s8GzmfSGqJl00oL39RIED85D135cDP/9TtRSBOZL7ureMoCz+
IvlwoPkmssmDmPrGS3B6AnPzRXR5mtYrZy1WL3BBIzM7CWJe8H8RELzqvC/Ndu5bMbBTka/YpMfX
eOWzIGo5G66dU2KiExXimC9urSMH/RxBt3nXauDt13rL8aDfDWhT4cG4P9APA7+wIRH1318AsEU9
orpMNp2ARXf3MZJrBMIDKU2sbV4QR+ho4c8izMviv+bpf/NSQ7/ilBN0/WlB7mahCP/L7dOiigbB
365cp/LZnTMq0aMKaHac9DTMIMRVpnEVw6le0an/mB3ZGH2tkAkCjGF0ekqAXV2ipJG9H9zvUPiq
0R4O/w13ZfYp/hldr0WH6NWDVgwKKKaYA6rg5QCnl+2G0QkW0k00kBwHmJV5XyUOhlbaIxAX36Q5
lVC39BFft2WTfERYzcKfxzCDU3Hzknnl15cYDuJNioq0q6iOiaTM3JTQ0Wk2GiBFVT6CyEc4y9an
5Y7iboFoD50few/PURrQiQR4rJ79DmsmqQ6FjKizJxjb7jGT9SOvVgDZlcnvznGgeRla4DrXOLGD
cVYNp0VKYo5cRLtpO/WD8cG87myey+8+6VPhjsQpB102BFLESo4VP6JVCZlrSJzqzeeeaVav9Bxh
DqM7Y9GEn8iLMlFBHUkAUpc8rtLmFiSKijuyu3OxvSdw0bQOdod4KJm43I44zGqj/WDF/7++ccUt
D8lQkWT5fHKrKG556Dji42Xj2lR7JgcFwRRw+CsxiPjbAXzuSCn4Q2+YhnlhZQJM3cxOrSLFqF/P
kXRqAae9/y4XtJDCv3m7ynlv+3gWtzi3fy2gV2c1qWofrUFPH90QV6fIJgMMWwqqfVe6XztGEiX+
Oe8bISblDspaFbMyUcPoNtB6T1dGZyvkrthOjbGjFVK3CAtY87DNLM9f9KpvfFlSDgVPTRspeH77
KqlshCyMZR6atY2fVewyOS5iZ4Ioq9i1Bqml33hOJUrqHxbMCLs0hY4nduB2Ql2gM8SWXrjMyrqR
YHNTt59CtLHEeUO0SyekSy97B6X6gD4nP87DnEbi07uI3L96V5EG38WVCROPjg0tucEwiAy2hUTn
AVfKOapPhuBdCSpu9kdOrUfgip+JBUEj+Z6y7wzjLl41PrjGnSII2FEc86+Mj2tKpMq1zqXqwONK
DXYLrCt4aNNkrM7Zd2Tgmzbvc4tp8aMBII7BwFRFEQu1PuirmePl0y5y20eNlGswBsebUfSOWEnb
3Hi8Z3ZX93juKhVrp56/CmfB9Ieiq2WbS2gjD0yTHg7Z+3+CMGC5VyIbkgMDf/3a/bDOrhfX4IHA
344ikWARxceuRHatTPwELh6EcAt7DlsXhB9z12t2wryVAdvUDHNUEDcXqZNRyQpIO1lVvACXLZQy
7xptg8BLhoKU2+g7gswjyt6kiZs0k9aTwuGFJVOaEse1yPPjMsu4opw6w3ebrN2eCjmwYUld1Zvz
pg49EmSokGGeAONZcdCTMjA+N6uLYDHgnPO7mgAweHs57w2+6cnFxU3ll/1aWPQc/swERTyUH+K0
4kZnORXZLX50jLJFBK8WuBJ7lYMD5NdgJyjrX167GF8MpB+WnVDSmJq5ZwmoeALhuZK6ciK1A6Xy
qTyb/3PmLOsT001a8p8nLLrnyUedI/I9M6dHB6eXu1EMPDV8BWBFOlVhJq7IjXD6kbIK0xPnLziR
D9aTzN8RLK8GA6UTmeV6+8yOJ1UuXb1iSYKrH/9z24n7J+BjudgXbaTo1aVBfXgc1FzgdKZbYRdU
pYJ5xsCGQ25dgQW/Wq8R6zQ0m7HUmf9yQJRk7JWmoLrlQmnfFtufKxWjkd5jEu6DukiffBOQY1mC
v6kmYKSBzNgUx22rIU0ULBLESc0xRSM7V/VoqbyvMT3oM1/aUElQaMgXo8FL4COvhLWq+VwcC9gY
/UTEFgSCLUi2T6XBrwUskLGp5qHHeiiWuEwqAEjwTEHU6b3a77XQ+y62rH317VFhWzTVA3CkTTZi
gj7w7CdLH/S4s/KSSJ40nO0ilED9VQIwnFCSiq1j8LMz8QDYL+qvpQJ90DfTdTlmsJXlMzdfk5od
mbSa59JB/Rs/Cti/JuVogjUU7ridtUyrdACoPn0vkK9ODIQikH1ZLR+SpjhshBUQl/zTqAr47WqN
gFxZU14QNwjaWJ8BOn0ny5lAeKPxEmTaDJdtOjCfTuC+DUTldnVEomoNeUatOkdGHWSLVJ4/2mrv
RpZeQkMgyAa8mT9Gf/gFRnYVWLH69nd46nmrR0qZBhv3Dmq2yiNJCg5fmpI2rf1HdOG/V9NEzcMS
5cxFwAVrL8O8zfN8gFHquwgawAIOihFnyY21uhAd/rnIhLb9N86whmPhobDhVkZ+QqYuj4GtsRgl
eAQ4S79wegLWA+8ptxG085+uUCAagbbxBbvTBBsy/AnyMjlCbBKD+GyKPYkeERwkpSji/c8D5VKz
Bsi+Fbw+TWc2aCGxzOFB5K+Bg4es/CYY+hI+swvQeGGMO9Aj5bA+V25M3qbkiAK983tqoTBj4TlP
WshTyuz4W3gyYyQQ0BbTljDlxVOjPtcb2lMRxdD0p8DnvrfC0pjHpIJG6lVEseIG3zECTs4XYKg1
oJBBuJDaYN337NUjzPmu3KiF3RS8A/z1h9W+R97x0DEx+/Go6M1bCrxQwBjkECI0F7gjBLlb0Dmu
9576syk42LL2Atnqei0GFljtoDcbBOnppIoxEDm8F5B1Jir+eEazobCLz7foM0PL92xrv4lZAB3d
txcqXk5PPHOxv+0YM3DydzDAGkwoMteoXmlVbUEWE5877/1GdPzT6O8ZOjlglEpPntf4VFHnqXOF
eHvPeMj/vFm79l6LrwyOFgVpKFn+H0uin6ltEbIK8b+3t4UWMgmkRa2mmR48iUqaaQ2DP5efuBzo
yhBR6uFypaR4Tm66pqJiwens5Kkhr2+CaOaTSr1/QCy/9xuJRoH4X9iGKUORL4ozjfIJip3KR4cr
oUcfemak8vRQqQ9tO8t8d8r9oI+uRvadKJkKbg/OBBOiDAkHxqPGJdgKtMIlxtEilhjm3TyT2GeC
FndljT/eMO0Z8XsQEUoevEBjcIL9e1C7nm2RGCKWD7EpEBnKOhHclN8IhE+p/X6FBrzAZg+3V+PN
Z97Yr3J2aH6vIDTBaXU58REnXy9apJ9sw8E9Ke26UxhaVldPwADCT58Z44dHWxfXlrVIQdLLj4Pk
tNqgooPc2EiXnn8R+qQ2NG4tnBla7F8yjh8idoYvyuJls9Rn2FCRofiKRH29z0Eg68ZmwDrCIWgv
wlnUctul0LWtmAIw8CrgmlPnbjqOZ6KGxyNN8q+fJhXBIZJ7HokI2CUeMGXymvATXb1/XUsfmIlz
Sx4Vdgn3S3Gz2A4BBuDufqZs4L69S/XB5pHjIR12Zdj03K8hyR1ciYGiPZfGkrsvEsuJ+erkO6YD
XbUPu9oaaY5sLPK0saqi6FH8dHWJhCy8GHlNNHT9wLfvefa3Pv3yjNpaprrdD1BCE8QEhibLl//6
y+cYISrjG1AD40//GmzZ0DjDGq3C6HkkX7n/UfQi+KURinDTu2EnL5swGneqVNY5bRVBW+iQvl9T
mCCj16fVAVIBUwgKKSdU5YpHvGiE18VOxET5ylLzEucvEUf9jbfMthyNZE7XVvn0/ITT4zi9LsbV
ECiy6ITa0Fiz6Hk5N4pYSlEKFU+sFCu5MT0NsrgSwdHriNArQ8tN/+vW1irunOWh0Lop/277OfaW
dXPKFGs9ufOumT8itnKUkgXi3hO+mp0v4P/iaVajSOmCsuso/Tc8AJmE4aGyxvrMhXmLCxkJCcn/
MsNNludEDwtnHGzvZxr+AtAx0996vIUhsNMUR7xIwR0FtqPOhrm1hEeAwUtpO2p4ULZJzwYgy/qj
XCg9WptH+GxlZVDY+/yGG2fmCSXns59HyXPo6TN2iytsFmWm9Kc3Xdhhg0xSu4FyhKHgvwtzG703
bBvjNLLTkMD3/AQGhy0b/2w9W0wHw+mf9D5C9XJX4yZ66LZQai8KrybGMT5AZYaqCiwXWeEr+8nr
ijuiUmXIQ1dbDazYDsoqBr4TlzalqlAFpu+1V9Gb4yk8zJ7/UOEM2VH8B4CtG9BpJSvSgSW0uijh
gbIGdn7ViDt99+CiUIBePk0H1d2pTsCaSmJq5sYQLbE1e/beAR2xo69p7VxrmQNnnYGPfTtvLtTf
w/VBObcIQPBMv90bzkBVmzn/31Vp69lzwPTLyl+r5IwhOQ/WzNNsaYKvIWQMZkitYoES/aYQR0G6
KzwkDYeCkKmz2dS+MowfWoa48CC2PF24oATLCwETrRV2DIZa6SlldQNDTDkdFRcFgO29X0xQCVzl
gCT4b/XKCQlhZQ5pvpK0SbZ+wbiN9RxcSAPYbxsJYW3P9rw7H0+y5nHxBBz5d1tCBWHlJfabg4Fg
HoHLlVdcdyXFUpa5zSpIVGOSY8DKJwSPwaxc/C6Tcri6/fx/G/sdsDyENV4VxhF5XzDWdaZmOv+6
j9KZXyc8/TvBz5wsXV6HTyrO3t0QYyoNpsagCflIdgBhX0ECyxLtBIHjT8HCSI79GvpJR2UFsUn4
c0KfYPxWevhnf5saOUhh1pwxVceq1xQ3uSfIC/vrUw4xfJaGfug7QyPOhcPAHjYYC5kxEIq4Etlu
p+hivvSHA/1XAPPNH18JcvDGKCYRNyS5YcKWfftd/qbGxgcFEk7pWQryT1yapTM3D2iAGBC+Ak8o
dcLxtLIkOI02nfjqh5sG16ig6imvyntiNo0OleJ3MbbzkyoEB+uyLGsAowXgxdPnw/imWrSn3PlA
x2ePrjizZqAQzczE0vjJhr1BEExQZ5t1jIwcxy9fBG7eDpRmBBN3YPLjwUVHaj6I40m7DZFfB6hb
fCwB4isJzs5Herthxriksl9yj2ky1Wqb+/YSHbFukznj59c+DJ6qx8l4Ty61OszPkzfRZw5leyZ/
3UKg3JJcRPvSLeoOay3V+KF9O6M3ytEzCw1aj/6Xa9okap8Cpitdap3/HemOm2njvRG3jvOi147t
yKAUYaEzjvXuujz4z6ZXSX/FmOFgT5DtubbmugKUmjzxucoIWCNPujfTqsgHRY+00YMolT6JGrVT
43pLW2+Y8rU0v/AIReqWLcwvXRcGS5D3ki9xK25lr8eSw9EPME36CK+ya9BmkPtFETc9TBukUCtF
+5pYlSpwiTHgmcWUzIB6nSWq7VGj7ey9ZjHWT0X2QQV52AQyzTyfEVm4Uxgsy56xpaSMnxR4g+dE
4BZGAbwUQ+80EbhzohKGHHGTR3x2pO6JTHWMsLwoLYufhi8v8iN5we5hu7XDCAYmzQ8/qfWg2wEd
E+TmzZdu4JNGQ3DYfTZyCZcECtcORnXfjIHqzR6RA0Z9cvyuEZY1ZVaMUlzXqMKHcm9dp2OlJ/fw
c2IXsVvro+I2SB1MNmSz+Yu5+YMasFkLYm737YjXi9JCuXJMXkv9WiC1vnOxNZx43YtLD4YJgXSh
Vb48LKmx5e4Ki4DL0WKdJQa6j8sVi7zd49PUMHu05nN8JbpVOnhe3sLj2MhNnyCm5ONRZQIHstKP
u1g1Aoyut1ofI/iMsw8gSec147v+xAQXieEjhyihLWqeMXhZK81DBXfEeQ/9Mt7xOUDa7CBvcnr7
NYIzihbWP5GZ4f18DtvqlTD9l4KVxobPwciXTjpMyJU1dDk7iwGIfmDBfdvPfH2pdX2jLvEjWoPR
uUlZNNsbhPGaAdQTDdE07VMTJkqh4+l4vdUFK5dZr28360Qd7bRRjjsqQsbolNE68nUDW0ohF3ei
ek7wI+wiKV3eOqIhQ3y6xdh/mJhxQG1azQh2ewmKJL1k9Wd/w2mZk81lYWpDWYX77AgGcWon5a6L
LjYAo68bpEI7P6+aE6F0ql46aIrjDpc0RJaVG4ynWz7dZ9tLOV+VyXHwJbi01zJ0my3nx2fCRy+A
IjcdQKRtAaQkbsfUqoB9CMwmp0ilCFWs/dqhLn6eaokob+ak97MJyloKQ7GDb9Y2jFMrBS9X+x8g
R1DMtZUlZ9sEYppNJb6dyuL32T7QKLnYR47nUMG5FQKThpAN4vOSuYkX0d2SDwEZFbL93zFYWZQ4
rb3jYQZ8TCITAFrVN9hxyxVt+7S6G+/LGLNr/dV9kfv2ExKZ225edtKnPh0gJa6rW52P/Sskoovk
mQ0emgRZsDMdoBpgZSaE0fnJZRmgKWiUuG9dPSRxAsoD0/ofQETbkMXk9fbAdobXtG+eUnxdpcJw
2J6nLHKPyf/iwU0vOKbpxh+J0xB4aNVl6XrDMP89CwqIPL5JHMpFvU9NjZp+JHTIQGK8rsXTAr73
hf/3NOIEA+A4e1XprsuAEC3IqYFakkMJDzKn1fGkUcKGyh8rtDjAGq/gQesf/D6gHrj84dRJl1CA
wW8GCPuv/IQf7KOs6A7yqMkML1Z9Ak92C96pV04msPb3rYFNw82ZaQ==
`pragma protect end_protected
