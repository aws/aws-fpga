`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
ShoFoWoA/JI+uhvjWOXcrR4Q02haKxR1eSydGnZIBi1MG9VKftWqUw9BYo4m4fFJSj9NQz5cuumw
E94gocn9S1olCWacBEopav/C8RP1ipgMxxdeAr/wqKQaRAz80oAt8Rv7P2tGxz6dApu4cE+Ith1O
//eMwSweBzaRetCYA6baLhlfR/SIbRyhVlCY7XIyenaq7Z6Drz3/W3upGwMOts0Yw0dZwp7k94jY
mYDjWQFT4KLtJX3l+vC1DhPf9O6DQ/0h59Ttm3zcjP27PyMA3SsPQSzL09A4o60YveIwl+7DBqce
0t3yU4YTj4dpfBd+mgcwinz3U7AZS1bcfTk48w==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
TUq+jOLEThVuNK+6En6bSDzSKwwXJ4pAuoH+hCVwZ+gp2iPEG1tJCilMk1BizAOYDK6JK3Hbmwxk
Aeqg5cqwvro/EjxEtBX4vskRMZijjaWgw5fxTOYr+LKlvhqpGIatVndXOqq1KjCUIsf9kga/P/40
KPiYZUb+GOuGz1Q4jL8=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
GQZNkRUZzULvXjRPYiiPuf7XpJJWPETZ0WoJ+ol5TWId/4Btv2vQZinhefNQFOxBAkuKTrKsCMJt
OQwnPLSZ5Iv77Ycfx6pW0ohFXf5apLdchi/eAEryOZpsNRQgKGpaF3Ei0ePjKhwYAgFS3NlSDgn7
13/oN91Akgbl45DXuPI=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3696)
`pragma protect data_block
Q7d9gm2gJhWSjnKcpkVkvJ1vGSZFWbMwz3VLF3l8H3B26ZBvNRqW4W/tBTnxJllzdXnOrX4H3rcJ
YiOPJZOxeLHnNI6CMuVKLdCl7qce769Tilhqa+O00nGrILqwh+hvK4PT5YIcZjpXv/KSs0tm5XV6
beAYk31g6GTn+EdQK0jzkMOCB4eqoGFVJ6anfoYJaOORhcjNmTpifxurHYE8MUBC4IHcurZUhrMx
wmGl4y+bqgB+EFbY0IkTEjidVZ/wfFX+K/RZgBGj0F/PjDxOGSe6eQHTbhTFESGLPyxz+6HMxZ7K
F85C9kiF0FdwtH7wVMtl9IDpSELeMmPnXRBefM6yQB3Wx+oNVA5KbcgfXOMGKn+fVlGtcy14P0tf
uUZcuiJ/j/9BqnzzgJz7E1VCmHuS7SWa48zxR+0bfdMveGkxqqwZxixxZ2dXFoc4cSHD6KLW7x1+
6dQkWESlZTt9c87MryVqqRirvRTqJYv/KigHHgAjXrxDBkB1vZodjvyQBHxcmDTLg0h7H0uwE6FT
KK9I3S3sJLXmE9hP02Ng/DCs5Gjk/fI2GzsSQaBDUQfYtJvsxZMlMj67J7LEzpcE9c1vK9KFHZjU
HOvBRedU/TH0M+fIWoTe5kZX4Dga+UOxTwMRPrJXhIu71CSbsfiIfqiistxjR101eWXYVAmUeXHE
kUaqk/CVtacGatmBw4DA8P3vq/l5F4T+Trmym1FoigZ42oyPlxgqPJhuHu0xPo/tmwaXCDnQkhXJ
EoAmzX6rdlN97pbngaqJ2EsHGsut6VKoj4C6fUisdOoDcxUgXtrPWZ7yZISHU7wUXAr+h0MVIVQ4
Fdk/hAtdQ+5J2g52iz2/6G9k7o8puONRdixTfey9McvtCzZKuYvB61a+A08tjeEm0iJbEtimK8sC
r09YWnbRoDHaYItUCPL7P9RxslBKIQFSIyNnRkRijwNrFB3+AUdeYesGk1403zaCB7qAyojdUMRS
6wHaLw94/PN927tKmJcbUahpGEWcSlr4VaNxp6XvR6E+qm/xxM6mU++GfOxzeo1pQbP1K9T25U34
fgjXFLBy6i7GibbFH1gtlqJ2w2rsbq4zF7/1tWOVNLCXEhDvP5yjGB9uRyR9hKBYgAos1j1ZZ8gh
kVTMcMTDt2f1Csos5ZIT7bDHPQiTnwn04eVho4RKXSrYfEoZWN6zHF/aN2OdKyxSfw0ZS8NYfewe
X0eKq/g29VrAG9gO80MTcxYdfJx9mq+yT23SvAKQQfkn7Kh8kY9yKyMUBFoHBkPiG+tufckKq5XF
6qTRc3nb7BZbDZcjhS+oZ69VJpNwHuiljsTvMkcvdAvGHCk++Xh9wPoKnqF+gvi9Np3RnRI1/QM6
nXPsg5NrXLqVjeWKovcSmGeIxFVt0BeQouY3eMJh5hVgn8CaqTeuqft+tx84T59cV4j8veIY7fhq
Kv/JNqmInoUOgJS65b+XBvq3GUN3LUbjmOisYH5FVWUcoJ0Yf3TqKQ7AnlFG6a5FE2xFhM0dJ4Zq
/aE8+ny2YCC+qauHxnLRZ1Cjz7tJJ1/2y7ycp6sVjGF9m5AY+km0tC55daxLtLBDQpQ9WfWu9oYr
JrESyrPb2tuoxjoAc3Ez7rEoubBFk+p9614/DEQUm5lsu8+Kvl17X5MsbacUPJlq1zzd+r8/0ZRb
LM/tvqt7aIeYb5S9etCBK6Eog7x0xMvKwbSF0DNFqf+fpERVNRjilqZCF7BNBVJ2akP/c8vhg7ky
WpRhiQSpKTsQCuDcpIlddBkqaQwYi4wvTe+Ob+arWgsrZ2tOzWWDs5sj+CPUoiBaqEes2ecgWl+3
d+xR5KYYAkdb8+zhrT6QATIRaFGe3ORtsytpBLVMJQWosQC4EDy+2miMm8hG03UfMaTfgEP//KhQ
9Uz7Q9UP8UrFq/Jrcl1nuRnLYX8YNemWuKybT2RBTefBnS1xHLIerAjbj7NWS0umNA3IDEKe6+v9
7RpgaN9jGNzi8kcsAsNMmRnmFIl/VpaP5ZSuqOGKUhrBJCm/IzqXp079IxfUnOwqMyhhk03utUzf
tSHknAtV/faCtFHaFnkZKiSOKm7CtHl+uVrUKUdrFbr9YUWr9OFtKJPkpoMNhw2CiJ0Co0gnQvDZ
dQmFtcdb95I+pWLmpB3iqxIihQ4MKkJIFiYxRYapK+9Tn4e0Mx6Er2ekq/jbABqsWQPVkO3C4g1z
sG+Y9FRE2PrPsOa6JfveYda2xE+bFIm/Zq8PR6UcLfx0MGxiWSFyEMREQXvEdfYmo0+MrRQgi8jL
50wYZ5NXhyBBpW/yliGVpxK5X69MG1gCibUphFiiD9f90//IutvDmjzAZtArTdvrfanT1GX39K9X
6ED9enxJrVHcLuohe5EU5CDrwiAjaRoErx+OuG4ak1DFrlskyhPbIW0jziLRmRNZfrO0xSCmAMJv
kbVb1Sh9+u2ucwp5RVECqN+D6l0zVViXkXeFrW0TmxAEu59yd12nnFSWNHQ4sezNB//7bAjchN+d
tvrl6TCRJ5cLgV1iOrrpS0tTLVWm0R2OlUFzLqchC585WlTMWgPXIperD2WHKMBzrb7v+NwppIMl
0HaCqsP9Crg6mOth1ow2wl6wJZmwToCmnSDIXQsKThyzYGankdE/qQpoPXPsc33JX2v3EiGa+P3A
px4NuLe/HmSu63JFAH8XgQN98J7oQsLapsresjq2z+H7TS0n/rDry6BepHC0Ru5pFzZ5PPFT5XCh
pICC4rGUEp4jw4iAWW5yP/WZ3xRbz3eia7GciDALQMH8zhGnY64BEAIo9C99ZC6DD+xTJlMhAEXB
1rH6U0hOcZO6ebjgzZy67oX2zOinSiLAoaNgQ23h8YLXAEr6eKBVxlWRk0C1jH3e5J9CeH4Njwau
PUcy8M/MJgax7XmDB/fjW6zDsuE8T5UwTd3NaqriosZpP6Y8JlIDfefYM72s/rZC6iwxFhVF6AX7
Ivzcmp0ADOHG8AlmNaqUEU5PyY9a0b2AfrnThBmMHsJJ9sPN0WpSSxv0/jRz7uBuk0VX/4n6GgLj
bG61kITZ6JvpwS2S+42vzmgW3KaeLgahTzTDbROAllztnvhjI4RJV2hII89KWH4tBQCJBWUrKBF4
pGf0b9k/ZQlSqGDP5nupltAT2Sd0n3QFDF6PzqO4pwh6i/Eu251WiC7WXWzd/g646IpIqyX433oX
u07WRmfplUNS7YWPXgo3knacbWth8IBV2zavybfJnEC+0gHbcIt9eh4K98n+UM0kHjAaCfd1eMEW
YZfHIeiBt+B8ucqwaCQfjXMHf29ZJRkRMIjc6qFYxTM6RSQ4BWh5GjzSY9CFfIFg0blFaRp2CK2P
3pg/ZLLE6S4kmWNFCy7SkglxmG8mSo3cn1FwxKK/jcS50G69qdxodml7GQb/xOfzSBs/akiLcdaR
KJ368f2/qnVVAmcPQlWHy6JzOKWc8ZjJuaKpQtN6HpzEtPkDlQELhUQVYTx68s6JvWfGWzvIpRnm
H6ZaX8kY3EXkK6op4Tqz6H9xoS8EXGc8eMbVMdTS9YEBX0qldaxkg5TE5j2lyPgVuEBFzhQ21TIu
bM8PCG5sfjeMZnKYKHHRq45w1yqQ6Yw1fslChHsYvlUy4IgxvU3ruCSZ8BU1XymJ5HSB8g2evszc
tVCTV1nICQxSoM3Sb7RqXaAg8hCD013fysY5KKhSQFEU5XDaayTZkbfKCryXCsFaxbkvWzHtdd0j
lh33wuC441xYwHXMHluddoFCFDQvz++Cez9zj7m1TmnCTh0CPTCAfXJOhLW5/1Hb3IweH4e/MtZW
8hiaVhiJHOZoom+/wHZrTKwMag23M1NQx5FGEvkMiDc1Ww06omqL05TzOMGZy0LdFOEnvf9XwpVL
CH3bGXKP2ZX5OciyAmd1LYn7BhIk0lJt/m5ZAW5AMOndl0LD5BNnDQteLsV2LM7WYKxdWncykrDH
YfTq/YRXu7SyabrGYnusuwL0L8sR63VQ+30gFnvheldqwWUDXiZDdXsD9/C6tZuBCcQmt9Xtyfm7
ewhfgHiH54xbCWs66FA27SpGIecCE8luy2nWwtb7ZK28E8ufVzlZeYNnt+A7hf7faC9KxoVrDvin
gbXt5Akhag+oO9qzN3ub50y3rN7ydUE3PK2Z03dFuwo/l8w7zEUqADh/oebr433enZ5vY8xtp7fl
drja1J/LjYaLC6YpLYEeWRZhy1KxlNTYQRNtxlKg7QjznuGRkoRrRFNprSy3pkUhQ7i1bVhcWo+h
sPmSIfMsk3ggL+GBtEDCVwa9E2/GAyffzO37qaT/pbI7fOkk0lGbdlApQgRpkAnXqTDITiW9cZcS
HlRvlybxGXPLYpSHAp3JZ3+3aOb1RtyY6p1H+hLOrAue3/hFZeicl/bBaH68EAlxXov9yjZPOIA6
/fCvCMglmDuzupusX4B1dzUUnYvfDvJkJB0DAAdeRGVxaIO7hBGi+li3Imoef08aX3+dg4vRknZG
gYZy30rcLfricQc3YUvyXJXDrDYhvo/vUt3G/jI+ShgqrN5SIKlmg3nYWSK30iqrxvAJJhUhJeO/
L6cjqpMeeEX1ra9mvVlrslKg59shDMd8TxXr3eNT3QyA5t1XRtllgSfUBZBalcc5bFBoCkekNuIA
T8X3vcB/RTn9OZIJRyIre6+n5G+RV4HhfwI7lOZ0WWl7MQvjKdC3ce/QCOClhDuEwJay02Cvg8qP
Nzn90JBtuo73CEmPD7rgN0UIZzGYKzhobDyNNMMzf2hncno1dow4PV/Tmo8Yh1crU397yPzsHUuR
yi1+0QkBD+vCaszTfbEx7wskj7K7GbHb7e+CWHCjPdvR7GZ8kxfsfmksOLn/wLPhzf2joqtcaKJb
7jjai4Fq7IZMllfPQRk+htUf1O3f/8NP6tYhiyfGDd2xtn+d8lQQJzem/sGmHdZ5
`pragma protect end_protected
