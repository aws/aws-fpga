// SHA: 43f4f449b937011c34848123159f70bd11b98098
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
I9Vw0IeC3pkT3VQuj597x37dNBljRwhfkSvLTmn+Ap3kHiImSKKpe1bJAano11WA1dBjd9vdqCn6
C7VF+EFvRNmBAZqLtn950T10W7ZA25FZyzmz2HQ7YHmrJf7EpIaxTv9NqDFIKvywsxwOvR4Icu71
MJyLy8qKx/r6O0Ywf13fw5F5J1DFCvdhP2NvOuaez+L2CcyIaXsrPQAO2I8X/8U/UPMW15/xr2E/
/IDdwCo1vhQdoJSBvOzxAdEDu+EK+SFqHG8XvPb3utlX7NExb9KJVqQrwFCzvmIBlhzuzd3IYGpk
xfqW6qXkf9U7QMpYn+k+hOgAYJMxp7PQOyovAg==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
up1uagoP908fZPvz4MEeeBgx6IGJjqA1xMActBrAi37uQeUZwUhMAUITC4QvKoo91HmKpyjDsuRk
8zy+U8R+p9fF/2Gb1Cl3hfu5Wb+H+cOvpWn9lATPSQ/YF7tBDJt9skGGJdV5XVh9C+otgdfCXStS
W7Gbzbr+53TWf7R3kG0=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
fivfhR2fk3nLuiCa/AC5/KdEMFuOtifOqGDAvTZ22vfsXa8EACXSnT3KLPkKCcPE8Z77naNseXpJ
yXd2gfxbbT0YaTsHi6NlBzw1yIVXTfQITJ6OceieAKfa0GliBVXqQxUz6yV039YTMVaXG1NwoJo9
bncGL0wJFoq2U7OMZS8=

`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
hG8HshecEfc3GNIkvwBRlLgQiErGX43Fb6rd6hP8FTTLxYrhvEz1ecNUwUPmg9n31obhDAtSMdj3
oiZfEIq13A==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5824)
`pragma protect data_block
hYFt8sbR/xCTYQ1+0wjJSehpWT6RzdCH6cry0nDfv8i6qZzumMC10sTUb9yh+3mY9fHkSD9NAUfg
p3uyhM4L/PLqQLrc93MXAZCZqZS5OxW+3OWhnuZ0ohyNwQTvcIHAVjHZ2LtZSVGNJN5GZhNG3HqT
ZZ/yvMBixlLlG7oqIBoQ7xIz8yAySgYn+Gtg5ZCZ9igS6iSw7sreWknhpYgoIOOtFWswKV1+7g0m
qHrX/7T7KdP04R775jEhIdBqC9VobxFv1zs3X5Fusf3cf9csNG8c9Q+fSU/07IZc9ADs+FQ6B2Q0
f4RXMSeM3WO7BWnNtny1RVEAqSvE20p7ybkavyQuDRH1jDiAWzZayKFx1MS+hr5KKeeW3JtPByaR
Ywigz3L1m3e4hN+T5xOYJhdrB0wvouGR9v3+URFPqOIfHFnTvm7RW3+q002hVxJJu88dxRu87OlJ
pzauV3R14kNABX+Go3gxjCTtgT+LXMQAP5pkZeTq/65wvUrDLbpxKATAgn1Hx9swh/Wnz0cDt4pU
n3W+giTepJIRWONanRZBcXF3OFZzO3E3P59e61F7ERivKbY3XHc3vqTUpfrlXdi6SLGu4naWMzZD
Q4AKX0x3fRHbSQtMoeXixurlFQkeZ6pEZ66NFdE1muGv5ek2MRN4li9gb7BFN4uTanxENSdoI3HD
eFHkJKzFlc8ABwyZNtr8kSDgu53DbhcsCEjSByuNE80wfIhrpVjR6XlLjp0uNMmsLQHPL5KtCBWZ
TUx+NWLxjK21n/a6GCdbmcPVWpP9VlaU4anfZfFRmqmALv9Hw4zJsBizwNSqcNoJ0SmCZ4nIbBAi
GA+d59KVVb48eXJtE+aTdcQW5WH6CI10kkQQu5s10YvoRgRclYEx4b08vOgEKqkeH60cYmcdy7db
Yi7Pprk94lg6aP/CAEGXcWw+y0tilEVOSjOQKx52YHt2jNRPZFEsWsT34RYMCQkuwze+I4KsDy3M
x78Qga3jg5APC0zSrHtAA6CEq7IGftgrA0z+YiazCB7pqFdPpWgHEwJPf6WenSdViRS6vyCZ2+ED
vuuGXA2+vmIPsE9ELqSGqmngQJUO/p9dAS6Ie7bWwZpAwJtG+T/NeMWPYX+ax2H4QCkcVXpA+XvB
B0a4vgCCWW5eRFc7WJ3jwgHV5NMXTLhmyytnGeQeCdgJcB++5P6N5O8SbCAnh1uaRaSDXENYeqG0
teHBoquBpN2LVo5fQ1rqI241Ib9CeGqVhRJ4LOi8wRv+lS1djJ14Dnmd24WkY42Q5tDGWn1ZD7I3
QJrjAoxH6Xcr44eL7cZbmIDUQUnV9jW4s0y417XGtnt/DBimT1dDF8a2WIOe9q889vCpP2pqHqAr
/0OaL5fReQ7PlAqdNnipuU9qaBrQ6Uf+25lYTmohl16hWSh0q/QmTWfsXefip3bnOwqdTDf9L7+K
h4EkYP3NVjt1H1KkI8IYEcwX6sy44zqK/vxMkfaYJwVBfI7spZxggm5+eWjstGKMGfj3GRBg5WyT
5tZHjQHqy9KFYk0adlZTjR3htdaPQjZWJ6W/f4JqoU+1ZMTl+rVV/Zc7Q6clrwA1nYieUxCq1T8g
45pcfIcafUgqgCia1opMBHy6829pLh24evxOI/BiMsMOCsmQb2RQ9asxdYLf1W71KodW7maeqwQE
SQ1MJbF7xaiFZ4JUpwEPK3MzoSA5XiY3cO9IxOW3aYcFAQgaRptWerysaGyQnh3eE5W7OrqjWeeq
zLdNH0zIBgBqkZ/LPqoB9Z/aMvC9Um5Xo3Vyo3vipnv7AeidwsWOUMZD7MxSVDHYH+3vzEXQnyrT
GgxINMzBFGL1Yt475kniS+3tSfqGbqglsBDWByZmQRs7X6XhsjWQ0PCzFnHv70NB2rsbj8DlN15w
YQ/val8PahT/AP9Zdati13jPawwTRu1IumaqgIkQIdvJXZ77wRPAkwX3g8gtnZ3glh3QbP8iO4Ih
Jo5cA8cnEABsgTI5R/IGAG3ntbyHXjEH8VLJDa8OcCtAw9p0tOd4yIx+E1aoil0/l5mJiD38hHxR
seEu+/XWYme6//g9nKATQNUHeW7jI1uOQMVIZe8H+sQ/gmdfy27atHRHf2WZ6/oy98r+xW4+hqLX
4h0qvmfBI6bKZTEixkaq/GdX/ruIDEEJWhryR3FwCoqMr1JlrGQuxYFVWsB0VHj3R29BXRdUj9O8
kIQeX0+oEZYnqllKbYgouY74+RwpXWqMceheEhWoyszbffx8Yvt06B1zUu+5gbX6QuaYX+pnpBa9
OmHpa8UaujPYwmRJ0PoyaK6b5UcQo7Y5nUKzOFzSDkp3o4QaaMVsf8craANgo7HPOHBgBvlgEhWl
JCjAQFq2ML6iHPa38QqEfoBQ1G/koRtsYiH4egn/2wVxPDMj/uNKhZhFRUPcO3kflJA5rRf3UODb
USIR8NalVEJwziwxJaudj6OklOuJmT/6kKU+AdQQ0FdMuW6/sJhFFhZCw7BbH49fZKVVpwWfs/DP
obw7zxKNLG8P4HJUl9F3QdxyoAitAmej5CK7iTnKW8Vk89Q71TLjmul+caPUpxdwDe8cQkfy0gW1
E1kpce0e/MsjxOkHNGOQkO2G4yfxmXVHNd2dYWm8MX8061PC9b0s47JxEYFthl1nl3HPW9QQY1NA
YHRLotj+8xA8YcGewKYCo8uTrQrxW3Cg9tAIIDxQiC2IjJcTrcy8/XQGX9XmQ99ZAecooAt5NxVC
0mZmCPywMzBx3HIcGmI10Nm9Oq4zOB9R/g2JfYx1Hv4dO3sjEganRmlYhErUa0RVpDp/EGlwaeWn
G1ix6ZOiELsk30iawFZ3FZuDyjOwOHGdcgBnF3nXVg3AR+RKDpXANBHDlc+VEJ4jk76KDqQyYcbF
LQAXTLyQ/7zjwunFYx0pT3DOy1qwyQdHWVuWsBl7RHkON8f1rqyX+YmQ2Ensl0JVyh2aTJmEae2l
pQO6tGaPkiZO4G5rnKg1lSvfZWuRkQAGVBFoF6+XHoPW+ovyhLpcayIDL/lUJWV6jvoO8CIL/J5/
4ufkznn++LWzbN33290wHua/bIrxoer5ET/kK8gHfUUcv7mfXKpftEKnD7cMq33gbzyCM0dfvTaB
rZeN7pnmb73MjpBfuK03vHCxu0c/XRz/S0ZBi7VOIgsqNmu+AOed8L10kLhBcPB/vFhMREgEc95A
WEf2uCg4EJGMztQSfUTyTawpHrCMil1YrE9NuDTgfuOVYBxFCB9m9MogZjIxdTh+dm00VWiW6ZPE
b6psc9bqN2vMg6mQGo3pYMill7EFgGDxAz1h4ItgTneRMV0BDs9VYV8iO7bUhIoBrmZImv/AmjRG
ZHex8z16Xy9zOdyDT5INvDgHJT0JNMHcFqQj2pllFlPGtwnHYDxlt0T6yqp9V0Y39Gu1pzBlw6IZ
gh0s+JalWqLy7MvfJADepCY7pk8q1hFgOknymx8mT2agf4+45L1ocnDSFmIH4omEqQNZzKD965Qt
vprPBKFi6wRzIhDZUI3n5W6r0IEJgD1l9EMy+ypgbRP5+3fMBKl7WRQfCx02gpM5Ye1Cng1gKcqT
bFBoZkj8+PyowETr8N+2icsRExAZmEqFls4Y6BtdIpIjQgkPtgAqjjoGjRUxPsjz731vToJm9NPa
jit8oKQMxVikftnosQu5AOxCnOVztnISOwDbonffccwQLceaE4o8AVpIRIMX2Pi1bHilV7qFypvm
f+d1xKIi3sHRBvmTtMVsJMVvwSk1DTI5lzyoZQyHNuc0La1VHUGHnfOJvf55fruiaF+jEXhtMlhP
XSfkWoLjR+dB+5m4GOPQvirF7YB2WombF9oh4/YEtfofY9wKrkrrrvQvt/PN+G7NSucDDfMDqm+d
PspkiA51/RZmBU3SjCRWTVERy3ny5gPLSbMMXgjS3elExfRxTvzBhWt31Uj7ZlmQxxFu6RPHysVL
tgzRkzlG4cScMK24dRLiENrwLUJYwE4tuzw5y3BNh3dfNOnMKPm6xq2crP+L5pRrDYFLS0V8MF+F
pq0KUk+B6m0pad+1kltDXFnOeH9GAcLaO3Ygbgij89kaSj+SiIfUQ68sbdLIEOJnXb2NxcLDmW+1
g/vYjxDU/HjYefYRBet/KLmngga8RPTer0QuUUUUQTR102nPY6cRq78GTbSc8ZKcHpyYMmlU4lcP
eVP5i9datG2H164FNzUuYUyMqdjeTMDu4/p19LVPfizZiM05i1yTLUvrK159FbNG6dXmnXmClpBq
S2gUlqL8ZM72vhdcsbHOOTOCZSwIlZBYKrQWsrh/8zeoK3y4hFHKtNvNhjeREHGmNoO+zCaMgpxr
306LJSI4R4DrfqQ7da+vXptVwlSuVVnttfKjM39AH4UsOQMhK1LS8BswSO0N1lbxnvqk7xVUm8fJ
YzDkM1HEl2rJkxCe9XqkDVvIl7h7WltE3x2NfQNWdg0drEdFOpLd8fzR6dGSlpp4pV2jOoP7nQi8
z6HH/BSz82wxYOs4dA+Td8WHPnGM4M7I+ZpLYEfsu48yz8eOLDxn+50emaFChnrSMPqhXpn4pMnu
+HqROB8Rts6IUjTJEnxWTS2FfzrStGkQ1IV3UwRunaufD1OXRxGB8M8cnXYb8DBQVoNIAGoacqdx
wAwf2wXmgLnsVFciK/q6/3vXrrEFk4bDw7xXd6Yo/tXhZmiVHVC1We9dEGWF/CJbn3MuVdkRNgZi
GUI9JA0lFwVzPVwvtCPfYeYukRCo7ibm37OJ66PYjSfR/T9EZBNiN6Hm2+g5FgQJ7yDl7rY+TOsL
Ck8r9u6/Ylb//94ySEybUzuvlfzf82wClCbcAgpIYJliCAfhhwm80R0uu8+roY2wiFukcK7ISgGm
XIFG1hCxcsLiA4jWqLE1PtSroBtUS7Kc0SKlYOjxDr6n74gIAqv1UwtUGwLrobl436yFskExboqs
odrQ5r5tapng4bKfXc3t4HHfF8/X7Qa8fapbuDMyGt6bKjm17/xnti+ajE2t2hyekCbfSNelof7e
VgRCFt2MtffSPJS/AO/MrSdON9+RuSyAzQoj/I6V0ohHEe1IFFzCp79d2JAEJ4bL/DW0SXvdsVpj
X0OHvJgQ9XFterqiw4WNFSgfogXePxHG47exm5c9WBmIfxSNDB8p1ZThYyeS1kGXhmnea4tK23aY
YcpBX+/YVajOlUEW++LCIy5Rdp3aTk4PIvUfpcc+8VVg1HzW8kkBkereO+tELXY8rEWvC/9Avek0
qlg1vZZXkZxRUJJtPqBZ/ePVPgFDOLzOPs54x6JDiC/9qp/JaAhnA413v18QTN1SD1zImdHcaGdS
1KHj073qgwk0bSgG2tHXJ2LI2R5JEp5YjJVR462YeOaTzNxDsSBOgXaluOrxQuP6J38dvjMY55SS
ZWSk66p1bufxLTcdiyv8aZnV88rKnc3uKC9WwZq+wD0CKuecS/oDumK4KqMk5jgPQrZyLlkbEYZ7
3o1FU7TyfZIpuSUBvZAaJm+Lw+/wmc7RUcESyVsfUFs3ZRCxraa51f4EIWwnzcHNchlgTmwHJZpr
bEoCFHFa2NR5iJ3rE3LfZ/bbZY2lUXmvtTMZ8Q5WW/DXVbxt3rwL4HpShsnV1UMoMfi77iIXLZYB
Z34xzDtt97V26/1Hy6XkJrANoFFWF5BbhqxMK9cY7Tr2GUltixf2ANn2nel2dhV6pysk0AYV2uuD
bsfLg/wLwPozEwOucTcYxjoUzAlXIG9BdTVUVrtaH0XcIV7LkS3HN1cVoSEI5/FuC3uJ4/2HYWPG
dF6fuVnv/5DgYPz7rd7K3Thm3gX5PVqZNAoB6WTX/ZlwWWqa1pQ+CQlKiagP4vKw+RiNHM/59Zj5
71WncGnX7qTTTe1jLNGbZ53f3PRaZ/A2aAlkBgvk48ScmVJ3SOWm8AAZJO/RYI9U8yzCRTWeFVwd
yEpBRMuX92Ee8aLgP4h071bD4YagvSKmgq48w93dCtVa9No+dP8Pk4T0/RbP2f4bPVNwvHCvWKgr
6SmczE8CX0SOZuO9wJEvdbZKD0tcFibtaDS7BtDGpgjz+xB/XtXKl/MnaItzS+tjz2vWtn4MZvHP
a8DY7ZK9HPOcTIB6lXwU04szxiYAEHl3AMG2xdvGEuTn8dXcQNPrEfuEM2Pdj090oLDeGY4AobI+
7a1olUVmSQ0lK51QeBNkDM8t6BoMsus8zKyaQXBGEc8u0RaJLkeToaZUyR08prlO6ajL3yEl1rtj
4D2Wp5dBUkJj7r4M73mWHjV8wut6+bRMy1KUXezu6tI2QtU2hjzPXAzji84OKzP7rDxK5IRJu8wR
PVLl2YyucjwzeOOI2xjwBgnFjhZKKTUZoJlw5hXBWjLCc/JRhG/nVhVsvlCGPhm2ao5eXO61y/dx
0oejxHjTNwYPr7P1FmoPeZCWCo78QQA/GG2iS/cABm71F1H937p+Q8pX94yAXNGhRyUudmi1uLHw
cByUjurlLhaElvlEIPM6x4ib30CabfL2IlX3YW3htz2K/C+yY2sC65OlNHXzcxEq7IRy+YrKkOEq
HOUuklU6M6dYW2ea7d4hTkOFJvBDfVmCFKLp8vvoNl8F/CVz6AP2kwLDFIzJA1kESIxOngbimG5O
hxvt8dZytdAOuXbXBBClg7PfbgmW4KX9KV0fkNoYxN+KPmd+VGShBhlEmp482W2wtWh3Tl1Y4xyq
I2sbVMhjNiiWIN84cKTm2/8yOdftm4I2OcaqWoWOaqaIPOHjYzXEm5A4tG0PwpBbsOjD0b4tBVPc
shUWbabgCOnwZ8x/YiaQ7N4zhe36lmJFxUMjjrbt/KX0J/BLdC+N+rk8FDk2mNkvvpABD+KUy0pg
UhkZ5H1V1XvEYooJVjCV4dVZ4qHrRtyMb6MR9lmnRekt+ZO8jWf/5eQR/NU2jaX2lLsyFLq3lsZx
Voz9FjZHYOZsLEYOCHvREqjAKxfq4JR8d0T5ktH6bOy41oLhGyuafsjA/N5bCGzOoPog5QDKI/fv
CIvv4Gqu5o+9j4SsqjrA0FPGlBqmvBCnI1oF2ECJKRUBsXz7GFJ7wThm+U8h/tAMzx8jKuO4ZbqF
iqQ4XXvAo2einweyWev0UHiepmRtOarPT+t21yhQRiEhsKTRMIREU75dvhxgpi50NNu3ITIIn3EA
46Z1jiYpIItNY1WG2oMGJMYrvkuQvR5X7IVLQkpVj6gI7HIn0BQGHLt8MTfQngdVusqn3D5o+8ga
2HXA1DXMcRhOhgNRNiGp/YiahEEBhdJaNkt0TmpcpS0zmbV7+cm+DB3xb1vQBGWCa2V5lSuCJjZT
9Xm8RuLRtKa9JLM5yGpdjLA6yuY6eP2RXu8cTXK1ochutqS11wm4F/e6u1pdJl28yUmfrV5ep4jh
d3D/OyxmD6RCPeJGEhIxEpzHvqLXS43eK1/8LUuW69S8XSkV/ga95XP/lTrQ4+jGnlRTyS5s1r5R
d9x6veZAS7zb19mjhoj71IQIxR0TdMUWZNVZSrXpPNP4wxVHq9XvFpXRk8LV2FGqNOhWwy3LqDZd
fK3Lzw1erlbTlWluMNONppy5Vrta8n/qbYTZT6meK+UprLspAS/QgZW3xfW4fe3eCZ5sfTheFG44
FPlC/3BvSbO/RkwaVazvlT1WR4jdjufvBu7hcS2FZv5LpNvRiFKUj4shljl4pEsupQ7Dvml21w0P
DN/3Qf0tq6NkvOMfn1ewp172pR/FjfIooqDzHBaAyhJpwMvnDtPdRiyJTDQDPf3vBSESM+zn7S1o
zKNHe9MWwLWOFQ==
`pragma protect end_protected
