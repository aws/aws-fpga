//------------------------------------
// Tie-Off Interrupts
//------------------------------------
  assign cl_sh_apppf_irq_req = 16'b0;

