../../../cl_dram_hbm_dma/verif/tests/test_clk_recipe.sv