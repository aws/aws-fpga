// =============================================================================
// Copyright 2016 Amazon.com, Inc. or its affiliates.
// All Rights Reserved Worldwide.
// Amazon Confidential information
// Restricted NDA Material
// =============================================================================

//--------------------------------------------------------------------------------
// Stats interface registers
//Register MAP
// 0x00 - GPIO 0 - read/write scratchpad
// 0x04 - GPIO 1 - read/write scratchpad
// 0x08 - DDR is ready status (bit 0)
// 0x0c - DDR reset (bit 0).  Set to drive reset to the DDR core.
// 0x10 - AXI Address - AXI Address for accessing DDR core (refer to Xilinx DDR specification - pg150)
// 0x14 - AXI Data - AXI Data access for accessing DDR core.  Read or write this register
//                   to read or write the Xilinx DDR controller registers.
// 0x20 - Write Words Low - Stats, number of words written (512-bit words).  Write to clear.  note is 64-bit counter
// 0x24 - Write Words High - Note can write either register to clear entire 64-bits
// 0x28 - Read Words Low - Stats, number of read words writen (512-bit words).  Write to clear
// 0x2c - Read Words High
//
// Interrupt Status0 - bit0: AXI-Lite interrupt from DDR core (refer to Xilinx DDR specification - pg150)


//--------------------------------------------------------------------------------

module sh_ddr #( parameter NUM_DDR = 3)
   (

   //---------------------------
   // Main clock/reset
   //---------------------------
   input clk,
   input rst_n,

   //--------------------------
   // DDR Physical Interface
   //--------------------------

// ------------------- DDR4 x72 RDIMM 2100 Interface A ----------------------------------
    input                CLK_300M_DIMM0_DP,
    input                CLK_300M_DIMM0_DN,
    output logic         M_A_ACT_N,
    output logic[16:0]   M_A_MA,
    output logic[1:0]    M_A_BA,
    output logic[1:0]    M_A_BG,
    output logic[0:0]    M_A_CKE,
    output logic[0:0]    M_A_ODT,
    output logic[0:0]    M_A_CS_N,
    output logic[0:0]    M_A_CLK_DN,
    output logic[0:0]    M_A_CLK_DP,
    output logic         RST_DIMM_A_N,
    output logic         M_A_PAR,
    inout  [63:0]        M_A_DQ,
    inout  [7:0]         M_A_ECC,
    inout  [17:0]        M_A_DQS_DP,
    inout  [17:0]        M_A_DQS_DN,

// ------------------- DDR4 x72 RDIMM 2100 Interface B ----------------------------------
    input                CLK_300M_DIMM1_DP,
    input                CLK_300M_DIMM1_DN,
    output logic         M_B_ACT_N,
    output logic[16:0]   M_B_MA,
    output logic[1:0]    M_B_BA,
    output logic[1:0]    M_B_BG,
    output logic[0:0]    M_B_CKE,
    output logic[0:0]    M_B_ODT,
    output logic[0:0]    M_B_CS_N,
    output logic[0:0]    M_B_CLK_DN,
    output logic[0:0]    M_B_CLK_DP,
    output logic         RST_DIMM_B_N,
    output logic         M_B_PAR,
    inout  [63:0]        M_B_DQ,
    inout  [7:0]         M_B_ECC,
    inout  [17:0]        M_B_DQS_DP,
    inout  [17:0]        M_B_DQS_DN,

// // ------------------- DDR4 x72 RDIMM 2100 Interface C ----------------------------------
//     input                CLK_300M_DIMM2_DP,
//     input                CLK_300M_DIMM2_DN,
//     output logic         M_C_ACT_N,
//     output logic[16:0]   M_C_MA,
//     output logic[1:0]    M_C_BA,
//     output logic[1:0]    M_C_BG,
//     output logic[0:0]    M_C_CKE,
//     output logic[0:0]    M_C_ODT,
//     output logic[0:0]    M_C_CS_N,
//     output logic[0:0]    M_C_CLK_DN,
//     output logic[0:0]    M_C_CLK_DP,
//     output logic         RST_DIMM_C_N,
//     output logic         M_C_PAR,
//     inout  [63:0]        M_C_DQ,
//     inout  [7:0]         M_C_ECC,
//     inout  [17:0]        M_C_DQS_DP,
//     inout  [17:0]        M_C_DQS_DN,

// ------------------- DDR4 x72 RDIMM 2100 Interface D ----------------------------------
    input                CLK_300M_DIMM3_DP,
    input                CLK_300M_DIMM3_DN,
    output logic         M_D_ACT_N,
    output logic[16:0]   M_D_MA,
    output logic[1:0]    M_D_BA,
    output logic[1:0]    M_D_BG,
    output logic[0:0]    M_D_CKE,
    output logic[0:0]    M_D_ODT,
    output logic[0:0]    M_D_CS_N,
    output logic[0:0]    M_D_CLK_DN,
    output logic[0:0]    M_D_CLK_DP,
    output logic         RST_DIMM_D_N,
    output logic         M_D_PAR,
    inout  [63:0]        M_D_DQ,
    inout  [7:0]         M_D_ECC,
    inout  [17:0]        M_D_DQS_DP,
    inout  [17:0]        M_D_DQS_DN,


   //------------------------------------------------------
   // DDR-4 Interface from CL (AXI-4)
   //------------------------------------------------------
   input[5:0] cl_sh_ddr_awid[NUM_DDR-1:0],
   input[63:0] cl_sh_ddr_awaddr[NUM_DDR-1:0],
   input[7:0] cl_sh_ddr_awlen[NUM_DDR-1:0],
   //input[10:0] cl_sh_ddr_awuser[NUM_DDR-1:0],
   input cl_sh_ddr_awvalid[NUM_DDR-1:0],
   output logic[NUM_DDR-1:0] sh_cl_ddr_awready,

   input[5:0] cl_sh_ddr_wid[NUM_DDR-1:0],
   input[511:0] cl_sh_ddr_wdata[NUM_DDR-1:0],
   input[63:0] cl_sh_ddr_wstrb[NUM_DDR-1:0],
   input[NUM_DDR-1:0] cl_sh_ddr_wlast,
   input[NUM_DDR-1:0] cl_sh_ddr_wvalid,
   output logic[NUM_DDR-1:0] sh_cl_ddr_wready,

   output logic[5:0] sh_cl_ddr_bid[NUM_DDR-1:0],
   output logic[1:0] sh_cl_ddr_bresp[NUM_DDR-1:0],
   output logic[NUM_DDR-1:0] sh_cl_ddr_bvalid,
   input[NUM_DDR-1:0] cl_sh_ddr_bready,

   input[5:0] cl_sh_ddr_arid[NUM_DDR-1:0],
   input[63:0] cl_sh_ddr_araddr[NUM_DDR-1:0],
   input[7:0] cl_sh_ddr_arlen[NUM_DDR-1:0],
   //input[10:0] cl_sh_ddr_aruser[NUM_DDR-1:0],
   input[NUM_DDR-1:0] cl_sh_ddr_arvalid,
   output logic[NUM_DDR-1:0] sh_cl_ddr_arready,

   output logic[5:0] sh_cl_ddr_rid[NUM_DDR-1:0],
   output logic[511:0] sh_cl_ddr_rdata[NUM_DDR-1:0],
   output logic[1:0] sh_cl_ddr_rresp[NUM_DDR-1:0],
   output logic[NUM_DDR-1:0] sh_cl_ddr_rlast,
   output logic[NUM_DDR-1:0] sh_cl_ddr_rvalid,
   input[NUM_DDR-1:0] cl_sh_ddr_rready,

   output logic[NUM_DDR-1:0] sh_cl_ddr_is_ready,

   input[7:0] sh_ddr_stat_addr[2:0],
   input[2:0] sh_ddr_stat_wr,
   input[2:0] sh_ddr_stat_rd,
   input[31:0] sh_ddr_stat_wdata[2:0],

   output logic[2:0] ddr_sh_stat_ack,
   output logic[31:0] ddr_sh_stat_rdata[2:0],
   output logic[7:0] ddr_sh_stat_int[2:0]
   );


`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Ptm+op+JUx/OyCnL+l866JDn9ep4ndGMpQpsNLdREDf1LvO9HbyWO3ZipvLdkPSuIU7vAaMhoK2V
ATeOYpFHMyEZ3dHYKpn2RG0iY+yVR7554qerHuoF0lZg/LvF3vXREmHTRHrfuflj3wCqMICz7S6I
Wi7KHbLeGrt4jKv6o4KhCoYFnb8gilUjMOGvrb9TlKfUP9qsACywH+OJ6KYWrPNgD1JbCbdN4kB1
0akR8nCCmewxIbvXmXakmEktDGm3JQDODce+jDDxN99KW/vUx5rdc6iJF77vD7hWb7pKpU/fPHCs
Tjf0RfHIDZhX5dez0gyzqyQxSHCMANYY/YTo8g==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
ZdpBzcBUivbK3ri/2isFi+muhXjpzvs36fdkJpcVLX5EN86AhAKGsCNh2SBDYrQDJZxseHQEQSLY
EqQ3q2LWYq0NitXLQrHPzEnyNHwRtgWym5G50Ppg9exXlOX9L8o8KaPX7bs1F1Rzy1hVxeZDLy14
sCW4lpaatswCUDuK0Fo=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
W6UYRTwB2bnhTprP+qRNFPorU0WSdAg1CIHhi4/e2YuWJC41OT8DHM6MIIx/RhaeFR//Ho8YqygX
nOGPjGIj3NM4JG6vI85f9KeFbQsCpeTBsGTMN12CGvQZVT4qiqB4lM7LBot4K8Wnf82fDpd+/Bbt
P+shG7OlGD8Rg4DkNZ4=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 35024)
`pragma protect data_block
wj5yO47cIsnl4n7r7hX7i6wJbgmNTu730Hj7hE2GAJSrF2Fh73UKtLppxdCDqI/NGEN8Gx/NtBSq
eQ/sf6/i9He9JFHmamFy1eD2io/b+hri5wxi+/BL92ZpJq7kdWWFqdOTwGGg0Jp2LDN7QyS2GztM
WnJMok0683VW/uDovSYMp8o/utGAXTmGbT1o3pd8QXw/ZoYdMX20frtLPfOO4z1hSZMRxUmBGlkH
PawV2ggjADwpsYauE/rXgJql4EyvAw4q5MU7vIIehBrLxiWiPKR4BsBDKNCmueAK8vPrjzuZOnMs
c++XEhfGidTl0g/94sa5KeunB0pVZjevO/UzaEIsiJtZRuu0l29zPW6S1k6rQU4HEdvCfAOC2g8D
cvWLyVIS/VCYgmAAtLwa5/M3qxtGn20OH+CiQnBj8Qzu06F7m6e7PiECA7EFg8x/q/uIXWPbmqXX
fqezs0nn6pAlCm/ajL2SZqG3TbHy2pZWok59QMypMXkiLebd6t4Qjz5xqjN1EwkN8anPJtyj+p1z
6yUHzbpScYqI+QlDGUXJ+lS4KukectlVVFBgYnQkgeQavY0v7TELjtWQTDU3xfvoeFfz8F11tzTk
f26dDPxJbk7YteckUpEYLZyiaU0pK6MUckPklj0Me4cy+6biyS53AgSJ6by0d36TceZAZxEXJiXi
HjQXKexmTHi0UitdyK6wfUS2Tva/HSpFkBfoEajzkzd2y6ecGP21z+TSiEGlspoHPwkhF+NihRTJ
9om03cFBx3bkSuC0AB1WtcN0Fjw7ljUOOxtYz2UIyiBzU/H3S5l4x8xQJ4R+9oOquMbdC9y1tT4q
abZy12UuBXoLYOmTftha4Juj4IbXmAzpI5y48dmHjXrPeuGpRW1bYQCbEXvroeHmzQyMyQIdDO/x
0gN4Kg9N7yf9XsenxVwUTXgmMjttWN/PBXzMHbKtexWnLJFFhSEPnTVEXIuU8xHugM0ElODw705e
M1t1K7LyWX7t0PomXdjQilyiob778SrMtNmt9zQA6Uy9bbQzZK7ZcOZve5cWuH8PCbizhSZViYjo
GgOxDNiLcFksNiUXxl/kdCixvptZt7UGr1oiep2W9WlIE6UkCRtr7vEg8/O2B54+PVEh+OfNh5X7
cdaM8E64FjILl71KQ8JRtQiKHbULmp4jvFTsEYMxqL2K83xaUmttNPN6IRi6BZKJlxKyEfl7MetM
92l+TG82slkBXbUyvRREgvglJoDWGP7DCbUH+Rkf/iYAlH0ugndZc7Y39vhVazyZWTXQ7QmSzzI3
pGzvPLlWTQpdXFlfhLiKlniNXsxznzzjJEe291NR0//IZcRSUPs+vS+Ctmqpdrr4b/NfvoLIVdIY
5L/vrmsqs6rw0H6b2fkJdy+nN3uLE+KdrsJHqSXdKxlPvaSvcLPDCiXlHAv+0+++9l5GM5ng92hx
drTSTnMCUn7SQc10xa+FdaQfMnk1X1p65iGXlBq4YFgO9wOpj6WBuEtdTpD+LGljeYA9eP2dS29m
OsmJnEZSXwdz3wzSpUi9b1qSNZrbjVv51Ci2/9jziAt9bivYOt++YQTr/4b24sZJMy+g+bqAOXZ2
GsvXHcteuru1VU87G3cVe0qgG4rgnB/6bOyukZj6823mRKhiizg4nzl794+J/FMXEE3nm1QtSyv0
SRlkYJ+zxaGKC0h3raomZLWZj02/rms7pc+8UuR2hzyFq5KezP8e1XSbuhjXb4uQ90ciH17PmBTG
A8qbJXdC5u/0c8Qp+JpHULb3y+Qlu0YoE8aYJzzZDimaYMi+qJy9vKuUT+bllbD5ZTrakay9+PyH
VYWKMx3JXKMt4+FFo7oz6UgnZC7G/RoyV+xelnH6FENt6b8IEQnGyXWNB3++E7AY2NGGqNKmtkp/
5v3TrbLa74kGpvVJr7JjR52bPhtf/+t1O7f25ZhpMwTdmB5pzK7TrWRlbpXOuJeMUlF9ZWcWYtu8
78keUVTvQM99Xn69qLMw6Jb4GsnmCuE9c/6kjD/K7ynHSuC876U9WU4UWITFp0wvoZFR6oefFjdZ
VRaZ07jBEpEmlLK8/zf1mevXo0F+BPEms/vqrJtKfAURWqLs/0IhGM93m/9Sw2dqkdUGb+2p2ykj
V7goKAh/vQvWursaJjxGekCOs7kMH6C87ubpiSue/KGG4y6pxPgI7v50RxpIPQhmKHsktpUcgkyL
KW0c34ixfHAAO5XFnMO17DCnNsPbzJ1Xn1z/KFjeOs64zSYwkAXooyd+pIZB6tRGiqQgrTxtD+Au
VZUaHFaO7NLeHCULta8wfiPhtYL9nbDntFrVlYu8UkHtCPpTBM9xAohM/3885+eDcmV0mxZlTzZx
Jqczq0zutG7fD8FFj4HkUvuGBM9wZs86nmCKxAQCl81I7vXaeP+rereUqxAz+/jHOIOTQGii2+DC
j+adcfaK+qgW2UF1cIWge3w097tKgkzUTXpkRA6PxrKvxoKVKJ78/qTYjrL84nQnHPZat19ntZod
EuXDmQRIC6knPjN4+AOcVp6RDgkcMcug/GPENMj5fr1OdtaQ2ulRatMxp0/ZK+Pt+AblDUz6zkMI
Df/vduQx4TBj8Akx0I4KK1M6+dK/++vGZWanTj09fNWIS30eNKNh4m0KiyoNoehOJHHub+5DkC7C
7IyKivlbZ3n6YKmMN4UNmeOslwgF26D53UHipTYG37k91YLobMGG4w4FKESe3dNidsBarmDsV+Qr
EYoJ+oUJhdUq0iS/rtUjEmENcxmmFZ4DSHIl27XwWi+J86y/agYSLNmpm9ivpGk2XKvuo0GDOlbI
Qb/nfdu0frBCqqTkZeqSbmTGQrQEBn2CiKf6j81VYBr4FVyUmvvfg4Isx9/DemUJ9Y0f5HvLEcK1
nTptJatOQY/vtb3O7DMcUpzrxhqsLoomZhx0JRM7Lr1xscTBBJtGiK4JA6uGg43igZmLDN77+tA1
2+tPQ7l3HnIO/hZC+oyoPpIqauvJsigfukf6GX9BQSIEtAJURGIHydRNmJk+aJqShDwU9ht0FJx7
zw8/6YlkNK8xvASfyi2iGHxpEAucc4PiiPsVvW1jUAVfoySAF1/kvoorBSNAqqXk1YgYEGu/KFS5
m641pRFlCFmLWu136r5FmDc2XNxlwNEIf4A45bVYsSKG6YWhy4dqpO7xZVPi4Z21L53aQo5wddIX
vgc816apfYQxFzzrZHWmdjKmxUseEy5ISuPXPadIcopgVHx+0cyXKyBTnnYOyOQlvJtVrTz6O3l/
K4IbWhy2y32Q3R7nQDMn/eAYwudat12TvaLzj7+5son+q7KMigTYv+w7Vn365ufnxCRBTyHan9Xl
sEpnM+FvrEQ0hf2C0FS5ZDBAKGGaBxbWeLjFj9Fm/euVLl2iuHrxQTtHFVfDoiSmqmMrE4uuGSa7
+Qplr8X2yzl1rNqQg7cOsgCFzEkdTpkr5WPujAPlOvWbmzCKk2Rf1sOckIR+zBfaszNTUOJ4D3KK
LOlUIXmgT4wmDOsccNMmA4dp6+TV6FqDex7JTy/ycoFFIPE22Feiq5hKr2M8E7sRu7OtkKPi/62K
+HDMoNzKnVwVZQsaV9TLWdMZlSy/LZHwb9KjQzO0Ez0WXFHGpRzltt6r6v1Zw/LjmDDuCPRbA6TU
mMCN/ghZaUW3IHqlxc+A8rkrfTIgujVOTbRkvILPFfb/Frb82sMgH+ThiMeVFvlqCfd222ucHHco
TwDmHa845IYpzDgy4V+AgYXdYYMDrSRvbLPN2SI1Pl6MM04ZGULimGhq4GGyLOd1Hm5ujswxns7j
kvCB0AcEwoQ7zNu9QyQxV7YxWv1+nr7ZjVpLnPaymFt5vh8vbed26uEVdzyE46Yk++KER5W62xO5
NEHQx6Ki942+cKDs8Of50yTP0YrS8o8RRkax3RmVHSTQ5SnrMPxVFBhJ1ZG/TzBaYCAx+gEEJWeT
apazMsrfSgUxyT7XND7Yb0RpUikoHK1bTV8SM6UBHyB3oCFUmKp2RNLkj86//H13YDDS28jta/9g
TEpx99Q0z1rn5PlbUraRD2HOYMq40O3KnzX0Ye+83smAfBOa/zpH4/DOj6P43bCFFO4CfgYzecjk
LpRjqapoB86vGuZhQiX/fBAaj51c0dHLG6qYq9fKV78DRebCBHOlmuKwowPl9JLix/qNWIEdT7TM
ybi3er5W0C5jrXoEtaE/ta7JDyszC+5jGxlemvDZ4cEy+lzQt8uEKvthVAWPg7Kol2QK/plDmEHf
CO89IyIkt8T7jVUNpK1Qp/enVZ+a7/RQtakQeZC8LXQvq02r9HMHoKnhUMRH9T4KFIIDoDKXlsjk
Xy4lP58vYg1tI44rHknOrTkwqQYuPtN1n3ILZy7VtwfS8NEdRo5R5etZ3Ln64ydTllErNzCFFubC
ve5zq6ukO2lDv345JvLqMQcgfhad+KccGYTB6uZ07BLXCqw9+UJjzWxQbgslqRv7+QX0zwGqlDf2
fKHO3kwcOjp3KVUSP7aNd7xFUz0oyEXOIOkbLEwhVnmK8hrSL0Hy4Z1Q2IBFUHWkFJ2gjjEg+LKZ
anqelKXcyLx0GJX7gCtZeiMxAVyZzq5FpGi2bXsWYUqUExMS2WeCyVZ7DNFC8WMjvsTQYvUyTiJk
OboKYktnzPyrr5lXTE5pDwnPJR7YFNUl2N/W0X61B1hl4hchVwB9C7sA/9i0kK0qv7Bcku3rphaf
nzDW4f5XuJ5RCmDVhYh7sW86XNV7RGUsigDWLfiq+nwv1owaiV/7JlIy/0zEkHtoclGrf3LQD1lK
aF8uP0zN5fiQSM3JbazbmJ4wOtccplxh773fXnnk/ZfIsQ5RMKsJn8Kw4rezHGp8Mlk4etDiO2u4
OdnJeeLhSGJPyEzzYR4jkW5CI8WkcsiJRTrI9LRaYUnFCuAcL8zrvswVps4d3yUoFYIHNh36v8Rh
9LJ4kIsp5iGwWyk6apWmkUj8letb3SDaRNGETlDwaRcoROKiAnNaX6Yr8FkE+xBFcwi++ymP13eO
3Kh0Cu9bmYxs27QycMosM+u4Cy0irdiptNVm2G4WBbPLUXU2Zwejt2/ZNxl6I3D3egtOyV2eU6sW
B58rjQOefFD6P3VqQpTFTRH87W7kt7bkt/64Hpc/NfeoFHyGlpjNDlYzpJKArnVGNtCQAynoJ238
ywQ+sUBfRf+BEtSjT+egABE9mnlJhMveprpC0f4rNF/hVZRdZXuWlziz+cKN2+FHOnnTw6grEHGS
YoC32xzAtQzv8qT736nBQOws8xyyKnvATMKz+fCzeMO2NN/wCnWbIt9UbpxEMGwXse7QSte3a5+T
4r9ELCFXxKysjWX7sPN0eD560G2bmmbyYwXdGQBd6T/itb/F8hPbu3qrGXP8JpJGMde01WVprmtS
hG9iLCC4LI3lvwkE3cnACx8bOgdgU4Vw7ClwBlydHaXDojMCoKjPBjkR+6xn+U5I/WylhTT33hyY
SlBWBndYauyLCVASV48YGLvolh2Eds08ZbJR5M7E9CqEm6dBsuBUjg46n3y4HslbawZVe7qnLPb8
GJg1nacC/YPq0ePBxdy3cZ4ThhfxKY/dii+mYGPStE7J9pSHsI3vQVNSjxWu19hwic4C2BhdVfMI
6KQkgz+o7XSGK2IESXHP5umD4zf3voA0CTqSEyzkaKhpH61QuqlLsrnXrVMtUrFzFbFgg/LvAA7S
I6+e6N67yYDyJxXuuWoDYOKO0r0jG2Cqyg624JkrNRmqsu37+VYsHjeckYE585XbeW189O3khTII
t5ELGdPefUm5JUtpMmBF+scDWr4vus2dgngMvtFzYcZqdOk2uNR1Mkd0lFat+HnDDu3lKt4uQhwZ
rQPCGI24Ezr3t3TPwmXXguwCSZg8GfI2R53tAnhw4H/qbgba+bCVQmS6jjkHZN4rnQWrJ1xAxgH3
p9NJmSYuzsgxXAO50HBf8qhdkktScdWQaQRoTiHDqdZLnju+MHna1MjPtH6s4bde1uDQmNTpctDD
oJ8T5P+EakY3I8TXfebp6JXb3GnZojqd0X+uCNAUP/k0pZIWdv8pJ2fIWvxakMiOVx5cBUrqCEAn
rPAwvi3VNvO0r1IGXIp+04I2wZOP9pnxRll73v+x3vkUT5unS7ImLdPbwOyBrc9bl1ejGvh1wKzo
1Fd+yt24D6KaGITrorH4qzz+++WIMZFtM77ZVfRA5FdVWtwdWx4CIhPskf63c0eWpKPyRTuVIGcV
i36sJiGJFu9fOS8+xa2dz7xkqEY5qvTt0D1zSRMhlNVB9n3cXj5h9IVsifEI0EJ/0LewP4j1W/7q
uEhOiqmLT5bt4ayLuHptbuZZ3x2Syine9wdNmncKMVRYdCuV64D6HsXURt9NULDMew45/WH0KtrB
QUDlcn5kWHP/9FyYM0/J8u0ySsumTpVsdfOxGM0jzYeiVF5dT9EtRI9TQdub0A/zTZUjuZMjAkKP
VXRxmNoi1mTERaE0+g/L1fqFQeMVcCirqIY9koVodmXPg/1U4ST7JSS4qQfcDF2goUXD1ro8UEkg
h0EBRJS3e0H778Pl9qKtFX/OMrbWAASE8U8aQnW84z4YpWWmDDM7YnLRzytecf7katOU55mIAYfF
QAqByFz3R4vni/vxLuFMP6fGyf1vDbScE9bxsknVAv+DrPditdirLVQqI/uMUizElf3Yq0tL81Yw
6nctwmVGjVSWbZIvoeg6rBDEgUhsXyG/qLHcwRH6NfkpX76x/dTI5zLpDC5JzH/DNNnub+I4vN7x
YrL7OVQFgJ7/DpdaL+9WKfEjuenyMJzv7R8U4SPMdoLs14rZOEeBjawmK9aoAGL+MpDz4L9td8Zg
Fij4DUfnj0TaZL8+ILGCUBmNX2TyTUx5nypm3EYPpNwYKIDDDSHjWSr0cB2GSotiIa3z0DxdMxVq
BKlVcCe1Az4qCNjqynh+2RMEyNO1up4apFfe0oqV9TQt578BP0hYUxWMKvOHAUFXfwF65lijtOXZ
rilUb1ZZAlhiC/Sai/3Tlb9VWf1mSFRREneZH+o0pKh37JdkXE7ot3lA7JihX7JR1LT+ZoTKoaT6
FSVQ3LbMEWb6GNGRdhHNJ9haQ5xsUwJk01ojEjVQRZ+nN3IwAg51VWZuxPWxilmx0WbtUyqzt1O7
ey58Tj+1Nyifb5lCgQ5YHymuzRIBABHzT1e9v6CZh5nxg4VEPcdWkxBEN82wE57htQQHfWjVXI2Q
eQBcqWjmQdJHHJCWfsOBLrZLtRbLjMIKyPcRQq4i9nGwWKnYS3D331pL9zi/S8VTR5ibUxrT8+tO
4SMxuweriI/jWbK0QzSUh40w6BRn3YZqys6KzULFeEYfUHSVPkT0vmebpWOPyavjoIPxxjwt31r4
G2NaVw3BqG1GwhctN94DpIU6sskSECNnKa9UR6WJ/G+MLutgzG7eKjmWDnqdLlOecHfiSP7vn+s6
cEOWvBLGdE2tV+nWAgqFbyRGWixw0sUnkY5IKL4mBqq5xBdgK8x9DQgXPMS0xyklFx8HOh15C9+q
tAfY4AT+VT1jK8e3F1uS/pzwTPkBZj3+jbGfunYuO2gExB8GHXfsA69Xt6nGMcpoOgQ7L82pMdY8
GEq56XMunXuoTXwaAdqRn5cZRFEPegSCJmV/dH9/ZFvHGqTn2xHjNlR1yh7T0hdPZvXYGmpBO3eM
7n9sEyl/iNac4IM9VC0gEydJtY1rqOWuCgC/hOOH9f1IMRpg3/yjVxfHaiDszX5ReKGcweTx3Spi
mX1WK8dxqynDAhFCHRfUiQLzsXWIG9GX6LXCCeQEMemBnsHvDgxmJ4ZWKLNoBK4Ko5SYHh4pO10a
GneR8UqcNGEOgcJx83upvHljHf63e/jHSesH3ol2WeiIS6+xXpTRjNzxM0a7eMKt7KUaSu30OBxl
lUet0KkkkG9PJj2Gxqc97+6jSYsrf9pbU3oB9Hw+JWFjO9A774BdX7vYZ/3o7v42plw49ex/RhEf
PU9xC7Q0ugY+oHcxhdMl1Q0q0Q3DicsMRcn8BqXxSsUFLRDrMGKokFDK2aZce92AndxeX/zu02Ka
1uFf7ixvbSCdnBWbThwhvxKY17dj8GXplJT7Pr0SlzG8LT5u5x6b+eq8Oao+gC1nqen09WHDGAvd
ZAcIrki18WpNVlDkCEeyzLAgCcOySyr/el3Wi4upSsTZDQKkzvPrhjujrlaNVps9xZogxW9JN/jG
GlTDuxQ5nk8I/y6d1mk/9Aln+uSy7PNK5KGRPuETuYKY7h4ZgIwFUgIAWr6oiJ064Q51wToYRur1
NTO/HUfM0xbGYJcN3HZB78JIPgPaLmPPSFruNZ/PeRYfDer9wAdOfw08kN/pRLcEVqd6sYWCgty1
sb+FTfdhFcqhqigtyB8pZRmtSn2CmJaaqV8rSBOd0eTZ6636UM5yqgVntqmvCg5BmbKByd91A9a3
+IcP7I+ScxG1FXAkZRlQUygHaTx6P0lrfOPXknGbqv8szybGtioCaLU3EelzkSzutM457kEJWZWi
MiRo/kJ+mpQz/f5gfgmt723DdOggNqzZ08z/dTjY587AYz7CMnb+HVPlWhd0/+VF4C6Ckahe6s81
d8HWN8p2msUmFaaIdqw+Dkdl67CM71MDY9siiwQ3sCREiShCJGAQcnVCPSU0LKf1xqW+GhXloeRG
VeCXKxlTqgWFu3QNsokcNrPNeAeLe/oz5IukMZiHF5RBDCkP5H540xvRiYE5YpcqYagXZ5iYgGny
fP8YTalxYhQeQ7w6Tx/wl8tycSrbb00sqg/CAMYx8qdh5BIp+gfPWoWbae0WwBBcRp764lhZv8fJ
q+dDmdLoJ9QYBM0TMQPNEe2Yq7Jkvk69GulJhz9o893Ce43SPItXe/aGVL4xp1mUQaJA3sygX6Y8
FAo/ShOOc1cH2OE9nAy06I7sT583MpkPObNNe20y/uWMRfjrcnGD2fo7GxbLEYPEGDh/Us+o7gf4
MneRSP/6NJ8A0Rd3wbb1zneN8t+vpQDefH1q8GeXXEiWxofGtt8CNtw7BQQCrXv+KA/oV59Y4XJC
4H56icR1i0iKVKmVvN1LvG7b4wcwcGy4JOHDbVOa2ipIJSFeZmAuzthzeQC/fGJBhV+2u4PzRzTk
cw4QEd3DubqYtBUmGhNc9YOAOYQcwHPxMf63N1PorK/ZNEsftx65fm3FVik4jLb6VUxoI+5juILV
FsWFfIvgifVrw8FmGnv/cKX7J/7UZIXVsSMpHGvae+Wp4PeAgZ3ySvM7tEqc96GLbIwVz0k8xsxJ
CHb8pPzpR+1xu+Yeaub9N6jfv7bpNp0jn3E35LjpKI6FnX2lXtWN2wXqy71JFXrs4MKG69uef20f
m8y8N0+GLWHSUpsbJRb0BVufOxWwXLsMtJ/p4V3YAx/v6O4tILWO/QI87VtfHpZG/CyaybLnGBIo
mY7CDie/duRwvyNhoNGxZ1ZwdA/6eeOo4vu87DjyHrglN6skv4qFWiVIaCPBuj3bnyvsNnz7CNB7
bbgKYQ3CHdLVFnWQstM5l+7FKXv5ffK8dukDEYfsxDOrX/KXEJdvuUnQpJc3vmqJANE5BQYQIyEU
lqf82svouNwk0A4l07QVkDghIQEYeFjVZU+wiQLrj/bW/qZVUBTmWD//9WmSdOAk1y24dEtyF+qv
tr1pJRWHuT2KHDbbu1gZwzGG+H9MNixvHKNfPaQaOde5CEPZ4RLO+RCEM8f8QN3a5p4ALpwL77Ji
JAZloC7i9t3nCBZYY+Aj7FFESkwKebWIe77TeBe2gD0ucPDgz8Dk0Fp7Byq+0pAHRN6keAociTYr
Mbr40NsURygMMVe0z3Y/CoHTvkIFrfkME8ir29yxNvIMFzpPKjQ5yOA6taVSjXhXp2ONN3pHev2X
hA5WuRin64G0y8m7C/gNg001GTFhbixjESHFsm3eZMhK/uA+TwOpbrDVpGtywMYAirY2blYzLkSu
uCNPa8cOPyD9bsAinwJiZfx5s/bZtY3sxZJI4ygPHRDFXe9u+xPM3cBs5xXDQT2pCU/6CPMCgyiL
Bv8HE7FVwAc19lLkG7hadcVxPMtbHR7hpLIO1biPVYkiDxquBufOUc8dBtlKLDg/R2krcB+Z4EFl
Rza6RPhOg0Scue5cVf+kxBr12bjFSFEN03caHBi6S7LyAf64lEgkHGKJ/kKYMPlSA13/Y3wcVzxD
KvOmB2DkbsLT3c3GFaD89sU0JpElAMv5LQMlTsPEbFqpMB2Kme3ZAYACu71Hhv5qBy2XuOru3acw
F8NnZtRVcdCFFWA4mMbMXYp6ernaq1ciTIxFZ1fSkKvW8NkK5hOo8nvaPXwi6tfWpqqwW0IpSWAh
hjJ+aJyT9vLPETc25uRTpl4MR8MVxxevbNg0SrduDHGD90OXJxmtMh1GxdP1nBm3X+2KgL3uFtnQ
QC8zdWau9Y4VFelerHkBcwAc5VSJZ2wQJ/2Q6frHIGRgBgQ+o8V4j0j0sq+aMVnvjf44dvn4O16W
uIIlCGIIwJddsNFIWPUAJYh5P1Kp0kc19MFMFnyosmjj0siEzR79YanmezzJ0NUMqGL0nfbtqEvo
KDYRWJa9R61iFA9xvGAvx+B9J5YPlx3iWVZwVciold18O6eYJhQwmFF6KHd0CPNjfn6qRhaHA1gy
JxUC+46Mmm/l9A9neUUm0m5gOK5rBjU59cx1JmsmWx7ZNJpat2uD3g0dGt55TchiyodxhrJPp6HP
otyI3ipKJ3tC16WkAiGEPbX3e/V2oR6/Klis3w35uMFXuEAu9XXzhxrIbBnhiR7/gjtsuDGJeXEq
lS/HmH7c9yyuH5coYMb1v1SX6dkw14UxwVE1PU1wejE3BpJo2422MKPD+rXtLXz+myexzzoLehym
Bobkr22gkV7ZPchHoth1DNkCLlWw8SLlE8HPvSrpRc7P5/21rvneKVVHDMFQfJEbDtOh1S8Cz3+q
fYusW3Ym1dPmq0IbaNMq6WHONxU/417CPciOb0+VbxPsJMW3rmt2rotNevhT4vsy8zeHxZIA2HK+
+dxHZ8zYhlVQkdRTAfAVOdLe+L0TsQNCAl48rR4tKCuQTJOizFp1osRqW00SoWYAfKfCPRw4cECr
f2T2kP+cxWg7cJXBgyCQNB/QGhAzGcdRPrKSTbEbd+GlsOlDYpcSJxfHbCLGYR7dJcmoeI06MVEl
Z/QQo+/9FyJJLU6BcTIaptPP3pOkamRuJgB3JyokTIFAzpm5PzZPL0B9rU6wOsdUXGJYlRrp+56H
NHO1zDloLKZqFCJaOzRF+Grae1gJeBXZebXmjMxyYkrz/GrXzxIVkzUezTC3j2o5+FSTUIbpJZoL
vpsTnbXLp3p5nKVYZp/K44dO6+HF/rn6XpUrYh5GAVFhr4Em/G+dURFaf8o22xQN3nuN/RbAgXmR
NEVqzZGzXoY/BJtCSuc/1oGqKFf9z6vJOPdKQq26uRf8h7f9oULFxHTP3NZeDr705Sb5wk0LDyGk
C4veSxB2d29vr9RdNdzPzvJT9qHiVnX3TkTGLTba+TtGDdW5ribjUb8iLgMU0ByRB9Bae/AN5aGY
0zS9tMSVz1irlIrlsW/geoCO0arg8T2NAWe5XdNjqSbInoaP2L4fGrQ4iW4Odo5SUzbKBQEaMD47
bLBS1MqG4m+BLz3gq2Qdi8aCnKZFRrVVIvBfOxdCeo3s1U9RqxcXg2YmBfIWEArKE2JcmySEUjdp
7ntekCJqQQsROtoCex/cLEyZkry1+vOoAHeACaYo5UhStLYecPrFTuODEUIENLxf40DsChvT0+Dq
lBHgJWjsUuRaafov0rnq/mZoPX7b5m75W7nr6vqz6BpzWzYSmEP9n+FnDJUl5kEnkoe6bMyXSH69
qeK2bDvmlOA17b+inp9AvxVCpIrhZ4iBbjlVI5Il7Pgj3f0dVNMONcF3Z+BkDpE0bJmqd4FqMffg
eVhmUBrcmxPfGBPLkSoBv7lTzNMqUgNrHalfFoXrAcdbJNcmy9kzuZW7IbwKskpdF8ZktOMxJJPL
AeuorbFuYosLJtJmO6GzoED43R61gJIh8Mrsn9+XZLUa6WOfOzqrJSS7J/K1f16y0EbEhK/BF+w6
8UjnmDsmtqLbWwKv71fxlni2HSmNxMyfxFie1P+TC4cm+lgpWJlnVMrM+O6o/YjV7dULRsEiw48e
Gkry2uC8WEbf22VBFAHLoRK+21zaFfVHzmIjoSG0TkNSLoCkRJj8iQ/f7CZ2sDUdOWdN4m/VGjYd
2E7w7L1DozRFHySejXI8LxEyDnABLT+iPMA5t5oO/BhIhcpu8P88macV4bym+HujLyaq1eUGEAkk
UPgKVe7B88rIex4tqgMCoXCogTF+j/wgnV9hgGcDktwTAqZ5J7vQcnRulrFL9CPCIcmc9tQCf3JA
awNcvIcVGIWX7E5SHF1kV2ZQ2CyCOQwpDQRCj9XvWlpbLmOdm+y3p+X6g/dO3RDIZyCjNNCLHCeC
SR9UUOEWZ5Him/cCOwMUELZwAcTK9tz8yRasPL6wP4Q3rjz6YBvvUPqwpd4Fa4A1DY4VD3IjH7MF
cO6Mm9cVdJ4D2fvgrR+Q4qUDj6Bqo64tAn8mgqco+JBIOdQ9CtGcAr1QcsvClpFdb//P91cU4vdL
Jed3aIqLWDb1dZYeiUYGbmdHeQdHhQHmOf6Lqzs0NJWkr/UapeshNxXUWb0ctbvO3R4vDebrA7cC
mqKPt9I6AdILx0tTStK7nGh24AE+gXoAu9E0OV7eV1GZfvyUMq6bLS57NFPEt8HUu6Xy9wTW96OL
oR+P2QjqyUUij8+beqWwv6gGrxuYk2Ncs+h7nlUi9PiMmvZ4blm4RLgy4WLKUx/Hcuyzxg8eqPXe
UwwCD9IsWSUIEWSH70pubMCxnLuGfIklnKGhqZJbGexdoAwMqNvuVjJK+wj8/EYt3Q11a4Qo01hS
YVdPrYTF5/CrW1AEJKb40aqZFDowtAuzzrYTTnO2fT7g33B01BJlBAdw6PvYEOBKhOocTXHEUgaY
9uAG37c+ygSpswE0Z/Im69PRl0RVb5VPuqe8XCVirIm6gdw7wUYZqbifZmEstM07UcSe2pAIS196
3G/dfCenUoUFYNs5Dsvc0s1UFyTdfTn1fvpeMNXwnjWEH0/edQBuZ2rbLmBMRjGQMI1VirPGDjnq
U7OSrgOnN/F5Y7ds4KuUapdY0RclfdZtzL/V4wNqNSd/nzJ171TuiERDeA3YTzHsBTVhjIorNUmB
sJmVANQp48PmX5VMVZrRXgIN2sZyD7A+CgFSV7jkKtn6G/jL8HO28ghbbm7RmYZjVd+AConXYBXT
JQWBLLzD3S3Qv26qTO03SSnjT3yYmYo1VdiiHFbQOIpYuBddyOk1fsvN/s4sNHprw45O2UuovAYb
Af2kfB6kjYPe0OIGm6ApAffcsKJF9GCnIUv9fa6YPAmPKGqbRbHheN9TSH7ESusdLSWvqBxXx4r+
Vh61QseKwDHyTOqJz4agvmwptJ3klh92FN8IhONUhHAcJKzPnRqJmbLFuM8hP5U2LKbL+NRg7k0z
6OlKrvsshyIchLdy45I3HOzwQZrfrjQVKkJJwaqgY4w926R0cflsypaHrPKDsw0U2Hh7DNVvVFSQ
R7BaR5bEEei8zWan2NvfOK/qV5p1bFjB2hXlkn/qdMzcji0mx8GKVoxC7JWPtTOpNe0Gv/nJoGxG
TSTtMscBDvFAsoi1dcO/EvmR0y8ohZTL9dznhm++f/C8YYtHnmmAY/tr4Je8JkspUKtIawiBCBBC
k30dCQlfo8wnR1ZpMJyCA15D3OxHBXaEPAxmfVtio4AoqfTx2lOnCJygw72lVMN6iBr6ZLSFRnfk
Mg6HkV2MjCELFzi3O1o2LrXr2JmH86n8skPRBTUhopGflSnhlKabMrgk9TK+fj0ajJTdguiJHGxm
C36Rysh8mi5r3nFSsB4j8hLLI+ZGx002wujH+GTCTQZAi41KhUt4UctD5bDQRR4A93pMwRoKV2/2
TqoURqdzBA4jTzgkdU8B2sn8gZCb0znL4HsB+i6Nrq1fqjZTYCi2vxzie4tbYN2ItMqKr/gmjtal
/zCP/XpC5e4SmvSV3vtmXkEPF4KSPwLsmk13yso80NZBiezJL/KwRjeFZEn9K7rocLolCtp4q1BE
fIENWcx6Yj66BpkxO9T4DnDYOhVZtWSWYtl7GlcQr/7TD11TD8rxLODTtbgk9pBapYXvSbCAKWz5
ZZSmTLJwb+AW27PxpW0/XnLdkpTsEUJrR5Ns9nYSKjX5PI4ItqjSAEnz/lZp0fAJ1aLwtWjU+iOW
diNrCV96U488Zq13LrBgY1xy+YZNhwPmoK9y9cnU0dxcw9jRVn9KgMLD5i7C82+AXj4U0XhFsAYl
V5Z2NRpSyM6elux3oR6cmqQgMccd0IbQvc3G8l+XnTxAbaL/pX65w/zxExJQB/LuEFvP8zMHf8JY
DNfwF3D2bOT/EszM4huOWFXjEWHeKuQQjuw6s3Ys7Wcvqh6PfbuvpNuEk0Y3j6lj6vaZC1THXJgm
HW5c7qyuDIProKo610K2U4ysNZkFS1jmgnv/uXgXl/fjUPD/piYIhmxX3yZ2X7VBs3ljMkjxKs1Y
2qGV/fZovlcfwpmq68RYoM2pnkm5G/GlM1caSTW2LCKjxMBfqUA66lnj59zSA4tHcozygN2ZXxGy
JrkfmWCxUSsrd4jX9nMHxyWvT3IUapKRJ3i4l5upWWNXf4D6yzg4K+KwzIwVND2gFd7NJASeCk4P
p4+ki0G6XJ/JMWzlBgBN+x4BbugGYtjZlka/Sc+l/i72s5tOZanitSNB+kUWO5Z+d1NOq6DmY9nm
/ecefvf8WSfJuP5Rx1aTJkwWp5yISO1DdrWICdyOsLx9DqdoR3pv3/yrpyKQx20qAxaLr0EDWSwI
ciZUISqyBDtnDJDSdPVtoeRCDKTp104YYS51pXVeNdtVOX0G/rokVNWjFTS4eEphf9OtOyzqUDXM
Nevso5UfQtEqBsjUIUpQLvwDDU9M5+FE1YtsCDWpRk504oOpphD+Y6P4I1jcPKWWYLWhl7xHOzIJ
gCl3m1tbJ+lXJOjAh6C1T9zSIEvA3ISSeeX0vRa8ckU/bbkrxF87T1irc0OeB6oVQ+FdYnU2AkJT
kxvYfj3ucIaZmnXrvAVRmLFRotVlipScFrwlWFmKx7+FrflO6CvNDzFl221nvVxQmsibfQODpQqM
ngVgjfdJMJ7Wy507GA3LMBI7gbaK8Yrihps/6eEV5SmWd73/f0Bayfs0LjgkA03dpsa4IqbvK2bs
2NnA0oxiKW0ptKguoq1jiz62J2BBhPaj3E0bR1W6AG7AKISBLIV666HRUXQPfhmSfUuwj1AzgRC1
Q2q5qs2T+oZPEUnZGkNhTM28L4W3PD3hDuMUG41Q0DJ5mj43xiAtpl96tCGSJyKfyTOPoYogyxrO
urzpIg1htPaX5z3vt9Lr9TN4aThpXSC1aufgey7S8Yj73qibk0COLBjkgq7Zk4ZNumZKVTuL3Hvf
7kp5kc3BE2cYBs3UBBPR8IZbeUMd8ZdbKqJQjxFVdCTQOf1Cqb77FjGHQ56cSDwVxcbWpK2nnHBf
wDR6d3AguFmqIxn0LGpHajQs8AZ/oDQ0I/vIdhde6QnKjkyjygRSPTCsbNkU59BvzhdhWZX9Ctqx
SdBY3leuFtqvo9M/IrXMSv8UNd9O+uKx+xPIgchr5rgzeBTa2RtyDvfgFnes0hloGYTjKib5Tg/L
5Gvh6ctbN9Pv3xYIkYI6kee+GUZmeYQqpMHAFnHAIJYoDq3P0TYCfzOSp+PEPCttnJp6GMZ5Z6/U
WMTtZXc5xhXWNKybJUMX3M3t9ZC6s/fA/tQPYJAyqD8XwCSgcrafHWTIuB0Kkf4nsrbgpZv56LAd
ZnUz1waqv85U/BMh0VhATeVmqRYWan2bKff87StZf5BQm88/5MxHG5pAXFXqbPmw1lVP7Iw4uIQD
nvCIbWZCPKN2hfBbOncfu8ekcw9bhB4lcYt3uDkvea3fHyKmxoOV+TG968qpUTA4jq8CPUP8lhZB
J6FxR4mDwm75i7+hLbS1dvh/jylUcizJrMCcSt3oQ6XJ5V9vCpzsKXvnrsfp/PRGNyInrhMaZiNe
EGTqZ7NfWMAY1aSPfqDL0l/iH0U5lDJbvn5nUX1Hb+2Mgj2fhZzcUOi/9tKQ7GT6PwzX5dM/8lRs
5qScWaDZt+lTZidgWleDH+9nmJtXL0tbvB3QXPAFNNzLJ7zIaI5vJV6iuPTJzaocGhAehED2fzHr
z3CdFYkcfbNQc2iDdlX7JvoxDwvkYHBys8zUNq5nqM01fkCVR9tigEPif3VX2j+pil2Fqkz2Y4+d
7iu8zL/8ysmNCm1U2t0gRgVIjShxNkT66RuN0gMKwvnl54MaDlIoLAFJFwT/Qc/2vCtVmsUT0f3g
3q9t82T6LZHWukyXji8umrQRK6/Jom3OWK2J7uKUrEQS2EFVyy3i+6mruNpUfkDVsptfuSbo84v/
0bJwK1ztoT3swm7Wl60WJcuZTooQ71seVZb7YABUMbpjyo1Yk0E+djl+syfF7WcXhW/1dAkEUKp/
4JOc7xjoSdTcp+zfPsUUOFp+0av55zjNOUBTS4ST4wAR8gg6q+I3/ekiWbNx92E7I+sVw3qHAfAi
0Sy75mYXbgzQpgSjHcjukErlsoOWn2sxHCzmMPcfMMU7yKB89IqLOGsZK6tW/OkuvDR4k683VXrx
4rfjOKAz6EcD6eboeFvDeI3S7gQAOFAdQnjr9sFK+SIsXpMSg9ADc2cm9HFSMYm1/sPNTz2uU4ps
ZOKt58zaTC3junUHKfrlDimbq4oH9gdCqW4mZH5H2nn550WE7Y+EMn0qK2N9t6NtFNfIAatfocx4
/mHwL+qVrkGCVrSiRceebsQLw0KwuG3FftVWFWMPRsd3mN0+T5qqc808GclDTb4BCsNWGU1zXhUF
6lgzK4oii0LJ0hVSl3M+83KuteWmXm+N4WR59n8qbTi7T7Yzf0Ju90D6HcgnYWeLuENpgEPEECHO
pi4pYbgZlDnKLb/degW04CGI4nPgHKpZssGkZ7pwxcyJgdpwLESJ6AxUugeArBkIlm70XYFXzBS7
IIsVl+VXwDb2cz3B9gLHYzqflHoK11C8B3WwoRBU6COeloeShJhf+esG3QwaI6pFQ02EpZ+2xZ2l
wVIGgTCb9y4qtMj1RMz0jRN1/zBoKfnNx/E1/C7X/3go8EC/Z5VKwAegzDevHFOpn6gTb0tqXFqb
8HgCoJubHCMcytO1Xa2zhCU+zF6poyMHXQdeMEa6BzQI1Ysy18IcVyk49sB0MtySxNhJJ43wpZ3I
0CohgCNr//JOIFOPSH+gPjadml9h9xrfOqrNPVk8a6UjzFlPaTNxrlxI+zmt+bo3cnM5vLzQ6Mp3
xVnLxfvRtLogv5JNJyPvzK/BIWW1ViF795W2og9YUUjeezygZ4RJGWdUzOqJuJNhJLJntGHpWndM
bB7VNyDNEmgixDtNHXIly55RecKZPE/PDOOznzPofcv4+FWlmyh2aB9zmRAuvGcm1TXBCZXfKrKD
45Vp6BG2UfUdLaKfY1iB3DtRlpsyFyI1OgYX2X38h3Wtw0KMC2SpDu/BK3PvBiuNn970uLnRxj3R
cFtAwqoP+97D3GPGsBCB3iAI9sPyWvUA7rtcB5iVwPrir4VxQCYJU0uNQtPBHD39/bEdWlg7tIKq
tpAtS/H5icTzBnXSJDn/TSPE08mr3JxyjeGwiNpZ14qAzaDLKpqGgoljn56A/fwtWHhUBmk35gy1
70uxL2ySZt4I6P/07vX9Jr0MhyIJAzTnQ7L+8bco2MCx7u87vN03y1HlJF7ZV3O0MGQSnbhdFLY+
oIkRARJFl5niyWDlILLQtET0klXycQ9iLO1tA1NdK6ityrd4AMR/RKOQhmpQm0+hJm/FOTQREdBO
Ri1fml5Xq7/EaYPS8CLa6cxO8jdKwdjCJsUc4yIlmLhx3KKYwgCz4YR9P5TNxACG8Xe71zc84x9Z
LtFF+TUTkNgc0Ii1U9w+XqPYJMekfSPyWZdePecEj0Fzia/sW1ylO5+DeWdjxQ1iDbo/y+OAgZna
c+pbDAwFtuqzoymLspKMZ3vaJ+Ap2Ch0YGWx0jQBLsRoHxZfLta36opBFgFuHokSASakg13slyY8
HeDalTH4F1MSLQyOvBPC7rgnhilcgrolR30d5XWybuWhYKgUjQx8Gk6gE4VVNYQbyEZDKtEXOPqF
M5pKimF0hdMdZIqYiyV+xNzmkRD0XqQihtkIf9T72p6C2iX50xauVufDLssDwsGR4clkp62FKOC9
X0NDmYC+4LTWGB9uMuvSbQbkb5JkhjJn9ucUxSrbvWj/geH+fFmueUD4HWAMRo7A3QJLoiSvjWy6
f5iBaK45iz5xJk0JQYe1b/0QR7hWOex/hdA44hP038zLWSUe20sdZMY+Xr7F4Tttv4fRKxxtWtFc
ujrPL0zAojxNS0JR1K5ebM9QJMgdIiSBOmT+h45cyYoopwDOSXj77Yu83ThgpNL+wqHMZRTH9p+7
bGMKPwwXcGyrgQ6GDgHkN+u0I1O1FPIdzTts3bL2pFYeqe4pjzphA8fhI78QiyCVqZhFsLi73Zmq
Ob66hVIOJs/68w5HgtQPkezBnX55/I13T6CedCrUfqOfpDY+9LjFH0C5wW6wUmoYwR/lMBi3lqH7
txJ6xcr0IHEWpmGwek+s/l0ySewCg1XYliUF3LDwel6bRzPDOwRTorTFbEzYX3zPRsV/tZupjvuA
a8+ztm14iwzg+uPC0VTXHaBAuaI9ezT5BbXNRoQbkTmu0ruwl73wWJYoYzl+Qfp/90w6TZ3EpUMF
6K5oQeviUh6UQ05fcB8mAE394gmzCP4qCfDENLSglnstEeG6rTXFIbth3yfwUVbOh2mxajFpBGpQ
etIMn/+Xs5R9daK1BS/4oTnLzagmVvVhIsvIWAhCoODCWwRv5uCKmTEgPwA97Yc+VLW4H+t0sjhk
E38CHKxRIkfd4maQ4gYEk7iI9HayC4visMI/I1XyfU5N9u1xwgzviBvACEnLSoz3Dv27gJ0tv8EW
VvFjkVpe/Dp71T7fDgnG6Yk82keOnUjI81KE+cjhS7p+qt3cbnZb+vCnAkgaG0/1ebIJ7T18Qn8/
XKg6qsGWpitrtsffqD8H4T9g6jXic40FCk46OnXOg+MDcYkFnvZvpOdjiN194mUfedAZm5VA/5eH
jWzSdUOUoAQtbB9BZBdt1FjzVhNaQB6UyaE59D3vMsghXO2VxmHzgJdClHobosumxAa8RPLXhGDr
UmyrgxU3H6R/iq0kSGXnek+163qGDDVbw5v8SYPMgKP3/HokZQYpPkRaPHrHQQxAxDNviP5gWmaN
tgRg9unSBEolG7iUc5dAOgFbjnh3futK5bL0rH/GDc18qpndcW0yzYM+puWQmzfAUF7PrQOm8lro
Ldiby78NjmqMKnnXK9Sn4uF90gTRt4qjSd68keZzIS+DpxyMgzD6BCbcfEPqbUPGRkquQWUxYmTA
LkpY7GhqraSW/XPHJ2nKjhSNIbPEiHNQNlZbvhI+x5g5/gCOVg3kQHsJtDXVW2mIms5YVsp33Lb9
Rbd8OJp4Wh6xiigWNA0RV198qcm4B6qgRX61TtznBpHM+4Q+gij2Jo7f2KxFxcv1/7qwHzg70gCs
zubUPDvQKoHTlMHXppm43IYfjb7xazIGDQpqg9o5OKXcve3TjW4SRNM9mHD2s7HXPXz4huTH6sQ0
HXkbXgo6MIs950qGMlAkBfkpLK+rsTyKWFBhlgEzn2G/Hnf/r/FgrsDr3xutEtvKCArUVOUGwlQA
NyAV+eXTWXV1EMzfSqmmZWcAsKk6qncVKz792AMwFyGfEViQTp3OhXwqAwEiH/CW/bKm4jSB5B++
03tDkE9EVNZgk69EOQ02bzuNUsia7IGLHmh6Dy7TtMyqL0Rn5zejW4aJqySxq85EnQ3haA8vJap/
OBZNouIa+eUwRIhMUi8YXsZF03lsKF7dI8m3FdBtppaN/qk9H3OW/eZXy8+c+zmesN8Oia0DRehU
RegB2neoORCeOM6nFSzxRdGUtNYMW2gd0uk+nUQ7Lg3Zg+ucp3Colma83hPGQHf8kRXOzhrfE8JU
dYi18qVCGAWAYSdLBBGmJePDK8qVlsM3+Kuryfj1edgzFM1OJvDfFgVUgabq2WwxiK9JmGbotuvq
3TmwZum3R+2+DE/oMZMFSC2AVmV2wr0edqtXgRVVJMeYPo6V5dJSMm/0Js9hsFFJZxOmx6TIsWYR
LKbguePw/JIiDAgrZnRh5/HxeyN0QiGsZjtS04vPQ+AMPDeeM5oau6ddkPYfNVE5LO+/S7uXcJcD
Zrf6DVjfYNmqtuXb/sqHHYudKd1HDx4g42DogSXdcoYPBmI5aRUjWdtlt52h4zIa9CBz7yKyDwFi
TUtReJ399MPAZhLhCdmvcs3AW3iHGGYGNCNoDstFhNnqgNYRFw7SMpvttiZlhk0KoaAHrbjjKBqO
SxzJhd1Qe7JAj8Q0D7v/EFKJ9L/A5hI0on2eGmwL6NYkAeJ6hiTwUZ2nbJhc/wd3na3VEq52QsMx
G0CgfesAnLQXvByXV6528WW5SjxHDxqdWYu71OkR++dgoLrVirs19qg6lARl/1g4ppmdO5qrmLGT
FX2i0X4XYWS3qxFX03sKCmP1Gk30HeXgdfG3GqvGYIv2NdhlaNRJidkRLBeL9m7aw53oYBHfbeEW
cs2zpl5hEX4Al8qtXrBVCEA48TRP/SigHEdmg3CY5OHo1pkKkpkLo3pzotOIU8HvoMWWIOZq3lYQ
C03xu44SRzlJVbPnvuQniP59k7RbytiO4FmHRCfu/yhpvFpad0FEOC82vzGEahPn5+LHGGDR7ea4
iQFovxAPaR/n+kjenrQ2vydRTmQex4xKPqftgO/FXcmvYQXd34BcAutrrclJd8QmCpF/dktlpbDn
1UAwGLtmU8PHMBqTfRSbP/54jumdgLlI9D3LEjtHWs3U8QbYrZy6Jeahq93p5mOH8Qsbeb4o2A6+
G3TOaSTXoPGtN8DAR5RNYgx7nBYOWstjISeFVSMK/70XUgY/XDsutHRvf4Orz3rpkA0lNk15pWUF
uCQD73JVfs3PrVtYAVh/2D7/cIVn3TXdHjfWXojPj/s6cHQh+qbM8r1wupRJXUEezJVZHTa75fTA
h7ttevjBspSXZ5X6d91DsGC+NQZFK5HnOPM3a3ZImAobrnj0O5TkhoPlC7LGl4BuzmtljYoNfkHS
FKY+Kuo7/wfFEJFUmfXd0bfZpAVRzPZak60nMUHXk1S9IthHzZwtajiXZFa0pcLgG4azXkrLE53V
MWln9JZzQOWpjbyo3GL40fo01D7BtBoVCar3zDqeKHW2GvttV4lLD/sOpmRs+BujIKdA/6Bg42cd
wiaLYJf/R1xPjHjIDyMdEqlCIgnuV9Y7qXf+9QBMO21odE9uHQz/cccfzJAiNGHjWT9kLXV+G0Ol
ckdWcjOF8R4pdvli+I0BGSufcfdthPzrRAkSZSqAlTFqCfQV/eoEFhIpsvs52a7S7Yte+R33YcYz
08FS4yiDFTq/KSck/HMYFDkWlD5Gcz4jus2EJXhAmeayqsq9W3AqN6srWiXp3IqTjU+2jpeDd8aJ
hTcBv2PS/Ov9s0SpwpJ7MDYS2yVPjIzxSManNY3iiSZkGCOG/bZVJuzwJ0/K4tU8qZ9X6+1VMdhD
C56joZSgEjTpmRTVBsxy/V9dRxI+MRC4zsWt6HioOq6veIY8AdWVa7HrVUPhg751QzVcgaqKlw4E
yvHhZWIyVW6B4ZQrFCkMqKDgRtYB4as6pLbsJXZe4MhaSrCyE6PrFWj/VlfVl4HsHEABCguUmvLF
PIz/LTdYX3+iAX02QsSA/QY5WuJ6EkljuFZNcMp+LvKnd8hGg7JgSzW0KD6KDvV1+S/2JQ//Ov14
bU/SEM5MztG7kKxmQaHuyHeg3nC2LLkkh9L/NlEjb73D247evcF9xH3wFoPxqtKcgU73vuVIZsDZ
u4tEZVt4EJHBPI5I6Rjn7cUhS9plnmiuXDT6zl/SCMSfXV78Dj/stgZ4qsuh1JyE0T2dOftpO0PS
SgLyRGbisdTO7ipwM92WLKjrrj21NJtSLIb24VW2gSor69dBWia8K0me2811rBYvIt8m+HSO4duu
ijzqKv8jTcsmXzlit/Qqfgoa3og9TlLs1zaErK0J2dEGGkpWMPFpd6GA3ksZM4C6BmDkIP/ueIKF
CPmmuctRdvPFlKLsefo6OvpqPECl6PgUPXi6CF7/UX9lL3Lpvm94gunY3VO6H6tmKxlgPi2pTuS1
oXCE2ZpfZdTGgDarOBYodDjBieE8wXUXeq384Yxmpha52w87Xg2jsJjUpCW9CBZWy5Cyg6C2Y3wt
5++MI/vahscqLMFzZbL32nX+PwGeTFZQslo+V4JxIGainuh0j9BwWWwugfYLkmt632B7nJl+L/oM
sJQH8jpzBYxbeQvmyT3T6kTU2pnslwjE61YdOIO9kPzs54EXlcpgsY8p4HIjsl45J5afg6vvUgTl
KRyi3zh2NAtOROGt7mMOydgmvUYa4ABD4T9LqDsrDlzUIUlDB2arq9OQL+SoAvDBnaZoMGnrXiBp
tkDrBHXEQQF2aDByogaD5e9xj9PusynoXpVkZON0jxVaOkLgcljRMF+PVkrDrfys+AnkFJZk2kbG
EYyXLXOMuTwWcvNujFEJ0wlbs0BiJUHTQ1H27SqWC2LUq+YQRZHy7ZxSPQwsLEEYb2wJemmjd7fm
1FN4/1LnJmVJwjJFfjp+jEwdJrLzSwsfgP0QEpK5gvJud60WidKN5xxO1nJt8UANNIALICFW+iqe
elf0hyHR5soc2zw2Pb+YJ1jz1JyZiG/fdQMEXT7BToKOHyW3J69AwqwJ0daFn7Mklto9OFKJrhtY
L2Hb986c+Hgf75X5Ti3/cfR/Ge5ID0poSGHIiaRFmK7yze+8Jnc8SBN3h9PnxL9Yj3FYyFle/LCK
G4fR6dYpnrYUsWSY4aS2LHFmWVQHUcyjAtA9XP4E9Ym6v0rX26MOvFhSSCrtJdGbaxT2ekL9DI6M
tNH2odNdIAc83FRO4GwuACP7t3WdrbJrl40dJTuGn3tL4hanvoTzHVxML/HCxASBsZ5CZnMzkZAz
7RFoQ1DojXrpbxx38TC2DamjmksNdNC1Y17d0GNRr8BqDh/BPUDAG0PHhUIBoWahsXZ1zGiOua30
xUO+E9/FJl2Fi2CmndkpS7EzV45G5FKiyT8yxucI+aIq5N15Ok5Qhk7crSlrGCGllVzJOCGwhD29
CHTL0+ArJpDtd9r1UrZI+7fv8UKG8JC/6kLwAM3seuIEHFEkWY0bbhu59QiOZ9st5sHGbh0MSqaJ
i7fEkulL2mvftIDwLj7LJmJDYnEh2F2WtC2Hllo3mjJOlob4axxUPhHz0PSaQQh386NPWhrPfZLT
cMGFRZpM8PruZ5Y8+MJRfjlfHcKTyZEMIk0wFmGHMfkNzwICVz/4Kuj6vHHdPTwtrYzLaujIxe6q
g1HLYioLT3eJwGy3ADfYg0DMFOfkhJBfKyTc7DCmJfEH8v4oOToIRPFZ2Hcubp/dZeY1/U59V1BZ
2qQ8+64j+hERpH20tivWBZfHJs65nmYpZAdmfQS+k1RZ56lfq7h/1bHt6vNsXMgiTZWkzcFQ1mYK
wAr8WRtrZmXyA4hwQ7usAkKaamWfKY5/KL3VtURAg1qau3flOnmcQdI1Myv76ujT4OBSdNhPaARg
+vNefzEsixv1VtnSU1edXUZrIYEz3bLe8V93orhVq4f5ElhNWB30k3ClLVyNDYl3X43lTT12UfI+
uopCFpaoqd9uY9LqzBAqs8AVPl33/G+G5m61z3MmbKaCEcCML5oEctY18Fpb2sXDfMC7XtdVRPiB
b6Kvqz1BoiOs5xnrFLldbr7PvFM2DIUVMbYJ0H/ydCVkDfjrtzxv3DdQ0wcf5llMHoHZWI2ZInXN
IYE/htJ/gdRl9w/8rQP6oA0liwFOJGQX2gbBtdqEHZu6/+4frFDmGYQyHENWvtrx2PEyafHZS3Z7
hc2a+9kP6/qeFE0k3Nird7I93htUfR1DgpTPLEgtfOkEDY3Gz9x/Cc+TIQMvrfxCskySXaHibtqa
mO56s4OJ9JUGoKsIADGKyfebSCBc44B5/cqAtngZJG3kAcDUmdD8uOpvvQVEndOy6gnKYx/hU/P3
R+nuYaqQaq3AfHrMcZpnebzeK0NasOkRygiN8sjfa3wE7TsNMfGqB/vBQun0MHX9Zzwe0MWHrW7E
WmWAFgG+OFocbtSFJ1WqTjl5+CLjC/RebtIUHQSIZhzHQSigoHrQ3rQFTG9qcySrKBKK9bA3drOc
mvnGh2+oGAoYipWhmlNrZvsWhcbqMDqstSRBfD/sdwleXUmlDTak53xMkI3zNGHWtgQXzVwUKjXe
2F7QblH4sOORTXlRy5Nc67Uq+zBZiriALZJ3XJh8XVcrWWTc/HyHG1zb9dxPXMZVVB/Qmwrwbd8W
vIZrIdArV/74CaCM3/0xxlcgk6Jt7SU7NQ7xgH62/lOo8d51HONAwktkZhLU5zKOeH/xPmmLH0jj
q0x8sKDrsiMnb4Iz4wLt2n8ywGF+/M+0x4lSX0vWwicGw2HLPp+sXPBVymc680ASfq4SwibPvWWr
Lqbeoy02RFpIt/XLfEMjGd/VIItJKyDRWD/yn5CoMy9Hk21Gad3WmllKHcP4M3QxO2b91+q7w/Br
M/uq4L8ASupfFAfMCdcmWTvat1PNr82sqBp6Nd2sULDy/ywviyWWEcjovvJNniorij/hfFKoKzrK
SkbCVfJlduyXAyfvPh7fcSaSCCtGOKtXHxZJPo719FedzLkTiTIMYpDQ1ae9vceNSbvUtt0WszvN
1kEdW20I1zOwXpOTQ/+bvhfMk+n154Kc1cWJckg8fwMa6pA+EDKiCWPsfwRKz2roiCp2JLbZrBmB
vmnEV1y7aa/AvRw5Km1yO3W5XY3nGKYl+bydzsbdCKU3wl7My7mcU+tG/+dCxSbVTvVNkncnhAW9
oY04fnd9m0LJJHViXsxljjroK86SA0NFC47juYBEQmJ2tHLVm4+vjoJtwEi/j+S/NGv25qL70jy9
S7U4p8L4jKMMi2WXtsTwAD6dpueNEq4s9ltdCtxh+pJNUtho7ZsuuGWJnoWLMeqwI9KHK2VQHsPh
fTQc6cA6dIHG6Y3zx3KfMpJUEV6zbNM6MpBOndvbTqEdHYIUCS7+u5JCP8O0GGL07gZu19TPFCJ/
Tq6y9JjZBoiXatH5WDX523GqduRe2z8OzUU2xxFeAGFq1NLPNnrbHkCDcBbjsHGebT4CyrlHEYW1
TD8Gu7MgrME+qyEh2+jLvV7kubJt4iOZIjxsdl4qulEWVy6Uo3bySnvp8NcX/xaiXrwczNVp0EKt
c3UWehDWvKlneemsfPqFxKguAtLFDacx7sHRKgKGvHl7oXnyS+7qTkWGqAcQ85VC5O8UvyD6z4FE
JeiBwNrh8iaHnaLy7p73SX/EUSXTVcqRJidasYUx5LBrDSN+y2DCR+iQ5ydg+gJVbXMwq6/In/LW
vm5a0tszvu1vN3KAhArBMWP+gFH4Vl/3QhhYRdObBx/n6Vujb/tb0wTCxctuPuB83eenHllGTWV+
1eDEkzZtWhHG167yKJHIGm5qhnYEfaMfjJe6zFxcgmjyYrlzFBY4kKuSX95JiIJPSFAFrBBF0HDn
IwZdunum6OR1P91TtF1T6oIxTvqrNUviBIAZ0sdJrJ9kjxZtw6TyroLfgXifzemHZeFGTEF7/57m
lyToShSiRBmnLRf8Gh+Xj4R1yxssyI/z5VjFVmrwGD2WPNd32a/vIWdnn+uTYUdu5X/zrGDIIeCa
DZblFPRbNOz7WJzmlfMjqEQ/1a8ndKUamYinrsJ1nLtxVoWRZxZl3YgjzC9grzj5Ri4v+5rqZ65i
dE152YOiElVfxR+MnlfVbdhH8Sm8tEhNfqEWi39IDMepptrrliu/zZfU+OVYaqDDaPoMOb00Iham
xRhFmFPtZWD9EUfbkLpytDcfQgkR174S3bn00RZlUrUijsWkeousBnOlVQ2IKuFUqjLvNvXROs7l
DjkxW9XsBKJxxpDan4mdOH6+Z3gpzJzrtwJsb5f7NnSYhAl4ZGznQpuPwCBJki9ly8tsvrt+gjGI
uZjssrxRiz8pfcMLbLVTHEu5Nx5KVS71VsxI2YKTfjBA77x/9i0LshFGK7uj0Oy5WgUt4qb0xs5d
8/op8Ck+0Z4CDANwKQkrLb84IEb4CtF4fygcDo+XvrlNYz+DvE5NVJH3mnGbg4J+6ROy3deWTzf7
IIhW7+kxFwgbYR0Xn0JYEHfyv2QV3lCWQlKh9KsZI3mZ31CJAjvNN53dpcFJf6spVUEsX6IJs76V
3sMdbNQtRX2/5rcaT75kJmjISh0t+jnZKroNZgjkvOFO+KBcjdv6/knKJ4yNu4qyqIr3L2Y3ER+L
IBYhtKEEaPUYeUdcdaQ+TJ/4rr89lNCy7VVB99sXPYPVDfPsyH4no9tl8JKtmU5wvwmlaNO7pVEQ
edgnHj07Gjntpc556ZHO4EWInUMflwaoOq3tJJveNtHBHgeF3e/kUHtyOTFcjp9km3VaJR8wTXD9
u8GYfBQljmgP9g64X+jVCnbTikCkBZZ1l1Fup9bVUuFHwfdPuAIf/UUtmXbCFwSiWAuDE5AuX6aS
Hn56TC6JQWXRVGgB7ts9gRwAu9Vk6rA70A6w1MQ2GfXw98CdnZpCDUrvSirwFRYtKtesW81Hi/lJ
jk/qfqYf+y3SJ8tb4+Qi+mVtmfXcjZiqnmlUiUjn1NgFamsvfWMc/gDnsYtN+GOAc/NT3h9BSXff
iR/lc1CryWOGXySdck8sChr9B/kDlbFSvNFjeKfT59F+Q2Ra9ls5nzJ4sPtkhVFPsVISMONdGI82
vtmFFk1cBcZc74wtrqu+mKVuTZNoJQMMsrjx5vSVxm0XVMVLpTJt3r0fGLkU1ph51lQH8IdvIR/n
CmAs7vRxID/ckb8DLCFTERbki0oXJvpqCJodM1jyZiYEkvPrah0JfDz4mdnBj1hDQU35pR5JUQLl
niOfbPP6pd+xUyj1MfYkNW1HljEcmTF4hUL4LVCm0X79mCSkHxP/lkXSy/IXvAadKsZETICBZDJl
mVRZJz9rX8fc5qF2nsw4xas1pDdQdlF3I0pBcCjoFwq0W1ux+oO4br0C7f+XB8gEO0J28CgrF9Yp
ip0q5AQoai2+qzV4RtrrSKirjBd0ajXgErN/bTbesjfSQv/2j0SK7OhK0gtpg8ji+U52RwDvfugE
E1UCKi4Go3zMqHPFpUkwSkf0PsXdj1yuCBCbE0wBypMuqaLcS6LJHIvQ6G3TNGYHENCuUp2625hn
7hT6Kc6nsq2c0WGCW/LFqJOgOyKZwXBgSv3J7HH+f9EToz0VaVgkAnX3UnlWXpL2GgD5qUg3AVU1
G8ov0oN9flD33MVIRA2d8qsfLft4fifcnxWIbH8azPy6kFYQac7MVwdqrUaaxEn8+3d9poFuM5Ng
HvPaNBOaq6jSUUnAjrkTncItiTx3X+dkyW7a4eb1JK7lhWROg/EXPRVGRPgIVFDTaK5/JUgRvqGq
9haBYJwM/i7AOJljhRJjYlgjN6WePec8FtKlqtQS5LkD+QCNGp/C7mUoQuCC5Nv8bT4dJCLdWXWf
/vanIGjVum3i1TriiJwBplAaVsoILaOv7fqgmgCB9qKFHyAmPLpduUmnFv/zoVkn3+CAQSWamke1
mRZEY2BpzBduyzyCrprtzxMHf3U7e3CiFqNxUFOLsjvcWe7UkjQrbsUmpHWdemPvj3BYdapJH6zh
2Zd39cH2b9IOyBGHfUDnS+IxnO1P3tiy1NMJrcP3Xqyych68GxCvdqhJa30WU3n+0cV6x9sUJKLU
fhd0R4oObRHUaGtQrC76a6WdsByIOoH1qaIHOUD8yRVuoVG1xfnJhuMMeiNaZ51Fkt8eU0YzHuo+
BAd/oKnYicL3cdlZi5T1vTenxoJdTrHE1RBJI2uVGZOZ04TFOQANmXEjFupVCUTewydmz4X6Ii/Z
VQH3MbjYcOGATmxgOeJ6XV1vaz1+1r7us+gN7uMYxJVpfD8hcsPZqIPSS10IyP+0T4FcEtss0P4D
jtyadxddTkeKw1h8c6hvejNvl6QR67FwmnNeonQx64WtQS+ULvxuSYeJ5LG3bk9UknJTuIsiFRgh
d9RXZOQR5IndKeB3L4gfkesLG+YmqRB5N9q12M8cooKE9TgljuUdeNfBS4sM1If6GKju8/iS5YrD
DVll8wgxYA2hvpsq+nkjWS241PLPapnO5KMQsb7hm8RQ9rnn26HxomJqe1rJgiBePFAY63n4jVtx
M1P/OzuhJPk9yhrnsqUin9fJFHrmYOE1hzgmqD59YgA5WMS2iHTaxSjcUQPqJ7MUoRVKOvkoNM5s
YdQVKw4dYUyM4F+w5kZ//r59jboN0y+ABLZAMiJ3KXgo3RaEdpAOJcBd2OLJ6+wz5TWGXRnEf47F
4TaGQpuPJ5qXxwoxOCVWhEJTxLnsJ66A37ukxjH6/hUR+76EQm78g4OAq8F2PrShOpgJ+GoSnsip
kSQAzf348kesNmJCe8XnFi6q0+55s799KdhxFCZ5MZYHTyNbZrdCNN+CWu0gOXcO4hY8U36vkcho
wSBdnC9kPIRHwfei2ib7fIcgeC0lfUXv0Sen2uaoh96d3ghcAH7jzn8qyv/uHQu5LdvZEu3hyPzf
4LF8cTEy1HI/dCxVTxMFsQhkz1Izvkp6wHQzZbxQwyJf4CJ8eTuw9aT+QSEDM17ci90/kGG3tOmU
mIYrI7bBvl8u/HoXJDFlt9zZDl99vOsnGTNjYWh6fenKrKFTs834W7jDQQ+iE27LuKIIqMyQPgKX
2bWgf8xW0BHqCxdfPf8/EnhaKo4O0+GXH0e9tk69q+z+gGNKNModDDtj5z5HvcQYAIO3lC4O87af
ybBCZu6IRjTSrYk2zTFNVUyjBNBkOkLsN2BgCXY671oY6UiIt9SbDVR6l/zy0YfDbT+9rdCuMPIx
iYouubo7cFJUqesyKsgi5mpjY4HWOmAQ1uvZps348IkijGj2mLlQucnrI7zdvxJdOz5MEkFFvU9U
M0i6x402kDjZ6FmBg9LmuRRDSdn7l2kdQ0RDK5YwdnJW6xC0dmi9qiTrTdTaSxjqHVimejB2Qds5
C/RFFp0QO43ARz/KPhwHlTRTTZVLjOWharZWR3LoKKPVqljNjYk2cvOF+n8Q9iragarkCQ8t1Q2W
h1k4JvedVdASY4THEbECb2hKaV5ZJXF88hfKPBEIsnDzQ9aonWgA/9Za2tlklfrbV1NQ+7JBvDb0
lQtyX0Iw0tGQLPEOLBceGKHetnYYyx4n9BS8i4Nw7nWQ9eiS60SnTUNo0SBN+7fgyz6YQgV5ia43
BAGenT49chRhNqfurgH/wam7yGu2TnhlvRmdrziiVlBK5Wc9Z9KDadavprF7qKjEo6dFeoMHDaxb
A6UcD2lDDqn4biQSyUbSxns1B7NqF9pgwTfLxzQ605ISa7SxEhp8uZuDMPW6UMuKk/gmDY8g19l2
6hdzZQM6tHXqH0n1ZlwKp56MRdiGaK1TWnDZcNy6hvqfO++iSP7DuJBLNKrl4uRQ0IJwLH90UWBQ
XjkHeZcubCm4R58wJHZjhe9QrH1oJXC+6Loaxb4bEZFL7A20YYzz8mDGXW2nA1m4Oo+tbyMXPJzL
UfN87h4l6V9Qq9L29sEXociJb8QLgDH0GiyuVPb3Uu0A0ToOVXJiKE+e5cM4P39CFuRKJaM0OJJm
UV4qgk67VeMRL7u7/H5VXvGXyijDtnpZVt2TrVsroC06eYBH1X+JX5M0QB+VYU3Movg7w0oyM81S
UXviSTUV3jQ6ng0RxJcn1D+wtisN2dY2hWcSRky+4kwUq1dVrb+rda2HxAlmpCrrUvSGtuWod4CK
Am5RU9RBzFsIFMa9xdtFDznifc61twGLx5S33DPSGuVsKKmwHaewZVpQHeLAW4GZAxEgUF7uaKU3
afVrExz8MorSvunbJFNEG6Fu8oe3pvQvlW08e820cYQo36Ux1M33u/3SeMb2/jOdGjewUDuTr2wU
ygcWQTh82NxpipxLnckMbfVl5rZqKURuWRz0S7Zgheuz0aI30jtnu6uBfD14mn1LHIZFI4IcaVYj
N8zhOsGzb6/0/8cQbBMCG4QcVMaAdb4jE5N/hXchyol7qWgTadw5ZKKEXBdZGXyE6OK7AAoOKJl8
OTip6g9qEmCK3GvkyZDNvwNtNEin8PMdoe+68q1M6xUZvFbPdK/9st3PKrhhyBxGIO+0nx7xQIW0
nmZpw5vudM2Eb/URo3ufzarkBQ9bhV2O7ZawKS0CTuVIa6HrQVVV5b3e0TWiq/f1dlxcrWRsFDD1
RcF2Bm10ymm6gtTTHzIu8I3su6ggNV+phlvvQIIlIZVsklgrKjtixgnjtgpIgq4rEU8+t1Jlncjh
QCOTBhUhPAngfBJhTcO9kxQzi1x6fRsx3Ih6RDs4+MV0iGxJ2ckm2iNJL7NOxvvFRkoy2NASh8ur
X7WWYT2gt+uISrXPCCU8t+sCmCVPVE6o85wjRr6wIU3kpIbliVD4koVO2SsPMlKQp6f3bV3366d+
qMeErVFvwlaP9plCMLh7+bJ+lkImK0ToqyvbMDupMeOR98GqJcsi9ZHZpSU5vAk15ugBcbq0fZCR
mZQ/zdkhUfCPlNezzP/251wylYR7PUnArrTwfEyk0AX8UGtLn1xUQ3NWqSdkCavjAQbpY3/Q+k3H
ESQQZvccXNro1+O34BWVg8RXK/1h3W6A5tP2eBjFq4ThINJ9VD5nXvlau2ORzGT1CpnmhKdgSvLf
KAeFlPiFqcGqyQd84gEpMLkyWJzPjd10rXQC3GGe60wEPz7GUFJ9TAfNCxkWHALcQB0y5kAHK6GN
hSYCdEG/u4K/yMqCus9wxbGJN2vHQ/Ot74SObb529nhiIRoEBAuZPJk85tcD6quX1d08B3yMOkO3
XVG7yKI70GEnl/e2HQ+BNbZ5oSlR35i44Rlh4URS1cERLw5V4jwvPW+ESoSW9aw6YpR/a2pLGLGi
0yiB9vm89nsEoQ6wqVG9124K9xESMPrNR3uU9bH1HFmwwC+Coj0il8wEMhn5lIh1nD8m8RLpgw07
5IR0kLmBrifW44UMxLrNJszMDKCKKbt9B7Skg/rKRZTGja0NNrzciuxSfOpcBjVaHH7FCi3xJQLS
gWH5fQqCdT8UuGD7QAmX23LCuzX7STzwCVZIK0kVqAlfx5ER3urT/JMXxE2tDQOiJoCe3RIESTFF
xoTQoHxZnat4BZacZmapqb3OF3ngK7eVq5bwbam7Oe//bXP5oxsC9RJUcbN5WQON1mlzPIzJjPBl
RNYzmEDDyovE7dA6+0ZvLJTI6k7r+qSeTTYF+PjpFGME6miqJ6PCnV+uciNZHkODdEANnK2X78dG
qmb3IaoFX9uq2ORIq/mnnbD9vaNkUwjr5EvqCNf5F2Kz783ctWXXprtUcKMBVXQKS1rsc5a6VgsI
+pRnqGE/37TG5iK767lAbIsZ98Qp/6WssdGL3t9rvQZv7HrHyvZvGA4L4ZrZ23bmjwmk9BoJH3gv
sLOEByshXSXGgh1qFh73lr4ZFjB18mUzy+BLVjQWF/5sKtM8BNxt+P0knXcflztg7rkyAK1KvNfB
dmMoiWRy3B06pWWp+cU5LRZh8FcFoMhwU/pMUyBwMLYkVKGjvQvex8bw3/SN4nyyHU05poMCxddi
LDVi5CtLvg8ISMHna4V5/Kx8HA0oR9xoCLBB2CKzTGeVYo0bK+4BUrSc85rse3jArfsxKCtTJYJK
u6sswuKNhWzgM6ytN+UoMmSGXxuIkfVpv8rGT2bY6V8rvZ2Lhxaaa78Qkow5eAdDF+jJv/r++eVK
m8aExEgYqZpVhkSMYgHWN2zrEqvV4YL10Jg5XbBxmYKwl3DXyo69p8oR8gZBNdNtt3gKyWNYqWoP
/oRVxLm/k5Q3/JqtFZK7EF61BagyWu7m6gLrPh/hloNpiTeUspO/lSfX7imKOOeq/paaCedSlm/Y
qu2t8QJs9t+or32zkIo2tUFa4loVl/wC8XB6PuKC43ZMmI0nry2zbXcKG9fzNkALwhlxGLezUOzy
UKZHGbT1xeeIRnVFCHt4ib3HxW3K3SXjWN0+z0ocW4z7g0PyEcMd0niBl+kJIrv0zYQlddT7iL4a
EG5NdM8NurS0Nea8Zmi9yn00FJW44FPXMv22M39MpWnZL46ybmz7glYPmCITw9NzNPl9X05rimKE
QdCGT0S6O8DSSh52YVRePLcsefnbSYogsQW4mvR7VueVGHDMlklBzlMC/AM9sB9xOGFsXGghGfJT
ilSeYpJAjAI3sIr38JZt4EcJVuO8LpZbl72Kx5cAIYi8iX6cd+HqqeDFiLr0AlGahFI6eMg9x1Cw
eo1iGL3tKkqKPCQhYEBDVdzTmwOXwWpsWY3k0xqU88WewHtt3XMsJT+4zUXw0Duf/QyU3d47uGfI
ZCZ8KiGXLxfu2v15PGcldPrYpP8y/ppUFvxsCxbzfApcOv73Jw68Ui6/wPNLZQvzvhEbCruLQW8y
pbrXhygNqekFir1EjNRSljE4exi7fSN6nRTMI4A5dtac5AckJKzDPiHpXO8bvz94ZiTT4o7gvJH8
8dloQEAptKhG4dbHunDj7eRPJtHqY442isZ3t4uvomhRDHM17VN8iu0ohcp5Zs8XZ8D8gdpDUgJ7
Ps8gyCCOrpe2TQOPwmxcXkKDn4aCEbXuvL5IrZBKOhnpuA5+rQYY4+DFNT0uvqpZWi99k5uG4gO1
2baRE8bWiE86vbbp1ggT+XWCD/g8bDCOQGu/w/CAuun7qBUP7e3x4kOT8UG4d3j0ZzKu07h1dkq2
AXF0bG74JzI41/Ze8Oe7mtaA1jgOw9od14ColYhUbD2HrDHbd1kANA5mo0z30e6TzxXm1+1L2Lsw
Dr24Ud4AGrTDi3IXnMVS1reKAXWXjg3BqQwTYgVr7z2QORiqtiPfwA8mE2khf40RFHq7rnefE3ij
D/XOfvWT7gMqSFaOQhCPb4j4VmP9BQ3fxZ3ov6OBTSnWDnPRxmdUUkr/yieXtLuJexMX+urDMzQB
IBA4tFEmA6fhNL8Mz/XAqwKXs6lkQ8d4/cgbIJ0wDOLD/NI93f1xBon1j/i4BYLGV3A0Ohh5ZshY
uVWM3McPvDuCc/1UdLON50GuPG02A4ZbewdruDa5RK9B1fp5V0cPKHzYLMU7faJufI1y6zCdvoSF
1f2jJEsHclASNU9ZXCOB3rhaysP3ve/MbJeyzH2myooJCxmBJbV5ZTyF9aqgBdQDMK6rLLFSGRcR
lJ/YF0ofhM97du7aTzIciOiSbEB2tIJRA0lO1Vd1eAqfNNyCpN3SZ2cCh60pij+sBDjFx7Pymmc1
3IRDZJcqnQRjhAO74NA8JZb4Ad6kUANc/hwCuWgpcsyJvbiTj5Ycpfg5PloHZnG+eVPHUjim3mXa
uFT8sSlTrivtJ4GdJ4FcPzg/vcyXPWC5biyxwpBFxw1Uux80poY3pWx/L31zu7/85FaodivqJHQO
oltU8lyBRx15hFy8Aamz4kerYwbWuoYrxq2GzEEjWVevtbgM349p8IkNT6+emQHc0Nw/fTUnzF6f
lpRMTjf3mIdRVbalzEQwowFjuE8PMpFBIJd9OZMGxkxpd0LcYBvMWIjPNS6xp+rWNDx/TO9YXq7W
5cYvfqAjXbBgJUJsvGBx7MYanZLLQKr3q7Qn32TvTWv/30O8h3E40mqC/ZCsDL6dYDXY2P7JEF6j
sPbTQCUA5ehs/Q+L+nzlRULdxts2hn9NJw9DUnkbytsAOp2iZfskZM3/j1tEpROBVtnnwTET1lSG
mI33weP+7gCbpWvdLmT0QmPRsi+1TlxYl6S+K3VULaAUFf0QCcMZF7PdHTRBm+rYaHdoJdBZ6cej
WZjJKs293ECerxbZe0CazPvKgugn+nXJiegM+ujjPqn7lE6v+aIectgHcuD1cbnA/8xzKE6rde17
YynEKHOOgPIulnJnoalM8Kk1wU9xR2qGRv1SNBe0L0a8gEkcPnal+zs5fwxDZBcE8Ha6O2S5rSHQ
RwK5uZK2sab3zXpmA5H7PkqKOxBUoMJea27gW8VD1dISMUWaOLWuldilF//JZmBwgrUT+ZRLiIFN
6Kh4WD1U2c2OWxI+f86J0KY007XHiv2XPLhphvd/AIUv4jZ+M205i5RmQQG9MDTUcHwlS1NSztFx
8WtTganL/j5pOgvShpF2liyhsxWALngdeLDi14jtE+2TTbh5EiE4vnqgzLUZ8lLvzTh+y0Bs1bzE
NtNRDRmZEKbbqUcyyFfGFipvkQ/iv/12dDcuAQW0EIm+oU4JOVMat/M30+RFzVvjAB4Z3vhuke/F
82rgs6wNokJLmWMwREaE+aue0wMNsNUtf54O9wBBxtuEdV4eZIRji/5PuUb/v0TKmbwFRP34Z2Qi
KPm5x4EyyQz/lJ9og1HmJsfmaaEzYUaJDGQh+BUp8G1qqE0DmsEwuP8tppTvShE0dUD0tc2+MEkz
lAz9fGfh8j9xsl/DTsv1RJ/8VkFX8gj1Mvk7V3xmrRccD25dQLQxuPjAlgNiZbag0MKb7il/OY/Q
hN6SW3cnv80KmfCpWyOfvO4tt0enmdq/b/TiGm58yItNiaF28gwRa39jMVZVTn3Ajxgl+yOARGEq
IE8/eUhSPsZxDIEp6tgN7Tb2l38Cc+mCdeIfsN38YZ1tqyKITF7ybgHPiR8OVUylP89BFrP3vtjL
GlL4bfvKDgGy3OLtnmC1ECnZyq0InagJvisT8x6mawPu4ngq3FzIGAShEEY00XVgG54WVVA3lXDW
D9zDp1+Jl4oenXquPA7fLf5H4cdY2hD5ELplINkMAfakF5gFfAsL8WiRlOIrtYAUJIUGoS4C3UPh
jrPkXpo1UNjhOEKZVu/7qlwhFye+dt0pBcMd3/Ct/aICFQN9FCjmlaz5kUN9HblsGdiOhElTxOUc
yqG4mnbIwm/9CT5E7E6EsWOwibpuMrX5qa3QvaOY8Ix3rkRFesouhr5Fm7EaA2qlY9LLWqa8wT47
LL19RJJfQ9q0Vi4d5WHxbZ2TKnju5mq73Puj640weQC4uRty220V9855g8s5RlUCDPtJc0bs8Zkp
WRfTiuyNaDSxOg6AT7gIv73e2NSTHfVpTmafDkuwnK3PUF8jCgkXyNED+ab4UOHVrsKAtkGiwNMq
rbEDVE9r/tIOH6lEXeiNlTgGyVKNhCEoxZ4sS7j1HVnRqDSnEXFvd5Vvc4kjhDjQTWlO03LdMXoZ
rl4qu91vLlsaQILKPsCvpsVZVvQWjg1h8L/nE2LBbTScD3LpkP2sI+Iz3EnZHGfd/POLaBPIXPON
9POISCaBCnUZhoLXvbJaOlUaFJlRopbyi8v42StG9MoYQVLcautUcL/REpN5JDzredASWYy2yKsI
iL00kuRGZJf+ROND1Kg7/ieG3Iui/Un6Xd7zRqL2Nt6vI8T1qWihS0nFX6v4wfByaP++Y5PYpoBd
qCT2J59VF9Qc5yjqDREi4w28Aa2tm/cPTsDJjj4K5RhH0w6kWbSyZjPZBP5bdERF5RTm8KUi9Dt3
mWdpAAYSZw466h9Yyan08oH9rkVsakTudR3B1ZIZVR/Kp0Y1Y90NYW7ML8qYOXOMtfMXRYy/JkRW
3g0bYgKWh7MxVVQA8c5Qy4av5x4R+yvbUS+VNB9oP3m7clBP0sgJan90aIu9/y7GF8RKl5e1E7Ph
3D2g9c/xNBpEw+TQZ+W5jpBjW9v81fHQ5k3qzjOib4L+EOWSHunLSLK3hio71leul93fGAKudU37
jTKZcQ8xTBHMdYrK2W9f00oae5V+Ypuv6yQhtadNV9tXTwvSB9X9NSYzLMVlwN6UHEM8ZI8O/X9f
S55O0KbFiQMtH3txqKMA8SYJ/kcYZj9GssCo5eX71hKGI4Xl7e9AtwG4alBCLukg8/hLESp9lReV
+eLN2+B6KjSGc50ZrRApaXXUuHVNmwBymdkCMzRhgs1C1dGuXWV5xWARkhkz9M1CFufmCV9p+1pa
qM6lbl9pODslpl9EAgzBam+HibTU8iw5qZU3SD3rRkBl5xjXdGp7Lm39c3ri30ndQHzhGQWO9eEG
cAu5uEQaiO6AmolQ8qUWVdt9XDZGFJnMKV9rxrICVlK5dmFbJIbwVXFMeUO6wdPydSg/y8wPrbQ5
uMvtPbkAU0qfTY2xfa/frMbS089/GSHfmafA00VEhmtoYk06/44tPmh0QTkKXCbjPuzXzAszmmWq
M928k6kivi5s5sn3OyGov6YovfQwg2X/rEAm3DXhIua8u62YP7hZQZWCJasZ2bhztvqW4kuNF3ly
4FNnjSxxnev54ZeVxi6sadtrynhgF+Zm6nQ4uv9UaqHmYXSca2UGYlCBcj/vUiFasjlLxHzjqmcr
nKSD5oPekX2hgC98zFZZ4mFM8ZWxO2BopShy6De77wS941g9ms7wCp1/509ANGOEhopt84eY9832
zFYzmqEXAYQsrv5Qh3nMXrze9/gIUTmAr5Z7EWwrLBfc49nQHEPhh0bJkm89Wy10IyyoNMOatUJg
Gsx3fXlzHlkwK4mC6wNqCkVZOdlYywrxZl0lDUxcroWNaqE5zt6aWqr8kwq2S756wwRJ+ahgXc9u
5oFCd0I2ldvEQ4v6pA0Ix+yel8jZ3Ejp+K6sikKr/7QV3QhpNeWs9H4SDN+nY0U+Yi5tkmkNPySl
iTCbB+Ccwu5FcaChTzaERLRJe4lVgcDAfr3xy+zo2CFX5gfn8zzpCe90fz8O1oyZk8Xx1bM5ooJU
Ppfu3VLraljTWednujwMiGer9Y7FkFv4xdrTF+daseE/7+HRaM5JnmGSIfQWLw3aw9zDFsSieIpS
zzts9pFu4OkToRico69IVO/dLYsqvaGMMWMjMMaG3G9RNBJArHj12Ccsp9UDepNF+Sx7G3VdHqsD
ys6Zqj0/Hq+C6eBk0ET8pso02PqlbWGELbY18kA6tVS6RBbH3Mf9qsitsNOnteh9ZoTh+UNJySaR
IDOhBQaZq4Gr2jfB1gzdiT6p8B7v/YCA+FWaNnWWaFd8Sl3h57jHvLdOfUO+uSgP9io82oAdyq8v
m2tHhiCODNGugXNkm7flIZpzlq0r6L8EWBkAKsa2gEDEnkhsj9zVfPIHPPuVzVjkCauwbgmMkwGN
gO1BYYGq8kmPtP6SD6KrInU8AdvVAnFMBRGd/nF+vua8nH2MH4owmYV7T2fW3imCTsNDEMcDxAMf
ssbIBJmPHpYmlp1BiCuGHnYA/DbQu9gZmHHWhlWacJullD7xukUffNxyY4dpQEQKo1p3zfJq2xD2
NAPBe3Wj0rodjmjaF2unnJzwptyFsWKjLysluhUDJaXJ8TR9jjq0PL7oBwWLqVm8Tz68WSzCF3p/
224MvO1wTO7pzEpRFJBqlN8/C537USXK5oMeUIPci3/yEUKWfpVgqRgviQ1kmTkFguvUsLCwWmNu
oLsT5yi/mzAEkl9Cq6mOIBqDoQbwjq617eIa8A1USfnHm2jO7c58XgNlecrWc8/Qd2EGvyhIqjYh
JZU/yUOeScBFC2g6hyCv08WJIwc7eYb7FnTgvBuYHtUlIbjRzsu3eZYzDW7tMjqD95QZ1Wq/ECAy
6te1mr1iiPidntSHsrvyOXC7OjJovNv4cG+CR+0UgV6ZipZvIqOjlaKWORmmtTVJTdak+rBvUvKC
d+ceGDdRLvH5j1ZjEHB1hSVOPG9kQFv6Gk30qK2QkqBtJyLc2dPt25+nYgB2GIyi7UlY6VcyLL+v
lbmmTeNjfZlqhCWuzEDshfqQQUlEszsItkcD3RqL1BWwt7TtF2LJjN4IN1op7N39QMhVCB1v1ypD
OPbkMaxVARbuTiWzCGq5ETYwP7vXydBXcNcJPeLgSEl9r7IYzyVcqD70QMe05fTU0mg6FLAUUE5b
NAfBzTQPRkRrEy4nYWn0KN0guA5nY5HebVtCALFX+smfyj4cYv87kG/K8kEixcTe/52K+OwoPAm9
1DffQeVg/RKkwhsN5A3IOjKLOtbUQg7lKG9Mpe3ByeTKOOcRZbKM49nfEZsWFf97wC6Va3cnEyVF
rJjPHvWr2tLD6R2cP3IRWrUH6/0EPNbj5PPYbFvL986jYjFjtjpim3J6qhj4Jx0E48Lqtw88pmFu
nyJjhbbXRXxNZTmY3Bxhsir46g7UxjIPtIxGjOS0cZLEr6xhgA8cRARPG4Ogk5DOHlCJx+jV332C
P/ckGX12KAA03EReCl/Hnax+gF57V6pIDAAJfTdTx8OjtolwApVY6qDUf4q6xWOWDCCEK6srKo27
5xZcOM4AmRINykK7xZsdS5PbJxQLM7wAaOb/hHcd/opjE3oVdGn4n7bOExo5b+Edl5/RJkIqgkbE
lroLLLrPahllJNcHtkKCthMltnmnY407qobW0/faF2wgJXxnyjGySTXLPvewFxeGbuE+KlKRzv2W
GlADw9jjGVB2DZOu6CS+ZlKg1wNzW01ieM/0o8HhYYZ3MXOLbMwZGTHFzo55xYJg2AhEll0VeVPO
z+RCzGeY6HuaFiuxhQemkCKeHh2oZMvFvlbPLdkoshSLkS3yfkaWYeOrZe9vdAv46WCY52hlNKgM
HHEnOA5+RAHV1xnoisdpozR1Cvh160yX0jv+mQGsRfCYLPom/Ll7XObwCOU8qW6J2Ns/kOJ+P2pM
gi3XDB8hSMbfLRKehDnmJpxw9Nuh0HPrUwTpslr7YAml6eBAxMy+HYZRGUWiH0XEA8lJaAfNQcxJ
5b9p+SLzkDuica+K+99dmO9s82RLTrTHsOlsP9uTERm3NrVBlgnNHLpBEjIvOSsbujRAKNExFHWC
VNMa7UR4ttVKtSy3ib5iiU9GA1Gyo3RVwAob/yAfM7skL7UkCKm8gG/s046xnyWcBhQbsQg0GnOP
dkFWN4PwsW2a8t5GfHR9dAvglTM/nXKJkDiIi8RHnIbw+S2emD+fL0Z4YJL0io1pcbIoLXGTuj5G
nn2T3w7bGUjCn3LocM6DX+T+NYb4GAVkXxpeKb8W7tZ24nwjZ31Jv8HuMau684ptrm9zOUWwSgJs
5e0rYFQexid5mHBClGTJstiyjaIy7J9BeFulnsIWpGBcnZs/3+jUWNsVObmPbwkPgtmVCEleL49s
FcnFJjI93hCd0qUxcEoRbC1bKLKb60PmhJa3ljjTp0YQtp1nlYZc1FSm9cYkBQRe5Ud0QfB8kQoF
YdXBGKyG2c2zCLzKbZLyjTYy/YNYbnOeXJ9ivRv+jP+iiqp0eSu3Pyg4MMxytSUq+ovR68PIQquT
5QDQc11g+MTtO3NUvaG53yPVUg75odRJgT8F0sSML3xj94RqmCiNp9Q7Zb2AtnS3PXLqWWcfu78v
X94f6GeyfODVz9RJavAH6Y3RWqq95dBVKQjbczKzAry5RcXBxIVWV3rX+WbWtCXRCiYzpxb2oTFO
9+XWgiLIOkGODM7io7GSWVTNeltRamNTVqLfd5K+0/iduZTv9A3JUmtbgUtQ53gtRfGcVzrmph1q
iav7ZVaJt+rQsV8CY5OZsD2v23Zv/hHIas8xvNjX1tu5g7QxRKD32Ge7PEfXG1f7JHTkzXCypTMB
X1ikT233ZJmUe9zhjArW4XReFsG6saVCSld1kjIOgWy0EEi7Dxitrguwni0t+0kf3Ex6ap1NK6TW
fKRSJsnqB+Il892GneOtqSlW7nMHGXlGu54m0HTOkwQCttWDOxJpcwL0wtU5Itds4Rtcc8zPKRrY
3Xg9dsFD0q5QgKcIXjcECFOJFzmSLfmfZ0IvnN5DqmJEXig0lbIDUsZmdZ0Q5pu7J4Fx2q1yh2Wm
9AqHS1P+gQuk63WFNqmFrvlPwG3s3Ee4EJoHwFQDpeuNn+p8+nweKjIQpAdT7QeBWmVDJmRRhTsK
YuFFDMec0xhP7gdrqDqCgz9lxl8KedEytV4rr3xUnz5zwoqmAjawNYG9vARB9JQpEyDOY1HcTRzf
WMoLWnKh9bkfaxRekg5hvpHDtbP/ncMo2BRJWwgvVfTywRBd7owCtM4xusVO/SPrMsoYcUhrVktA
ytwNe2U0o48GWJO+G+O7ZoQ5XoI4r8Gi7TRz8oYcgAsSc67+YF4pCb4ZcstOkqhhjgnWySb5j1gk
S5q96OcUblRMOS1Ho5dUsIlbpqrFggkka30vCJcBPh4x8pSWm2Imq+DCxw0XRGQNtGAycB1LuiMk
cYhQCUgdBS81Zqrb3fr7hoC7QHeAhnIu2O/YHqp4U4bKZNesgve15bF+8SkYKUqalpv5NCnrxwSc
gmF55qe5UNX9w3D4fHWI8a79o3DguYzSdSDigRf8oD0Tq7UA98CIh6kwvNgopsqA4DhT4JajV2+5
E4/evzNsE5mWPBY6Lm9R1+tPZtbbM6S3VTM2huqOEq89yEl4PocXJxIlW1PPF97QNtuNJb99Zk7Y
G6F6dSe4nTZf8nlJgs85KfiJS5piINK1Spblc5shXhGU4hieQApLhFBoX8JtNgeOYsuAKTIbgGuQ
H1gaE3+/onPn97BV7Pl0K+OyO/aLMC9esIHF6WHeYUeyba0RiEW9Lc27Y/3sVRVqUwh6ucVb31JW
Y0roZBuRPH95hLQEleuWz7WsrQztRWBbaaOPMseIHOfj/7Btj128jeKdKST9ITwAmuEWXknH9La+
bDLG/LmL1jbf0BfwP5EEm9i/ZteKHOstTwGp/TR/Y3d1oDTxZe/MCqY1k+2ypTkTsrLG/ak32Xtw
kK+b5A0o+S8LAgcoDUucx4JRYbfEUCBzJJta30e82D+TVA04Up/Wne8mWc1GIVq/DanLCgco+A6U
ysGdBSThPIE8fbeDnVjawxjZynNklyWICwnVBAUTQMhzYUMNKqgdtY/v1nUaSzR/VKeYH9wTmy9o
wVpYUwWg0jnNueK7lDncuA2YVa252oknxwekne7zikM8hhk0sIypeNyu4oOKqeXKccQSeRp6tEOj
7gCmdXZOHJcd+aAw4uXBq+R8/gAVTRiuCTGGh5LTYWbGi2vNiIqolc1W1vPwk8JGYJyioBFV1Fg5
YEEul5wCH8QJnDNnHOzSDoM8AtrPL5a1n12e0EgypNo2GMnbB4F3ZSAMUQVYLC36TMD2yei8TlEO
dohd7bFV448N33mXkPXiKC28KhS3jK/Og0Ycm1JPZ3jHWJUm2zlaj/z31xPFbz2Vrl+nKGCSwtn7
D9Xqm2UINsgL0zkxnHdhhxBTx6ck7yjkK+sDEe+nfu9ciEXvRWMhTNdNdxBtfuZ7VQd+iqENdQra
OzQvPLC11TsO7C8izGgJ+eolqA2X3u8V546JGTXtrKViAr726VnFZ2yvftRVKAtIt83A6UvVPrZ4
3cKqfumm7ZCX54aXQXuQnU1IA4kfODijDheQ8Yk/SVzdsLFI9NGSVpDh6U4S6QsP35cesMnxNpDB
DPb6INyqGXj2n7Ws3fL2KOnF1gbKo714zdyTym7oYEOVzKORNOW+C/smI8edgOhkW1IeVF4jZmbg
sKSStEOZ0CkiERio0Hd7hwMXp2rc2fPdKYHebli4kJAVL/CaeW3yYHBHqBWNIn3Nct62zQCmh7E6
aJTOUzC+lOAVXVqHHLRESda2PKdoi5KIz/SqA5l+3ZPxtsxOh5madiJ4xMw6PkP0uIK3Vnh/6SrH
hSuGekcLIVJrGqtOYykNfXoTx2d2Xb4/qxxToQR4LFAmk8GThOjOXjjxr0gJ4Tmfj7XT3rkH0FTu
pfZ+DkUmLlZxVvDEYtzA6fcw+IgxC+wPTgBMgeO0+AEpxIfG8CoWvg/uQ4OVAhd3TmvjGhyNRRLM
y60Y8Q5e4XV6R6hg+53/rhUrIpUG0Vcgh1gJcyoEZLp/Ha1muuhiJBosCJ8CQto0F+R06wxxJHsk
QOG+pD1zV42VXT/GRTPJjhbgY1AdM+cug4Sh9xTtsbGn7u8WLk7/ZgMH0JNq8jZ+PRcWgw5I+kzl
RGzD8nbm1qAmVTRhh7Ac03mn6RFjFbrq4gSLfCSiFvEXu9lf7emyh2JQztp57sUSOvO/oE3IrLlH
Oz6ASPsw1vsqABZWCzBXUCFjJu3W6G8L2Pf0JQ8X7igx6JCiIq2VEDFKWqDTtmcLjnNQdZpP9Ejq
SMq7X5/xQUAnRD/OTitGrV1j4WogATtvh0XEtUHXliwEqjW3eLbiXBM3+ErNP/uNT2nhWNMqbXnm
gGJyhnC5mC3QulUUrNjEt84EfoMLB6M0nCR1pc6v0rgGFqZ3hIR6FuU2fnVLqK1bBl6TRD2C9WIx
VqIT+cmO6bjLgCnshFtEqyITpGGYHxxA9LjVBXenQMLutTqtiOVV7mOrFwhDN4JYGmLZB9j9w7jI
n2mXOlZy9CwooBilgJe7ka5SlV4rRAt/hbal9lBeuaKg2RBjXR0ZC7MEq14BfyhkOVVS6fanGMTF
W9uRAPZvIQkW3DzKMdKCYXRrB8uFH9MeNwt0ubjEEdqhutb8WRHAq22jllfd2SXac1TUC2iFxmr2
XLGAnrgMmicdJp+mfLR81dSPYtE1lkPi0zm7rtePYTc26s/segZtQk80xtuacQS8XjvdSC186cU7
dpkFo4v0sdR9A7InpM3IJ2Nk4M2ixgGK0Hp9k2mAIqQvog3izbubT7ZH5+2/I7bWOkwqrFrAtUmJ
vRpg65N8WQNb/CRMQ2VHhxBUjlm218DaCzcoQDclmQbPlcs24so+cakTng+mPCQXvqiXJ8spj8nE
vhXvHQw/KDAP1vn6TjMPuMzWECpE5HnHME21yGtkOcxbda00FDgMiMw/dv4Jm7YVwbGahq+5ZHgd
fb5vRt0PN/VGPYzg5VUo8A5MJ+to6BZFqYfcc73HI2SbfD+a2cEuDEl+FKdx5muFApAZDJoWWsGB
v124Owqs3cz6Y+5bpaWzwRhkfS6vZs/2Mk6fXtxyH7qfM0A3vJyHb7+S4EABqIeozwEEMA0I9/d5
3o9t4iC+7vHbWDl69li6BsBwKOrIHorog/PnAYXlpbWHNJpAZM/tsEgioiqBcVwSXrWQZE1ac0sD
ih/uWnQPbQ2iQcrAXCmwk7Edozbl/7Y8nDLlVFfmEgqInSED4K7WtTnWL5ZXICIH6xyIM2pGoJv3
MCLPDYh7FOgcXlXRA9BZiDDBSpJ9Ep9pDLKJMTxKDfwNfM9F6+cmjxu9rbMCjnTqX+m21AhT9bPN
69zEaGdBQq27jXSHcxML98wVCMXpQZvlLls4dPwWZg330zS8WDJIolrCL5jP+3xwGoO/c0au0e39
yL/NNGiep6DEMCQgjzG6eTa8nL8l6FbkI4GkwMzOgCYW3Mvnz0P/EI0KfJRu6yABr1DLyYB1ITxx
1pTH4Q3X8QoGKiWx3uC4GL67GZsHCL+0fOavppSezuvCynvbgMfbNMpTRhYM7ZocCUohHlrSOFzB
pmoVxKF6vEL1RTJgDU+ZC6/8seRgZP7VT9ANcGfUrnErgWUkU6V2z9GEOBgCw0ifqtQkx+kNEePx
gS0wy1u0OhoF3E9Aru0kvvcL/ELoYIyLLEMK7dHuXfVhy1mmOcsp+Znpk9EpP6SAhivG9ptX5H9Z
jhRcufAVXP8fOWzI+kYhxqoDVaxsELuOu2t4xFL6RsdoG4Dxkk0pL7cc6v76eA2aF3uoloeBPw0L
abGVKI8kxQDvNNrUCNg4e9QNw17HR36i650DhhvOeEdmEItE29YVlNRipJvnsjVB+FBJgmENK/31
mUAQuZpXLxrv3WQQs5+tm7pqOgXtaokLfhxovF5fbgFtuZZQtN44MVarWJr9ZLBCTRdMXryIbtCu
gZQJwVmBHQpDkeOkIMeuYo7sYsrpDSvc/vReScUM+fjTVk6oPbtONkaByWUioesxM+zhBHiXgrl3
eaXtuW3alJe00TP4KR/IUML9WaDpuimImvlp5Jamz07Aj6S6U6Du81okfBdVfYzTPNauTccdH5Sk
yfycGcLelRQlyB0ZUioVzuWHHrt4ZMxX5sIFrNNxx9ZN+rYcKdltn6cPt0V4p3NJtchzT29MYgUj
7Q4mbPE0HtUZJb950S8S/NIGLssQMY9i2+HDjSm9heesaB0CDQm4mfAapCL2jc7/P1m7sO6zF/MR
5QwRrN/yKC8r8Vr1Dnx+FXCpextl+MI1RaFyBV6irLXTDpeddX7iMJ2c4pAstGr/vsypQiU8QfT0
cpe3GzbRwTsjf7Bxd/5s2u2tL7Xz25mF11lhO1jALk269+I+e5nqyK9opx5W9psewsGqr4Rr2BZ0
ovIM/7mm3F4sHyd7gFRqe1deVCiSnFIAmyNBOWoFVd79wIKnNOoFALMAi/P1xgzFN4quleI3neI7
vJ+mhTwtao8EixWkot9NDg3Lobc23+MAIosm6E4DFKaFu1QWqVB9n5QfmAmZp35TxDyXGeAQCK26
VyJ6SmKuON1PGpiDfjAynqpQJjNi7MNmPxp7rwgJe5cYul3sYemNPx+HBYPRBsr1qhT0Wlk2oAGh
je1XjLK0j+yi8I0uLSWQ4E5vUbtD0pAc4IoHuPrydvOJ0mtCxTEX4jnl/AtY/m5kpi2izRV/nxvD
kdfNRh673cxX8jB338SbyA80dq/mAJ0NH43cx0BFQvCfLFu69Hqw2Z+tu7OU5nJRS8Hhl5iZ75WN
neNo5KHGhsNdaPCzkLG/RHkE7bbZRez7MDKCVwKAoKMHkFv3CIzcnyBDxdC1lAOQLIVNb3V6EeCm
LZJu7Ks5HtT6Wa9C8Y+pTcuf62TbrdNdMGlQDI1EgwTJnfr3hNPZ2KZx9D7Q2DcMFxHEAlIRFkRE
Ftufo8OzVXm46KzNDxVyME4MUBAamAAFASR6CLcmc/uRusStG9L0mjLFA+GXqmUAE2/zDot/kVol
XwRS9HVXJZV4FdWlwfWezgBKvA/HuqGFduiXM6k295X4+2y8fH7Uf2BodMkbB2YwkXzhIe1KnidM
N44Ov9/jTsObj/FPFnNwtlWK6lb4YN0moLLDyovT+sVfR9np2KMktxmWxORGFw1cBF4Bwu2mZjAm
kYwceWDVDNWfsDp/iOa7Ogw+Yjsq1fbHD5RVnOekBSr2mzgVFt60fDHsVG8NmewICu9N2/Btd+id
mjktLA/D/AkJwD5Xp2Ej9ulXAyd8ccK8uv7RAYjMBesc1WmlneiyH50l/GkU64a9sTz7TWrlED1i
lIOIOukUeH24o8m7L8SaAM9QzKkQ9vvaOdmpWUnvq3wj1b55QTya3KEXzqgB2DZuxQQfxpxGRfrz
ZYTZHLX3ZAIYfczmXeapq6ACwns0VKCR6wROigqB8b4ek38/2CBrDSWQSk3fszkPlYBqALMVKJIw
dUGcHgx7R/4uqQ79QJglKlz2m15CSTJDGrBu2PZqVegDa9JPEEam9U8BZVICsOvVlFhF4y3X8C3l
ebjog5TLXcgXKBK/Gwg43Qf9Yw/eifTkNpbMurqzErf3lJtz4BnaIsKIuNgrYzk8PlIKI8l0XTfE
q5a02dEE4n+4XwIN+JBDcTXujJffj/SfO7DwWWSpQs5XRPb77rjKuOA+8vPLdDNR1cqwOyWgEvyB
sM+MOp0xN81OV6XgWeS9DnzzaWjK6xGn/n+7q/uhabWh+QTbP/DOb/Yz4XjKvN7lvHb/wX6YrVgA
+RgkNeQc2hqCjBFLSBLz8/8i5klB0nwlEqPvBVxv3rSvn09ArOXntnsIDr2/z5toVFT2I/KppyN7
7n35XU9l0UsBKZXKLsa1+rjzD1SA/1YiOVjGTuwrEOgvuAN1G6fwDfEAaTGVeHHH/J4YSjM3g/kl
R0asGdEWeEBhBtbt8KUaUr/BzgPzA8T5RRjJZDgylaKHoJ36+0mHke7aaHsqHG+bl9+UjFaZavf7
G7V9n+cehrjO3Ei3Q14DwcHWOIIVHDsGq4v1usiwGAkk/JfB/DVOhvElZsk/p0wk0FDhlSrohYG5
Gn5MVyjYY6XnWRqVTU49OzLolr7tFOqjobmndWu8oYub4bxXttUJdBkgKMGw+nRRs83G7GQvTwL2
044DAMOBAoXJ4VmiByddhyJ8H9YALAv4vpisBNdToQeu7Y3hlL7o8IC2gIWbadlpE0b7Ql+45Pt7
DtxiOFYgDzFZVYEt+CmAKSb8GbHfhfgnirsBJbwEDZxID3eyjY1oOGCZQvXbKBdk24PCmmeMl3cI
SUSO/NSNfa20JFq6Bv3+aIvKx36lcypp3DHhZoP1BthfeKzeepKA7GUPWuwZV4XPPGsHfjQSRs9X
FbfK/Yg+4+5Tcvb4/z+s+9oTsYNjdBFOBAHmocdGU/M2MdINm+6j5ynUJiaKbanpU5Kl9msElIV4
JGzA+8UVWbYGmmeuaT/W+F52fGG4c92J+Irq3ArNTAaHGNT7NbbC9eW/gUxpfqhn2ggSZqrBWKek
p+32FqjtPXHcoe4YSDpu7QuQXMNGY3uEoOfpONBzPBh8OQBlqF5yOA2gWq/D+30QvASHYCh65dUu
5auto2DaYiJH7TI+5SY6SHemTEY8qftbTxpnOcBUMmmXoo4k6jzL3erXmHi2eNNmwi8R6vDpAb+H
3/bAvL0Uid2Z5b1hLSFAvI13MIFo/sbJrRo=
`pragma protect end_protected


endmodule
