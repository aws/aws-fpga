// =============================================================================
// Copyright 2016 Amazon.com, Inc. or its affiliates.
// All Rights Reserved Worldwide.
// Amazon Confidential information
// Restricted NDA Material
// =============================================================================

//--------------------------------------------------------------------------------
// Stats interface registers
//Register MAP
// 0x00 - GPIO 0 - read/write scratchpad
// 0x04 - GPIO 1 - read/write scratchpad
// 0x08 - DDR is ready status (bit 0)
// 0x0c - DDR reset (bit 0).  Set to drive reset to the DDR core.
// 0x10 - AXI Address - AXI Address for accessing DDR core (refer to Xilinx DDR specification - pg150)
// 0x14 - AXI Data - AXI Data access for accessing DDR core.  Read or write this register
//                   to read or write the Xilinx DDR controller registers.
// 0x20 - Write Words Low - Stats, number of words written (512-bit words).  Write to clear.  note is 64-bit counter
// 0x24 - Write Words High - Note can write either register to clear entire 64-bits
// 0x28 - Read Words Low - Stats, number of read words writen (512-bit words).  Write to clear
// 0x2c - Read Words High
// 0x30 - Self Refresh Request - Request self refresh to the core
// 0x34 - Self Refresh Ack (read only) - Self refresh ack from the core
// 0x38 - Restore/Skip - Drive these signals to the core
//          0 - Restore
//          1 - Skip Mem Init
//          2 - Restore Complete
// 0x3c - DBG Out - Save/restore debug out (??not sure what is on this)
// 0x4c - XSDB Select - Drive select to the core for save/restore operation
// 0x50 - XSDB Addr - Drive  address to core for save/restore operation
// 0x54 - XSDB Data  - Drive data to core for save/restore operation.  Read/write to this register triggers
//                   a save/restore access to the core (with XSDB Addr setup at offset 0x50).
//
// Interrupt Status0 - bit0: AXI-Lite interrupt from DDR core (refer to Xilinx DDR specification - pg150)


//--------------------------------------------------------------------------------

module sh_ddr #( parameter DDR_A_PRESENT = 1,
                 parameter DDR_B_PRESENT = 1,
                 parameter DDR_D_PRESENT = 1,
                 parameter DDR_A_IO = 1,           //When not Present to include IO buffers
                 parameter DDR_D_IO = 1)           //When not Present to include IO buffers
   (

   //---------------------------
   // Main clock/reset
   //---------------------------
   input clk,
   input rst_n,

   input stat_clk,                           //Stats interface clock
   input stat_rst_n,

   //--------------------------
   // DDR Physical Interface
   //--------------------------

// ------------------- DDR4 x72 RDIMM 2100 Interface A ----------------------------------
    input                CLK_300M_DIMM0_DP,
    input                CLK_300M_DIMM0_DN,
    output logic         M_A_ACT_N,
    output logic[16:0]   M_A_MA,
    output logic[1:0]    M_A_BA,
    output logic[1:0]    M_A_BG,
    output logic[0:0]    M_A_CKE,
    output logic[0:0]    M_A_ODT,
    output logic[0:0]    M_A_CS_N,
    output logic[0:0]    M_A_CLK_DN,
    output logic[0:0]    M_A_CLK_DP,
    output logic         RST_DIMM_A_N,
    output logic         M_A_PAR,
    inout  [63:0]        M_A_DQ,
    inout  [7:0]         M_A_ECC,
    inout  [17:0]        M_A_DQS_DP,
    inout  [17:0]        M_A_DQS_DN,
    output logic cl_RST_DIMM_A_N,

// ------------------- DDR4 x72 RDIMM 2100 Interface B ----------------------------------
    input                CLK_300M_DIMM1_DP,
    input                CLK_300M_DIMM1_DN,
    output logic         M_B_ACT_N,
    output logic[16:0]   M_B_MA,
    output logic[1:0]    M_B_BA,
    output logic[1:0]    M_B_BG,
    output logic[0:0]    M_B_CKE,
    output logic[0:0]    M_B_ODT,
    output logic[0:0]    M_B_CS_N,
    output logic[0:0]    M_B_CLK_DN,
    output logic[0:0]    M_B_CLK_DP,
    output logic         RST_DIMM_B_N,
    output logic         M_B_PAR,
    inout  [63:0]        M_B_DQ,
    inout  [7:0]         M_B_ECC,
    inout  [17:0]        M_B_DQS_DP,
    inout  [17:0]        M_B_DQS_DN,
    output logic cl_RST_DIMM_B_N,

// ------------------- DDR4 x72 RDIMM 2100 Interface D ----------------------------------
    input                CLK_300M_DIMM3_DP,
    input                CLK_300M_DIMM3_DN,
    output logic         M_D_ACT_N,
    output logic[16:0]   M_D_MA,
    output logic[1:0]    M_D_BA,
    output logic[1:0]    M_D_BG,
    output logic[0:0]    M_D_CKE,
    output logic[0:0]    M_D_ODT,
    output logic[0:0]    M_D_CS_N,
    output logic[0:0]    M_D_CLK_DN,
    output logic[0:0]    M_D_CLK_DP,
    output logic         RST_DIMM_D_N,
    output logic         M_D_PAR,
    inout  [63:0]        M_D_DQ,
    inout  [7:0]         M_D_ECC,
    inout  [17:0]        M_D_DQS_DP,
    inout  [17:0]        M_D_DQS_DN,
    output logic cl_RST_DIMM_D_N,


   //------------------------------------------------------
   // DDR-4 Interface from CL (AXI-4)
   //------------------------------------------------------
   input[15:0] cl_sh_ddr_awid[2:0],
   input[63:0] cl_sh_ddr_awaddr[2:0],
   input[7:0] cl_sh_ddr_awlen[2:0],
   //input[10:0] cl_sh_ddr_awuser[2:0],
   input cl_sh_ddr_awvalid[2:0],
   output logic[2:0] sh_cl_ddr_awready,

   input[15:0] cl_sh_ddr_wid[2:0],
   input[511:0] cl_sh_ddr_wdata[2:0],
   input[63:0] cl_sh_ddr_wstrb[2:0],
   input[2:0] cl_sh_ddr_wlast,
   input[2:0] cl_sh_ddr_wvalid,
   output logic[2:0] sh_cl_ddr_wready,

   output logic[15:0] sh_cl_ddr_bid[2:0],
   output logic[1:0] sh_cl_ddr_bresp[2:0],
   output logic[2:0] sh_cl_ddr_bvalid,
   input[2:0] cl_sh_ddr_bready,

   input[15:0] cl_sh_ddr_arid[2:0],
   input[63:0] cl_sh_ddr_araddr[2:0],
   input[7:0] cl_sh_ddr_arlen[2:0],
   //input[10:0] cl_sh_ddr_aruser[2:0],
   input[2:0] cl_sh_ddr_arvalid,
   output logic[2:0] sh_cl_ddr_arready,

   output logic[15:0] sh_cl_ddr_rid[2:0],
   output logic[511:0] sh_cl_ddr_rdata[2:0],
   output logic[1:0] sh_cl_ddr_rresp[2:0],
   output logic[2:0] sh_cl_ddr_rlast,
   output logic[2:0] sh_cl_ddr_rvalid,
   input[2:0] cl_sh_ddr_rready,

   output logic[2:0] sh_cl_ddr_is_ready,

   input[7:0] sh_ddr_stat_addr0,
   input sh_ddr_stat_wr0,
   input sh_ddr_stat_rd0,
   input[31:0] sh_ddr_stat_wdata0,

   output logic ddr_sh_stat_ack0,
   output logic[31:0] ddr_sh_stat_rdata0,
   output logic[7:0] ddr_sh_stat_int0,

   input[7:0] sh_ddr_stat_addr1,
   input sh_ddr_stat_wr1,
   input sh_ddr_stat_rd1,
   input[31:0] sh_ddr_stat_wdata1,

   output logic ddr_sh_stat_ack1,
   output logic[31:0] ddr_sh_stat_rdata1,
   output logic[7:0] ddr_sh_stat_int1,

   input[7:0] sh_ddr_stat_addr2,
   input sh_ddr_stat_wr2,
   input sh_ddr_stat_rd2,
   input[31:0] sh_ddr_stat_wdata2,

   output logic ddr_sh_stat_ack2,
   output logic[31:0] ddr_sh_stat_rdata2,
   output logic[7:0] ddr_sh_stat_int2



   );


`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
c8JKX9BNuDkb0ZrKkm6zlqZbqBHWdLr5ISC8ZlprccNdL9pHd0Yh7ebdlRbHk6LTCwoB3O4/fVm+
EYNT9LSDt9vjOmGOfmj0TWBV5dmzyMs+JlvIoOcYY94j4YFE+p+2+JslI77c/7768ib8m9/EiZ69
LQwB1CCaj/3gUG1Sg74s7mhuyUSGQtdKbj3vZRAULdOwXr1sKP2wT/pnUK44unEOzvvPTPt6vR0w
9Xd+K1vu8Cn+9NEQpjxJUeZsNTMdMUGi+c7QdrQmHHE5aIjoOLfCDoWxSNkYJG8ZX3UhF5nFUs+z
NV2pmhZdMfEwbTHVtxRpZK4EnPzqehqpZXz0mA==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
t14SX8Isth9t1rc1FIhl+ir9dhyRef1D370Rpg7VPZA4/p34OvTByV+KBTmm7LZ82MdsNM7AdDCf
ORA4inSnuT1Vjtrp4xs6u+xV64KF2k1Cs4Abcd5lCQnrkwL2Dquh79rSX7svqbynF7qB8R5mWhso
dwOO58vdAiN5C2x8dGQ=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
XLlQJTxpQdotSPNgUhjGkPekYsR9yu0x8V1BzK1XW5KY6wl2jX734DedoeRWWv2oBoeVW1EA0bzE
2v2GtJzYgdONIosoZwnWGJTvib/aj3XXayM8UnQ3EJZ2Xd2LEwCzkzwAsOcKfpQFrFyuiuCscdg2
tJRldsG+mk4Z5ENfI9o=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 48064)
`pragma protect data_block
pSjZ/QzpFJD5U8URGzSZ+oxuLM9JxBh6HdhVbTKUm/gklJ7AaecylDeASvgwCogDoai5NetNPTz1
rPvkYtad4todvVv8dyl7nvTew1vMg+YKErmYMoOGbSPTzrSP/mmT+VsBAKwkbhDOwA76YT1HRPQu
cjFd4iQT4XrH0hBiv9G3wat1TL3G2M+l8Q0cMJvS5LNyLTbQi+1m+HjnVwoYpf5T4+iD/hVVFjTY
A/TdjXDDTHczmStiweFZQNnRiin2Y6kL6pyVkN2vj431i1Xgtg0dpLbG+axBlocVDqUWS+1rwHcZ
i4aUEtx7IjeZLpSXg/CNbDJbF9Yzl532SPQzpY1801/wjPfeFO5/fQzlcxtgtremqAerV6u1uWJO
NjtL/mDXaRU0tBspG5UF0DWHqHzWK8alUgvvy4SxtWTBeSb0IgFheFJhaZXx+IadnGtS4WywjE+v
TY//K94or2PkHK/jwBHpxJzKKBO3qymskh2gHSEGGwOy8eya08DcJpfqK9TnCziNU32ClDmvSMCK
Zdzu8ypUtNO6+ZSqFKfkzUx3PQL3FjVkh5OGxWIRA5MAX6gfNqFjt6fXTwlbk7qeqEx1aUoSoaVQ
krsZ0MYynLmOzc+b0YdhYm1NHNfsloTiRKFfDL37LsGtdS1LjmnKZ8Gv8Gf6EKXHVZVC4zrNkOU/
ynNA0LXUEk3pC5vf5KtIRpFWbYQpzrYzS0f11hMzS6DKYWFo0zvPJT/igp8LidKtRO4E6RBSHQmY
FB7rwUewAZh/u7+k/+IbcNTiOFVR8HQ0/VF4mFSWBPhtKaEVG5xTPZs5+i7ynnBvaNiPVd8ERi7p
jn7jz7Sqc9Se6G+jJY+rkI6oFBWPaNimxDcHzWG9Y8ujXfJgx0K3Jp2BNohz19+p3rR+Umg24G9m
b1je294k5XehSiTvNRI91I9R4aEdYCaFSJHDlFLPkPV8EL2AMGvD2aNKt6ZqXJSJWmBaPCD+4YH1
0msg6onij8N0Lf6YpxdMSXVpPFqb92LmLYo1orYFfBgdNvoAucj+FlBAZ5L6AKxnudoFZLTQyI5F
Dwhrp4Ms/Wvag+IV4L59/hjoDnxZlnfl2nMii73/+zSyPI/rUFUeemGj0UKiNSPk9zgv2WUhlEKp
QIcZFaR8UE9VbRmeUVp6eLWMJinn7gR+HESteZufIMndocBtUy4VzNx8ZemXw+MssCP6ZjOrQGb1
6rYP3kfF6pFmQyc8OvkdaCJiOi+o/TbBxiJDkHWLRiXBS/+dGf/lo+g2ksvULDxDN1VNkquse0tQ
wmx32YE28rCQ1lqVMeu1L4BgFhIoEbeutxj44kGxfvXv7jUVOU78IQRYnil05LklJkm2I0+Q3dGt
GNJuC/S632U7K77wvNo+9kKbNa679lmacrivOcUP4g3wGxy7e5RbwKXST0b7xV67VU68JOQsKS07
wisFYS0BQk8YQPRgZOZWyUGsKIrBf2NuQJt5Zx/j46bKYn/vwcBwDAD9dkzdu/RoUQEzA016G4B/
Pg5exOIqxc/ycLY0Pz7u+J6rR6+F62JODDoQUwfivD7dpwXAh1NurysEqYNGCKRB4V9mZBBgrC5p
iy0iN9pPvoIRAR5JQVXWQsHOfLV15vFGozXhC00C0+1kBFpfZ8yqH9HovQFtP8lCmvk7cZ+8hYen
qI+EErt+P9nrmWfJurXj+uJgYAhIqa75w1Sk27FtcNruaonEno4+vYoMMmaUzlrDVodpHd3/OHl1
vZFpix8mioqty9UU0iGot4nvzp4HyHFexcowrMs28STGMRLqYEHmHZabvqA2kNUnJkGWSSWqFSNF
4JTSqYUvDSO8GQi2vDCm19U48yt2MPz28OXFj3fC82/Kh+YVFEtzR9kGndVs7DxPdDgmNumjZM7C
3PQCOwd9QHNMt1jdR0ttTszWC/tuvE7SwUFMH8QMNGeIH9JVauMT7t4GEmQ3AfzB0ZulSC4l1nBc
FjEcEr/rpFCBf7FdhQPa+4ui0CZTwxBmU453/vcecJmv4wrah/boOm0+bxI+ZJymaBDT0b/RLZaJ
3xVMDjqo2Vl/Vuk+p99WRTVRXBgPnGLQgK/hd2Z8ha7LDCKj+q9t7b48FHioR1VA36FZTln8kKdf
eBR50dd1YBuqp91fX7YtydgdeoTc7uFZZKp8lVq9yZxQsaYzLXIAeyJ73PauwiI7qUTSFwSzEUYT
WYDk+TrdD9nQl9j417wbxinhf+EhujweBarkN5SUYCYuNEpRQ1B7FQatVsnVHzv6HiUu58DCdbnC
B/eVlQJWY5fw2ct1AaOvsjsxHn7OuUu/mUIXb8ppsRK80bdPwgYgt20BE560f16qjI6Uiy+5M/Ml
yi0W/DLgyTqEXTyPk73J8EKfqBnpPMRzt/URaN2MxzWoRmIjoC8w7uMmlVDYqgdCQUI2PaMZ5ay/
KDZVufua9bEmZvgffB+wLxvpeMd7B0x+hRd9JXdYo0Ak2HdqGeEma58kwhPMVgb0nWIVY/yKe7bA
pLbclJ16AKQEW63Ulo0jFPea+KPXH8d0gWEkWCaIXAbqthOYnBdF5evlJByQ0xnc0t9+zm/6BNoi
jjW7BAe6tGWjQOJLRQ4SFhiHxagfY0aQSNVxVxXyxUoPhnn9MeSifAaQvqcHLzQwEkZP/rin1dX/
iDvNn7GzdVlfqr7wKFT74mqCDPWz+x2AF4IW8PT5bLQ/kBV4bsf5d8dp5guOVPh3u2xv6uBDmQph
+HediAgVpCCC5IpYnWBg5f9XmKZdFCIq61KLsZWbkhi08MyHCmaBg2sWS/Ptk5V4UtyjXDj9Eitt
eOXUaj3UifcTIT5pXMrK3kZ7etW6JORnn/2tjK0B281E5vUKj92dyqfKpxX3dYux3OZffrca8Zla
sYXOjHxoi3bne884XlYx8CiDH1SpKgf34v70dwv+c4QOfRTpDxwAonvIJbqSc6I9DkfQ8njk+OI6
jYpfDe/XtAu9GBM6NEnNgR+b6b7c4wtGoqBmvr98jP8pe+rPBdTorbbvEGeuaWRMkiP7CjWya4uz
PT+3wjeb8Xixd27QUhxvG8x8bRmIp52Oa3MeTnrvUfukpj+9ArgRthj3gsO9WGfn5xnIi8N2Vfov
EbLAraWju7bkJq9vlO0nEpi+eZVBF2WRu3YPk2sQcA7cfxuGb1Bacu2QjO0ue666OOvHFd/pnZTr
0b+mXmIlhJ31BEvhX6pwr+yn1NluRvcE4pR7cipyaFD81gdQcoVaOg5NMKTb67R3D1bnb4aN++Vu
kHePtNImL6Irf+o1Ix2THgiH91DQbX4G4JkYbf/ZgLkWfhb4JR4dAcGz6vLN+FuXZbc/QJ+sKDAV
SEmn4NdhtVbCXp+pGK1RPYOyxM6fwsYmQmqPJMRL9/kQl54geGA56nt938fivcsC47skx3/lZEf+
yNtTkCXcGv5TvzPyF1NF7UdC/x7tKv37+uupQKXKSUcjoe5mJ3I88wJMk/WeFBIRFOvlXe1oIyt5
NF9v3wcGLIfWLAknAjeqK19hKnyFdmrrl78KpB2YVGvb7vJJSE58zXdYaZ+U7IbIvsVURcrQ5NRx
8SWXycBqM6iFFf1pW2xLaF5LYphht+WsSHD3Cgmvs0lBVwRcyhi9MDRQPeRsy3cd7YnMkaC9T7A3
jI4n6O9JGdJ8SwUJmSCNa9n750mGWBi8Mwyp6sBJrKJosMIsizMuT3eBZJ7ye/1cVVPVyNFxTDFH
rmR7HY3JDx8DAZ/lKxZFeDp7Rk5y4zPhIVfcyzuXXvQc2sIFSiJoeRieVy+8rAyv/owErFETmMAZ
w3FEiUwIVSsSZM07ofkQ/BVsBQAKxOF9ugOE1yuKWkLTczwG73n3w3I6Yi2zZ5HunFvpHeVelYJi
SejkK/Ku3JXmKXKGuvOPWrksbkHb+wXjYcZ/Mo1xgahNLKOA8hfxmKTVfI9shHTZcJGHRtlYu0G5
VfRhk4DwPoRJBRYn7SCgCCM2cLDqGTbVi7fkaoTBxxAm6ax0L82/TM1fI2AqfCidGAKtcajyuWjb
YhY6+X9jAYKVGjo4VSnhjAPjLEyPEoKCE6E5c3RA16PUqGL+DpgXll9a1FBzMtTC9XGe84IKb5wF
/zpm7is/cj5ZUGIhmGHRB9GMWnCOEAbWOPvikuIia5eWDYeEsTKrPUd7rJ9SUpFTMlYo80LUoTqC
r84lMxcaERE8CSyiy72aTXgbmGrIsGHQdIxb3bbFu6CnJIcLxILUU46U/SboRbfnNoVZ2t1gR35F
Ee/BGyaiD5XtLF0dwT5uc/CxrahtOFwnI4s2VWTW/VOCPAjtFO7NxV2mbFfoJlzzCOcqyP/DTbeg
8i8KK/XnriEVkfp9ZpsA/9oc5tUS3cCDxZ6Z0GxGXJs+T3H1y7MwsUMV3PbtetE0Xil0Y1cZ014a
WZcniVCUzYATR/IMjYyc0/FqxPoymvgVyswGQYfPlLqxpDr4H7BNNa7sLsTbgqC9Zi7mzHstHpUF
FCS/lQmtNjQspVDFH/v4zvqzRraIZEsgJvFbzkv7KgW5jI/ZuGR+tzO0z7jyW5KQTQX9fcbPiE8M
udaf1bZB0oOkQbnz7MFE/golMtN5hYb4EpS5/HOKlMFpxhWfP4COXCb07ZzPFc1OJYIWmr59JQP6
oteZwYX701Mk0ivEOE6ATj96bwC7b9SlwiMS6p8NiOXQqYxEPAg4yFlgazwOSpYtjA1DSqdewl9J
5xRxRpKQqq2aLwi5Aoi1u9xHE9ALZ8aLICp1odUE/hS72wvZjMThxhaTWIupJ4SguhLIJO1bNyR3
6TKzBwv0UOorHLGvjcmI70sWGr2t4bupQsinlpWBbLZYTTcSIGOkSktzt56DKeL89CrAucV8j4ch
VmVLIBGne4jkfoAKxjV1qoP7r0Fho6vSHIdMlHICdrCpUmTTy7m6zxQUfuJS7qIrEvH4zoK9uZY9
Bxv8uDPhk/y29zIqZoqbQdW1yZA8VVrse404PnueLNYuV3Qc1nVlc/nX/AuuNeBIWgVHFDgz7O5q
i+KS7Ec8XYBemn89q87WM1TfuEB4jxc4qDkThOX2FURckIcYWQsiWkL6xVjkVvcSStejiGOEi3Kv
xswy4CCaOWXbDJRos1OE+/jWe5s9Jy2V+BC59Cja7qaBdP4kA6jmXSQxbGPSHy5e9bId1AlhvykE
BwrnGV4aOYitbKr+s/vpIDEqtwKtsHjBN91gwqHklbcFeNRvR+PVasyfgr+RT8AXeY3f9wUKTwHw
TYhI0biu4D9A2YEMeRvtyfE1uj0RTGO0D5uICBplLnboeNZZXK8km8nI4KdZyzXbVCEinIdzv6VQ
fNf5ee9AszTgXIzMWuGNOH4SmhB5WnkY2XvEKekS6GQ8Iv0R6gFVZUEdOJA5eMOLFCCKRKcDhTEW
q4Htza5Z8vN0EqbPIuOb3IBAk//N4xuUGLpIhoWRFLgfgAQkBrTnokKaYoZIFfpdKmye7n6XPtcV
okd17H7BSfl28mRXI/9WLRaTF68anLv+MaZ2qvF5Gu53TbRBRGqVV7ht9Am3/PrPyI7gJaohyfC/
yu6jyX7/bvq5MIiyv2lYan05Btia7AlyZ82461K/6JnVzQinPkEjoUqzSDSKiKKr8lhjLXa4hk6s
ndIqsAJ3lGXaQ9hOntlrBGRUYF3lz3H2yDmh4fbw69WpMpzBRz5CmSMZ6VZ7fx5FYzkJ7y8dGUMJ
vFXwA8xR+H6kH51sGDlr0sj5k9b2934rLDbKxExFca7/0KIFfsuRLh1vlYxofPKa69qNx4W5M7QN
lH6pSjprnFkpMScv7UiRi3xVndO+OVC0aPel+SR5tiNJeaeySLcRhe2x9x4ecg80iMR6blwIyPRT
Ah8mLcS3gdhdG887dKVn2mw7eQ7JnACjIyEQ3ZnvPTTTgbEstebejHVA1AheUSd1/0GvH8hFhjaV
J5zJ0z9Rv56Bg/Z4gFc4+oVXQ8wpsaeUGNytUYS2azjrfAsW3yh0cLACzvaITB1xdEsXjZtBytGI
kudxi4vvdi71MVq+wG9W9NML+/JUKQUcxqkphlyAyHEeVObv1ZI1prnyVXc9yugeidXnYIM7j0nb
0B75009X+hD+x/BZdGwo6uzFsUa2eklRRnjkS/vmbveKb1rou8lPwvzxhMhDxp5VmYWiw+6Qha0i
UBVBJuayRX9vI3XtU3EIFxnhrRcwdZlH2yaDRxj59znnZmFz4QRF5s+Up4OtgH3Af/He0JeZYDIW
jvnCDJF59czelntcdrdt43fMWnWyim+gq7p+BFHNaijLoX5Ttj6XxMPsBeuojF/4owHKMf0a3ao9
Slv73vIn/J1GdaO9nWGW3zh4JCjIPhh4r9J5yX7rwnnjyoAoN/U84BdM1xw2gFDXwzgGdBvo2XAl
cuPXz93O/N7kDMYe9o8sjQYC8D80Bhrq1Orxz3V+bSCpHaBCNH0JAvOihQdNX7O1Pg6ArIFbmPiz
0Gxuq2xlPNMWLWflzcLAOhPqnSWxnsw/zxsZXNGSGSdidFR0y1ICNV+vqv9xTXUbIK3evAmoMzZd
YtBGygbk7n64RDCyQB0ytrpQQhAKjtXByWNRkuQGqBne+Zw7Ql9WendKpNSOJQVWLREl4T1btmrY
mhOeerJpIXA/APzK2tAZswiLMnCuc4IbtXMNT4tprjl8Id3na2FYgiLoMX5/HDa3p97UUWX1L/AN
NLb5qfz45w7MKh6GnXXHPlJngLcTsB/8QBbtEz6+Cs4Z4IvKfBcOdjtuIbzvo0AZdq7B93bm0226
ek04bpUP4cR4t/eozFW8LaF0vL68zJ+6skoyK6xBgZF0qSzd6wmzW+KpmBqmS4PqfEW7z9/X8Qx3
7LEAT30dy/HPeLdC04zrNd3QE2AbcuY/Xx7oU4BE0MwcngBG+XXy8cqjNa6Grl302h7zK9aazVTH
7G6IPbMvmFcZBxcLMSSjAJfz73V1GJBc4MWzJ//olMHAFYbTvTBNmVgK7gvwC1WELCvtHav4p/ZR
Vyu837HMFBsiVoEHUgEWP+ywKp1+F49XKpySQDTOvbD4Q9ELvUxV8hH5tCxGopUwMrY19pSCCe/e
5de1XtPet2jggW3Tib6xOq2KeMTZrrvMDgtZ51vGu7fLLlvNJ6vX1PhKNydzU8tYulPFAD7yl9mH
JpfRLyrpL4E8vge8NfVRwJ90/cJ+wceIm+0h80pFl0WxMds0nQ3aggzNmhKXcs4bjGQuWuWwjY11
U3/llA4rHGI02hn2V1Po/vLRxcmHmwLcdy9PuDM1CtgOvvPLcANgno2kXDMb/kWzC142wKyMKDn6
uPg3yx5qs0IrAlDtOy/dVDPBN+4F9kblDywuCBtkxvQa4xFKMl9tKmxzuzuSh7HuIFMlBYswZBb6
4XZV/IibX3IKEMkqNtkR6Wn2IPFZNLXpbbVKwrjwznrm4B95WOuhA6/zBKzz3UzGvND8jl4JZteg
74tIhGtQlTuBn3xwO+j4H5TECcgMCGa1i6h52RS2QophhHMG46LqWTaHGYkVXZAEBrpra6+MfCSA
iALpzdzOXh55tNHOY/8BkZxLSInl4OTVib2WkAOGcyFhDARUfXgwG0vFjGXFOL/2EADaAX7O/JEW
XyjMg7mn4iao8z0bSNSOrHIX0NoPqUGAwr34TY0s5QBbIBdecSAdcFNCfJIDW8kpqLUJqICqjFml
t8SlRFtouRszAHLF/0UR3UEqJh8iGJQHc5hy/o/tU7FRXBx212kWLNtfJ5wNu2OE4pLa9tKi2jsg
BsZG69FVRcbeORhQzsgdpqFCdgeO0rANTiqlyeGXMeW4BOV359mBXgbr3oQxQt5y8Ckl9V7y1kuj
vmV2BgVaNYjdLtCAxweIrgkxtWJdmyeyiwBT8aOCy8EQBd+IaAixWLKV3Uo5bkFHH3owyh0dyuJA
qtRHLE4Dw66OlrB/fv0SC4jAdaQA054tTqlTeVwcvWg3LlBB9lOePCLn7kK8D0uQ2HDQOF4DE0D/
MJSfj9tuPiN8GjGNsB0WsZ3lSNI7Ja7AH7ZSqxhnBs4Qeezc2Z6pB/0ANgplfEg/fCn9Dd/rcFfr
1ajjgFhXbQoSf/iHHWIX+arojjAPorZPloSEI7eyxzMG15R/WMZuIMUzN+yjFF1NA+Irh1JTKppy
Ikf91NTPg0/N49PJkt5fFptbOYI+LCeNYLw0DmB+u68wfhaOsqDE+EgTefStF8t+xE2OwvPGSjjO
8/t9GkrHnGSAefmhtAgUB0QosQCrRebnjhmLcBJ1IOUlitquU/T+ZFDJSEUcVpMX4QB8r5Py14VA
UIB1l4pibEHGOPs+NQwALQUBDbFxcLrNt1rPoaKKE5q9G+vbLxXoQ4qQZX8Or16PJcfufVXxIffr
VnYrD3U31/ogr+QoS+pCTqMVZxngUH3AY3fOr8yoMx6eS/5KEZwbRch3QBPWBQAU8fo8CDoCDHkk
OO28D4Kbv2xAXO/h7oXzdABlQoa/ijR41vdcB5ReFhL2e1hfRBUvjoapcf/Ddx7+ja3xHbtr4u2d
ntvYxdOaaFobvnAXtf9EjugMWgKvGOOnmr1YQhZTaPmSUBz4WHJHfJGpnjVZMlFLalLtLEjI1cvg
ua47dqGPcPQ/fjaW7FXH2jpGF3HWMN0FzdkmJMD1kH01C67GyX4nFDRP75miXApAVlYKQVahPJEI
5zjX1Y86FzZ1spBFI4NIj/ut48CxDuZ8rF7we8DU/DB0RabBD31Vpgo7IZX0tokpSaOFHVdaRPLj
mKn74uCnBxaK36uSm4tmjn+MD1KW6PjEz9Zz3z4ZgkrXFkCMVwmHRvFkWyBWX+xloM189mds8G7l
fuKvX+UFBiImdg8weCFLYuXPC7zP1nTB9Tr+KeL+Xh3Puq3XuHKO+s2w84LmQJziZv9CZ7JSndBB
yKOsKoarU6r4g9zWIU0i+QdI6iiz9DVwQx9H2EEKR0tn1ILZJJaTeBrik3j5LMuqBs2Th7Jijweq
hYyYxKhjf4M2kUhGSqJx1r9BQwGfdh23ysYjBtjuSfrWxQ1zSyeq6mDJ0S+Iy1CxdKHa324IxRuH
t9FTffRvRrs/RyhsKyCiDVXxWHTJuS4PnlMdBTH+I251+ccMedPrrVENSlQRarXrqtIHiN73hsLd
pLEOGTAfKF6ICIQi1mQQ+Eg1Dy9XNT+dXPtdkTIEhJu3Yv+CmFXhcTO+a/+IojseaBkzKdDb2t2T
znQbxHZJWhQICpviLEhoX5C1yxW93GRo7wB0q3RW73xuDrS4AduDla3ZdeS3Qj4giLpFMsxh+e8h
W/3MuoxKRUlq+9aELFcxGPI2zshnykBbw05XOKyMB91jsQlKAwpShv3sSSAOjzNVQQtGoG14+Lyp
S5KUBCms/0lgTNS0g7DISjE197ixAHXYCjZkUTnmR/pfgFE4YQoNkeeOJ8iUCS3b1P3zTE7owR8g
TzUgNBMvsRJj4tAx6WRLoGvZJBS15keA4/pQ6fP/leQtyZM/bn3mXIk2reaEXLKpMG1SzxNUGf0G
Y637pD82sTGJoHdxrhPIDMuO8C6AHrpH58IDH5VdOaEealdLv/m0eHZJlG3gfyd3AYAE7HOiKoqp
awb2GZOibQ9cqPI7V7EqBLElXt5pLPsMHhz3RGdNwCiH+GnReSrVYKlXEHGryZeOaVvajpg3H06P
dfjunShghTiNx4C+0Zw4NQMUQnlLfczQGgbR1ZdF0LkbQmrir7JhYEq+ZDVlrktRRBi2EQCwhD0e
LLyJXdmhtULF7h/AJELklYJ3ptAmXZtiDnklndn3sn+oWm0kplW/3sjmsjI4t7ZgX86Lw+1S8hfS
2055GpPJn1m9TfaZNVqtDMEwiP7S87tvrP9uWHhgtJ+iDdn/Ayym8hOTmcdQRgyMuo5jp3WX3Aqj
eOp6p9xSABSy+SCsj3Zr04bvdejvtyr9lu7kiWkYo0q5sDkAPEGzmT6kyIFcUGN0gWr4Ei+q/O/D
xcOf0sXbcHLYxrDgSXjmdtvo4mJgxZqYZZCpgeeK1FV5X604GljxBvTfKn/+U9FXcinc7SWv6n2y
/KKilO4P3KGAnzlBeE8xE2Az57hDa0orVLREE9AM+QGviMcW3W3Ah2Z6tzDXr+RwnUF+yzaTzPeJ
f0iOJofqdYMohGZ9tykK74wfbz310Sk0UK0pCPdbY9m4gfBrt7KYH7Q2p2cY+lryJHzfYGZR+O4T
CG6QbtJ7n7dXELDvjcR22k8NmpUqMVdbNbHxrbR2JBfSRenUp/e8V2dSsoa4dPdgO8peYJ8bazEm
QaIjq5kw7FN1kNd4OfxqFtdoQJzlFZ0keaE8KPQz4qo5hQwWn/Hgurv6y7QsqAGTGWAKr4lrwe+g
jshZi5QJiSnyfj3JMG3D+u3HRJVbx+BXFORndv/g8zcdhVgrFLXazJrK7/zM2BJZ0W3R6iJo1V3Z
qV8uPVFg+HA1wK0vumeLAY+on+8kKTmGPFIjQV0a7/aQmIdgjFa9KSTIEsMY9UaWCGc5iRne/Iba
dTgS4W6AYn2kfjK1MEFqfq74R9HNppv6teljiVSqYUCS3yM8H6MlfE7eYRvdR0HLaopGYvvwBtHU
VIw2FRDSQUCzb9jRHh9h18HEQEi/aI54OKbIlDdrsFOefhZhIPAhStMSCAtF8tJ1xll34tQ9S50i
kEMnuZhKLn5oGrGHDKBV5hXgLK4rNoIkgJ3wNCp92ptCdKibyOSOjGJuzXcnGm+0hKGj0nDMZyZL
97mWxet+CHJGv0T7n62fHzLDCkB0W79A6k2UotK+C/e8K4iZ64v2GPjYk5YdVTWbZ9p2BNAxbEg1
rxgd8cqJUe8Gcl86ssipWRJipkUvDe1q5FD7msOk6+sFJ7gAq16OLxKinVW9uPQ3qk5HBJT+nVU/
mkaRUiCI8p9KkXoG0o4HeuUx3KEVBoMm1tbyrrmcHA+8H67CgIRtodLaRXm32yXceyBrcsjZSfBo
L5vwx7qY2yghR8P8SXnbKhVPg5GH4mPAkiJt3bmjPYroEqQ23cIsGQKnvhTYfqkVSRDwLMb4R9LP
ycLRXyxLyh9DxU3spt1QHb08FcOaYZDfS4xXV0+9ONCas62YRbZk/SoMH+8eVTV18pTqMZ1ytq39
5R9czNLDT518abW7eDrioEhjaMezkJeQZxmrqsMb2EY4WnE3RuPN3Al5B8QW2U6J417onk0/36lV
6MRCp/1H2RJQceJoBAJeNIKukP2v2jlYKfpRF0gYCqPs7irBfBytdAiLsvZtN+bk0VnulE7EZMox
FyWx13K/4nmHlZDrf36H5m23rs7vAHofn10Q4M0Q+kbrUu2upc4puHZo39zGSclGwGGRmAlAFwWN
fbl/vjX6ZaUX2yElZEy3XMtr8WFPyaIMIqSeycPWlAr7avpfIglBoVYNTbmSoUAIGnuLFUTjQihW
is1Rqak/Fb3t0ubP4IgdWE4B464twE2JaTyGzc8LAgwbdUzp4D6+xXi/WillyhHB+lBFks1HFG/T
JzoUIVNE94j9VRpgwCC+x2RFIv3c/LgJUJpd8lqoJA8H9y161PcWbZExZW8QaAbgum54dGeYwyTJ
pml6CV11uM3kcVMpYfWvVfBhV9cCORkVwsT+dj+jICngGv8GApq4NK97+B1IgeAJ/tNp3U55sA9I
f1oxkWBrG5fqnLiMHDmJYY+jYvIHfw9wp3xxiYC/LPMbkgv3WsyLQ4X9WaBHqMdjmZnSrCkS2HeP
x9I8XVr/+4W8bWi6PC9v7nR2xtGcj4EiE2ZCl/R+3g4BHwxUSQhTdidqhZrNlzA+IG6ufrQVSdD0
yeXNZ3PfUDwQPmChAIxAlxa9QVioCo+DfQs8b8WpUJwxMHDWyqFD4MwwRN2+rwJGkDHCx6ulSKM5
Aoe87ebIJaPNgBRSVuXK4lab+NSAnjE3rVPJSuHO7FuUOpDj5DFCQjiK0UMCCMFdy7MwuMvwxK27
GzCdKzunjNe5v3zO8vbCis/hRy7kALcWK4Fw24AGWtADsQxHUBD64Y1ypiKdQxhtPnh+/RACxDFq
//wZyFE7UTh6y55sV5S6PtX9z6HyEgTbQuP+JROgfjIEE180jRXsgsWJ6meBosqdCaFKZXqxNVxS
hvo3l5hC2uvqpKzyUlLRl/393mCPlRsviyOVvNJ9ExdooKSIq781HeTbTolC1y8wUBd70LgtXjq6
lOAYwSOlGEfR1FGXYc5I+2MceIRhVjIasx62tca88FI5H9iAF5KVm68PEGd8xPNo3l2J+uxxWO6Y
vggcq9i9PU2FMRh7h9N/oXKsyJn8nMNv84n9wEEOFo3Zn9/caSTGz5NPz1O3pZIrWm2mJZ7V/caM
uQacwdhxbuLNUefoq84wY/xXosYuKFQ8IuQPJ4oYze2bL3Bggfv0xbKyxQY8QbrqZVdaFXmZBmqh
gu7ZMSkByhYrhTpipMtqEFhRpH6ZSbuR/IGR770KbzpIvRu9GjS/nVXlcBCpUYslzunz1/X5TCEE
X75YFx1LBK2vuvVGY50rvaeiea/iH9g89Cy91YsOVuxtk8z5Qf5iEul5oqkfDBZJB7q7G0jCtD5b
/Qy+U2gNqyNZUV4htVnPChTCgUtL+1qhuUziCv16uDa8OFPfGWPugOxrKwPLI9P5HT5G1lqGJArO
nKsFTvwMnRRN8/R+kPZlXNWMxzmgR3q9auw1Eqy/Fb8PMlVmhx3JIyMjYZaqA033wraXvOgEr3+3
q4qDaxOYErZXLB5krXl8IEN2ykNehYXGkVqqT53F3k18914jp7HZYIF/pWq5UqQJnzhjq/ajJ2cn
Kt5CKHc9VFrIZmMU14tLPKxtLG2KeAxSQjzNBzVrMBwW3q6OJw5X1ssMK3S4CNXGruCy6d1oXVvC
lEtqdXl52gTqBoFsCSSR5SPzKeyCVs5tUm25uGeGfAqSwgbBxpPvDarpTe5AC19EnJgAk4hhA08m
cz0YFXgntzz6sPXxddvjVrtXnCB+lCm5CbK9u+rbhkHCVxgSQwnPYs2PXD3WEacavlb4Wkof3Ju8
iN8kfbZYFZY+SjfUA2oftNG96djJeaZeAjD1NZSRgpBn2bCWkIbVky1Rh8utwCO4UWcqpeEzYj79
h8VRgmTZu6tkzxobEAr9q9coTYySEwmCcbck2yjz6XSq5J0tDaos/NnDCOKdPkL4iZ8ybkGnCFGh
JhyFOow18Vo9UOiBjDTQngV0x34qoMooItmMgGV7zIy+5XzpT1XqWDkc0i0zlJQ0pkX88pRqGqIc
oGVsxTL+aL3jNYJK/NtVLhL0TyujEVdBs32tO77Ftc4pK5oMGU8vTXe5pkJnCAWXkQvm46dMjCQg
Ob5kZn9YbnDC0pGat73QZIFeltBGWbsnFkLfY/C28ApQcYm29W4QJwYXN8LihKpAIKT9Vm4DHTK2
NrZxZYA3b5U5GYKsOSYeOkZJajtDEe38FoUEMAyMZ/n0fskZ7IiisM2NFrqb17AoOTL6GS/FoS5a
w/IJR94YLor+8ZzBQ+ZBapWlgvKw9ZkLTyegg9XnWoK4xm49rNKdtxn8C1T36vc+wg3JdZx0Eq3x
6bLQq63cXJS7LTZuuB9neemQEnEEC+5SzYJni+ZJEuYyLBFXPwghV78GRRPtqB/FlThcNuDpAZN5
R+Zy+Pb3FPaZ+IBkC/VPA2KeF3u+epyfFZ/SuUuZyaPlg8rtQdijKnmXwtNnJgfKyXwoDZp1DIcT
5En1wC2E9tQD0q2VIaUG0qNlAJyWfptbfuKVOVeaAoWLwOuhBXV+zp+xdT3r0cjfhq+irybb7AE1
f8HLb6wzrXhQ3KaIB0Ag5Atwivx8PCsImIfZX3XEECTjk/v2+3bzUo4a48fSeLSPcSJjIy9q8Uec
HDJ5iY0Xwfh3x5BI6Q/VGWj/jsmjUE0TuF4iODqUWd0IsrC8ULNoCq6CxoXW9p08YkOMSQjSFXeq
uKrocDIIm+z+qInfQBYrX9UU5R/pfxWe68sgSefgFV8ZcbCX468VTLZnK7HijCUcRFPhvjhcPyjn
O9X7hVyb/bs9J7PPe4ImZSgf3MRQwdyNdXK02MD6j/baUdEUEwYhVVl83TvxuJjkaCBWxGTGUrn3
YBCPLE7Q8+e0udN3VGE9ETjTMwAI8D7xpe5rxgNGN9lMmH+jxjJ2ZZ3QcviqgSvqAAsFOHF6ldt8
ymmIiGgwA1cu0q2L9fC5Zs3RLpsMZ/4TSIPPjwNzhzPs+o3aiiDLmi1YMjspNW0XS/21h3hSY0pp
j1K4upYTjV7tb1hWf9VaKLfwa8Jq//4f+aCjUsCAMaKh/xI4cqYNZSUorHZlDrShgX7VLoE1ICva
mHoMzS4fEsGowTgyEPEeqooX6iyjqKpiZSpXDL0rq8CBV8MNr3hJ5xdrYCwkGNChFQTBv+iSpmAW
0/2yziq9EbkSRvSp79fzL2W1tMJvstPtSZPaodhUeG7vH8N9JEeLfNhF8NtBbD7w1+ch3Keq+Fe5
j4WLgyZC3lB+sR51IlUZ7kkSQUJ3sQWWPR5Esd+cAFnY+x0vLjvzUVwxm0Ux+uQ3nPRWlOVlM7Jg
uJKznAN+LbISUCb3Dmrze3aR2wbNTZwNDcPAkpQjzWCS79FUblSWgWQxxa8twAIn6Ulx/E42AjpZ
G/eUSJl/lKQSnC/9rBhyr/Ls/9nUEWmQvrvFF2tG4zvxZUSGM8g8qU8j1a6ByH6ByHwUrwCZdDqo
GrUrQ/liwZkbFh6hbxjXXjuKKUHG6jI6tlnPik2CmPbD7DqbVXKFYOLd0vOko9psc61YqdzahGDQ
VGqHq6tPzJsz7ZrDSWaCvrZ40ppjx9rHVXLNolXV2/QxZMZDORZTJo5EcrpU/BTiaW/sEJYTQNCl
l9EXvX7CWMi3HSELWHxqcP1WnZsw+Irwedk8nG7HqQ6ipiE5jBiwbo0YPNujYvliD6ClRRW7984J
cumY8eIhcxUR1hoa2k8XV7YtCxswiM+7IpUqlKTXC5DG0P5SDGUvoFiH98LmpW+T2luVtg8Q20/D
yAcJHiHea8CpeghgtfEehyKCpJ3ZSGxgnrP4gSQciSTrvWq0OR49gxmTkmJd4N7+HBmtL9aDoquW
TKEQG4TyxXApaHM5pyRchpnbPz0ThHjy2mzgC0XiQWkIcgZvmL0Ro3p7XZjdct8PAUig9tm5URWt
shKDPlq9KuF8KgR/V+uCl0Jk7HwYpKXDV4GWaEDckct9rzfWJrvxEjXUZ9I4SDZuzQDbbC60o1t6
+SEzqYIzmHfc5YwNOowtrg+wZ/3fHcHjI/UpA7qr/TMKs9/CCm2JvQHcCKKcoDd+faIbjND7U5Rs
UV6pnCMtoDv7at9WsUoOGAW6mmIrTK0zfLlKp6jczSeg6KGwBl/lMgGYol45bUEbxobgUIKUoxyp
0supzmcj6O/eM+nJvwb6TYox8ZWFvQLBZF9I8F9tnYDzJZ04OY67PCQyrQ1X7aJngi8QwrwOA0J9
1VEXx06iACtNg79e9l558nsb2OTQPY57QWNljJ05XO1k9U7VMkeE2Y4y0UnnoNw1T0XoB7pLaNe/
/4G3C7JuK+NBUAraX24KIKbP3zO0li7m9VOxlccuSznTUlb/r2rAe19uRhBmPvnKc41IXQf3Va8R
HZMaG3/XJUNnuK+UkWEAN/vN2IW7+9090BRrcp16Zc7GYrEg5bnOlc3dNdsL5K0X5+WKRi+OEclw
a2VxznzVn3mQqpQRxsD1lYjC0M9fzwPW7VwDw0Q2BwPhLmBqRAlSvMlkkZtDEvLsllAYpcZ/IDsl
d8Kzol40SUznUerhIPs4e2aW4ZmfEloPbwcJif4mlVd2rRnpfbZnixA4hFWWFhiVm3XD4Qzb71lM
l7clBjX170ejZYzTnqsA/BvocZ2qVrSSZkIfiaCQh1F29Xg/qTRSdD6rQBRsVmFWRNI3rG8dkydl
XdkCSFjSjhec/UHCBmHgb7R729zriniUQPSNmi0U1r6GEQ3vbFY8P2aHMcFBchbdn20WWPW1sStu
VYq4yL2LVtCc0micC7MOoh32Xj/wZDYwRupavmBJLnwwMvUKJnUXMed+vsq++IlP4LEZW2HpceDH
RItTQxUwHUnU/XKMJDB1uA6pr9VtmAjlHieTfKF62Kw2JsZS/5KTrc6yV/C8ywXPUcg7mokooiaq
pHKkf2xEhb5aAplPiBz+QN2qHxi9ZVyPWxvUxxBuphZ4lomTHSIxyV3psMiDgk44w33Dr73EyrYy
lm8rOtiL/I//CfXVVp9C2yMR7Zy7plMDdQqXqyZuixU+JfudKyhSVdWfhdWPTdODxMDfP9G4xV8a
SqXsAfkakrslMaF0F0uO5TQkpKZKzXnqlczkA3FPVqXjDpt9tTGKBbHRAbLWQpLebo6pMrOxBSTg
Ws5RXHk3lGpxOaYH+y60I8CzoiDJ8R8mBitKcjGlw2dfxFhtFcySWkGyWC0TRbcKzQncZSsht/ka
dgkrbbw5EERB9WiSqqotNtk+RwuP04RYBOi9av3ZRx8+abi5UvOUN7QBEixndYAXS5aTpu10T3He
cBqZsow+SJGCpOP7SFdAjF26uLKFTrSBLNa3MteOIE0nVqR1NkwYPhwtNFOExc0Ckrr6ygWMRJCj
9mZI9FulYBKavBNAimK73QOX+Rr8cUkjuZWw43cFYqJOrpnwTsuHRqUANsja3xtJ3LwJz79pjtzu
20Ez+eRm56vj+uTwhpmEA843Ql4gWup8y+TjSyhc06vqrF54zeyjkHM6N1dwzoLo/mXmp/bHTH1I
7fRPGpI3M5ns3X/dR0vhAvispurEj+0dQvkfBgvB5s3NxIPyxrYb/Fmxr4BmUBEcEmUPoTweN3C5
8mM/QjcIWx0hEyxxA3ejtY7I5fHp4ifzkl5xNLEceOHE4U18BvPtbjlss2rYYtlPv7bV6wRKz/4S
1NymPPISV8ngbyMNI+8tGuAF6nKL4YrtawZxJlBDJylfwZD8XZsvvABl73fbulYJg2+s7zKyUpDz
F+Md7NoRmsHdq9gjBoE5Z5a2qkOLoJ/Wss4Eajds9WFli16udrfI8a2CW7GWPvVm0SEPlSHX7xLQ
78teXo22imut5dVdujQJ7mGouNiFbPsgJRPUll79dbXIX+y0TVDZhRj+kEiFDBc5O1sm4HUjE1p3
ioJNGEX/afAjGPhyKl/nsXHmXCmQ3dTeIbq8zfweRjmgrukX+yj/o/5a2EGs2c7Zve5g3hW1ixIF
dZ7E2w6Y0DD5muUnEF1efsrPI7LaVsB6fH51S/a+qI9s78ijT1VmqXSbyoFgcCrUrnLFW8UIuMgd
ZuhEjLWK6HaqJQnhJbp4HOS9il6UEyG5d4VetSWItFSRckwylOAslGg1qkVeVhZIcWYg2/+PVz2K
NqVSl385Oq5gYThhHAMkGz3okpYCYxMGMsYibKPwaFPHNTSMuhmXZeh/oUXvyDV5xWQxgP6Gpb0A
U0uJn4q+msElHhHRwLowPtl7AgHYh3i9klSn4Fz2ycIH4h32P021zKP5NVIU4d2Zpav3HFLPd3MQ
rA0qoZjutQwZZdNbrZ8Z83wwElTeVWWRVJ3Ntr2fheDlOq528RW28F/s7/ALqHRPZ8I8lUx9ZEto
7+haCK0HsZPNrdKVZ34HfN5HhvM1YmYSChQkNcrqapg9ZNUP3LHUz3bbjID9Hlo9nAJWysP88adj
YrKIocaopvBncwPBrW3+yUgzuHs4Ug6AxHNe5lkn/HcGlXya71g+XcrrXNNtZocCN4XfJyXu+r6K
FWFbB9b9KKRlBzYua0WJw9rT8rNGE2Hc+PJl50a0zpMNYDET0McIcqHjtCvamgWExh8R2Eoyn7R7
/MY1mtE8m3za89Z+MeVMX05+E641Y513HeOpTCv1Gbq7aZa3UWzWItcelEJvZfG7Y6Kk0DsvGn7F
h2ZE/BVWFGQVFmB31P0n7PksULOex4nKFNvjsITEXIp2bjVLHaGtvnKsRnPrciF89xwzqNQZstP2
yDSASCbR39p4ftJU7yutpeUQ07OimbjDrzXNn5z5h1t4aTNsTouGRAm/Rz6M+Z//EjyduMCAtTiC
ROd5043NYxcc55lwqxIfpV7lhbSGoTSZ9qZcvGYpDiqDDFwFd3gnxaQEzXAekx1ZWYDL8npqPY5a
91anMwTCFoPQAUQBtACvPFvYz9v2P+Rp5nX/Qc3MVdSbJZgt/tI3r2n7W4Y4aDtR8j9jy6C/PPAb
UhwtcZd413oqDkT8TKOFgUHz4j7QZrYZ9pHFKYtN3V5pnlftbqpvxkcLwMI0j6RTCfprFt/ApgPr
5RpHPiEMptC5Z/Y6gaULwRbJCx0ZQoQ8nCqzBP8+BQRJ7qUmL0PFFgk1AP9/pMRAVzaOWIUBue6e
52s0ZKJFw93EKnodHLRVRPfCgVJtob2gSPg7t7rVxuGKmKuUkHUBymia8pNF4/CeBWHmpf22pxN5
KP/JcSkDRCCncm2bIMU4mlKnbiOETorZhdpMl6OfsRocK+KbuXdDdepN///11eFHi0v2t+8p49Ht
eFURAsCQoQNtgVDNijdWXMcpuAVEUd5ch82vJy6ZOW1LuqvVnEMe/o22xuWN+NKp6ZxZdasIrdkD
hn0WYw5uvaf8UsmSzoZbdg2O3sJlYVYsjrtmIYNCPfR23bIR0hPMWdVATSkkHpIbRKRzOIFtKZit
I2tIxjVUay9ul+lv0tGQcP7+1JwS72rbV7N0UGwcWppoSTnEzbeznYNF2K3Yw0bWlh6GZm1ADE2G
QavAbcPhA13qxhg2ODPp+5nomZ+ebrG/xFERFmSlqbybE8JuK8zKQoXcXa2K+vAOH5xaduUbgN71
0QuwqXEnQMNyiRb5lSIzwNkfp8b2KSJ0rjhtk+lMV+Q/AYH1f/CAmujY34xh+uh0xuYrZ9sr7f+T
LWL/+VujtguU+kIlZhLU5vFs84uEXL50jnEIACcliErj3o0/Mr95AGfD35ZsSWppjbOAr30oujBJ
M3K+T+2gkeez4mcccWJidyuPtrYINl3vZVrmo6lI2sb+sPg7caD0teEFb1KuOI8kS2MrcQDCbkED
6oDTaYoWNQcOfBX0botK2sLSDaDKJHlLcZ/lY59TFFoBqx0duVhNpGv4DyN6VDaGHyrxwPQi+MtH
pt2w4WeyRIjJQg++KnsR0bGzQfrJvP4wc2HrsBShF951tPQyjlCgwGES0vE5ZoI3S5P6D+xrXo5k
GXV1P/2QWd6SHzAGyPBG5Bn7WpXCn37YNTRrNlfhXuSPgsJ2SS3WUHCfqDI3DfAHpck4vMw0sSBo
+0VWUIuu0JXvjNH+NFU5CLRXbLJKM9io+Tha3OG9J+M6IL9ob4IwxoUz20UhN5k1SDpDiU2u3AXH
OCqPnYbTZcOKFRrbFhiHaivUsO91zvvFLih9rZ/cfQvnFmjeqY1dnlftwHL03LP5xbeHUiMUstjn
2Yv3GqR7EtFv7fFO2zZyKAh/w65zHfaKf4JLwOCdPvqacMZrnPSkTWLLkfFbpU63g+EsBXbFHQ6r
7Wewqk6si1rUuRune8SUBkWelZ+thpyE8vuz+5bev9Oc1g40chXGxzdzHSd+EtgvT4QWKsouiQUd
/YoSqbt9sqdeToQEV7P6vMb56JJUdU0g7s+xXW1TPsGLUCAeDf2yOxXir9FpugzqSpGkEISlBffG
eCBy1Gzhe/zs+4OjkqzP565W6IDfm05CHEeW8WEem/zrzZLao/7rCn+DT4P1bQBNiVVxMjlKCnbm
7JMWgfk3Ietdg3mfq7BnG3m2mVJ6vjdYcvUYln6BX+7kcMypnTERcV1B5S8BFFRSbSkskeJSSX4V
CfFCC/Ue8K8ajSFpqy1/8+4yrCoiJCL0BesifCEvGnrC1wYcLZ6CzHHuUiQNp8xE6R0BvMozYO0G
WmpxQW/5LD94lZQ809a0kgkMLyJnZPxvgjms6jRpEiCb+f8jzTP/ektkP7VEZa49B9SaCmePi8f6
nIWuna3JdxOEKtdYwGvmYANhyKnQTTDgsSiSOgnrTYGm7XTbxYaikUo+AfZa5Vp6EUoaaTw2bYrQ
jGtnyov5DTVMgkVBHnOMJFjmEb+ekhkRo/zmzh72PtYpTcm9YkTxLu4avsP9qrq9pffdlmKOnjVJ
prn51DhUBIVqQzlyJwV+a7ngYnVYjfw71LXtnUvhrmEUdSMsOJKa45mhzaUXSE1C7hxN6/BfnhrY
lWzPC/sCI9t3tK5hEip8UHtp2Sl4+j6xq4OjUtn44j/lrSQq5lb2sByqiNUXceC9gBKHXfo5n/X/
H72Lr8iPUUqx4tR33uLaPdPsTjkB2qDL4NvjDeyzAPTGu1DMv/bx6M2aPYAHySsPfIA/TCPyuNZV
92R93qTD+6NmQEGNgUwi7v0fXoVlgu0TU34uEW0RezYHfhUpXEevmdYsBZhXBVmJB6GmvxORxkCP
u0GXaNoIlTz1UWFEdl2trtjekZckgOBfzsFLTdfc+75fBqMSY3VLdRnNIewQ/2px60MC7oCQTpFK
7mVt4MGQSNgG2d+LQMi+bz/EUfhocS+4124QLI/bQoXjmnWfrbREUsRKvXYaV3Ka2TDWa9QItHe3
lW4kF66BShX59Aw28aS3SlF4wd8xkrQzTwdUsTJu0pmGyNz7gl6n44BRXZvkuNg+z1jpyFIjFa+n
idZsnMG44d/yL4A3WFVeeLL/0mMrbr+xqktxhCtWpsRAg8QNzEnImnjPKL80qYTbjD2tDOsXdRCp
n5cHdA44j67wuOI9z5vkCRhslKZ9LH7ddqgN7tyU/v4xROzKKKqgbVwSKmKzJryLPonAvONSPfVB
jWvH0HtaV60OmDFpOZI4HtKTGKdm4HE+RL1PCJLa6Z+hulsGuoyO8C/DaZjQKa50S2a5LLoCJ4Gz
yP4Hrh2dfn03XHD+7qV5jYtJlim4UzKkSOPEXh+jSGj/+YSHEJ6A4jxL+pnq/V7r5gyfTSg+P7Ew
MEOKfYEcDH22+yF3fpq55QDn4sLTNFXp8qP9a8ZqKlbpCU6vjYqYng68BxVBYgnLlHVohnZgMWVv
zQuQfxTaOs8kBidSJGV0EOtNvvQMmTIMY2vJtfopqqdW8L/2wx8XtWa4gL2iZSyGmxPadE6ZFMFH
MuaozeHCGsz3jCkajZeeaUp2UXVcX09UODcIKkSs0Q8dgz4HxTkTVXhJjIHXd+5DmHEkdPwbtrKV
ktoeB/Xz0O5Xls3A0oyGC9admEZmJSbZXfalX8TsuwQEsEaFm7CwDciToDJW1yJJH1Q4bol8ZF9f
MVMUB/6kAvD92WxyG0Qfh3/plNaSRcNzZNIvtWNHt2pRh/NOcDpUF5YSkGSFTRClttqzuedTSpkt
oziYSbhFzwNQOGOPuhkQCozGxB0vUmE8aOhA/v5JQJh7211hUcgi7lDkyBUWnr3Rp4WtJtYPOy61
w4JantXkizQWUcb/ATzf7UxURoN0jJCQxGfwVc5Qh/D4iOUdsn2CqCEDGCn16s+4Hijextngm1vK
4fwMy7XWnflRE7ZKxzrAuzfB18xkFz1lkt3nyz2Hi8BC7X9JrMDbBoFfrqYbNVc9CdLLnqukn7zQ
iiqtZxt2WmaqX93ASLY64sEZjD1sFuh0NBI0TwlFppdpMaU0QPSaA9SLDxTt0XTom2QjwBJX0dO7
1ql25avecsUV0GGwB9rThaigmdlldVlGfItF+4kiiBp0jBy0eUqRvUIEllj2xuDuHNyftZxwapJl
VPJ74yfKUXyR7bUZHbPVWL1Rp2p4dsPFVY9Cq137a5aoUATa5Jravuu3W6mGr57WpUK2UgeADBzk
Rge8alC6/oQ63IMwRZjPNElfaPxvleiu4ySB2p78uf97Y/yO+j1xkGSxza9WBnBVgU9Qjy29EL+A
IXtIDNAOeyqmP/80S0z+nZppt6oFfTUfh8MS7UQK8Aq8W5J+NdoZVkuc6F3v18DbH48x4ku1vfl9
8zITXzpEuKf+RzTiRnK54RUTlIEo4q2HOVtlLbuY+Xjxsg648IbYRiwQTQCfnHgYBgSt8A0eebE0
jFhvKY5vY/w0jXDBFXS3Nxd7hbfEY/9IouXBwN7FGqBX4efRZ3LfrnJTr8utMEEV4JSzN8/P6p50
ZJASZnYs54MR6eHEf++t0NS2QJx0B9/GYF9bp8CAwRywFuEHDIQ0uVS9fb/NV9RCrCLS9jNIERFm
5zfZX1TjVhxm1M6Rkly72abOyfjdIWLUCtpqEGFkNL/AZH9w4SsxaP2aaId5GN49OX6OQrscWZcq
/SXK7WO8V6yojeFjeKlMoLfKAbWUNhKY05lPHhHPBOAVDfk6nGJ9MhNmEN4TV1Hj7NNrA1/xBIuf
CoIe8aPwAidUSprWOv6TsC4cO6PeR7aSC1RikeOATuov8n7L+xL1PEpHEIlFzemXFXRgfIhlBoG9
PlXbb06C2vkuh7ra+oiu/rTG7bP7/ygaNbrwUD7OK4tnelMx6fIHXnHvc842vlEDgfhGSbNFZLen
N5qKAnW6mKZICzxjbkIm2j50AbDoRb5mwMOUefwcVmcKOeMEsE7cqgA29Huay7WojjC6uzxvbLYz
jMQ7uU08UAJ2HSm6NO2qXn07E5z95rV7ElDW2gZlpfh3k7BJZruzu1OasqirKszipXWFBy+rcfUi
fPoy1QD21kPVS1m3r/+S35gVUmfq7FBEmTOCFm2XYn1dzRXHy0aPOwZzyfLHmkG8b6SVUJhlQNG6
tYQXDaLR033djrvpdMk6OfMqXqKsBW+R3BfGfKZNc4lrkkPgS+zg63Ykqjnc7UnoFy4vTTkCGXuF
Y1F9m/oiKIvYtlAWiaigbVPRP9Q1xRdBV/8+Nnjeta8TzWO7kNMJ4qtdzLWQ4KEz8QVgUbmG4aCV
8aOTPvwoFESMBrXW1HN37YjhjtpijO39eOqT8ZHnRU2qsk46fu/ct/yb5OHb/Lx1IDoQWIFuPHjC
2b3bcRV2BRiU2V/X1xNpxvANQVu+c1BVWuU8s4vC1v4o2Z9PuO24GQM57gRiaEHpaxSRL29qNVmT
C5PztI60tFa9fD/Ct+vTl0tO92Dzj+WkDItHhsW7kmLy2rgQHSgCCou3GLMoZsDaUJvFXz8ogDH3
UCgv4RIQh97iltMMu6QJNMd8J5FQWqqgT50GaqkSzekIYdP0mnOYBdk58re2CWiO6wVtEpsSUNZ7
zjoN32F9cgzKxyhHsrx024WMqlys0GwU3mU1GUudGgP5wMTg5uFCFwfWGPWW31OTqVF0OZA1Lj6x
mxJlSmAaNE5sIUV7YlbL41GxAO+lFzZuVe5xH7uxJntCVgKqvwDDQVQ5qdADqtGYL7hPL57Am/Rh
1+dNCmIdpSW/0yJ9EHlpqIBS14nW9WEeTyGSCvHR6ijDI5JNxwfemm3KLJu9zEDU8ETpRyxhA4OQ
prjP6HKnumOWfFWppyETyLq9eEzdU7BlUg9+wj6jD7tc6TzLqSsV+XIBdQVOQipTFvsvZrTI04df
UpBU30kkVwfvwmObjcGIA9wvC0hBo+A/CngV2VxtBheAjGdSHqaK9XsYL0+Xeqyb2WVCzFpapFPs
XdX8lj7VsUcAbf2ASzJ0g39rtA+6e0fVB+T+XbC93fAwC6837SlfE+J4/xFzytajNKWpDZyHmDUA
cJ2uOp6+ZxunEsSeFKSS1Q6PHdIcmtlN0b1LDqVbmNgWOqraG/flSYHyzw2mCHwwwOmWdz4mDhXJ
BN6lxDhYt0P3Mh1NtdFcpW02v0dQCpyHK2isO+5N9hp2AmqrOWv4ZrHc2Wp1/MAvSmkZ6UqVk/Ld
s4yaYVcE1wtHbJ7MOCsdW1h5+LGntLa+qG3wCKT10wxVUP6qdipXxZsPiSzHuagOSABZNvEn8r3o
YqzYxAw95tDqDnVG76sPYQwp0PpZ6OqBwMynEFUzAH0xufBWOdRz1vLj3BAbAr9f45wQkfvUUHOZ
2G3rsOkyAR/8DrfGSlyJU9UMufW/9UgMrRR8nDJ4JolbNN/xQlY+OglQ0DfrACO8UlH4PiQ1wB2t
9SyXvOZG4ein+fPj92+04rw7cVMkQx6FKrIdZePJA05XAYK12CrnlSBU+6dbu5I3or/Uhs29AIDA
m/J5B8yDnwLtfWyd5thr0DIvWf3z2x7XPBl9rEQ64AE0lqcKnl6yYqxBwi6cQ05llB5yt+oWg0Sm
gH2flh5Gptkib2XP7XQ+SjHhCF+BhX3+st3RkPZbs51fW1xdUuB88GGLS2anmsSqG+0ybwhzHHdX
pOT2EAiJfBYIXoH0QKmzowXsfUxoAk0kq+BHaBmeD6H0vb3xIVMrZynZK137xhAzBVt/WCGgnkaP
ylhof6VJZTjoNSDJ7U6ff6IHBUceHQZHDNxdkqf/jb/km9wKbf6ArMvDJjj7kvfFoN9Hajk9OP46
vTZHByZfhjkLyut2925sUQ11de0do6DpbUKXMBRh2hYmZ/JzsvQ0Aa741TafF1daKHgpev7MHd51
weuj73+s7blU26bk2iFQD5PNlZGW/K6dkpL6O1WCr7QD1joXlVWxSDfEU6lxcBgQxU/8eLl1Qy9k
H7K8lKjFbl8pIizXXCuZAw1QEQsnPaDBgVhFKGQ5oIms+r1LZKX19S7WWKmBBHjLyMDygRYyxsbV
aFLMmM95nTfSOirGgScypnlh2pfr0f0qB02fR/b/ZgCzBmZdgbJ5L/uRPA6v5igUW31F1Gn53tk2
NCDM0ukC5Fd01mQvfnHvLjFyHX2JhVNc0cfzVZjYyoYefkxUfYIDV/Dv/u2kaPR3mDYY2aeJOpOx
jC2k7HAQh2l3h8qYK7XcLgxivVMV1SK6HlDOcbCvhywO1zmbNlBgYrRTRRAxoBcZGhSV0sLSFQk9
XpC5ZW0bMjDwZXprnX1nZuQTVusYn1iLO5ur2kKhFKHZB5ZAepBmw98cEEsqZvjrl8vpkqiTk1Nh
u815PJ9meYtOm2ofmWh1RopOguL7HGyz2FRWwVsHXPTA/t73tLXHAxJ54jzNBX0kJwcfVYvr2afp
nFNGgW9Vs/tbl+pnhEwA5OZEkTxe5/riWz5AeNRAhV4kmWqkvym5GvTFLL+hSIKcMkfPW8J7q+6w
ePqnm/mxaCcDHUoTWZo9xKEUn+0HiTAcElRCRzaruJKDj2+F+4hc8SkUAGU/+DF+tT2aqNaJ041d
sTWueYaKVnE6XQFPg6DQJaTjvwDo+qilzc8SP+EoSyglyESfJs8YPkavIxP/2Z6lkSKGIEnWkwgn
xMLmoN7Ww1ecmFKwCZvx6NjTJQslXjbIOPcoJGRvjRRYZoPKGW/DWwWh/KXnT4uhbiiz15jh5j7T
JivAF/PGTNn66nihBbFUg9jwCnPeAVqdvPxeLet09MM+oIYI/tTM6yNz+HvU+qBthuKG0SBq1WfY
XFOC0M7cQ4/G7u2niwNfvC5mmFM/N0fJRoPQ2QTlQUG349jrMD+eGFLFolmE6OlfD8eVGP1rmbo+
/sGX8OVOof7S9pvpOo3/xqTMLE1micJUXx9Ph3X9rrih7F6MBxmFuGbVINK6bEes8OaSR1Dh/AK+
pDH+mUPvP9uif/FfH9sCfacmGjHWf9Mgn+DudHJ0vdmIiz1CT7dg13+5H4A0TVuvfVfhD51KIX49
DaXELwxMCTtVo4Ik+1V7RVbQiv6Ov8iK8TQgUDQqukHNcIjOZ+NABEZ+NHX7hE9ujBezc47fTAgx
Msnc//WElLOINutUSfx2kOPGu/Vf5y0sj7UT3/Rw8O63kxNoa7HiM2C/bUgglGdNmvKiwqw5YKHk
stmtOj0lCe/yngM2zkLbjTbOyEklPsalVhKwvDRAh6ASbR/CBxAjjPqT1tY89ZErCoc82PPQrC0v
R/eXkuMpR0qxGy1ilsrRDa4TuWOIyE9rVJSC70QSBYxNYfRKwj0df/6P8Oe9peufQbyKBzTxqYRL
ww5XBzc00o4TAUG59KDZOqMa/XLlHN+t2kMdCPGs1P13n+dLgQtTKlK4EgQewLhTH3+F9Bj9tSeG
2lVkedAKMxYgnugMO0fuAi1gf8rFApDTgUz8+xCLk3+kSD86SdlmYRjhbhkA1rwRH02DpDHv0QUC
pJA1yp7BTLY8aAR+IhTHNq1wRulYxvYsitiEFGl8htz0IoxyCeUZKAacfq3H5ObAn34KEaTTptoY
oVz4n2ehJKR/k8NjvBTYq7yDUPr8dv/aKRY7xcClsueADwCNqaxJnwvA1kZnyNO3PdOjBJHzNEZ2
2RkX7HKHQqu0RCAlONM/gugg5h5GLQs6712nobl0TlPPTdIB76j+Jfx97TuNA8lll1fKlqSIj56a
zghXRCc/sn2ldXl3rNVSw8YsNljQAS7tMaZftJ4vTp6qW4+v9jiWNhV1ADqqVBZcuMdK9o+aNYe+
WpjGM282ecglzps1mzOgD6WXH+Y1+KIN2MuHOQzFuwHSMmldAuqt3txyLakCfYXr3UQVRoYVueJl
AtqL95hpf3kByagq/Q9ODq4vPrVPJ+2wPsaMIAxhSq0BXJPI7LwJMAD7UzGxYtX1q2/sKvfWXkds
dtcIUa+vGyTeEE+xzc9ZYsoyfziUCHYfJcMZm9yIdHBO4+a3yi4lcw7rirjce/AFCVgM4Zku+w6P
zFjT7Anfer1elS5IdtWNaKIN1MiyTDqWOJy9E53HdKpS5vf2lXTmf6hCbD2dlG6ufn+FWizO8b1w
XRJCI1uDVpB8ofWkVIZH2NbirO2cFN+KSTiE8x+palFjMVJKL/hRSsVbzmuub097bY167BlxWgxK
mRAhmaAjrWwpE6qmvMBsjIY5T5YL76mKiPRWXWRcbsLues3g73J5GOPnbXPon+WkAnPCXgH9xneA
IKi4HvCqqx6K5R17p9sER0eVFmyX4l3F/B7AfvFI4QnuRD8nexJSJJAI6u98UwZzuB29KnmGT2fU
wBTUWM+d5eY64nhOV/udi2Pom/FDk+Wh0Nh3KYRAlFz2c7OIvfaInnJNHbTls1T4e7ZAaT0E6630
QKZ0cL/Ul6R+rxAXt9qoFyUb0b/baySy3HNt8bHq6AdiBkJetvWOUzfvs6GAoxuwcYIOnQtvC4mg
Ga82I0uaMcVtZKjVRGe9PZ7aZDXk/tnsMwdcCPB55s6TYYciAs7UERA/3bDrZh9ywk2ublpl+qmo
Uf3Fd+fANJahZTgu+rZqqzYmPykKI3xIcMqSlEhBSkTw4afhgtvLLoB4/ILhlXpkFs7MNjXvkI0f
gg2iCUhQO2FHs+gL/o13KVfcdnTrLza7MH44g9AGuErSgOZ16zpXFsKkxRnBdaCbTew3/6vPOQQE
lFQFvq0IL3xsJBCXq0//K+kAKXHrXpXIBn95gZgXfHx0pifi6aOnQhrNJaR2AkRhScR5E9aa2FhR
+29qHSLS5lA2nLgqLkfab9uiHwsSfFAM/FsvT4RuO2/li6gpvqCwM/zIwyH+N74O0ChD4osYwE+G
JBq/UJliGGZGiHYegc8bDDyGIduZTzm3rcA+0JYw7ksbOqIH20euf6YjIAhwTBVgh5WHw+TwZpg5
TmQJm7+h0QHuB8c2+a/l9E2zUw1tDhNJApzWJapREwaWAPGSu4RxRzL2LXg6QMiBSfMgg0qU2/Ky
kaJ2Phy8oVA0MBzEU+hNNPadvNYffS+i4HjKxvOO7ov5GppMZGxGq/MWHKCxn8hKI5WqalWFaZT6
N1yWgOUUcQT17Lvnk18q7miirK3RjyhIWg/ji5kW8uvdIx7A0dG5gSpdZsmdJ5Xflf0S3UEelcx+
k+Kl0ciaMroaEvu4sIz7ot2/KbLSDiWnq8V5vIBQbDAaLKrRZW+o0/3FxpMpyWj5Ao8kj5toYZlg
pMPEMv3l1G92BUrBMq3UALTaM898YYclR8XbmZ51e5aIH1ah9FHqvA2cuGd7UNktvVsbBW5MO/6C
On6XkYe3910cJLzfxIs7UY/qh81+fK54uMx70FkneIvkdfLOPpeU9g5tkmb86ceclQmyu9h82Pf0
1pyI9iNm/qiaotn/RpkHYlRPIyWywV3F2MF2n97q1TbvpYYglQQc/AVXikot9LdkTs5izb3WjHjv
JsBR+pyPOGYufrn9p9zzJ2JycmO0TMBfbD5CQFIv8+R2gX255nXRPsDEx90EOhvkqBbdpix9fQlx
CTIzVIzcWodOOEY/HmMhlBdheqrmVpv14BuMAVxWx6e+rDVYVScnixt5u43eH4nRZ/bCkbn0kxAm
HtlzUqh5odIit5+SVenVi0XsatMonUCMEJPd9ldnkBklUAmTEOp7EJf+O7fnfsRQUDsMFGnDl7CC
yxZg2XGEmuarwQm1UcnAfKjgEkuPDq6WPj0lt7Z2YZYEVoovvPdA5s/o43vb5N48Xdhw0Wd++sUG
UbMIZSd8ep8hR5K2X0z1wxKCN+8QBVXnAiRA8+i9JXuuUhx5A69gF+nx4QTFRbge8bJrzM88C4Wc
DFgFhhA2vx9vl1xpIQ0tZZ7SDmXJlu35sVGTipQ+PchUdlhbzhmyoO1TGqe6JTbiSUjP3eBDW3O3
7wr3j5p/1eRgcM3j0AbNf+2zlEPwZ58W+EOb6+qLkXLSohztYwkhZG4h6JiQinMfEi8AlpExRlLY
YQx3sEN8zpVtNm1IhDUyrna0VdO8Io9twSZamN2hOLvEpZyHjyXnZt7HGKRamVaXmLoXAYJD7zbq
BmXaftQE5dv2hhf/xgorKib7saMuoq7kTZr4fco07TKjEALtgUxpLhbao7Y3j3Pfu6INg2xrruEj
LgUZrizKejSC/3HHljhmBpVf4avQKXhIpS6RRDDmNp+EAm0EpHGqOGviB9+XKDNdFLsD/iEJYOnC
LFachMKO8tW5IrzRlAzR1WRJrivpM+mfx+GAx+iJTdCjFgs6vQU4fFF6ortScmwmp2766Lbhs5cD
0b7R4IpfcfzfLG94AMR9eIWVYstaGarTmNMzHefEsyhO0zDDh4zYQE6OcEPUL9ar+RWCaeWnSUMO
3lpx6FuFeYjzUT30Wp9OB44ZXkBMjg6Ro1gjYGiAZznnzr95rNK0/yicpD39VuHTxUf3n9LfXpSW
Mw/ndn7lsAFI9nWTmI38dZ/Pn90EKQcBVZmFKfs6OZdnZhCq2ZUfHTzeA2y+F2wPrBqqO+F0Z5WV
3a16V4RUMUm2N0fj7e3x79r9CGyW/Gpr53R5c2bWChgWIsLoGIsJ0VwCGHYyyFlo/Ii2hRj7kRWj
apLNyeyeQDvnmGQPRUONIFEEIPSaTO9MkCBlkgpyuvY1TDJUOSbLaZK4qUOVJHI2Lrux8nekmkJ0
o8GVDksSXpwa4ekvgQoRe4noHm+90x1jlSC3t5ArTwiqCn5g+YxlHKJeH2RhSYyJ0OnRVQ9N3Nn9
ZG0dKCnsmGmLOsUEj0BJUtg3CbkZgdl99EySOKIfk4MjdaPhTHKzouZJNC6dghmCyzv50+oxB6fu
aZsBtj0FKYT9f1jwb6ZPVhjf8hZMFLERW+zC031CJaV/jA1s0xClvWo+K8UtLcr67F0DH9Yk2dTS
bvxmC4O5DvIya8+YYmL82mmyCUM+B07tlW+Y+1HQjG5/MTu8W80+AFYH2gY4rTLZT4Zz4ea+oQSF
fa+MIMMmq+Su3QCvqqwX0Gr4KKD2tiu0Unjv7jBbWI3oN+E8ZDMlkLHyXjGkHusduZ85bwnBmGpD
o6MNLl5TeWtxIiSJowmw9mySBavTCLETJPJdugn/BpOQqhnivyvlznzNJymhI+S/LEQyJhAHFwRY
TKi4hXEWtvdzvmTPnTy491v3m7x5xUVZ4QJeh9VoTZZnkHu86bKcgdaFO7wTBGoGsk9+khRAIo6s
n8bKlpem/Mnt3JjSLguWoqUebvpPNWItrx+hLFxFEIOpDsMaQDUVg5Z01vWPffuIgIFQMFQf39NA
2pnqOAgzWVMXaZl9iLDYVVuyY4s20ZcXeXVKi6mvVnTfC9WAlDmlqeliT56689lA3Ax6qT3gOzQD
a9uIRiBRbhg9nL7njsmHlDe+C4zlkpuV0F2xlNUqIdnA3Ps8s+0R/9Uhv0URIEXynwfEP++EQUqG
gqbPgbYS1kqSLzBhRtKAqC2GX4tX/V/xaez8y4zl2j8238OQc9x+l5T8uAJWDFrJ78gmDSm4a08q
mtgDq3lu0ZPoxGgdmm70WP047PSMy07am1BTjz/D90LCcTFvqQAYiTupJxsQpEzWBoAsDAi7trOj
G+GK4r7CpXeL1b9DMsvn2jDpweytJJba94ZdvLjod00AlV9pZBFR7ScOtJZmMteBfaW3lMXP4ImW
6TcErLX+dJNfA9SkGcm+r6ng5Er9tvnp28HhliurQPhNjRmDHjw91XoQep2XC3OFgUARb7JXRi6c
ejCLIEipZgJ4UuH4MDEnHzMzlmnk9abSpBMek51SHiLC1Wb4mpwI6m+11FMdN/T/m7v72CkcDNmn
QpWu94NYCFeewpLMhP5oOGraT0Xz6Cv33ixBpkSf63ZbLJzfsC1fe0YYWFqa9PvEWIwWvXMOyYsT
CFsQwyTHgFX16hq1p8phAjT9xEWgisCeB6IJnXyBDw0toUgpS0j8RTHqzlIZIHBx1KlvrNwKa+LU
nE/eJRQifvQ5LI6/97EbWw26BG7kiORk0SDhcqBdcV7FTL5em7g4Aroi9kG3r2UyQIj9b/jPxf/R
IU0EYysaV+wBY5DCTIb5oCyAldoJt8nkHHyz656aLEaW8PWAreiZaqnqhEdzAue6S2d7KtR0ev70
IdquSIzAr0qx7fcPY2QLel3ijiAC0LbY0Fqc1Y2qOy0BXGBGjuiJFWJcfYNPjZfwWbJbXlTQbAwG
0zmKdJOLTymHttwFqi8t92LTDtx3G4DrF6nfd2p4MOyHM+4fbiqtDh6RdMczIslJ+GmxNb0HN+Ig
llH7ZSyTU62Ks2MAPXFJVmkMmxB2dO+BClQY/9xNhD5/yFfbMsWEres72cMvvIrPC7SxlTsk3yZp
qVDzOZ24VpG9+vi+TJyP16ufMiEYI17FSpyr4x6B5Y4k8lTya5UO429ea4lluN7q4eBywHrxjUW7
fggD8DwzIC6tlEwgGH8l/T4HKAOZgcEwpOM3RenogB7KZKuLb0oiGlaQcVf4GxjTliwHHiJl4rhF
gYD+miKGuUgX8s4YzrmlWNHfaX9pYmKzCuSbjEm6wh0boXWqWsCrh2EbyuNIiJotDEsvF3PBSPU0
2lWR3QCRDXMrR3Xi85FaZW+YLh5hliFc/p4MC29BOBCnWePS/EV4hPJlZHRl/in4g9j8nXGCXLMq
5yJF4fIwGq4C/dXUL4CP919ZM6XVnKo5WJf9Tv+4x/e4T9PKDW3MfF4SSkVoYyhU17oGJWcbXbct
dfsGJDGNdldgmhQwheoX7IiCOD2XPxPZaPo7HE9GJrWHHmuVTBE9DNVowrARfvLYLpaAqnwoG1Xo
TxAafeQhqn0H+1K/bu3ht/WTE9fGNAlHPs5pG/raXTAvRGXqs+j/QCDuzzmPKmjRrMZY8LL3ikkP
16eav4OnsQb5/sxvaqxrSkAhZUdR86ewWVkEyIBW9eNIniOSM46UFaAJWtTSgvDBTmFp2GtHmNe1
eFc9V2wf5/19uUuqIhqg0MQzdhLlqmCCTZE4okd/xYMydFdHG4ZD5khAN7Dsg9Vkf7G+8B7jZ1rB
mrifaJ8Ysoq8DtVOwz59snkAhdhMAnp5idkesMwe/RqmTFTuRcNBVYPV0XWX1McJl4ajs+ZxPz+4
LhibI1bfahtW7iqxfteQIvsQkwdjSRcYmnOkgj+fWyUezR9XZL7WA3n7qJIYv9CVX86bT6NRKzkl
XTK2Cek/7rqdiPrVx0QLYFKhb/3SfP6l/e6X5v06a9LY9yXDMqSii7kXNojwvnTJwyDbOkEpY5ux
dhlYQ8xUJG9vobMfKFpjV9yDQaQS9IkdK0Hm8eMuCVUgNYc1XfCKr2ufHE8fJOvliXFUhy1INWjZ
rrlROz6eW/nz2wq4X/ZSliRp9VDR/uFvUNzmHldh0RKuUJGd8234F+tdIUUSK6h8RMlKyefXYjR6
fAIzeodKIQ2uAB0swHpjyPpUNrniZnwWmb6SSzHjJXcTor0grhf5gja+1f/RcdqbF2G7Tbg9/Jw6
Zt4YuMN7h2aFjFk/1CHuo5nFdMGZqqc23GH+434qCU3Og3ukdaOOJ6SYfLBZFVtirJvWawmrnqkC
wIVdQNHYRCW3t+ZF8GR2nBwm82ycdloFzi7NrVEtBt0w2hriQOE2zi6XAWLWv5o5DeUKRZHbyf0i
f2Uyir/49aYvfV12Er48jX0ih6vaoRmKbLYjwOFUpQ/OFIYX33BWFGzxRGqG23V1ei5R2DCif6QC
4MBPMYnCvAnFuGxhEENfCRF4hNZTunhOYiE7s55/t9f0FWXHzRyH5g3byc6AynaztOkwzRwiDzFJ
UW8SnVe4pmkPnpLUp4QORv+FnvsO1k2cOOXwWws5MiadYzvkvaQwVgtdz6nDjNoaob9/Y7t/gR76
dqKHnO4xRn+MtNsugqbLgcLXN6BFdqBAgY0VbodwUf5QbV3pod3DGI+0ufK/yK6AoiXT37bnFDCt
XRe/4JkBtGpfUwTJGOoc+UASKi0VYguCfvjRadOP97vFEwDtSzshxLJCOBBfFXjb6E4CbVFKHaPi
waI991yPWjG8w1NseI6tVsRYDKE7L09vTjUWTvO81ihfPLwOdPkeOEoZHgNE8mwh90RdWff/qMtD
15kVqSjJZGHObu0EcthylEakFuLwtgcxvg6VVJKJT/Dl6KslJuh3Y2jIFlorHskTEtLjqqrdVfED
8lC19J6XjNyjEXMl+bKffR4KNIqQueANhCsItlLYd2yMtJtOcvwcieGwvds8kc6MPqJrbYZ4SqUI
vj+OV0/fDHdBqkGX7dcjGYqD+6jpmmoxBVSZoQJUBzgb6c6IxQ9AdXOJHaV2EUE2ceqrLiVYGhyz
cKvpZKFVx7m2xJYVvZCGqu2jX5CqU65KKd2CUoRS+ChcHyXlhMBBQ4mHETsqCX+cJHPwUbX6T7Xr
JID+/9sV8jYpsvey1RTWwI7JZ6/NzNgSigpzAKtqQQ/PjtDV/gRVt6G8U6fLRNigNYE7dCtaF2sf
yfDNgSBXwG126DVwfBr+vhJQMEOsMbejyFZmJSD0h0X+H14haE46ei5E/vWu1Krd6i0yp6pRKY9u
uwWxfa4rBbdamxHgLOzH9bp+dGccy1yVxzPLeOpm+Q3yq19kd/eVJu2+ZhQRk4jeNmCEOFdDUX/o
xZDtHrQudWtag+zHnehPdlGMlVJjNu8VdmiHN32HWvlGs2IfuzU3CBKpqy1buwIY1Yk1FUB3yxbi
RNQDjsgDEBTLsMYy4GQ+yu4PrvSJ9BzBIDRBxI0DwSIZAKhWaUtDLnbaFZTJDT5ImvbdiQACkql5
+B8BP/+FY71BrJLtYxaq7kCYAv6t3dWB1CewpElN/HwP0ikoeIpkePGI70rK6Y+T1XqNjy9mVFEh
0f2RF/8Aqifm/JipqiVT6Bb4U7kTcCJByISjNbkzNeVUaA39t3PtTbGtLwJ9S9NXQTPTqdurWzz2
7I8L1z8hzn+M0YFtl8yBeDkACNRkZp7z497z48AcrmSjE4LKwVVLXgboNZ/sngz7kG++i4z13Ue/
s7G+UgsPpEX9oTJV00SOw49Qi7a/6EzVvL2leHyBuqFTWgEOrRZJ1AOS8I1HSPF1CBbI0emteDdr
20dKSnEUiiyXz4LO/PAQqBPrZmhuVb1OUH4p+xVBeGkADlExFyou4NXgOxoYLXnwUqEBvShp5ife
Z8QwbQIwp3Yh0pyx5BsyeBhfoNjTloIRXVSVWmmUiVi1VHbJ3cfYVnlGahtuGVfnZ8ad3NvO7kiC
6KTvK9gKKwBrgpMD41pcegt0KuCWPRdAJVPh5SPaRGPCnV/xe41UHC4Vqzofu+5uZk1LrkwZIM24
S4C7HDoPg/NUGng1/2M2IrKRJuceovWUA4psOE5biaqcFLxActRE9RrZFHzoiQlKDRwqfv2/4Bw0
DCAA+PGm4POEYRB6glekjUx0Z0gIrTfoi2urlR7t63IjRq7kpXJKy+ww3j0m33fpz6JNIugK55b7
reKWDSBfTW9Lsdnq+4xpowgNiJZEATLkxd8vOpMbo3PdQbzh+QW/GH2tkFq2283g7UiDS42JvxQ+
7b2yzeaYNmU1xrP6kf+TYTnkX0F1jcAXvBLmrANspdSsrdDwQy/cfGqi6nEO/nBjnOSg+07x6kPi
OEpqUrzTBvvEHlMoWwbRWgAcx3p/mX7I92HvQPLcyU/fDRFwGBOebgY1ZZ2TzZAJdEiIcDpfeoq4
RpwGoPWke5I9x2JDFNlBeSjP9ErXJtS+C9udk7evlkAZyN9hVE41B2GOLk02I+oBuU9AM7rPluQE
wlBS4oJB/Lt1M3mkHfrB+jZnBH23gR/xS2iXl6U2Ywq1I8D6OphCgM/lvMtVxUcSB/lBxK9baqTB
SSzC5PYpdYjBbcqZS6LuHNxRwkjoZKb2N57dfpv3f/4NblYM8/K/xold0pSAB/IJNIDLlaHOGY90
EYA7X3FYCo53Q5zXB0lwnsZ4WH/1rzSnLWCQjd77ml1K04ftTMsd3iKDsdSxvUuUwxScAwDY/4DD
KgYX8jRobAgoGPhqSSvsROQYIZyzI6v7sm6ae8VehHLxYWKe5lLORZ7bp8MmibwYtEBc7NBbGtS5
3rDx4MR0UT98MwBowQ060u0CeEURYZCMmnnWy7QDrBgHSt7/QnAJ96rxeftAwH0guJbAsS1aAKqE
m0f/a+qkDGhYy3sfbge4VVr2xfuB66l0o1UbNQmI8J+fxOWZP529B2aJ+P/onF1aoMl4RkQgsJvR
skJY7KiitcZmtap2SXn8+DcvecfAN2D5eILbPSfxNm754SeyDjFIpY3C+D+4NFzdE0V6saA1w9VL
HDEm8aefJvcdS8bokJZHRywNw+MvBzv67DDmPxWKkHNk6OUlb5Zmc6u3V/qlsyMabWRvhrCHIQWG
7H8DYu2gLPe3b3tO49rBzb4NMJO7SvKC4WrqWF78D0k9mKwwIyq8JZnbte5Jf1btUP/his7MSoPx
Wkoq4xH3NCL3K9e14ImMUUUBjNmkb848rV4FfAfFUAr0DMyNUv5C0dVz2cqIhvtyKWBYOUpm6jN6
LDVbxQDOOvjgJjhKzPURa3DrWUSYHcSkBEh8YhHifBQwIZE90gKoGt8LOeFdUE+AS1gCsoc0RQLf
S/BF7cefrczeKMqB7ABOxWfT7Pss1pjjkiAeQdKQ1jUpIAxBvsMElXlsf9iGC7oebuQ3M4CJfTS3
jU9ElEhZa8136/WmxtMQRuTMyhcBJBUM9GZ5AKEG+y6gZ4WS5AMxrGLs9npMfYHmk+URR23A77EN
tFAT6F2FenTSKePpiUoz5bEsTTevq5uSocrwTCTXOYxLulsaO2/mirX4jp2+1IIWDD/9gsjhl4cG
6bgNvnZ88tNqG0S4BkIYeMql6RJwLCaJOYTnZF/mDgDejP5fqqWMj9pu6oskUtwpjLRWhKA8MXrD
rLhrzr1MsHKH70ijjDGlMk6I5XWwSoc9SD4iUO3NITFAePi20hZClOEYVo9swuzsXEsS1oiq7hft
y9CG5EXyzVC94Ehl+t1BXSKyGaF+qB9tc/jFSzQyhsl8VygbIMH42JiSn6NzH7xPirHD+gssilng
aidmiBX/nky/5nakswmDkI1zGSUqIaARV8PfgXBkS5NgQhv/24EcG7pJ1GxGVVhTKjTylKVzb8Zv
VqUuHUtMK7deSGH+QlaMBknNyjBJ3DgNurfpZ3H9vV0tvhdfk77fLl3gh+Gk0vrZVh8eRfofg2bG
1mcwWdap/UUaElJYGBQ+lPkGFRqMhe7Pm9Bi/WMgr8Alx4DzqqywDYm9T1ohSkLMbhpibhrA2ggW
ZGPGuFCt+esOdJgIZa1UMFSdFtUk1r82v2isAvodlWO4na1RXC/xsr/QjtAFuyo3LzutMnsw2cqS
vJ32GA97LW9Ly2MtVt0ANvTEsJNmms3mmoz/mqTP2/+qy1m0CTlzKaQfeibFgnMGg1uKlqJP1cgN
IfKt2O9qIrSz8+UXm1HPWV7SHkppANWc7e9VYlVSKvdEQINZUgKRFA2JOqSTy3N70Q+jYWTQuCXf
uW3L+F2s5JniRD5e4lmJAnZH/7QRpLKzBhpDs0UOZiRARCbjvHDkOO+PixTTO9m3NMwYQA+iYYPX
+yGSHBez91di1y3ks5b6SKa8DTe/yCSTKcdveY4oUgpCXYJuVv2S4BvTystv1M4xGrjD0tjwDJt/
wBpvZL+QdjFN8IT3O38ZQxkCSF2fjTYjKe4KZxMH2Xh2u5BYEUkQw6X10raXa9FjsgIz6Qk0oS+d
b3uSqaKdBTQerLnRU8eybGUsCkpG2wjZkcQTzlbcwnDBs4IZyxOEKfKtgCYQL36g6uQ1QmJohPDq
H/jkH2tOZyAemsnNtZp38+QEOUcmdpe6uJjnH9M6r5k5ZgFQlfuwWKBtMdwWW6qGNoiA0CkzABr3
J2UOGvG5yrNcENMV5UGzjh6A6Tdq8hgypvgQyBJxhWObBr3D2ojIx6UCgQbf1oJ6ygfNG6iFm6D6
LH61cOsDMFq+ps/Gvgje7Tg1X87c8JUcSRps7fpgqI2iDLn5L0rKGe+ZdPo1k76wsxB0+3z5uIQW
f8eVkTs8MOqCddOGAW8aISyEcg0U5Lzm490YwP7yICYaGUCpBCctoDrAGEI4gJALrX8/A2HS/eOo
eR/kfzlvd5hX34S5ljK3bi4U3mXD/AV0+IycdJgyfYcN9k19+UjdRRlwkX+U7C23hkSOaTNQDBen
W6UoRfHh2FqykDAtlVA1c1bEPj/7xNiNYNpLuGP0Zycdc1KKfB0+PYXXPDaVtGahb/Mt0UH7gtH2
GIy7pp8lhwu43bLWgbukEv4UsMOMLODnhQpaTjZBwc5k1hBshgz7DYspPTIJSGvB3zzTI5KXJ2wH
c6tGYG11aW6zFKJc3nGEk2RhTVio2kWvtCzoHVoeuFeMwOzffIAK01TGokwCF4uTXoALGSSgkDYp
iXUSTa3uucssjAeSsJL3n7lIeJdB/s8HwxXYiZTUMi20/zFxcaby67O0lIyJf8TN09qqPBTOelY3
Kjtxk5aOZ3uhxRlkqDUwJBLuEfoyDHCiTCT87N4HBMsFSXp4+LqJ/BrhQuUcWLqURXUSOTKPe29S
MTSmp6CdEbzK8UkpzpXQJV+iFJtlsPebCRc4W0vbnJCnNXXYLzto8Sukj2qpkdQDu/awZjJEv6F0
pA0kqnslb8zsMFYiBxaLMx+b4C3n1wAezvD9tSJOGa0ZnO6JeTffrDewBl3LbnILW2k+zPhTtnDn
qCJ26I1ofZhod9GcWkLpdSwKOn6ZkheLPyqTGL39Z6GmimQLt+TPjaklCzsQiebt0SEZTYqUFvpS
5Zp1eY4acwBZABQRR9de2UUoRujaJXDV6bDc8faKBBPwUeSI1kzQAhatN4jLlgQqzfL4RjjACEoE
4X7ru3nMnax8lTsvkmrA4bu9UIs6jbmRiXEgQtKiA4IT8memRNASOPWnZe0gjlNWFfFg9OUrZ7e+
drgSxBwRB4HWslYIm0fe99WuI2pixak+t/Fwirrvkelum//BgLQSleGOmOXXWjYbJaDyEwHZi0kH
iXqPP+TKvXgcJGropoUAn6z6ADheMFsh6dMeUbKy9IfELXvPcpfAWUk2ISc84y170M8zrfJiJ3xz
IX6LGNkC0WUAuc2Sq9EJM5+SQO6Mp+oT2jBHwjhJyERBr5stVXa+aXXZf4JCqwx0JLkzmjDxKwkY
Fodh7TLGBjP3WLrNvR6tQXnuhGH7OWSoB+/ujTEKhycuiDoNCIvGFOxhP0a1cgKDgsJ648MqX815
IrfnOqgljo2M2hIjfCQ51eN6UBpnfgEToZmQSYyLkk1MIj2OeahGK6rYgNXU4h4Sygm0cg4XwguZ
6lfVqTOu1BkYGJxAfnJrHbsnWq9BHbqVMdxTTNQo2x363aAsgHeshpwy/3EP6OJmXkeSKl85p1vL
WRCY7+ihspppEIXnA8tehslwelwetM4bX2EkVKTvQVQWgpDpQSYvXnBd/n2H/7EJqFAM/gtYgyKw
qkFnmPdkwKTooFULwAFr7EZF/zirNzfyCIpOQzgfN5G2/igqCOgiS40nnPulR23DHVLefNTuHg3e
UTPoG9DV98M01SdYEOm+0fAvA1mCOYz/e8Cphhm1zKxxiQWn6N6uQZpqE2+tRK8Usrc/LWCyXtlW
1d/UggMIg3xiCt3eIIxNG2E8XBxTB/7RDIy9CFFmPr+QwCeEGEmZMHz+UydrtnVpoBWMSrdFz92J
1XHoPWp2lAqFvXQBp0dySF6aZIoNtzDfzhO++zoM4eT0HCnV0LKHNF0tfzPm0ELd0kq7dgtWicF3
UvzStkgmvQN0Oz9hHLC8gnLZtVCfwLKPyLXQLfBHwvIqzgTWz8VfOyHQaL4ZX+SK6swtcIkakHRQ
q/rbqlRavRxmytJlO4Gae8X6MCLSDlirkQzjq2AS5ABWIoPomP5erWRFEzAKdh8Z0LNeoWzVDCh/
LlMpAESsY+7eVOYxsK9C0gpb9pN2zbZJRaF4RLrQd1CLthfBb5WClV7QGe9cnkCkyR/QslxZa8xW
oBdQIrXqfFjBLAQY6QPxiB2EK5ShuBfDHqoISDglJzRSB5VZNyBIR3y2XOEJ0THlkon8Otz58fMy
up6DrvVNx4hetEFXF6d3QMYYg6kxD7s7J4cd0bxICnekxMZVNe9tf6qbbWuoYv6u6DHlY8DPoMiW
e4sYYFoRRdlyHjnWZB/lIE1vA7SSBkxI1odd8kEEJj849wJU4ZxFRnwrmz/T8st/fkfly4M1wAy5
eUPORb1nPcdX+xbAnPPIsZZgV4JsAeDAmk6812NtQ/6c2F5ZgC0o7mQ2+Tzogx7FWJwgKDuA9GLC
v223sgqAsAt7nZXfaEESlY190bV1W/vXZYa4mMTuSMv6IrMRINSOKVTg4zogTIq6Jq34k4AE7QlZ
hdhxhOE4wU7LhchOcWlYwWkNtaACcz9Mi9GjQnloJmPiKW4AAtCc2ur4xCUUE0yo0BSh+pruY3nx
XGfvWolss6+0jMQci66AzbwZB0wEC3hy1N1SUcl4oMC4D+PCO40qDIk76HNSgPzhydW7LH1oUksD
O2P+hbiv4UoO/WeE8XlOYEdj3XL54hy5vtYuNKqzDM3FIaiGQC4IS6xZcJZmGMS77OTCAusXTID3
J8GQmwA2av+9LsmUOaiCM7pmdbaw2m7um4H9aBYL+SDtQManaR/lbrpzr+5g1tIboZjEppV80bbe
lk9hcrxuUYjaop5LP8sScn/6vVMSTafyvE2R3uGm4SeLV9/q/bNqXsHkpfygj2EDz967kdPCRkNQ
zv6x/bv53i0aklZV3GdwgxXWlyH+a0/8fYEQgzjLMo/gVCpY5WwvdDfZp9CushVYjBp/20jx1Gy9
jR5elgZ9hZvZ3gkRT6Yhm6cD50bJhCc2/aUpOCjmDhGTmKU1E9Jp/Y6vX2HpV9hLJzqAdK/f3bX4
/rIySk7BtXsIuY/S237L1gJdfiDWmoaLcVho/ZqlRb88DOiEPAfkwztxTEsZv+OLDlBDvbb6e4g3
6w1GHlyT1zQgbAso+pwTwuPe8+o30eLly9ZBU4zp3PLkR94GfCzl/dDx7RZBffkfIA97mer3fJFI
Swy13Rs2/jY5Oa99nHBAR9IMKWxmA2n+IFdgUs8D9hZ+eS6JOSvx8CgY0fR5bIgGKt9YF/iWqXQ+
RhX2kKVcKmqRozVIsfQaVbvo2gzFE7ufvC8lJenqe6ElbVplHabZEUXmEXzLuwI9At/pzgE8OS0Y
oYK3vBSZEj1jEK8g6dt1vvJRSEDnN1jr2bWiAW2oTYSNAk3qqY7N+3D05Bphep7pY1/DPWBZkfbR
HgB1thkQhnl2+kA8tbUM/IpwLbG6kUq2CYqEtoFiau3nMVN6RnWFypkUL3EXhKAV3qMqh6ThTsFP
CCNm6TyjarYrESwQjJPEV2Cy5bLWHGsJHv2wK1CooviQyL2ss0X74kD0kS/0N9cmSskbV1ZKrLka
MvdxIEVAp73YNL+OCFkxB2EI0+VwVJX7E/xdJHtBkTFZGLwLzUjHNLqpBz16ebQaGfKOsRR3mA/f
6kAD3ao9BwUyCA+X69BfkZFgV7QN/T4b5fUGicFPTXxRNKUpfxOvVgDh8hJZrWuYWtze1tm+x6+5
aXa6RcQDYRtqU5btoGiaG2+UqEpAKGj2nSw5GjiFZ1A6scZydsvDlSdVqKQbbXT+T4FvQEbi0U19
9xjHF0l9jdIEXG8/mjSwKb2H/VkbCs/yef8Vv3iXyJquKJrnNB0ctRBPz3e75E7UnUhjrvSFoN+r
Zc2VD2+Ew4QrvgEb6bLCecfwd9PryS+IXjb/wpAAw2XmwDe6ZbuRHSvXHGKhBep4R2zERMs2Nm7m
67QWrV7VBlzmDrpgtNIqfj/GClPdYSbF+K2HaUcF0xQ/srqXttZ+cl4AqpuFw/LAGaCOcKC9HoLY
YS1mifp5VYNxJgZOfFZBZzkdnm5ErrWO2JPHv2j6MuIZxxcu7qVX4r4UCkIDtf8me6/LLM9Tbadd
sSZxtOymDIq0eRr9L9V/tdPU2zz5aIAFKkVMf8SSsVzq9IzVs9PbT51ZNa09jbDOgzjrLJIl5eO6
lweupHM06g5MqD6AOnB2ROwEMaSGO03yw5HSyqQwR1/rgSPoekBrW0rUBy61xtCyahGnNmxRvSy+
fH0L/r43hwKVG9BS25aMdr45Cu4+n5THv/FT3v4ccXQWBzi+R3BaWS+b4A1iJRox+rIc9/OToLne
VbuO005HOc7r90IS62A8VO90tFeMiufUlVvunva3nhB4xKzC4JRwGcSPhyHMcc+7sGzF5PdI+S+t
w0I2GGiGF4U/QsmYK1gzkgZT1hvZOuYXsZojzHSuduhAaOztpjWYSD7o+nIrzPKCBa9WTkO6k6yo
FendotnhXHHXexHfIuphUOQk4kX3cWeFSD0lXBGzGwbLq93+cAHCu5nsTSbgqzY3iwv0l+LfdAUp
prezeHNvrKxo3ySeSgUGGxBz2LM3p9JCxwnkq9h4XwtR3+RtQAA54PRVTcYKmjtihu/tSc28QxLO
clBV4GHyOW0rrSShKIMxCIMdazrD+jgE21szf1mA0i68cPmJjMHHPW1EAVCQ4HQvPfoPMxpOfD7j
tPN7ctjR5UpiuC2zYYPiwjZ8dKRMXbFio7ESXyHQ3FPBnv4GDxKTspOGxiIpUFb/TvFT2+aruL7M
58Syu54cHoFGLgDtg+okZMecpby7gcDDG14tagzJpd1ffPqKR0+FeHEEFjv1LLspTlzXCst9RMew
C8AQljNcRjIOq3tGWYTl8kYiwbRos8HgGHukAmhK7deE8/TF8OeWsr7G1S0zu29rJlWCxOAMb6Of
JRVKOHOaFhVsrAoP8mCUiOkLD24EssRGVcUqMKswhoUqofRTCbJSNwRZNztmIC5IYWAqJc1l99lS
y12STcWhgEj1131x/nfCFBe+kdmrEPbq36SFbLRfKKu5TYMV4nnYYC3XKHmhzWZiHfsmNvs2i2uj
dPPncwbmUQDsO+HhisRV/nAE+xWpFZbIelNab7psG12M0DBqMEAfw9lKv1vjc/Rw7fXQpGaSU9U+
0SUaWXCdOsIQ0ndI+qo5zbyVQxs8EXVvgJWGxEKEY5w1ZPjhu/qq9379pSuIgGmrRTZXm2LuXCCS
eVf53rV2QKcS1rNzNlFhLTJxKr4mn68bodhIuO6kytos2DWtZDoXm09SqdgeQpXa1oJDPDMUf9DF
y1PVHnCPZiznOa7+jptoXhvbgtBw2My5dTHejHCnloty0unCu9k6pw+vJtbx2gupn0yRMA/Rle65
G1MB8524VyMrZgy6aaRPc+8pqA7qCbJJLsH89E0Ynqn9sRLCI3JcqcRSAzdn1c4tpf1+D6A7tbY4
sgHHY7fUE7mUi6XIurbCaaYkxKezX4kasho/NfwifrKT0MRW/j3CTHa2F8CsClDWbPU12AlgPUC+
OXtfUAGrfM5zF/FVVQ21ETfieoJ/ZoLn7VHCngGzoUhZGHH6fc4qhpSl8xrRdnqQ1RtNbwq8dF9L
szhLb4XxIouiykYPvxUzNldoUDqw6lrDHVQgr7XtzIdLZE9rfYsH4VGTZsZmK8Vaw9yhlfQ5NdbS
4dq74dsNihcV9aq1HV7cFmJaucLnj+7rvyGF6YzYUUQBELWdq+agAmc3diq/nxx4ni4EXnk8TLxw
Ptlz5aLyFtgsHmjVtjPoQL8l4zA2wD/GGiww3fUWxHCP/fUK521fJKxrdPtDrXddyDeKtOKEUbMj
OgB0A6loQT8qaRCbeKPYQG33MVGTiLn9RNQymYZRh6o7RfL/qSNgJHDiZPLb8c8ABxMSfDnzBXlv
q8fM/MYB/QXvGcZ+X6uM3w1Jy8e9kO0FXB5K3vU4TyEqYpK831EpGhqoGw99cXBBYLMBfmGiOLin
OCS6HuaBXeunFfZJD1QzWNRJg5EyY/OCH2KKaFwuQWV6+8NRJaNHjU73QFro08k21Uuo5PoySrPk
sxxxIXeZNKj4e2YvqtpQlZohKT9X6CXiluJlxtiOg/stLvGYeyV1uDzBroVr6uclHQ+koawTCvYH
+GwDPFDo4+2If1S8wCpFppLMw3CKYveH/Foo1ngubHoI8wxbjKy8yX3V5rOuIp58eV7pd1Dhm8Eo
dtJfkuiy4SsLjt7uM9viHNhVUagB0zaLpAe3Gez6xBaG6/sH5535qzM1VtYP0UiuRg72IvTTfjXL
lHLk6S0/pXyAeNH1vnjD+gEEYGREOde9Gd2AYVEhGcz7TA7WOd1P+inP6hTt7KmJLYYBcjgwMPbn
5EJZSP/Z4FhrkovYz1/RH33nm29+ju6fnJ+kxx9+6W8QKehmA57NeDg627RVAOXBReOYagPbHGyQ
SpgRELq4TnKQVVUfMq48A6kM43gZLFSa2Hq+rA9VjlZhW15Kzi4/nnav6CVcIkz5XM3kE2x5WSdR
wHrKk0Oyt4ZJmRpKd7pxsNhKj14rA41anRy9juoF6v8P/TVEdFTat6NSoQFPW0jPJA9SS0GLMz/+
r9/lHmsh/Av41XDNckKlMhQTTv0lVB1k/M4b70dh2ViiISYcISb5b3heRJQ4rvH8822wWwDsBYgR
GZ38wrEyEAAXC7Etx4KM0rev4gIdTD0sXfQnRZjfC2PhNxBh2c1w0gFZp2ZiUTawfPuneu3EsmE+
xqlmjhmwDQlMvXsUAKax+fOFtaj4/JLklQRqGGlitfKqm7br76wUptZ+k2vqzOhElCY40vctgW6z
NHnr2DIWA6H8F0m3pOANZCDfoOnrVH0C2nQuVZO49+abAPwc6cNDp/b+8zIwfZY4ShG7O7kawz+O
abSMrT+Bv8QUKfWeslf1aTlO7fxQCfx67b24iVdNjDf1ldQFTIFaAvYGd5QFkIEraEcP6C5XurfA
1tK3+kZVystOpVWa11QL8sRackkC++/bu7GoaJnxFbheQpGunD/LZ2FtlHHgKuB1TU49cG4Ap9YB
mP0nL6Fisxg+e7iS1a7lqCGw3niB7g3X4DrIO04iyVkG25MVBhtgsiyqy+q7vzPs5zuwP6VdoYdJ
jSCiInsCbIvUIvA6lMWmLdnXwsj3BF/jWNA/d+2d5k4auqQMARQ3flIjQych+lQ1+kT8Jrsr/hfB
70C7G1zgQvgjRnrk/1UltrWsWhabjPi4e66nb/5662wfwgdPArETBUTJIR5zyBSzlPhKLbZlnaFd
xoSrzrzr0/OhEH9SgCTyO5XlV0/YqbFuS4TG5KwMUbxJSE+qBKSf1jjBGGbBTQHvgVzbL8DglyiQ
9pzQNj8G7KyILg6mkc+FCm2vo6TwhBhVA59wziXBXrhuZxGZigHpeus4fcwL2wQYcy3pc2PNVqpX
5HSxPb/DbiFBuC2nJA855Sb1ZozT+EYAm/FObHy2FQG4X5WdeX5ZSRjcF9xu9/zrGI8OVV5dZ1HU
HSpUDBJ6wZ6hJD6p1VyQ/WlAxi+uPNsucw29kQrxp4vsvBAaiq7pYjdP709qBU5E3KbaukjvCs+P
7UJRdzKRRnTOvO9ZMVkKHdSGEqw55F2uygUFU8lFBxclj6pNouRbMTvEiFb3gqKsmrlsVjDEtyUX
ORbNZdGk6Tb7Yfj3wGPi83kkGaQC9u/GTb0dGgCX8k5GXRy8tPBbIOfjTdJMKDYAi5V64vLJE+dq
/uZOYBZxxHXpcGoCiGJjUxUQNhDfwYoz789C91LP28vRvAoxqtkMEoIIWmqI7CA44b9Q2dY4vApE
ELFwTdj3UuGGjlUTCYPWPJHbvtwbNXF05w90psHdeu4w8QPKfBhDg3Jz+RDEtzet5JC15zFdUxs6
efdeyx+WGBTV1bGDVvlPPEOI7kxjOmk1DDv9JLMh0W7rtolJ1ShENu8xIl0ug8p34S4LEJPT0lXM
54suyt+kqVEt5XjiZNTPgNtjKJBdLQWWpEstCI+VuFbqMZQVQnvDr2e6QQJm1/WJbwC06uDoiR78
dFU6M+EINZmBv9i0bYAPWxzztYSo55L6ZsEDqz6iseb+7TJBX+jpN9GXGIY1k2WgaBZismhOL2GM
l8xvU2qudninbI7WCUSWB4NduRF8grHVgfciJc4sQJUoquvPjhTUyqFQbpDunxcsXWYKPai8zBd8
Lv2DyJEfl1uv/ABEAq8skel1d75lej8Y/61Lmhjw7yv+2C1BVRZr3wJXHCVY8x558de8CISLHHop
9lxJ5/j/oH9cGonYSMkp0PkRQJDu0xjdDcLL+kc8BkQGLas2Y73DIuc+2teulVnLqnZMfLdulPf4
+des9wZTStBsEy4zacGUDkSSfL8KCQQ0jU6Vm17zBi4R4ZjizM3cMD8axbzrzAmdgG1GSHQ1KTA4
1jpgNKsjqrrWy8bSgWL1vYjhTcDsh138BH6e840MJhumk43syE+qOXsPfjNeJafubbxgyB3F1TQ1
yiyzDg1ucPoDXuxI0Q/Ril/3cTAw0K0/oCEEd0nxgT+ytXGG8tnwh74w3MiCrn7CZp94Cn+uve4k
A1uJ4e6pjQSfnvdDW8B48MjpWDsrhYCYmcR1Um26bsr6WEkj28yDYbtiHAQgpvjLIsXZsuall5w5
R0S9/ZSTgwZU0jyd3d4c0jF7b7Jb78rML5JL11cQX0Jd8Y5bMQ1yI1HaKZWscO+Ljef5iqQyoGmw
p5ZaITAcPEGHwq/Uj0ydKEDun3hG690jSvl4jJomzBN9YHa0lo3+htA0NIujktZKvKzwFXTFlzlN
TIElJTguKBX2vUo9osmfmAXzTXSjFdpjJ41YqStl60DSpqEXQ6cPbcrqxIi8I6Iq4TzA66mLTFBw
64Or8Iu49QM2ftQwGMQopETTgc+YmCTuaDqJE3fRR1FXRMthUFadrVbeXek8vxffMT+edmG35CJZ
gJp6HBL7bdWcFvtTZGL4x23j4KcXUcpR4phcHdC44d+QanomFTplsPNT36Yw5ExvLtWTA/4AT1Q2
LGLxUwzoymytMPlKpttAU1oUn6zAJ2BrCTMJsReXwauU0uBrK2NY9uG5flJcoPjpuxgDYMdJzvv/
GDle3l/4eRQU8lh48F3eJYUlkTUk0pxthB2g6m2Y6hIkPGG8bfxp9smENo3xbRg5c2zJocGMFaiE
mgcmpPBAJAOPMjuV3MDIi8UHXo24D1bDjmIEQEHbEW8NzRpxDrN5EbQknACgjuetwIqtHi/L3p25
04c2tcGNp76IapVas52F5lwimREhSXzUO7IdBIv/tp+Xfl/pIfUZelkW9UpX3DHADcd+Y2jxp68G
1BaTF8jJ3z+iZEnejMGtcqX1UGpVkxEFgt8WObLzB9hQGvx694gOz93HdR9IAKpXfbdBSGqryYrN
66g02m7s9gdwJmGgeWiID5IlSpf6zNbbsjeIHC40wq0HQ1hzdCjJ7aQzqJ27nsCF/CopOpN5pqm0
t9bWoe/sthPzC/6uuZBz9VRE5s8PwCl/LhMBAnOzjCK2DT3Pv+0pOF6KCyLC2h2ESOv5NvR3xLEo
Xl/3S/XdNSFuEWqY6BMHodTd0RKF5yrv5kBlMmv7GY554Xwv7W4rPHlemTjzsP+iHppqZURZsru3
y45vkggmK+iZ8ZX6Si+0ESpqhmnFayEHXNYv2Y+a94X98fJ6bQCfRfnhjaFY9H1gzfTx/OARLWbm
0HqMainKgLqOw2Qttggkkpi+hlGGpvk2RWGK2BEuJOvXdf7kuEzWE/WvLjatnLES/95i48z918M6
uUQ2+eDjvcGptYP0hbVwckUjvhsXNDf1fkUVz5YUNVHRqwzxrB8Gz8lfDopkSGlg0w/icTpxYbxX
Z+Em3EdKIynliaQceLz8p01mhtWzso3wbK8L/dJPwXg+9OklYM0USzdCnaB5tZQospvD+YjlXlFA
fGgJxU8WtDd/qD9HekEttq/dIPzOeJd4mzOVFZmXBXXKg0shihMczvmbe8YDwz6z9bIRIPIlXklv
NVNkWeHrCOZLS2zQMJNDosxLnnWh7KwDLY3YmAgkVprYLWmjRhGDjQ1gWAIaVvQI/3T5jzcPWA++
7Bjry4p+cA6n7iClgAHtpFotjX3glM6SVtN06X1yMoJKlFTXb2VfvWE/O8L5eoeUN26B6B0IAa3f
zfiuxLD4Lr+Shk5vZ0W98uZ7y+oTXcaL3HRj1AQZKM8oAnmc0o2WOWuBz1VPR1VnG1M7N46GWDm/
DWPQ2hXtT1vMcIEHs9ANtG2It2cODC3CoItdxAsmnCQaGW4uEtmus5PSwb2T/OVJ8ObO/L0vcqMt
bhd4bFME7i8xdpnQHCRdoQjmHgDqm2Q8biTk1v2k0sNYA9UClzfirYsCrBUpHMLsKzjMsy8vzjDH
RVXAVuWnpljkalSKm2zhJ2oIGDJIXdqnIUdgKIi6PK2/LAXeFtcuZO1U5npQD40tiFTV3G1Egm17
q5bB4wz0PkgYShUb0ZWZAaEH8ADkrSUc1D9LqEXcPxlWyDu0kWZiCzcLv2ARlLsICTfHShvV1Yst
w/f3lnsGjP+ik/Zp1tp5AXTzOteB0FwGAjpD2OCzV+el/03NN4pNdhOyUT5/gmnx3x05rpkcK6eL
dQi8aYIQaac9+Yzk2buPprPoToi9IZwFvBNlzjPyoBY/03seJyeIC6TkdwKqZARHY7X+Dj86WK27
o4+WDcHN8OIEipz2YQC0BXEyjzvlsJaoMUhMWtp6vZ+63HNRp5Kx6AUUlFEchzGaKi9wpi7LlQAR
qq2v2oyz6cqOXpdKSmLGAG0tKob3/YPOnKqTxghCHdy8IAYtyklpwP2Xko4IpzLtpXmahFkETNLM
+UyiNo8RaScDyUtUJn0GbNW24zkC99nbAwaBcw5t5sGU/ucE3MyRzG8Q53pqphn+w8lGgBMV2art
6jXOPl9lJlE7kL5khKgQ2xPQGnqWzyFMlrThPgqzE8Dvw7asEc9hjaFx2atLcv8SPE3sg78qcbSP
56QgIbkt3KjdGp14fZ0Z0oFd1B/mU8zHZ1sfeAxq4TKxpd/RsnKMwIzrVt1UeigVflXo5kKBf7Gp
ar56evfL7wMdVmTWxbLnazj5z8qslfovGB36XQZjH9hG8xjPw1moCs5HMD0RX9nCdHRDfgI4Dz1L
1/D/EbVZmmBqmigf5Y9dIKkSCUwRZgNgBL3URpbsWSMxiZrlKiLi/PLGbvUA7BKKWXpQ283vma4K
jw+/mD4RrNsmLhuI5GcFgoMBb+46yOMpEzcS1mDAOpHDglmTZmECfooaUNKiSHM7oIx46k8VsCKH
V623a1glck+s+ZOWZFRclfXgNVq5OrVC4+21npDAtTZfxv67uuU1eTg7EF0jIdibNSJhE85oi1aR
1n/6b0emCryWvTLxKvBub6zOrftFRz5aVgCdJmKx3PyMEGa1yqXpMsLQCK6IFFkCkts4AbQJxcAZ
jWiMCO4I2rq8tBQtJcUmMUwvAO4sD5h20rBHe7B3QO8WeQsDnZJC7rAya2CuGaVCtrsgoSnwLeN4
OwNNR9GHPdBpqJICjEgjXwTCdmjDfnUDgGZ8zFX/Sp6Qc3qyVUFPzgS9nPTkAmWM/b+Lg7p1zdF6
JmEZfRhvakI4cB0rx4DiwgIbBRGnDwhqBOLUyFw+BPgidML5pFVAyIl52PEnhe3bDcShZy3Am+Ci
Ie9d7iqELR/Ekh7lozG8LFuzZLIs8SPqI8eTw3J3ABYjz5JKHj5HtX5CCzKMcVuKg68PFuzI6Ufv
kqmHltEuHpSz96q5bgJ8GlaJJCSy1+fOq/9wQr0R1r9z7OijmPfzXZ8q/OCHKAVLkVqJdMQuzNhJ
DtX+BqpYnVrZE9rBb3W5TyK7MXST+A6Q9rp9LAZtw3qMk0xNYpnqddKxS4And3Fi3BFYDbvhH/Uq
88UDr2O977HUjSBMseMbGQb+w5+ASnJy+Xb3aPEC+sGCNhZuJPXn1rDqtlcxhc+lkGepRhZjT2wa
xpYFLVE2B5HliTbYwT3gKxF7sOc3MCEzKfIVC1UhZzWK/Y/Agkfjj5w2DssKdrjJMtn2i2bXRQYw
R29sZda0ghxZMPY+ei1EBqNbp52by1mY1vLFq3edIT+8v6oJsiGeilOkBnXd6k+27Qaw5PKW38bp
TUfXF8XEEF8yZJVwCb+avMTsqhh9u9tM68a3O8SRki8S9ADS5++0QACzOzSNoAxWQQhPqZZTBfos
HpGCJi0r+JtfY4VjOjkGvDOaqgHlAKN9GxHtFfQ7bm0Xk5vsSBJBZunPxxRntGEGvI7vX13YZH34
lEAlapT/lWDuwX9Gk7fkf4wgupmjcUvB9mGXOnpPARWXhYwdxr+5pAzk/oYI66CZQ6jcLzu36o5Y
DWcnhrlCQ9WbiX/d2SfvhgpqogKMkq58veiTY7OB3waZSgHI5iJCHCZcAC69XlbbCto/NmCjWE+x
buxRO9Wcv2E8S0rkNAADmXfeBb8K2Bi4najfdVPUdf6vk7sbW8TBoQtaokgJVck6VGQKfPJYkUoG
NB3jXSVdQhxdLPNP/3xSgcBVVATWOPG8Y5+BDoFLq3doBskUikaPiPhtvba0G2o+4p7vtp0hCSTF
FcAYZYkN60Iqx2njfxSoj0q0WWUCCrEstebzjmRixugRC2Su41W35xafT7RRIuKe5oarFb6ZwJvj
3AWxAwmhQiVVGb84Lbclx8ZSojxKkm1JAbxiBXgB3clM7WfrjEl/Op3l/0JZaQ+kP3YPQM3u1Hdv
qS/kGQqQS12G20yOFJ8Te/Z2It1NLmZW8T5YH4W6kVFxgwshuPbxcXiVEUZIfG0YpgiAqJmCgvmG
aYwXetcKQ3g9R4y9tb3w7Wx5EMf7Rddm4dRcNKIjIVRdBJ7bUyCFE8Ml4aYKPnBzbjbvFeuvGFMV
5XbD/oJj/RX21gvTlmEym7yj18nTKAXZN9h5VhfRsw9YgqIcZZYWCJmVBnIrNYfAEPITDReI8STa
78v390aZgroCrPUZwSdTUq7tx6G2WOgXXa97ut68Pr/kZ34vFhI/N6SfZVaGn/j+9+BBUiRqUzwY
Hsn+OhsmsjvC5vg1wn7wwf94vBFW6beBs9vhrq4sHHWLeoHlHzeK7sMwFlVDr6NYuaxVFt3cbRLo
1OwDR2MQLVbElA+OA8ztVBawcKP1ypouIUy8pSDzT7rXKy4jMzCPMJIfG9TgN11il6Zyr7SmxxhB
K9XWxgmVnSS3RtcPA/svME1u0eAVm0O006JDPw5sOGP7uFLCA6Ane3VBiAhrc2E27qXIm8ZLObiV
Gd2hL6q/by9oyzJXCOscLbsI9tYsmmNxXWXSCSNSwgbF1C3L+xxnA0sHVVXaFArpyTSS80Ucx3+0
vz25YHDFkw4fIVyhRGhIHLE2IdqIIcDEH2OyMAw26kkeg+HOdv4MIyZb0cVQz23ZCngRc89yX7Sv
1w/gR7jUlU/EtMqMY6mZLtbxsMuxb9/sks2dyysVkDIOr0euLUiRJ+fNp8NVBFKqXRlPSC7kU8sQ
u77cP/JOCNs3EW54hc7qBwtMyCBa3qCl650nDQE+kttRXs/Xrp/WJPVTdSXVJA52vnNYOYNMz9Zb
17N5FM10wuY2lfuhHyHbXszz5Sna6+MQBTJA8Vbgu/2rPnhoVLmUqAAcAf0e3hUzM3GXQDhpcZeZ
fYhY6DMSZuuSSuIie8kGiWafx9NRe14dp6HAmNaEKNHd1usXhxWRRbO20LX+6EZiFwSvtt9hM/Ae
hKmvKBTW7oDzURk0OJJmxTlg3RtGa48+JN+dDnMOSt9kZSNMOEosATGDcDKBgma8YdeJ8DUjUDYK
mEjUdnp6ia+omvIqyfSacNonbsPL0a+8WSwFN4o9OJMWgKdLUEPRKaPj4z7JDE4G04cTA29Lp1D3
VOXKWD5fTnORUk39S7s+hcy6UCCSX0yHw/p+cLwMOP6GVdnJo1QQ4nFraYjOhJLin3KWS1DqXy9U
2tJnhoNceQgtFfk3kt0T0bjVvPocJMR1vQYCxENLtKRWzdrLnNc5f0apCul9jkUd9s9EpX3CgSjv
0Jn115n87iFv5AxPx83LJ+CTQwXBOTDkzUpZwtOfF4B4YX7NYXjnMtxS9N4dmj7aWpzIqhgwY4IL
AhSV7AnKv0785x3wa/JKqMvLKNBGFAIcGY1owOq3SZnhPloStnjYoH6V35Rda03tDCtCnzXoh4Ie
P1BSH5+neILEimaMqeb0COUznxgoQTsMgzg+hY+BX18ro1j9V2sXk7ddmqZhwt9uX3vKbM6OwUp5
9UfF3k1NShCJJuRt0tcqmyRcRnA1W0+xLHSf6llrLZsqwNaMMX11QeCofFZej60uf0A5rnKsTP6r
pNcQvTTg0N9dVX5dObgOpGDpZG1+UKRiehjb+4M638GKxeXs+NChq70yu3gQXpCy1uPVL2dEzEeR
9igP/WjNQvtwlc/WvpoJ5jC9TUT6RA6G/5NouzQEg8XxWeyuihKMth2othEHKNP/yApTGDTTh8gi
dB5icUzTNMS9J3bv3qCt5+THiWFZcyhZpWGTO8/DvhvOb8FeRCTcuniKAVD1QxhMFHTUwxOtjI47
xAB0aI+nr0b4RhsImSzR9nZWxvfieHz6CB+sNOHSvOrNSOMWIxBRRvoHsPRMSZeJef6CTnZsanZ3
1VsaEQ3ROMGTB8yzSHEQO1Ru4SjHg1EUB9KBworjR/RQ87PFqkf6xcYVaMdfSwsPSsmTJ9nGpqsg
p2/vLucGYSlpom2zvRqIYwGOX5LG2SLFHn77qTMbcfVWm7uXUNTDt8c/8W9KGIS3GZs7myWqypD/
oCq37d8A2c+LQgFs3wSNCCZY9wD2vL1cdeGWmphTuxrne9bHqBD7IUB0K9mJn+zfrWPYtgRsHPOf
lT8cAqVcSMSerADhcI8QQW4s3Qmwtr3q7QY1PB5jX98X+vQ5Ko2XrFidaOQoCaeaBBXALowfzubG
eqZsx/uswacj/gx9eLCzZ9blnJxrkQ/hf0c/rWsykWcyC3EE5umP5fmz3O3TVntDi7Vbf65VFnLS
XCZeZGumz4tMnE/VQuBv9rOTn3AlJpJZ6nPslcwloBsVTFKnvcTFuKEzVEiWmbD8SmizJpheJN1Q
Z+hyqOT2vZpbNRDnbezvqWJ17R3zAeH+895yjVRYq/xjfkaPmYdfG/9kho3wLNBiCGcFo3tYsiH5
YTq2rxaG92RS7FUS11hHLfBfC3fT2FK96cnwWk8mh6hENgXAEZ/6KWT/0ip7zxhL5Oa7q9IXfkIg
3qE2etF5d/6eFxbCSUY31pBPq1eRDgOfossnTLlSgx22MuV9r9syLegRBQVNzJ9dxsae3CkpvOVZ
HaQi7qnVP2PcCxyVGU1CiyMynBbEcR/97Cuoa5oum6WZuUPPdwu0gKhqAyzKCX5eQGBTTUGYqfyg
9IErRX2OsNMoNvmJAAjlV7NPagdZKjq46qlHWiQbUklhQJEjv+HaFV4WEEZdoXycEZGb67PFYFg0
9RwMFwm1dTA9dBHEiVkN1Zs/ym/+kcEZ6JuBobN/j0dqfgzAJdgLRou/pvI1XTx1rRKpmGSzDb0C
5XS9A6ImUf9qeZDmEaesWXMJdXU1Dm1NCeSjBEEXeZSsh036t6e9SOzf5b39Ne7TkhZPMSfdUHbC
/BivD5SS2uDQRdsu/SRrL4+SC4b0sgcZ1OIAaqi09fpnXTZZn4gTPuSV+y/jpsFFyGRLIdIc2pP6
glzb9vE8XvzAPniN4J0B+1ydrkqFTQyQM+3WCaHA52S+PyWWlEEaJ6aEhiHkU/a1WnbtNJGzJ6EK
rFJBSi+lScMbU7l7xOHXB0y0v3LBGegzsJ6n9yk/LC5GS3Klp3a3S07IyGAeqy3PD0x0b3Hh+kN5
0ySmpwyhzguhDK4FLXD9dPdEKPU7C8GW47FXpZ6YazaPr6o6FaDfeSwWD++646ItUgLD1MnW8aeb
A+Cba2PdoGGouIfwYXVe6Dl+zI4LECphudHmu3uKdGvmBQx2hhTSGPTWuv0mhaFY/yLEqqYvwho5
9jyH6yBTU6LBavNyPhxFvr4jANqMhasmQM8/n62Hudn/kGd6DKYDFarZ3EUnVlX9jBOT0scPHNGs
Ii0v59HHw57eI1k7OibawMp3b7/+f9jLF0bfvIIL/n6ITY6uXYtmIUdnyWqcWVGekc43K/YI5cSP
fLbU0zHBuKgfTrzbRUIl8cmp2/3lKbhTj1OU9w7OSrYJQPMBmNM3X6/eFwGVMTh1e92ieBVQhGBH
UG8xezaaDgKfW93MwTdWiZyiPaybNuaRahB++nMFOTpbHGIpNxkt0xDZP5vcN9uTvvU5uqIvyZy7
SeX4fslROj/eJmqLKTqxsghK1lseAfBzkE518fQMS5AzGHFH+xiyWeaWjdQx237fcnGEWyHjA4UZ
ojflDoCwxsTIm3xW4twOSGWNkm/m1OIln9o+tFLFwZRH/WD1Zo/51YNgdbDMVYE7cOk/HaG/6j6O
YsWo+dc5TOqkWWeqV6U5wgdNmcT+HJrRhVhBh8b0pFK3PMNwpFkQJ6sUD+rn9x0deX56Zr61nve+
CJnkhm3vHRGWvPlcJIKiitnM0cd9kkRUx5vWNZ4UX4xAgvPLeMd5ViVuJ+DH+XAYiwsgo+QkyQwg
jCFH8tnuwKegAV4V0ppdMy8V1B7feOJ1BmhDTC2ubZIvOrx1/HGoS513oyRgpDz5lIkrCsOEsnnh
3eOjemVHfGifUC95ZnlU8V2sstwvwF9Rfowzbxlk4WeRLb0W9wn1mmF4WyYOlZlbGviDRH9lIgZp
GOBqCKqLu/rDKlJRkcqgz5gdpIx0IQXXmHrYvovutwDS9R1PR2hsZNQnB5ncB4CGzPPxkoUlxFht
Xyvog/w7AQ2A4STreyIp4Tt14zn8GW4zLKFg2gTneSo1wfRAfhTN1fK3XSxIcpuT3rnsDknYvgFk
oerSiWPIUTbUKA15N1OaR5uXz20hV7OSgr2EkfeDUiTj6yEhaWg1CY3nfGam3kzhahE3ZMtxhHeQ
cIe/thRp0r5NZ8/jAtztTC8d3EUIXBnArRO1wiEdYaeOv340XCqBFtI6PMch5iJyUOlm9EI35AZx
f/bReVTAoIWWBvaeJvUV0yYgNyU0OsuRZjJJ62CkWVvKHRmHglTUsmoNMr+7FWyak+7+OkX7RYTz
O6d0mqgIItLPugks3yyVBXHHQ0Z4tMa1RxMrePFqvVqNiNjnfUCojkzSm8C0BWTeQ9BC4GsKyxX4
qis8du6GV9xekPk2LFN/MpuVG4gR9znb3LEtgV1P70cuXVERzSkKM2iUSYCF8TSnAjuF3eZbtsWI
65ULFiKQ+tesmuaUDbKJ6hKXFUCzURmNqsTEcfNaCZ8DqRQ/52OC/NJyCwpr/hKPlTdHZH1e6jsM
rgSFFgpKbMkxDik64PkYv4vXdseA5+X37rABR2cNfhINiEWYSphEppiqnciDpAIimqzQvIVELN6U
/cvjInRhZDZJALANoG5WzgJtc/3oaauyVai9k+pgY6co6TJp6R/Zj6Tjv9sbRU5NZsVxbwxp6/JA
z7Jg5T2p0Yj+u03wBDP0iTGUz96o5L+6/Gx3+7Jl3AzQYr/o84eKsvW3eTuJyfpyUwYcC0h5VnDJ
uy0fb/sHGr/Q5qO4k4hEz/3iLvos+qQ0XxaZB3yLe5MGztP3MmwhuYWkKAdPj4yhupcZBIiQYsOK
hTookoRHEBGghtzaHPIy1v9F59eemqWJ3OY7zO5gDN7yqJkso73O/eNa3xr4fm/LYgdwwtOiWDMG
mdF1oaBKICWLhaJGWtLNGNl2W15zXB1WXKBu3nroz3NtDua40xfaPb9N9pQE3H1T028XeY0EaTOn
sFwsgfOxOLXm7mPopru3ZXKoA/936qga4lOqsVu12DxlkobKhfUg78dWbWj7ovAsawkzmrI8Np4V
OmAQHgu0829hUsas2HqyUIRydEH2hdgKRnCxgjoSy7m9+Hz4BqUvusXNDUP/PE7O0TVQkAe60cuw
XE7FpAtIhCYcbAwkYtQsrCLQdZZ11JHaMe/rsa06x/c/1hHhVqVAekl1EVEPH7fm91iPVuuyIQkz
XIHnyat0+BSiW0EfhR3jNMRMbEaoZBi3pGgEp9TyoCpDUGOfi7cFKZXo/rGkMSZLm5THvUOiYIAz
7B8G9TugiEErGjNssBq6j6aYzEb2sCSLs0qijcH/cQ9O9aUFcXobNqREUTyMv1RrpwwRbT1Emu5Y
RR1RDqkXTtiZbrm5fupc5GxxGN9Nm4+7OfvAZ4lObai3HRtraFJNHxsmsqFgs+y19GqjfboRf2vQ
H1rV9HmvXelXGz05EEeE+p2OvEBPjq713UWu2EO7NHYnn/oR6bBKSPP1ENNDhmujy0fSr3ijdPY2
q9uWwB27mfY5aAjXJYT+IkXa7vFOAqNyqMzrPEj0h+BUY+QQBHXDxzpEwtejQ4TGaBx5ZiZnp/9O
1TyP2JT11BEU0nmToumFrwWKIGaG04v3cEP1zWbs6S7k2M0g3WeELU8pBR1ndpsAm3i46ck7Onb/
viHMFWuL+PeH19Vw/8ovjbn6KYPxqM99oP2LWABjuBrjkDKmUYxb5vBkwhOc8arxprAtGV3dfDxh
7yB9Nd4LLWWW+PuNHN7Z62wXFQ2WmNRR8QN++D2LTReJ4FFR8+25k/UJcVdA9hc8YrvVvmKR0JWe
8TzU3v5422KBsvwKyEbiAAP7g/S7jT+Dv0+jMDeLlE/5eaQIlzN9wUN9k3YKhfez5NXdvubmTnrr
TxnNrviX8o7FbJrj72YPbeubiqXZ9VZaM4WAMzdXf/DXMvZWsdZHHkZCymKhBZddkZShytxIojd8
b9ppgEg/oyH0Qkgz0Mr8EX7P75cQH572/D/isLT3lyz+FgJSHZj1/YMKqOQu40bxd15P7OyFiK5F
Wx7Vsl7wT6Yba6lOR98xcY/CcxwsC6AzPDzf61a0xhgygRVgOWU2fiMGBldPpBIAhKodBIXLYnjB
ACrF9s3iW6ePVj/k3rlpToRFT3X6kUb9mb8xplZUqKSWFqLwOSnuNUMmrFDDThp2xAXAg4+eAxT6
Pkui/uXna0DcrbldF9O8qWiwG2+M7mA9CNB7Bn4CcvY7T6fUixUqKduBWFQoEgp/9zU6gPWb0yK8
QFzE3E6j/6dYXLGWH5v4IvhwrvYtPcvjlASfzQ9OTYBJfz/Wc7eOGisTCBUnH8t6lhy3cXBDKKWF
d/o5g+m5/ZcMawnl/mRKcBtuRB4UDQrIDRHqTk/IE+82DSHwwJebPZfCue4qX+yj7DQXcT7DyC2k
HRNHIRArxIB+WSWn/ujM1xlN70E2zA82Ddm1LQQmmgJE1R/8UZAGVThElgQbHcSEbNXQDQxkwCeo
D7XedKUfQwcGF8Lm2oUHaOBuqQsAjmgWcreU/ardilckpVsj1UzlPYW+n1D3CL8yZ6VG16R8CGJh
opkLlurjhnwPCtcIJfM9vYEiRiFw7jQItCRDZWNNF4G5P68CDT9pw+culCKDJAkc//x1VxEipx16
0zdwanEacerl473O7+tUdjyghv8UsSqs7HC5/dxeigypOESCDrnQnxdIz0mbKXt1s4PHgl8ypO77
/tyWpbrdcZP+T3RpmxNTHxo4dH5NCcyLkYa1IZHEHWA6+HXk8hUoPlEFRPbPAr6THDTNxUq7GEXq
ZFXZt62a4CIgpoEsQbLQP35rJ0aX4PvCucAmtRXcUmNfP59xB36hr81F1if8ImEWeESV839yUGW0
nMKCT/QLk/DlN0TxIQTnhhFw1DkhruLPr6llXyEwirNU2q3JW8fdpzt/RS3G9wmLv+EGXRY21PjE
vRrMma3MSPZTW+1xWYcqkNTGzkhcw5W84jW7gUMkUk2rnsIkcP2B/NQxB5K7S4e+Oejv6XEuzfK8
Ayu30UzbmxIRh8QtfgW4q4kFsBZ7L+Mgp7mepVsV1guNrze8EnOsddQFCdF0PFQMo4Qx3JlTEjXR
NWdjTpuV25VyP+GSIEnb6JIR8LEY0gvmKTK6zJdGtcHi9ABPeY2F3WwXuYdvEA8oIbZXtaKB7c6Y
WJd8LmsmP+yHBsQ+E/Jd1NNmL8XT1IZ7by1zs3JhrKsffN21jYpMMIvZEUwQCafN4oFJolsvQQc4
sfQVPmJ3TZthlysYUKTEhjANP3UNun7Fg5oi9LSwjNzG6WBkQZbzQp956H08efE8cpujKMfZDHIU
5AuYghO1inOakzOo1qSp9JV8JuGQs5QslE2O5IFDxjgm0Ir+VCiyAVmqNH4WXPi2mWzAPNWT1Raw
PmhWBZINYvQU/22sVyYfpblkF1E1PiWEJuvnftp4HnglpPQuuewYuzUjtEcFK4AyfKk/gwY9feTJ
IzkCX9gJdyXx3+eJSH2zWM58VCvGCMTC0HtEKiGb8V4bzn7lN80CT+4YZ87B+I8j8wbcFUZhRiaP
hRWY/WzV48nhRwRPdHtdTrmffkKphEpnaMclBIIYPt+QXg8+JVPJk98jvSb2raXLQi6Ry8ST6NX0
IPFXtUN5uXSQPlzum0027GDok2VXzUjHDzziSjfu9YvGFVTw6pdIr40dCXSZ/1xx070XdYYWsH8c
atg9+pn4AoqGLlIyFL+wJUoAinT5Ie+0NXP5TzgUuz1oLsV61AAp6B9zamMuiv1Rgr4wVzR9HfEx
v5LBS0DVbVDhcg/2Bc62lkg60uXWUt7MNhWalzQxP8Am4a2ljyYHANsApu8ueaadNeoNw9EVLTBV
rNjwSoXnE05NHtOHlzttz1TMU5rwuJPksY+frnwdd4MHwkn67Rb0bVl1IXWljxUTKJ+paM3MAnM4
+TZK9bt+4Qn7CGoIQ82ZlrOwllRGjfMhxh1hqAPrFPmbUb8kdLwi7VVCx0c3dmpnZvyVM5mYvaLU
1YoyqoWbqODo8SBGWptg16duUCSytIQd9KRUtiBY5l7OgRxY3aC5cfoX6v/Z2ldYQ21TCjny1S4Z
SWnRI1itngDi7/Uj38Zs91i5+jDQFJJcYLswXywTLpJpuEaykmV0kQ4bLSyzSOA4ihHY4ACN9flI
gh+urlDJ5tXVh7nI5F0f5lUDMG/SuQc2CYs1xAH8W8peO3QS4KNJpl0Wlncc6Rf9WGa4VZ0CELAZ
nShoFV2fvJ5xF9p2FxpOBcX21lrS7aHK+G9VHAorE0/WdQQ+KLmew+P238yoFvSXy3yVZlhNMLF4
7tiG1H3zgQiJAWoqSOrf2yWH1zyY1J6QvT4Hf5QudLcLWibhv/nCZbtmXyWwiyikjwUktSfnQp+V
kmR3+Nzja/jDwzdFPRCzH6RPvOo91/l8Rd+Yv/VE668cF8RmjZZ3epyFcf6YNJTxbfoJmSPnN5rT
voRM7cAjO84dGtcAU0ewpLgsCI5Kh66Hr+7JjGS5uynOUPXN0y1PRP5abiN2hX9mClx/D7FVt92E
VUaEnfoZYcGdYqWBmGb2/KiCzdloh3r9R0ae5g/4JZjoKdES5FxmAs+BzaLVdiAq29fthcAtD+MN
7/IJwdMh2P9OFCxMqLRbV7t8uF4ZjsKJzR0Bcx2PAA8nXIUdmlM4UJ2MTnWLSmdzqRfd06gUj8SA
fhN7HSjMqtncsHlbzjY1az51A4m3eu7yXIEGCkN7mpRApUKrqSHMFJsgbmZHjO/JpWt5IeBA8fHl
G7CCpTBOk7wFAf1+0af3h798QO3zlmdD8wGNIUVFn6Cba5uib0PIo6fLJVTndOonnbePF3l6zryB
KAP1MehruR/4n01xezO1UQQR9h2Uvg+Br/ea4FsH4wZFyF9J/jTGybPP21PGipeJvsOswhEY5zzM
voXqn1SwtZ4tKi4ROJ8l2i4QfQ0k2qNDDGUsoJGIpUV0H8sCmkpzdFS+uqSr23rPkdVe3J3k9ibd
eQ57JS7A48RyBkMfNTdAvORQOI6JQQ0QAY6zeiW/JZofV6fB7xA/cb8boPOgHP4adH5mPurwf+E9
WiiNxYxr57e6/Ejkpv64AMqK9mYznj1FWbLR3Accl8bJYK7xV9gY2rSHtwD7CgaveLJ/EFw9O2eY
+xfqY2Daa0DqFl1jVVVFjO3HKJm3Z0gkL5dg2WlbJg7kH9+JPfXxqKcFp14DqHpWqNjhAZDKrk5n
Irvq0lt9PbWljQ8vNvNE0uKCJS83/dhcET//65EgQHpn8cZym26hTOxK4S0tAOx5n0XMPCwzVtyj
sLAPMZM8h8DOgR50RcrBDJT7HrnSi+/Pcm1v4HJYRAB4Tq3Egcr+MU6nxNgYRtWVAMExGsWkZb4Q
PwbQuCMqCH/dCjVEuUiFN1gz8XBgvC9cLhqR36tVisV4XONRXifL+yfEmtiQeRo7rwNQ8flXLl9N
UGIsefApdrmr4/CaIc/sehsjOhLOhspzpJ22TI0oxSarvykADiXXlNrIfaelYY6RzU65NT+x0O/C
AyOGPTIkihYOIVg0nQDJmCeWorKlzVWUGyM9/upGt2umAlOHUthNTzWmLxc7iJzdrf4LdZAt5IZB
xu+DGLd73OWFOEwSonr8MN5j0sqU2NOKBCpCHZcKji4tTFZopdCPae4164/QNlCusVm7nTEk8M91
oDc9NNisRkY7YdbvLsITvSASle9dT1HpHiH53oWf8MGLpkPBke1TCUfb3TWXh68W9flw442IEajv
Mw2nSNwLSHK8fV/FVIEIk5/5Xj2LXGBxSBtH2N+EFLg5C2W40u4IelZT4gVtuzhlaPPP+As2IFkC
3uQNzmcmAdb6Vhs9s8xvX8aBDGycBTTqQ6fEwGU5+h2co9OyTThQ/QJXJwISBWS1L4BF/chNVbYv
c9nZf8+tmubS5CwlJhJq3f2W2+vShV655hcJ+/bXE2iQQh2WqLZOUFHfVGF2rZBWGtCqx1Qvm5Zg
+2Peto/EXzFG1lmF4u940S6218K4ySLFQvlLMNjS8DllRvzBpErawlmR2HOkAA1b5zh5ZC5IXDJn
G87FwP1KTxMnsNEtzbBZpuVFYqpeO2mPLM0qQeWilkuOd1ID3VAr/1KRYzhPwNzEqE9m1RSzbMXM
7a8GZVChXDEwNYeW8MFs1seE4HkbaGd3PYx47T/4EbA93wHZbzc3rIEt5p0PqlN8ntVnaLWrhBUm
iZEW8vle08IqRaWcZ+fTIe3s/qKr0hCz9OnwnIWfJ/tksoPoG3ZHpAaa2M3FjzQ+Wr9MpgL2Fo8Z
0FDBTJVOKArce4UChjgutDLVTaz/W846B0Ry3tzgSjaBXqLL+y8ckWhAg0uZsz7A+FsmY2PxpI54
MC/HrV3X+VWcYhwu73AZ8ozZo7exVLmhuIvVoX1eZyYiwbI709aoVcysa1FLNE0a64IwBHYWeyoC
Csoxye+iu3f/HERxfnwUxwrJ78jXNbFjdiWVCM4s/LNZuN0svEs2BQ4zz0oqoew+Lm/tD3rNZAAH
S6ZXTyS3S5HKPQejmzJ8rf96WbS61sUp28gqpVCDFnN90+F5v/7AKA+/yvo4WYWTa3jqdGD0TqiP
MN389pRy6Z3nNa+fwJhytlf6c5FcmsMU5wuI1ThEVZhm+wlh5J9bwIr0XYiAkX2soHR6HOkX6ni9
ZUJcBhs6pqz/wW23wfAfWz4Ew3Rab7ozAk2LYVya9MRGmHeBxsQGOBupMOsPeqLg7EU+2B/BmieG
yWxP+0yj5J/9UtyM0PJu0Rcjgo4isXC1+U2lfyuzbOcBklZuTll8tCBXZsBRXoBn3VY/aZFwUz/h
RGSzWRNTF8Rmmr+avwRWtEwxrm8I8JMGVdnMOk2zVj9uTnEgXCg7Uh8GqnD+YZQg79iSLy4mEgaF
2lSWIg8aecLdA0G5CVw1qjvbtloCU1uC6sFVfXaheI5VVybEHMoX3j02DUWpbf+B/UqrR0kT0+eX
qHCu2BQN166+xs/xnhsuzLZ5LEE8WrdksT32omKoHYsw2WW6g2K6n+IGiMJ8RBxYtLxU4RRAGTS5
xfIPQ2tVWvsh/mG4QeQ3p83/mppthOQHl110mV7JHOZ6efxEoRh3vzH+TTwh1zTwmcozfDvdLmK/
BVjmdxV7nrWDOYkQh8EGGNT+terBrRoQmubr5irRUNKsdEViBBm7EH9A/nLFMda4DQCmLX6oiN2I
joCIioA4a6+C9bBo4tKNNchYvqcXkTtlhE0LJ2gA1yobI0HkyUHWjNBQeuffcvwdOHwfPuS9mFf2
GnULs7MqgUwvJKpvxNGPmH3w5XFXiM8EYIZL2HIxgeBnw6gOn2hQ1zJNl8VaL6dPKXzfmi9gKDCx
VJll1TyDPBhbRyoPrsdwnfpg+FFX5253s27u5nSvLkBfnJk0o2RKMtq6DQRs6KjDjHPoyXA+5U2F
tt3nvYWpiON91xDogcKct/1qCA7ctD6rwaMa5R4i1U91e3mGv7toiSCkmx7MVP6yhU9F8HbW/mJY
6woyN2KVGosSy0LRItvDERsJbEzaFg6yg5llt6urdJZKi/5r6daYpu6Vvd/xQw7+3REcUFegrcIZ
U4mGb+ZmPgTq4GAC6d8QNmWZekr2NZwRCG4qnqt7Za3rAU7lTtImJ7h141lRHBT4Il7Tph8+NACe
CynTrAEBPYgLry7nq1yhMbylvjoVX/x7AIOHOuAlY24AtwcXaA+fyBDPLZPvyYlQVaxErrRXhIVA
JlplW7vBJ1YIJiO22oJM8UgpWn/VgCUQ9TeGdtkqqvvJED8kPO+tT1pZtTGzho/eYP1t0gowcinE
C9O0S71lXD34U7N+7VKuaLDJNIoegcemvo8jG0mX58DZvpFWFdM+pPKGUp8TzBo2b5ROnBGMjgNb
zkXf5Jv/Lhqtr5aMgWntCqrFkQ6RM3BQI0VRJutDFqkNoTBMXnaUFANO9Lsiqdjy1MEGp4U5Rb7x
rLQ5tOfyf8BEis4AFPGLK2kdRI7Xzgb+sd5GcfNWCF9RRhyi+7jSGP6IGBpnW0wLLfSjmd5Ko8bn
I8NaC/hf7I8Mj0FJs7Xv1S738n3TEf9in1EPT12qRtdGJeFQ45VQlPccQ+lcMqHconp3aPtjeIwi
BDOJEpzXjyn11QrGmS+jPx4DOAxfJaDlILJJOqKxQK7b3HKLXH+wW3fUwkllt2bAdp5RckbwT7DV
uP0PXFxEEQzZCONnoLtswTpA/xZ2Su3yE42BtkC/WeHdNFYqoKlpto2UjEN3QkAiq2Fs8tyfikNX
PDyLJqQfhILXHjpzN2bthzFqgHlOTV2uxbKyOKgKVy3VlC021Du/M2RX9vhDzcolwXeQsqSNn/Fn
CrFhbTZT1d/ga098rOdlGwSEsI6C9zHf8PrsQiLR7eYa36QGGU/nq1fOYGYVy45jFmIpycTpLTAF
tQ4dg2G83enaNWL3hoSzA4vCLeS0sXT8Ph/Y0ezGVljnAvfzUHlfNQZ1bsUgO23Ul/C8mGItuFF3
uA1m4tpULL4Mp/lWU+fn/rvDLiFGXhQaueBEwAYA98419TQzrVgvN9yJqx2mLKLJq9LboAJ2z0iO
d+IHrJkxx/7H2yB8LM//ElBADNhG1KWGnufH5TJvc5WeDV9rbse8zjyx2SBfY2dQAjLt8lDYylDw
TlDoqj1xO9r+GsSF9iCPykCnK66jhPs+hBX5UVm63OhLgtYpzZQubKe5FTmxKMkgVGDjHO2OpLCH
sszsqCPjTbB3O5DqA1oC42clxDno5e0Ga7Y5FxGO5YYwNtnXQ3rhQCuU5FjfIzbkPCSRupf5UL2d
PYXRra2CZFZ2xTfkPlPt6SlASWkvp9p79OXS/S/kgoh42mDSGLoODpDafPY2v/AUmTTU1WUuCe7T
QPLNInMT5NHt0xKBSUIEP+/ZBsJF0ITC0l/nK8YlwFih9A2ippLC/nEkYKsf2hkZnTCguCoQKhcS
DMcppM9zBIu8WTRY1szHPePTXMFa0m0jzhlcSjAT72Nx9L99H4+QeAp95l4UZPTDS0D6zRyrGO6G
h+WBsUXTRTHoh67nD32g249mKqCt/c5iufwi5ay+7VGnefn0EMj5J6EbasPmSO2sGmiCOJTpoUvH
tp05+mCMgn2+eFZVx00FKIUPYQdva3glqgLr+ctUgunzO9O1RidAMlwJkCZcHS6hc97WqEQH93jA
E+nteAElQhQ5J5cNyuFVHuaoCWJcdpNGRHsUxwCTkPMRCQXVrhBuf4TLYZ9u6yIaLsg+pu8vKBmz
TPEbt+EMBcz0dkj4oyuGpG34a9j7yQXHxO+BLlasGsppkLYXw4NDWpFQCQWBmqWmIPpFgjYHghuH
4Ev0zUOh0Ac3ueQfb3k6TijEvcF0tBW4ZiVGCNbgpm73eA48ZFou7gyQnW6hc0T+KxJHZkhx2gX+
CgVVEbjNS8UJNKEvFsc+LjDzLHtkCFEdlp7O+5DFQJDc91LCq1Q0QVOU6QNScnBSVUji6wBCC+pH
zlySIevqvBbO/mf3os1euA2SogIMaUANe1xloG6tspN/PdvTqIkHSkg1hdq46/Zb3yAb458IH0sL
QEO/PwsZQoJCElCwjvhHaAx8ttj95omkzLikUO///leucEPfVsb2TizyqHTuQfkFgfc54YpSdwFg
hZuGwPhADQ/OboaNN+rmcCA9TbsMf7httW+D+RDX3VfEN0QhTJ/GXB1ofL42tluHw1rEYx9gLt/n
Wmc7UtTlBbIXt7Nm9LTtLvND5rAY5Yd83CsUUP98cImaWZaRRzAFr/TqfXT8EFAjjpRAsQwYftWv
vasy5x8vhttfIqSyJLA99K4K0dKuz8N7OySk+RGeNbcoEIjXAivtGpNs+I63BGUb6QBuVNsilkYI
4eRy896lr04DUelh3agxo+NRDbwVd0qRHl5/cyiMbNAM3XnNW/BeKPsUGaqOm6vhJQw0TrA1+Brh
tRfJJ9hFDlk6y+67JIrfZqt8gwStPdW6ecRzXq+TkmpJt+PKqrz/GZBisSMWlXbv5WQixNcWYWgq
Bo4hYI/Ha7lkUfwhL501/U1OlQyEP2I/brFUrzOvIWX7HnjEC4Hg0pSNQqsvdzA8IS0MXb1v9edx
EjiKmyu/OFx/GngTXAbfaO7ZTjfdWvdQQqi2z72TlpSCHf4AWX8l5gY26vkh2ZPW3BmuX3IM9wmC
odsbRd62o1moXdB34Bwj7TGOq8td8THX51K0+NVEh2uV/mA1k+Vdxa/aD6e5IPurnhVx1mcP1Mz6
CsUYiJlMs9mew3aqyyclLN9TweznJ0mUfGBCmR2tJE0qhdQdQveVuh6IWac65MAnZO9tg2dkbnUK
W1wNYwd4VUu1IkETTMKGiEdL3HWL3QDA5JwIWpoVU6k7P2gaFrZ550CD7qXEd4okBDhUY++k8q05
99Rj7JZGgEQghj0BZ2ktsQ+bc7800PpFgn465Ja0ze3pbSZKjDAZTHWwzXtbUwaiGCywvFwfcodA
QXIyIKdMWA6vwlzvadyHEabLNd2w85S51X8rXfBxUkmsDcJJLlcksy7t8O0YfnAVQDpN2awGv0JN
LFYZ6NvHcHIdDhzhPupP8tdC5+ACPY4+rnWBXP2Ui6w1t86HuAlfPfcx4sWE/VmVikqI2M4W2YEQ
Wu1GkHN2ShbJSWEjOaNQdAPS+8wLLqRZHD+iYpCBosBUBdU74iP7l05y/zkJL41s33wJUh4zZgq9
jdzTo8h3fWEYULlh3sVU3OA562b3q+eIGhb9eax999yjNMzZrJJX6U/jh5WXub9ZNejqO6He7bmX
bllNonIG0ggOfzxd6g==
`pragma protect end_protected


endmodule
