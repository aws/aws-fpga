../../../cl_dram_hbm_dma/verif/tests/cl_dram_hbm_dma_utils.svh