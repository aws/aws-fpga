`ifndef CL_TEMPLATE_DEFINES
`define CL_TEMPLATE_DEFINES

  // Put module name of the CL design here. This is used to instantiate in top.sv
  `define CL_NAME CL_TEMPLATE

`endif
