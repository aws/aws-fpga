`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
llGzHlLmxjnydZAk/ysliPuLS5mPcUH2rLDBuQigGk3nbVOeDhQ0qzgycSNsx9OevMccHEj6f88Y
VWa9askX5ruwyRJ8LUfsrGQfky6LgFlOzthfOleu3BKlVdmPrrheSKsqp4skeJ6gtafazHuWewD2
USWBWNW4BWDOVtQ1BjURLzULtcIR5rzYgcLG/zxy3iUJ6pz1pC9fC+UW4ZvSvx4Gu/3GDulTPkeJ
uV+2MM97Mq/PoEH1jTRvokqsP8WMwM27bUAJAK/kBAwZ24urZLsCvozWK79CvgAM3uBdLOWUMRd4
4HKJgM9+Zl/LCXOj90F2GeTl6rbysTF8R7QT1A==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
zp9cqO3X0WO30+20SahZk+ERVHg6VEUX0RAjgqGoL37Yy8M/OiCPfAZh62OgRIWG0QQQwaLHGXfe
ltyxmCvnaBi3fkoN/U1WamFcby10nSXYq5c4he2N8KjNPK13QeYBRg+V/343CJ9/KM1UrYF5aTQj
NBy5cS3pGd7IfJxLiok=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
aKD8OFYKPPZhWVxZK7crrpAGuxx43clwHCRix7rgnWP6GCiCl5Q8/xcjtyHFGd2A8Q0a+UX3qUc8
uaE++wefuHP5+KnyQmtelRmG/1ZGlSXltzOWb8P0fBwl6cemcyTHulRQZf58buf3i/FTDiej7vPy
OeMyk8Vtfgo49BfL+yI=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2672)
`pragma protect data_block
+//UvX3jMBUeXxZEUboZ209fpApbc1XQHC9oWOsigoy730M3bYBmq5uCFL56ylQ1CzOMYGlrnROP
slujwuewXPPUGeSPlADAa2opHVbVOuBFD3CgMnVIay/OJnwYIbeUI89r7OPRhwoDgRhJC5EPZWjV
KFkOGks+kWDx6sw0nU4UgqNjijnh37Jyerk6wCIXTXfpqmrrcoiyflxPW44PNhhGhU+/R/TORIN3
LnFlCJVXOdftD847ABCLngP1tgGAKoVVNRbY2xxLx60IuWCSjqYCSqSle5aFOdRiYHWTU1PZm2sl
U08SqcyDgRdGwG1a+3we33R6yj3Tf7t/W2NcghzkRgynMwkJKbHZi9DFOCgxZmSFt7a3Te44B+9d
QoeLcV3rV0OD+pBzNEZr0jVCWUcYwWzr4n+56kIiN9QSrM8ZF6wy+CdNWIzVnhy9YERWIGnraKbV
Sc30rsij4OB48ZaD527gvnEcyLK5CF0ZZa/ci2nm0uMXhqStAsCT+5ezE1E0O+i6ykid+B5rN2v+
ufzRBkkbxfWW+9HkckS+doObkC9TLukBptm45P6VZa+NWQd/kHjpY6lY17E/bngATdZWWQPaOWc7
eb9HLJwwgjnkT62yk+P/qVl6CJGoZ+WM11cU51BpS6VR1CJXKwtUtXMMXoAIZx2yOfq+OHXJi7KE
6Wk+B2LKysfO3CGf5aKO17zhHgGbA5+/1LION9qR7lKgTHMqUjSeKr4K/GTyRiY0VZ8oNGHCIYUZ
HVbhubyQCIZYg+a1PsNkPJbPvSlQ4AhshmWBuBi1g+9mAZw0jWytq0/0sAG0Y8euoLe+D55U9pMz
C+RWvSXZ1NLPG4Xz/vEXadJU87NqcHhqWAhOKR7r9h1cPL9UD/I7mwnXL4KACrQIkhp8W+4sbiRN
gVvcfOIxs0/f8K+S1G0Zc/GNAEkuf7H67YSAntv/zFtmDs8Anf5JByDEKwXYo/Kahz+5NCid04ox
oDP2BdN2DTRVbt3dEgGISvd2QjP/Au5I9NSWRHtaBcd6XTB7St4r9hJWvJ3uoL/EEdo/y9MqeuRa
Nj64l6ZQDXeaeJe2P7iO7/WMXqqVdNh+1H+CxNKyP/AGdby99TelCDlgxE+mCygTFSXHhtjiQqAx
X1kDtP3YPT46jDGxSrM7AT+pGOg2Vh37IcYvQQh5iwU7ScDYLSnAJfzbik47cwHuOUX9CeiW8nPp
+YF095Uqn2SU652bT0om1+VjFFrVR1AayyO2x7jasL0H9Le46D7a/0Rp5BNpIFgBhHEqD+e9dcyy
ii9uWst0I59nSLcT+YbJqzwPGn3BTTwQy6IoMnvdFHSI9riQDz5HFcVL+784z95y6H5+V1eIhyGl
uBMEvSj5CZrRGjq9Kz1InAM9FCYs6uVsgMTnpEuHjeE6/5MRNPCGGBNifnyWm3evqFa7XMjWQVNB
owYINXuDxSC9DVRMInd7A+SgzScgzSbE87yeUvF/8LYtJ2JIG0qOk+r3nR2R5PJxA1IEOOVGY1uE
jMY2tP4IxTKuuIhb3Pt+42e2WB/thQdECh457vJR17GhITtahAc3HPURoXYCwAbsxKak6l0Q7tIg
bqjQwSSvVh0SFVRjMPY7HhR5qgL6NDikcaXS6t7wCvJD6xaBhetTbiMGkVMTzP9bc098o6NsASiL
G9TRIs9IkyPnmBGUCz3PIszIcVB0pMbMyIMSFdlk1Ovyy6mTjmKvCrh2r0G6v22jqPxB+WH7scSt
oGoAYkTbTfQJzTzqrp/r8Vv1b636dULaA7gSF1DpSMezq7hAVlY7S+exfCYwXpOtgjqOwdZ03D2o
ovXb+IfVcPOiI5PYZ3JCc09r5+IvrNU6cpRgQ5Jgt1KszddkIjCK43jV5+i/RCj6CcW+Mzm/n/BE
5aBrDpwtMB+80wdS7QTNKgCe7P5Xhqa9yREIjHeWWMK7h2JalGWJdbPgjfYq3/lKLNs0wflVxXQk
moId0lG0ZEKkrR4AZ210zKRU6TQPfOXXJzImJ2qqth6V7T6kvpV4+0QFSajpr2hOI9jJcwYJBWMF
bD8zunXzqwUBZ/xdXhQP6gNDohNXXxbfn/jUFgFwR5jTJGYB1xfSugjs1vSUgcwBYYN2f0/K4IYY
7zDeKKENoQq0G7X+oi9D5UNaW5/ZGgJnquqev+ilywO2pBE7cBUkcENa5ehxxR2fvzVdanO4vFp5
R9GWTpKGKE9zaORTMdlB9vcwnyfg8UKI7XxjKhQq5pszZcP1qkOwb/jQPkS/SJRt2Y2yqvOelRuG
oJfqvxVrWOxQOltNxhyQ5UU2ttJ4VBl2yGYSm4xPqri3Q/buTRUIM4wQyWM9/ZzVCmAFxohNRRfO
3d82pZooIjiWziOqrZIPz13QF6XDE1ljq3R4m8o8ZHY5yrLMJsVFr6osAi7M5w/fqiClrdXHCfNJ
y7+yA8t0nNT61qho7GW8KQeLgeO73Cd6CwDjtA92gJRZRtxREUuLF4R1UF1jnS7+1bhJwam8rjus
Zb4xzrR8nKMEPuWBdWDBGmV3FgTn5AY4wkKHZPg4MJMAbXMs72RWYOReY7YFe7WSHQx+2TdQ3lB1
u1K4Upup/g0GtY0+1iHvlZS6EGcp9vlLPrlgzUprzuUo8kM/K/79abqb/ea14foW9BLSAuwgD3Z/
5XJjjjyVBXuSa+DXwiUxz+4225J1GiZzoLM5FCo67H0InqKU+73qUrDzevPpedF/3m92x42B53il
NkvePCj9TCoccTkkRS8Kb18bLXExmD9cMcaDv6hCWfQCltK80pfTkWx8/yNQCu73hzV1bcay5EKW
SidMUp1LV+x71tw4nydFJ9FtB5yBJntrPwaBO/uH+H4FGjAYb3cC9awZfyiaSEUWfj2cvG/17ezZ
jkwN/DlahCjdzlYvKlvZcYyX+PNNjFK6JAz1sLORIqvdZDWKutVy/NfSKJO+H90yljx6pOoRN6zy
EdPIsoEa5qnc5vku2yrETNisiMSgvXZeSp2SDQp/5KtfJFiSOg688smqcb5cgXzk/J0JzUctxFyb
kTyUo8oIG5ZkFeN5KrVYMClAKJJFxKd1kH2dgk/KDbq6YgbP0Mwh6gPO/Ci1ylTwSz51HalsbNqN
F0mbIS5NUgTrz7BBynqj3PpwGN/LrI2XR22c6cxrwCxXJUm3B5ZiBzdKHZQDrOhKPLnD0McKSsWN
HaKigYILkRmzc7u0sDwLt3WjfaWczpd2rEepVJPU4EQdXEIU8eMFgiki3Go/J3rj3ez9500njGFv
/FcSaOl9XZ3RNkPVJmhUXwFUrolqXEXqPmJYocc3tO48bXt+STL4CHpBUXxRn917Vqs4OBbp2FkC
GOA5yo2zHhcfAGcJIK3B7FFIxKBnML4294CwdUPalKNw4NsTZUS3oWDCH+4A6OCMktPgAuEnUt7K
KOlgWU3e88dYaO1/1ZYpVydTYcTIvUO+RXAujdJVPU2XRVdjqgytMuKFIwqsXCtD8K+n5kPyafIF
AfmOFWbLBc3bURoPqZ6rLr+3in8RamFayWBw9gZlnYuuiC3hX+NTF782uARh5N4saj4=
`pragma protect end_protected
