`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2016_05", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
rNMubEMaLbjnMIX9QN5TN/lMnoGIjbNK8YQQX1d28oacd5osi0sb89brEVK/7nmjzIQuu+dt3+fG
dtxIcQkcIDPEURPaHEdvKIgBGUMSL7giVxQ+WFA/nQRVziaAONG20XMFKDJH1pgnRglq5+JAgqjE
XS6kZW3g5q1FlxYNDl+1cPVHitBsTS7FAt3QvCgBRfvW/u4fOQ5Base5kEsyO577LLktE8JWYS3P
d539ceIt7W9EWa1pIl45STPWGT4lh4OX51UtiNuvOZTvlvWS0YglH14UcjuYk8LTtUQkWyb8tHO1
lgzmAoKnSzuJQRkecukCNlKGUd0iTkJj/HiCXQ==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
VJHIn/4IrWqGj0vqDUA3fAdVd2oAuw/BWcXO8bVexXLDKEyTAyt2+CNq0r3nr7eFZJ1lTMfisvoW
hNKtPbiPdBBjyFD23yd9do728D4YDv/bYZJtLuqa0FOYq/EMCPBEePJo6MqJVsijM4z8Vs/20/7a
ci9cgS/wuuLjWEnqJsk=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
c4rTbdyriJRELGCJ9ZFtBNQiJstRjbRhsw8m/S9KHJvcxcz32KE/H5F+Xtrdet753ydxD+K/HwJt
B9IaQBZwk580UO4xzqq+EtlyqmS1D+eZAzGUHYdkAJ1HycjsKGPHVMP4J7TV3ydjdDuw3UfJWyMI
lMBl1YwagQrrnSGGIP0=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3504)
`pragma protect data_block
xKMyvbI4QEWAS4f/8KWXvSasc5tnZN/Zs/9PDQ4AkMIMiWg49Lho/XtDzN6oaHKnWYL8RBKAfW9n
ah6KFKipqAN7M9+D6OtkEq7UgBAqv8PnD1qg+VNsJ/ZysjmOkceI2lk5ssrDv4iptEZNOBX4aN8u
Hc+Lk/Alm+70vgqRfpbKMFuBO25LBHUoIsCEebrgol3fIJHwVmQaI40NL/fqVJX2UDZR2k+uthsa
tbaIBP5m0hgx5WAWXIUhHu6lh1o8ZlioZU3850JaAdnutMCmIx48D5vDu3tXy1yylVgKEfU/PZy4
JV6aZTFw1GFGPBvoXZgxZI3DtzyRZWMz2NtWzSg5EcNDSBHPi8OGRglZXgdktWblS75qwm/cMxr8
BJpoDjdU9EQdRiAefYFCmiUxQuVIbJTghQX1ek0MKLnH+YqUpLABFC6XHuwV7OhqoShyktQd2YZx
B3hF+V+tGvMOSh15wEw29v9Z6eSVzJBB7hys4nXQC4ZwnWyZNTAJhTJNGfis3V54C26gIfeUc8Zh
qz3YW1oH7CUIEA5wtEMuW4GgxVfuzn/2ABtTMUNNAgOepyOpNQHB5h3jRd9GMkUHUpiAsVpwj8Xs
r3sK1WZ8f5ofauUR6nS0GZ4KUAqbMUsOvgMwg+Dj7PQL5CkTCtLg05GF4VH2KGW2oF6GzlCvFi+i
L1Dyo+Z+rkbfshWiRlPhzCB3bQBjVST0YMJ8HHMr6PZdNDEcF58UI9iThBOv6v9HSQK6pahT35BY
3aHMoImTY6NTHRQQfEd0FFAG3IhaHvPiLynBmk9J9QuG2MR6LtXn8anXyJZwLaUuivgr3s/MXRaa
ycuTVBhkoZotqoKqho0VhbaEfEW0Z7LveojufyzXXauFd5NxiHvtY7ZVyZnEBAGEETnL49xio7CF
AmZuhyxBO+cfkDVlkzb3js/+VbhK4PiBgn6ibnP6B40ywl962uxX9TkQQD6tbD10OypJx2Q4QZkK
O1XAloy0dPRCob/FaVI6PbWUSCgt+21wIjkYySz38ByvJSABqYsiVWM0hYqHV105AKQhjf9i70Er
QhbJLsiRN6k+PA2GiSXIXWV9GymINUan7DhQKekA8aqmyufjgthA+BKgCp4t9ozciCwIai6bDPjq
Xi83NNIbYzzVnVptVpvyVkIyxvH0HDzJsH/NiWNinQaoe+13O1gZWkFycVQv2uft/LOeBUDNeR8i
kouSGHMlmTZPTy4LewKKkQkZzaxxEkaJpyEFUuRRPJDnbNjGx5liBXYHI85jFPnQ+chihoI9MdnO
+TvQl1YqwBPpBKP4Zu/p1ldVDFFVc9g6BlMT5Z3gj2j6KSGqPMK4lVfA+4772Q0P0XmtIC28rR7i
4Bn4r1OnQW9pJe/Dh9xYgSmIgWeGJRI1Potrtymhm0vErSIxx2gDUzuK3RxLWgTkOw1d2vnze7Zx
r4U3o/PAUo3ak4obdm+qFYW0mBhpxkdYoU1JDUj286zIajUfN+W08Jofzys0Q0xtalZcL6ZrPw5k
WLrd4XC8Btj1UIp87CoDXwtWohucRW0LZ5/47/oG9vqxsAwCiLVTF3huRPBglNJxUh/j+X4+0Xo1
DqR7pgFSUwapJT9Fd+o68A+NCTIxP+sMxgJd5rU40glx/IATieSB6kL2CH4xHDOmTSJa1FTzc4/F
19bg00dXhoPfvm+kpmKNMUhzxtE1LZSyHJK4qeZg0E1z0S4Ok3K3srN6jaMe+1e1KpiFTcGiSrL8
iP0mzq93kPffrKv8Enfw/UrEUtcwusv+IhYtapmVNCgR6LUdBtwkKail/3W2CmPeBdb784F9uaVh
djgdkP0FwScMqaAeHMoEaSWp+K4elWzvO2i+qaTUOtn0L2kXJ4KcRfMBvOAyRUc8oxG/7SxgBl9C
wXHi6gGmaiAvdL/mKjgMAlsBef9ODNW1zc/qiZ8xGJ0wIqNLsFRrGEEYKVSZ7VjiOKGbR0dKLyVi
eGKljlpYQVW97NK9A3I6+gQ6ysal0kIn11RfIK99uc9rDLGK8GMR47tKCvcbL+UzA9woXJURMcOQ
NcUBG/knF75RVqWRix6/Gt+NRSUTTWWlywMREFii8o6YMEWdY4HpjmsCaulhd+uCljaqoYAGTWwl
J2r9OQcqgVDOp4LzM/sL/LVpLOUAGnceEj8PbtxQOwyDvs1e53NsVUJ8Qm+b9kmmgbkjNZwVZWtm
OIRHjBYRDdDv9/LE+kZ7rDl9Mew7M7pTJ/atSeR4LTA1LFSqoIof2EFZrqonsliG11nW3+YVRKX+
dIzNzafkugRJ4O9+Odt6fA337pc9Dpk9sBIlYahGqqZxsu9qDRlFO8+6E8qnf1rvWR4DiodJeJnl
eHHFk1/z/sYv+9ZgwnI8KbUtlsseh61Y+vRwi0rq8tQwAEN2FhJCKoshWz+FyCglEtCd4Qfh4Wdc
EXppylw2eJ7QTx4Vf3a+IddLps7gsgQlmwXE6NE1juibVDpDuKi1m8gfbRwNCM/Ghbt4QV+ENDBJ
xnkMcvDaK2mwcdYeJtnqPIp0KGBcI4ePcodzpbol9XV5+2lhndz1hZ+w3dz6a7HuDiXH1q+kXrID
36yJ4AULHatEU3sIYc48BLT1j6e78kqpYsbmGYVs7HczXXipJDnEXn44bOlKB9KOCmltIc4gnetH
PAg5zHf8KAnye1FmJzjowuF0WwfaSAvAeh5xM1xOTE/WAbcakQUh2ezWcWcBgQUO7wFQsZIz2vkZ
ujUVObD4vByqPGHudzvreB8A/eBciKgPEmkp1/sfPARuw6Wu4t+VxiUHWKi1cwBI8G+6+953RhbB
DRwHOY7WUVxWDvHCRc0LzZ6FemAjpwm+Zy6UIp9AXfI+nKXzQUhlJ6m2zsYMt1Ut51MBCGtnjeqc
xy5dB46scCQlIxoqCUv5NwtstB9Oie/DLE34W36sQUf2JpGVdFFa+Pvr0Sa/DEvFAhYRe65vI2Fx
MF6LzBNNK71zlZMeay82vrbkyDLiGmFsjJGs1otEwGIq9b8gTR1jk3UJ1/1LOIhKYn3K3gFqMVCS
ok72lITlkZQwAECZl0AP8644PjSrx+gPE4eZ2WFRcsw/DqoSBavX3aRkRfCUL9Pe5R5BhJhrCPcM
edoDT5kYpwW0hJh8ZVdD1t5Z7EeMxlGLd1MPyvVtblKuMYtqDEDWIkX8eveEIJ5R3hQvSaj/Vq8T
Cxq7eoFPdtZ78VFF6zKE+s57tx2TixIKkYUtj9DcnXqvO8C13muG9V6g7C6m/V3gBWL1ZzVrCbGp
xdQfOhGC6DQknvhR4u7/ZCtUH+v36792ZU5F7EpI+6mGmpBCmwgYUR5q/CWEFFC3lfKeSpby7NcL
72w/e2DWiAxAe2pgw8gmWhcOqIDJNcYJJbaWGaImNp7sQcnVfTomT3757Ew+pQIs5RbNxuJgNND9
tAlOVDiX9XfTSALsFkgoiH8I2r6wL9MYY5UkSyvQ/8QVR/Zax6Uxg+BOFe1VDVDrkNqnBtPrgBSq
VRhHd1CUkVMU7Bys3huoEooOSP5MPzI4ibVrxR0jLZXF9AJri1/NtJIUs9EqKOViwr9uCubUpGcD
9lXMjF/XgN74Pycg0Z2mMJ7n1OD8f5+r6SsuOekVKcq1S//3BmGM2HzFUSa3EzGWuqn8EsBeSf+N
dVSzDaIcTCTij/Wg8qDXBf1MscczD64hT4795/AhEki4EjlYz7CFh55qUXUA4o2vlm83dA9QuSWn
I14fvy1npGZ8+5lJL3EEH46Rf5hzUJk1DN/kzlXhVVBCl5i0fy+p5NO8Lg7c7LZmACMhUlG2FSDv
3Ja4AWtjtbhnsAOA+cpaoIhlrIWTEGgBRR4tWN8duymIMrA17J5nOatjaEGyLv/tG90t239pzLo5
PfiJVL4rZry10vvubJn3WZGYOWclta1V03vWaKEraM+rA1eLvFeG1jA8SamrA0MQhH//LbekCjvf
wcG8UU+rFpEr1MjPW8lnPY+uqdQdS0cgEZHOV3z6C0qnLxUK8BvCqpQcSl0sFqrp15dWmukA/+DQ
9paCgTvvHk57mB51qiB4UCgN87FM+Rt2lLAQWnUi2bKEW6lQn5RUAXISjqhsU7LFntRVg88fs18K
FSMm+E0Ge62FgEbwbgReghs9JC1ZP7s+hQoyzx1PItU3e2WNg7YI4EcXk0E2yMOS8/fEb3k1Wtlk
VCsRNMpNoq7D1P+3lohD1ujIhD3Ekpi4vm44qY6EQFUU5j4NbfdmSPEx2J1XgZE26/Ml7eKqYSVx
vZpYT9IfSVm5iX1Xa5npVcm3/g9kIUuaXe8doxNrQx/4QSjXz3SE3JqO24Xi/sAzzgqhBJD1pQZR
yYOBYalbDth503Acaj9DKYfIOcjzuOZ6dOICWxqrSctcqVEdEstt+TCkBPWczw2g3pXh3Xf/2sBX
/qSR2F04KxVO0ssx+ifxNv9U88xdshY1NGV6jkaVc2RCIFd4L/KP+tgQfi2sDtPsAkNwq/g1hodX
P/tDc5IoVixJk4MQhZBS1rcUd9RsgwvJsvAzOedjN+ru++hRf3DGtHVrvLQfkmQqmQ4bOM8T326r
VTSTEbVa8MJf/Va0diWyYaBrSoGyyscyDsdyynDDowWZUAMFOGp0cZQU29V7TWHBLKhBAMaHDdYn
gVrIvkmYdn/P4eMzGJQNUQgdYhlXAQx2yOrh
`pragma protect end_protected
