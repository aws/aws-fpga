`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
llwd395QfRJWTfSPDCrAHuhWWTPniQWFOW8UR8u/W64JpK5hkB+w4Zz+P+YJU8egvPWFRyxeg9rI
iTpER5gxbVnLHytn03ybFyjCvfA+2AELYRkwBC0UCMd+sTF+FpgENl/OYE+66EXlKF23YvKa/44P
6R+q9BD3TUOXIqgc9OglvBgliH+RY7lt42Ek3aa98GGQmO/1KYBZKOEfjhR7H7hQiAKCvvE1y/AO
XmkRWc+WsIcx6N7WV0etnoQW4A1iaws+PSJLSsu3ybVfz8LLbN5mVY0XwK3CPqBZTOh707GTC1mF
joBwUQpUFiCvonSceSxefeo+2drqyMJcOtEqZQ==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
VlNbiMjL/1fAkSFeVBcX+zeIQ21vBpLlfbcqZmvsgh/fvHC7XkwaDOrO4h3bg/GoSXVm4idORYBO
V6wa0lZJPf8KDwmL4SQAWVC3vNlt51N8OnuAQml8JK595NmsFABLVBwcwzoDwKIBHZpOeanEOi5Z
+LJST2U2ZAD01p9I4vU=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
UJqvVCIjAT2LkpODpdV3VCIVWaPQasV+bAsRSczmzn6hwW+9V77u33bupAXaMkNQQRfQTkFtQBKx
pXyhYz8/g3N2mjwP6EoViMddGQrcgP6uco+xVPq1tv3v5rRC/nTdK6XNRSLBJyIHWQQxNY85rzw7
0xxALMwY9w/Sy2zS6EU=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12128)
`pragma protect data_block
iJJhL47M0d6KM61F0qW30DwbflFCrOSZQ8N/ufPKYgzyj9lvPo/1uYIfYukeJc12bwFXFaLclCqA
UMx6r2PmVyFWie7U3mw6EdGsWgc3TeF9C1OAZUE86+1k0CL0DfSOGd8w1scHxl7ah1AfaYz3FfWk
tVATYIVV+rtTRVAdwJ1WGSgs1VewQS3MwiWWwhTFOFO/FDLOtQe0xgOl5QOQOZWBD5VsZUbUjifF
TlwHav8cEOHJija6652DHKu+XiQYf0E0W/JCbfpI2eCMkJZJYfFtyZGgT4RuxwFjVKdkvF0tOD/g
K4VOboCDBlNiZ9OkNbEK6X4E7ND7rzz0XuDrQIO55XsuapZQN0ABCB/r5c+y+9hIqjPatSygqywl
peuHzQooMs2RZq7WkZGnamvhq4BzYdP1Y2kDNvJgWInQy4OggJ3UJU3IxWBPd537SVl6g/qYk8/X
uEmN2SmijL+EVfJt2QxYY+68nfCN/R9jT2W9baR4Ii+b3ppR6yXiEhPnNENmjNLfjOYK71sF5Fq1
fEpL4viskhLWFtrhDq8MHvO2A1dt0Z1MbHUGJ8MRpj5YCkqiDQory97C1krXMdvYeyzbYdgc8Vu4
MYmk8ToW24O3rOSsCLBuHDczuQdHRXZ/nDiKvFOY8iaM0VV3pznQIBCho9pQJST/a0OIzLCpwQNC
UvEsfvMMq7gzcJPfj+0ydrTu0A+Hz8GShhh6SqaZJj++UBf2KkuSUYnKlC3xl8iNlHqZ12P/DoNn
tms3QcVh36BBi7g383R1eQ4pTJoW3sFU8cK2ymo5Q7FWC1xUDFSptJmT73K0MO/buo9l4BL+kjVV
szonbq3tFZ5OAZ9Ey825tfMbdEWpVluIuwQbb/5l0e1n2/tF6tOwn+JRyZVVPIViA3Le/5topZFx
8Sdhgp0gPj+hb6PEDPqadfFc3iZFpCMH0CKqypuCFrhv/suCuOwJCNR+QCWs+FSn8mDDWXmS6Ef/
enT9FEBh8nOtdQOE6SgZnPYEF7qToLvc02ZFIIOWn9Swi4uo4YSPKi/UkVxnLkviTOMSAaxJLkOm
CKjP2wq+fY/+jH4Z1EHSq46tdKluwbhXr3nNgRKH3KqmTgF/+e6EBpwIRw6LeNkQIiB9s/bQ+Qjr
UAaSgKPQjJGYO593MRHjKJRy8CjX+zzJmLk2epfEC5RNrfNxYA6DoUvWDmp/7dRt1vDiCHTb/IfW
TtGOhq1kpW2g5Tu/o+pndGXNPJm8yOKhWc/pqT9n/LTMsnC5v/jiOunzz6Ve5QQSlBARAld4ap/D
M7VBb0tceOBF6beDIx6jhPYJKc2Tfo1sGcodhbjJ95yQgJWYnHG7TlNl144Nwe9yjfHzNiUvuw57
etVyZQ+HatyyvRMssq79tL0JD8ea+VkQrdY4DnprdFL90QKphGJUB3rlSuegp3g3hVutuN7p/Pzd
J8cLvLHvahU2YnGbjiZVGz1Y2TgP5rX9fzOgoZGGFzPKmf0tCjyq1tUyJm8WtiakGV8D0ybhhWmS
yNKNN59GV7rgRfO6BkMcMGppbkihHn/07HY0IY5WldkCL74JZ9nfK49UIS6LEzC127q0WAUlZiAg
EPAXcjxyQHcips3OuFXi/OMnEY7QiWslCSIQ6yYPRr0/aK1tnUcPF5FWzuKMGKcf8RKqkCJw4TR2
fw5KNvf+plZgHJlmsuO78eRpUZmVwBBLxz30Ff4Vm1PS5YbDgg1rHN+AYljri5rbsfQphgi9UA/u
ULJAJ9QdtSA+uBx1Zmz7i6cb8Or1XkB7nX/Ho1Jbb9Fjlitx1xngAW6Gnu4co/2VdSM2IF0pF6Bl
jcCcSIpXlGe9snb9Zmhy/OBQBm+2OID+HEmpEJjIbK1HWg1dadOQnOTjmc/kxEbyx8kjAXrGUrFJ
y50E+LHySJZOr+ninf/ijIIIONHKiG5nNNwpeoORQJbhVMox6SPclQycuo6NQl7R/NLKIJqUeWTq
h84Q+SqsqvCBIZGE88IrP1WQYGUiVMAg0HhM8/QXVh24A/s1mOPApcD7KJxzGyc0WtZmiB5J/JRH
II4+LFdwxLrwLF/Rt/OaE+vWpo+nhDO5ZYSRvYb35O79F8izwdgW/h0kAue9kDSjFUTb+oEzwFXO
YoziVrzKeJ0kWs2YM2wrlv1tlH4JiUG0DIolZO3arpeZxVfZ6UVmDUTGvu4RxSD9eymO6Iqbf8/s
T8mZElYwIvvXwcPaJz5+1Ip3u6tIEtk4qa2V/bO4IzxfFCGHg7HEUzovohot4ywt4UB4ExpJ/Xa9
a6uFkImQb8TDw3e2lcmWLR9UbwH11V4gass9t9CLuw42hlxPol+FS/gSFQtdPey6cdiEdo/2j/Oa
VuNaB5k62iNfzbYODEYEPsNEoyNSfA58/hsfcATdkFoewzdSsTTBtLUHin/CcDRToDusqwmSY4EK
6Rd/Ku1he9RKhPMjh5jZIOckZivYPcPPN0Y3qFEfd2oEJxRcdZ+JALjlHWMLKbw0U69IiNo4bL6s
20RphahdubWcxATr3rCXtt4++8vMe6nv7R3MSvkH6H2nxjVFqNvl7QSTOvKMRI+/OMqz3GGf2R3u
0+YGmKwIb547F8HpTM3TSLbewMjy3lGNflabbdMoRoVVzSTLkaoCjmV3LTFC1/ngco924W9hk7JR
1pS1sNqfdIVq82a1IWVnP5PxInXJ/vy2AywI0iHQ9FJZuKkYIPN5jCAk/WKJfnG2dnCiP2R15Teu
V7bdfiWJF2r70CCiBC89zbfifADDzRaVfnrxjEWclJG4oegyuWnoIg9UTHvexYizXeuSy5cM6qZY
3ZOEUWg8p6DBXllD1U3St7Oaq0qTrLWK80TaZOz10N5dfB3eUDEMAYKvvyL8LIxZ6YioWtkFQ+/t
N+3l5+NbHOQGDbj52ErLI3idKqt/REBGZJbgizHLx0qzsKCbV25HtpPscN0JSEARTb+dPp/aRJbC
TQdaSCG206zE2hqBHYdESSD4zmVxS7UeWffGIzDgOcls4TOLE6xlACa69jKnNwLKGzp5zMsLTTwR
YxRcxafFpwfMl5dBuH0teOzy5gSAISeRPMxMA/Je4LgOcjMB6wnJGqdWIQCGDxKSW2A9UK8OWWxb
A6gyGxmPZVpTUeZ/A4YShmi9Pv9duQyT7HropuL3gpKrhPYl0dFv5o3LTWrmHMT03A4vB8eHN9B6
yVVWQDkesi2635Lc4/liy9EpH8gMjcfMo6QE/IVoQmDI/bp/6lZ33UCltGy0e94Lu87rYwLmKesf
wR+HISU4QKSV7clrkTXQR7ey22Ybhy+MyOwC8NHqHBwx5WKd9xUYbEx8npxH0W9/rv8pxSnRIuwm
3pLTogmE5r7+iAVKbu2hru5ozsKt4fzR4SWwgZSlyQRku8Wt6cETSnEopKIOTJBN6+i9tOxUtwzP
ABOoXKT9bXj6/2Mk3RDdfPbe9NDuGYnoxIVQn8/b2leWIFwWS3U3eS+xUFjAmWxpg0+uj4pJANV/
JfcnsX0QQg9HjZ39VyCJzQN15PTCno+jzooPRhXll6gE/m6//E7UuR0pKlI1S8cZ8rz8cbI4W6Fv
cXgsDX2zNsk2of3ZZFNE5pOmBQChMMp5UhhX1jBRzroK18B/0ZulmBLptj0ClHtwPWnmi/59GT3I
n2eZEmVkvR8X9OYUgUmUvm6Svd09nb97Wpsa7Smk0NR+BcF76zupgN81UfYp6PsOWRxTBda98dqb
3RTbhM/slDVMxtoQ4uCp0UlnuRaSeOn4uGQqXVqy51lKlmK/3pflEBLpJoOSlIAlReLTGwzliDSh
BXH3DmuLl1fW06DY8n4clhFJr2vFA/ndy8b6Wj3JAZsyWlrzNHRm8//0SCWP/45MIhFsTn7cxPo2
v80R+V45KCYOz/RC+1eYo6oSdfVTWGmqvI84TsSGHDH44GmzieVfE78a6YO+HJ+oq5csqGlJ2+Ng
1ru8DY6yxONlesmWyyh2+mdPbQRCvGMawy1fe3pR4ewz9WNsp9C2raOB29EfvUvNcMxOLRo03qaq
5Tg9ZBnO2j08XJWk3iCG7nF3RA5f5l6QlxdSqX5PQvwnnKVHJpI11YAZOsReIe5ZJsj3pUBfOiyJ
emOvtQrakRyE+RrCWJnYxaq2ItBLCTBLx8hSqaua6BmWNJAZ7SFT8v2ttAV2CN8ZUciDKRTi0yME
rUIvYsXCHaAKDlo4ozfMK3OvbnAw/OLdcUY07Ax2LN75S9oZHU0ILRGNewiO9FwYzrhwi67excuu
I31+BAbUAQGIwdqWPjDAO/9zoJfYWEPbspWWGQpisEbJHqJ9HLUCoe/cE3nnnUdjrFl/bit/ivF3
7RGDtt8e7Eb/l9xTdFmiwcHR5rCpzpg1PYnZ/kX4auXTRJtjXQ+GLuktp/yEIH0LnzZhMck/+nE/
U2zuE3YkQoFZlk4eBLpNOp3tE7GeR0Ht3DetGTk2K3+oTnza1JZgeO5hz9rHrUiz5R0xWifv9kp6
ZRvcjOGwubSeS5ChKNNxh1Ty+02zDhEK9LHve5cqRoj9JnWVj5NxHHgU1IhgyzyHPOa2w8u+mNGA
uuPlT2tEtnrN+UgEfFX1hAFdAnBz1qfXAVf4D9oDMroVSmup5WSoXdCKpCglXwMlUfvRMM+wMcc2
9McltAVWp8HA6w7rKhMEhD+kNQcuvqmdbdeZdMGeuI3iyTv66DbQy59wp42T6wY/wVpONKn+3HyJ
UCtyhPozWi2ROXpNP9ZZURjHnI7JHRGuyGfZ20l+ETkFvBsR2eTb/XburzO+DCR7EAmZcF2mzwrR
sWpBI7GNfsKQBfY1ga0wrrIWoekafSuvHS+QMtgM5UZpNFW6Dxgg7f0zC41m6GH0AsQ/HN3khIJP
hW4gvcJfkiymCo8yEzKjh95NsN4+x5TNTsO7Z4Ghjq4+dimnIh4MRJPfxDEJTYsX9Da95z1f5g77
yAQpv/I11JqR61EWUXri3tGvlJQR/v3p+lHsHk+EEmGepbm+GRfgVPGoOD30w6ZjylaEkiQepIr1
oWlT76Y7S6iUl6+/D2PV+Xr2xcc+XmbIXK9T9MAMbbvS7uUCwqWusFfAzi/mDVu9hoKu4c3I/u3S
hic1PDfNsN5w6bQPPuYCQiVxMCCP60qAXvcQVylHDNQljZq3UE8wDYWK/FEJBwNXIK47cuYIAD1g
QYyLh0pOTSe+fppZcSh9hsRvSgBNl9u4aA06wS2nP+9F3y1NTlEM8z218ZKfNvnWAj8neOxf7rDW
IIqMR0iwrz9AhrZpoaJc1DajmAFlJu6Ei0PI/uSWbuUwtw5sfDjvIAE2xwFqHC482H3duygHP6VE
Z6sBGYQMwtddFmhxxhzpQrKtuDrOxL8oS5vBn4NGG6gvFDd95tHofsyDusmUSEX902TkLyROIel0
3XCrf5lbbfsGZpnQD0m+8PoK8lm7H8LqkBDY+1Eum04TFQHSvrEbQXykwFhQxM4Jnqhw8QJX8uz+
Id9F9jasy/cDoh/C8uxBHL1lAtJ+JpvmZIqIbd638emKQpfgVJNcni7h2FYGvM7H98P2JQ9oKp07
/0fFhVgCR8v9lbyEP9VjGdyz4TBeDYBECiD/xbqah9yNobhYk+GsdbX22j1ywVk8gN7Icy8vh1eo
Fg4MEsV4U8hkEfkeTw0tZyQWyFL2JEad5KSXYpJMisodOnEflX1NN30myywKkQpbK16zDWneVNRn
NEL8GkmXRsNo8ygofrd5rcIDQ0cZ+lbNx6HzRallwq3C2Uj4IGUJ6P3jHnSwZwnKstwq5lWlXaOP
rVinHjHaYC20IP0ykoFP0+x6DyINXBv52+0NALZLbRzgjty4i96bOeCeKSz1LxQfossDilib4lZs
/iUY8CgdfBJLPMVpVwB/+u8bB5MT24UDJiVIHJvcW8HOzUq+2LMaguM0ag8ZBkYZx/IRuLNlFzCg
vHJw7IJHRGRWHp28PBhUhBCiMi5+MM+wgyGb41SjOWBzKTbzJYnbFdIW8srksVu7vgHLBA9efrfy
D0Car847hfanU/tJexkw0xzPn44A7ByZJfw/IiesKe/aAqebMutYSq9XjlVvkvzsA6yLRWgRylDM
itfoghY5ACUlUkPQMzdkMITkR2ilPZr/X0p4bh41DeNSavs2E4gh8StbnsfsX8is9mOk2/T26deN
2AlZnHQpylZ7ua/gDKQt3coAWtc+A1At/Y3IUdEAopzMwvHS8828h8GV+yQYL75LEwuc7T6rOCFP
XaU0Jeet3RB/SUqHVMdsEbZBCCoONLSUzAOmNMazDWaelNVG1zCSTyvYM1+GitnHtDjAL200F4Hb
m2PGYSw93HUWOQLlWHyGY7MQrK058Fauoc9mpy178nMvYa/YnfPWSTQQQOMvCGXtjk6rIGH9I0kp
sS7GvpI8KLbQ2H+IoYarsKjeiAPF+Y4DDwS0NlKPSuuImRxHU51TAx+wy6xegANilx3Qb/txE/pU
01x3F+ag984NW7Px6+V4RFZMzHdWrT3iYfcDfX7FcUOlqXxi0/eancS641ZPjQBq8zK1AVn+2RlI
j4+5qrXByQh7PUmjeh54D1HH6+SRBzRje3FzlmIoU0MUfzf1zjdDqieE3l7eCYUvbjVI+XWl4Sao
tdSDgF6bxxliZgtlYYgeywVBtfnb4NC2dEKoU/OuTH+7SNqvaKS/+tg4RELedkd/oq4MWwvnLvUA
2jTr926fNuBzyFJ3fZLezacDYPSPjffCxz3PtJgBdImoeyp8ru+ayYTfjA3lH6ajkb+H+RsLyvz5
I4PntUuNxfisHqzNFa70l1s+YG78Su33GgST5E34lssoV4I7Y6L6e5JDTFMv4M4nXbGxMmUt5mcW
aXJMU6ftwNT3eDHBA7/DAFoSTZAKA9XtT+AZWZmKeq6A00A6dSx5X/du6zlEeX9dxQtKKd1qf0lT
i9ogG+iCJlA/Hm62W9R3KCz/SgOuYOires9YeqLO2ecNo7XC85pgvaEugjm24Z73lmqcPUD3ZJ70
6igHjXUFfM+V7G8D4Mt6mULcAt97YBZrCMyXj6t6Rm9kuz8+jpEgwfH39xIm6VUSbzZc1C9gPz03
egKrsquZ4+0l6gv9bXzDOFY686sWGN+BC7VnQMeisvlkVYGJGu8AWcUYAwX8QGRvUxeX8lmuEl7O
nfYLh7HSSPoiXnEdB+QM9/SjfEq8gaV7BFWIJfXtTK2sk3SxkFNofGoqjGdVc62t5R//TrzPS35P
0HAmG/ikZCFtoyQm7dBiICPRXC+P0tBXI6d6wlEqH8KHioP+C3kyT7wPvTcdFuUJKF1bI69xJD8/
dJeSZ4KplV25PuKmv3OnHxqX9DY/PQlZOCJOafEc4ELLQkYVsq6XlkUa+NZ64AoxUhkXiSUr4qOn
0R2wQ1VcmqG0JKKyL+tT/zVDNCtIa9+xj+CCJflVWyn3hAg0rAu/thWBS/i4L9B6oESsD5eTb2B5
y1Wmcn20z68fES2iuhnPVVqZIoy21YiQiWYC8fJ44xV8eXE1PDf76q/zHOEh2Mr01gj2DHHp7MeM
RNkfEIQVGxKBmxcWPupO+BeyJ5qFKZ4dHtc8MLA0N0+tSKhG2jUVeUn8mFAb9rOPI4jtEi26CPE3
hx2Zip6OA5SgpPiWXFOolCxkQzEpZ7AF+7udDNSn3dFGE69MyveI79EBBhywhyRk7d8GAEQ+OReR
O8gC8bt5NSCx3uByy6BeCivQ6fHdSZpOTTrCRmNjy1CX/CqRjijkF0x/6jkzLXhqSgXvFjWlngdD
ZZPX7e3VYfrlLaE5I7wPdOI4c4JgC8UmNQ+v2qkYKTUbXmfhcwVqSBaSYM9TY6TrPp64veu+LuYO
zOh5cT9iTkKyqWUVx90voYEsJWiNLEsB/tQJ8ATBBNZZMjFZ7RVc4m9CvmvBZpSSnkW4it0cVaPQ
mSBCMa6qDEFOz+5B7znCwZ6odzqSA8Elc3TbTX+ui436z8RfzD+14lpgm5Dub2V1fLwF+5HFPWYQ
WiZz2RUizmokIuDHmslbfDq+vYDrBcV1cbZp4LFuwKgPaha+4HJpDyTJ0EXXqhMxXUDAAKom8Pbe
WDhrrD/ygDUfliL1SKbBkokgqzAawLAwJysJtBkxIBVx72eSVy3BL6Nd46rNHIwKioDcqTMxB32L
7hgUVrpOlV+TM8EdcLCKyfXYmVKLffqWP5d4NedTlRW0EWPCff5BuMNEw5+Qp8z21sJo3XCXPY0H
6eQkUKoeSgi83mm8qGfiWgn5Oyn+otoNsttrOe2xEHzK0olhc+0nHJPtFFNps/hauuak8UEl22Q3
9sNmZZxyh0r//bcTSneKKfwYepji+VamWLLMKKhSB7bp1c4FwLL5UDm98DY2nzrJnKtC0t9Mi3s7
csbxIS7eczbIIIPDt9DGgT4aTZj1s1b4RqLnBXBIptcbHuiwCkjB0wvabOR62Y9/LrTpH6tLYVQK
iaWMp//9qOIoI7yMs5O2cJQMdkSISvOBbYbuZSRrhM/h+pBEpK7VunQ1+fhGb9cqM6XdhoGba2t7
XaEDs8bkQQbn7mCo2ybsEvfUF7Wy2sVTuQMJwSYO5sLHXdXRU+G5Gx4jmoOSOZKwyKNjFwrp/GrY
Et+J7WFTNV/bHCpmRowEZ2XS3WZIH8+xnNISxMR3ox8ovTU4ZDcoyYDcETmgDC/HGFDAWNAIKraI
FMfNsZVT4ghRuqrefZg7oy/VR7mdLFuktBENxL2e9Fqqln+9mjtNT1xTw6PUhkEwjfZL0n+6IF71
YdMaByF0V+I279fkO1Vikl4fxR1xybcXo1R3F0069BCyzPpOie0pb2/lTM6W8x44qCFL7UVZL/ia
AAbYuWsJhKtFigcr3Yjjahi+8JA62DWY8JruNvBD3OaFKBu9iPb4kaoocPr7GnsTFcDqMj6wgrOh
+hsOJ0elE+uGyf+noO7A3p80bIHQ6sM0YsKmmryZRcqzakWwFn4cWnWbBIfOQkaww9NxCZAFOM+M
KMkBT8c5G93UzJiB5lIwCoWGCUcdIBOcrafeUS2EB0rHr9xrLSERu7gkb1iMuNbmJP6MIBLIc4fi
Wp28AqYZss21CDT/GcFmRPL8b6WC86qLXxTyvw/Twq7E7ksk6XSiLm4AAI4wZQx0+E/4O6HpzhIt
+0N6pIv0M1Lg1QtcQYwngsbkXWcM47PZo25QF5uyR5goMvlKW/lK3mOTAv96c9yWhkb6ivxsNRTc
wggqJcDv6S94qRuQgW2TNddCh1u7LHW4XDB+LMTK0nWem5+OBPkXhPeLjtYuktZFYa1LdCTU72ys
GVciMNCg67N99Vti0MZyo3KWxxRcBDMESRxtN2aj/2LSQ4PZVIxmUJSfwpHwKc7GXvhT21Hs+A6o
F3bLtwbJrJK8EKHUTmMIrw2bJwcwrbqWGMGdzsGxXZau+vq4CK/RCEDd+BSz8tNO/E6CZzzVJnIY
jpK74ysWphEXTvR1u+5eUaEltS+8uoPJhro/jFdJRBXAqjAS6vJH51z43GOZEY5I9emTg0zCSGqB
3q7QNkoJ23l2DHhulWVcf8KxnxolXdl9RgPBOc/PIbIAv1vinuTV7kIYg7zs+B1kbgYZd0Knh5lA
NIog107Di0YZpouUJiS5N6BdufTsNOQal1N8k0lAnp9wKd8fL1GTPW3ElSvzrefollRQQ+H9/IxX
0IN+sPtUA2L6KplUAbppvWniCg+uFHIoSxpQICU34z/0O1AmK/FfgXuzDcTYQCpRTXj9uDRyw5Nl
+OPfz37TPALhv4KsSjTtQDY0pT5cXWZc3tlSFOS8JMz9UfOXjG7cdHn4+9wPAv+pPOMwV0IA2gxN
pPQl3uyHeprMF8Gwe36mq5brXooNZaH/NLWGHYg3GvVFqfYJDCemDFd/UGvlYQR/lS6sZyUiO0Z+
5XCmezfBUxfiLKk4jbXT1dX/IvSxpNeEZWxK52F6ucPF9UvsBV/yN7/kDX+gcZ+XAXl9NbPdp7nH
ujAE0iNuCnDBgu+XZUv3Zk40NEbVT0JQId7PgLY76+slJCITbvSu7mZHetQN2nwMK0T+XYMmwSMq
W5r7tZh2HmLrbnp8L01YIXqm0e0pNnC/VX1z3AWEciddVlDP3t2aC16JcEMTujtwpJRVeiCGKvtD
3TH+l94TZVYcnyAPFxfLi/XBD1leb8sX/0ibTd3ocldEdwWluIUYYg5tdnANmTqh+kIHoBbYvI7e
Y5DCQ+PYdT2vHnfGI/LrpKY8br/+O/EgfPN/vkA62seGTL0A/aFmyvWHpkbcwGqDt+33M23EvpIx
79W7D9rfRkD7v9xW7+v0aZHFIt9yOLN+AC0cqjjehBJnoWwR+PVXH1bgBdyYj5DO9GIFKO0dKnBt
zNwuNWrOuFfuvEwUAGSOsqJGSFddwc7us/N5f/yqSdPjJRnmTglvUMtQtCxHt88TUT92Q7w+t6eQ
O+sdKB4qvNBFHb6GeRNpBbxBKIzH3Hl/2ziMnZtrsbfOTXNTRKhu68DOcXnv1RXbbYfP800CN8Gm
29dVW+1LIomgO8V4fbZXi0XI7woNoPP2gkqg5zKuC54lnX0/YBJ23EFgZdmie/wJ+yq6DVWyZ/f8
eXLJqvtohf0Q7EgdXKx3+9rQ0yjIMOoPgxroOtBu2/VrmK1EZNBxMBN5q1qzkt6MCVWFYigR2KBR
diH+4ekHESB29EVCDbjrTzcHRnfnMn8Xc3TLtMRx9h2E3bgp+TLiHBXimn0k3xAw828HC48y1t+C
eiyGKcxzXbxjSNwyxI0XseOZnLBeNKpYLVD+frhtXjhcZd1cf81LhWxLUJQBfndofqioohO4UoaV
etr33VxCRD1PhfOgQiUDIIbhhqEOpV9FfCHhfDqtVO0u4FKT09PuS45YBm9cjUu4LOz/wgsFHknN
1k+gsxfGbuiVr07g2KAP12aVFMuLaZtkr7O6jDFsJcoa6uKHaBGwteh5hT+pKqGivsOj3+3RSU+0
krdRQbTx6dxGedARfRspo757bi38o9qhH5DoxmTkgmXdxmjhNcB4NGa2nd8zqxvU2z+LngMf3zYn
Y1dqld/HQKCw3TxYGzzmHjLJr++CMsWqWq+mC2bXULU920rPQlgIg81kv47K4VxyZPERLBlKC7Cu
8M0pkDlj2alv9NYtz0B6nIKpEwthojUE27LHgISlfPJQnTjQgPXTuS+SRND0XLXi9IBa0TDsC6tY
EeiM2fqkqDfaxeBuAlgZXnpIj8ToTMhmo7npOrPPnqg6FwoB8DpzO6Ja5UaKCPObhfNhu04r4wQG
40IYDCBN1raPYpHOPHbar0XNnqXzSi944zQY0H4IjuemxhNsYwIcpKYmFDibNDziWb9HRgOkpLca
mZyA5M0yfm48hvKJ+RB+J62OYDG/rog+U+3UnTI8pCborxBkXgFbIhZH+Zi2RIoR1Busy3/re3LL
aOnEPBvKb3e73LE7USLjrtsBcffjDG4eQHde+eaAPc+ViaPRIgWTMOjbkTSckrh3wL6BCgMPJQM/
0xRw6jPIaNk3LDCbbe1Y+kv3d3P/Q7Rza4K5PHVZ4pGR7TXkJKvRbR6LZENgyrv/tyyF0er7Upf4
C39JiahLOBcCKtF9XIpbeEIn6cK7VY9RyM8nLWK9hQXjEmNOeqJH61HShd9dyCyTKEuiBQIUQiff
A/GuzB1+UbZ9VnWSoDXvUxJV0xiyvSTSz6cZMhGKIAQUaXFX9Lb7JBfdCAsO+0uitTqMEj0Cn5C8
o9CpB+zdK08VrSQWq9O1HuDs2PqF+yA9xtTaqBC23H4ImS8zzjl5bas9K6luIqocIbJ6AtJaoGAN
fJpQhYoEnM80N/GgVmXq98Xowkp+AvmcxzdSWPhAqJBMhkHnUaelxOjsByeWhmdr1hph8mbsKaZX
HVJFjG0MqJHpmYfXrgRvr2NSZ3c0808twou7AkpfLxkkx8U1vRxhrtCkaeMK8SsdVPWJg0cyMdEn
Ug4rz+9zPsIJ2om8dvNa14OARW3GRpoMAfN41N6XEVpmFyCJtsslqoXoSeTWv66flXsHxt5F1B/U
89hReIl8+fO3NibbbUSMzwTrA5gEZ7m6Ft60x1rylpOpOxQWfDtmrB/Ie+zPRs3UAjgR5F5GyZ+T
Ut4TdNp3IS2Glgfy8JweLmFi/YhZn2Xt9HA8YEce5XcrdM6xrp+FGpVgRcyXViTtXxI3LOaV0Ide
jBUwNUdbgkv5VOh8UMjAjI19k4XEFaTWtJI4VuOQhIrn0tg4tHHL8svk+/PPPkfW7HguMQVKrcMs
mzqYZb3M1mbgNF/fVFfOft+9pCgcPwonvq7t2u9iYy9mopCKjtoGbmi6UJpM8JJGmKsHZTZSoblr
5EYPFZAvSpXRH0lN69e2AfbcxAKCUpn/sZINUnFG5D/qua/ajF7B7G1nmFqpPS3YB6Gr22p6dbXw
MnRwW/S1hFm68nTkv4hS/KfR+vbvRqfaYLbVag6C2Xurb0Njsc2OFM99NoDWgaLyEuHpcCpXTeRa
j5QE4TDHEoMy1P3xAsCPxeJNize5j1ArQCweGi8Dh0kdpVY1TtTAkehxLi6ko0Lh4oPTyCKKvGSx
mGfFFvZOcCzjISNSf1huEiGup3Hkos4T7TgP1Us9XbdO5kRMLtfgoa8GLzIDsx6TcLqssotFrAsT
c/2g5yIgqs1Td4LvC90ryW0GxBOnDC9XrwEF07jziWefSYYeyJHjeXNcUbIfftkTPnBti/yksDmq
cERqTIBhxTk2ZbiPiCB+so+eKm4xElW8R+U+xy9x2TbO5GGRlPvz1P6gziA7BugjASxBM4Iy1dub
2xAUemCFhwKYHF+YaikSUT8irlGmOyVdP+9qtgOZJ185y5LnKVk4K2zV6/7yVGrWlGn1i2l0kJPx
rlXrJ58h8dgtv9U66cbz4/+PlxAbKz0jEVOG4zqVcyLOr9GNaL79CGrt4vIzb1G0XC/BLyZMeYR1
S6KXBjpr+96eCiRLHniYksuEK1MlHRd+Tzq+m7w0kXUsFwfxG9/L7PwfR1p7jGk0Glp8FW+hBjC6
jcTAIh3lyF+AWVSuu+FjgjIpKW4tAoUdpxODMKxxyBhl6GUG+A0Ok3fQ0bOwttVaT7wJxptsZN0C
ykn6yaA+bEo3MLhGUm2I5ttQkq3ciwXNdb//JG+XjQv+6RwT0OLKRKVUQ7ZXkCYOZNVh6u0UXsM7
OD1Gst1elDn2kOWr1Addmi6JF+dhZ/qUEJuP/7MFPaKn7ViX1vJ1LuuBk08664MukEbxNFtgMKrC
FF1/yr712zuecJXQycGOuD6VKnUDL+3SyaeO0Wl0//SsopkgbsvK+hP6vqxuN5gQMh0/BFH/KBHR
Eo/GA5cJ+hhqlhxZiuqh2bxff3Wb4QXIHgvdrN+YgKzqQxEhpbaPOVNlOZs9uFSWjMNOY3F7oeJl
ijH9QtcP5vmuspSoGU00MJXJDwOL1Nvp7dwtB2mD1qabqWm3K7/eCvvgl0cxo6XC33vspM1Jfa5Z
wSY0Y1btL+dlG0TSJKijSnx3PyOzC2a67pv880HivaokJvA3OrNy3cFOpXCxIQa2BAWvJofybYFY
+Qsk9jceLk/M26bu1n2yhdhcruG+TI9G/xIa3N1bIB8wbnCI/PMvrLjJb+3Ksy4QL3Y/mbUo8LFl
pZtgKifSSc3OzBl8TsS5rnJ5bGmMNXjAHz24OkdGHNo08SP/3dDXzOuzXsqqTwKmU1j9WK+E0HsL
X7w6eMBvO4UIyBrHdED67GMGN9b7y0/bBp12M4S9GeVJ2XpGR5x2UmXkTPINeAtiPs0kGDCyGQ8d
7h3cnVQOBMd4sSWEzsRT3WQf53IBzzH81xYqEZVAtnMiTkrRb3FAx8c9+jGoOy9SKeq3mgrBxOa5
zAohDSTB+EwAHyiA6a29uYmGexpUC9yXoalAgJRusQ16XenF8uIeVEh9ETlODcemzjZpmZDPZoQi
6SZHd22IzvwePnZpHyLxpkGTnSyJjb1kw2R1gU+9sUzJNiib8R4E3KOPFpXSHZGx4/Z58fzjPTSo
yxH7Biwt4Xgc03RyRYymAm0pSFy1m/jkmGl8TPlEnZpMAILIJKlhG/Rk+FL42msbop3pWS0oQu+W
LSiRJ7bKL6/4ogW34Mdh1Tsy/t92WxuieMCf2HTcZ0l8yoneJykUhP+tt+DKuedft5uEG9fxI0e9
5Kd+e3k+l+ohFJeWKA0ZNsX+j1gN38c9j0hQKxByEPviash1c1PhnG87IMuuCeXmdXkbhfqkPPo6
N4SX1zxPiI7Sduxbc2bZ5au8VBD+pZsZMvucOMP+6dfmchiLY8v20DWeA9+ShCo52PF5Z5uy+WpD
jJCQpHzaNdByT9Z/6DxI37lJZURnGVq4OY5uQqt4JvTWcU+AeR3BDo5hYM87cFRonCchRIG22/Yk
ZHJYe3CmYObdN24RqGTJERCaIGuroxaYL9E0ZKhEM+xCCZ/wVMApZjheJ4F4f/Lpc1CnJtMcMasN
MjHlqe7FVzSE4iV+uEoIrBgvZVZjIJ3Ho6STEBVtftodp2HJPXlnB6U8zwNpGZAVUYU3STiXuXRh
7PbNsZXwM5DqR0qeNlnYmxS0sGyGIuAnnHyzkYblx/cOi1axR528eKmrgpjD2bEo9+hNZPQPCZ1O
SCFXOvhBBTctfKDl1/iKzsQbKkHFcrPF7t9nbcMbIynGEk3PVGMdcdnfTeCrOYc9HByPyrdRVZCS
G8JILJUUPSjVW1HhzEBnuRPdp3qyXM/TiasggY3FOIPGDpOWUhL6eyvThhlFohgQLS1JzB5NLeZA
CSn9R7TFcpze74/cwOU26zyTcQz159bRz7TzMIII/YRkjSySzwuDss4PfikyQvnRXoqXHjiFTxmY
VeirPstCFvYd8r4iPOSwWjZ0XgaGvQnr9CmmKz7mCttIfGso5O2/pTTDnX+yFhBQCQmyKG8q1rdU
d8Cm4tOyuDAQstZCZDUkd/c+sgLcMau/4CycbU1hho9cVfCuZaGocq+5KqV1JFQVZuQGcM+M2vcU
nXLXfOkFdGGfvJ+AJXlB92UCl2lXmq8vqWoYbSX7yDfEZDcOECmSphVaXgr6YEAx7NZdQ1cXDEKd
Wv3uKx0XdLeO7gN0PILfnSqVOlftd0egoSeZ8FWeiEv2IkwsBWJeLy9SM3fJp9azKPqXM4kcjAFg
83VqVc2KcWGAL9IphDRC3g16v6YpOb72YLgEb2QD+bxazH5hAIddwRFE4ANx0kBXYB+fyngZ3Wo3
2z7UrOOREQN7gIqqIWQuVijGIHzy6JLNiUPg/Q888eYqcz2h+5ZYQeUQJlcLOfm2IzNnIYegX8Rt
OEN3jG/42JMPw782FHHYzmdKEexqRR8tRRLzWqL9V3mVvlA3cgJIJoigBScSyO5nj+1RwhdY4igb
qsL0lsEaWjcr5+FiaHN9SAS4vIzk1ahJlo0+eItx3HKN3BPMJyXOTLiJteW36wwSiixbgk8vZ1L+
SSOYnQrD+FYKdAQB4j8w9jMaaEnstDA8KblmBnpFv0JXqmpTUFqehqI1kLml6wMdmxnVfbwf5qrF
RmKiNFUiozTQ+rlxmo1lD+GKhTZb82fozFMQLwzhqEnzJ2H2PgVnlOr3Z9HMk+MkXHnC2lius+kr
p8z+dZGWOzKDXNQKaSy6MhL8B2LVyu0qy11+aXvmXSJWXEVpHWUi46kuq8API4JmuTKIwF/BhEqd
d8A5+OrlfooLCgHQZkfQvWJ8YWUNom3cYvNuVSW6oJ23v+3GNagZqQalz4hb4A17ovFoTg9OVI44
IydGspVQLdHTg69zch/awjk8J7C1BzMsTgK7d15j61SaCopdHS24IdkBe3wgfRD5VHRErVUpFlzq
vUGCjQuHhZm7ISwmm0jv6Jt37NLFSvuCAcpM0UBDPpsgCX1ivZWpDT0JsNCUsIvM13fcQGz4lycS
KxV+3sj5TOyQPuX1xZFArO8SYukNiZVlcqAuNtfpZwzfpdzkVUt8+8WJMSYF0pMKgTgECHd2/XUE
oPPs55ip5YDTLHzskoFerMXn56UgPbn2LT8RU5xnPCBaLuiqoYEgg50sWFAdKFZeTU+ZMRs6IUbU
l4qf/pMIllyEK/3uHvilVDdnaIrzGno4KITBv0Enw0NeRasuR91JyTqfC3423367LCnhvyRVZxnv
aig4WQ2A0vcXy5uXPio3zK5u2MC701flLUZHCAsPEI7kf7T9AQApo7PZaSU=
`pragma protect end_protected
