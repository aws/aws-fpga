`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
CPJpGocSV6UwckyUGcP22ZpRrWKPgp0krAmn8MmPkXwl0b1+zQtBK1dBGRSXaiAaK6vph/4CerOK
hlWROjzkr4KZ2oWEWfEpo3+KEyDAUIdifSevkf0hYGuBDPII1/tdSnzIAbA1vu+KGYCQV9q8W7E6
K4yzTZgyFFabavqSQGjSVSCVsXJqS4X41EWLh00s3LqtY/4z1a3N4skHUwfqADuJKFgJSGpOUpyM
aTndiC/9FLsDmHa1EUDPbCyGBLsSbBuwAoCjTduGbXNoVzSHsK4tkP2h6U4VuwDwdJfLZDlIUjyi
8vlDhvJS7+TmYWxIK6jjwOo8mHky6bPdA9Q5Sg==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
T8hz0x6V6LMAFKq2+ujkb1bAjCrQFi0vZcG6Zl5VfO8xUw1DHfZmsWKCpDUiAVT4gBHdljyUJKAM
bNiIwzWXAyfMNwsp2wor3F8xrct5ADRMCRtJuWSDLF2/UDNaF38tKFuZzwtM4e/jsZ6OGZ7aOPUf
OlSFP/Y00u0P4Zxdz/U=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
LIYGP+Jz1fjWvA7DU4J2bYpPtWCsCH9GyTfR3Jy7zmaMMgXj2Ovp+egqiKlhIz3JlarauDzEzcb3
VmS35041lgljEwzBf3AVIJEDFglM00vhtcUso45V0emsy6RDAPmlVWOq9Q8L/eoOFBrcLwuvK2D0
v1w0MIHY/3N6ZbNhCyg=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1120)
`pragma protect data_block
3J7eI1nvax0I9RlDuK/caQ0+NUlr0l/x02zTKiYqjr9YyJCQXDSQnA1A/kD18ffk9kleP2ldrL3R
sqigHoNQUEZ1RyZ91g6Q2LJUecXA2k3BpvnozVbV+JsBL49lJKtQNcTVXqbfYlOMw/pSiaUPDqat
M/iwCVhOxnwsnwb7sseMmBE180JEV8YcYCEtDH3Jha8+Yb0vv7HkAlnZZXM2tW6vvKhyuKVxNOr9
zb6kQR0TV6aA+j7vb/9T/c8e51A0TdmdnqWrIYkJumwdYMkgFcqDBWtAWNtLRpHtLe2gcZvLXNDj
+WxkpkYU5AybPbU0LsLJrdNB5lJSnQk4H2PdDDfI2uLK2dSd9d1i1I8LzwsTVROv5jx4uWDr+g4s
jt5MMRxY6vqkyyn2jERyidXgEdSwGjcKYCyZrgmpCQs93AqJile7X0vrJMdv4WqLRC3PH+WRMrtv
nhdUWGj5X5LDoIQye4fiFQTVQtmhoq8hZVJVtP+SEQgkk9WFzcEA+k5Is9sbp9CHYPayFuZ/ttuC
isBKBUanp3znDcAZoD8vt5Sez5rMYrYeL1QLo7NpsGYOa31kRW13WYAeWJax3wyUEpZmuPxsmIt+
bMoT8h1KWVQl7TUq/OddVEsO7B0eISf8dhSoqo4PhgSBI/9VUTQbgMNQKal/iRgzG358RrlqlXsR
DJ8xxjUuE6YfBHGMnxs8uNnifSAbn5+rnKJSyB+o1dQQJEgrsh6qTOdL9PUrw9ZMiB338SNpAS9V
4B+L9/qhAemtoV1So99qoFszF3TYiYsG14EiJAkXgYb2zxCdS1XABBa5oKPS7nVuZx37OQhXS8jP
/OY8xzbycVbvasHmtlnPq0ZlaU+K/ghjwdEAoNWm/hzzWmq6tBKl+Ib4j7hdhlnrRic8jZBmran2
rluq8ZZTpxbuZVimxYplDVdeV6Ox6J/Ry7fDjaCO1SxgsdQzUbAG7V/8+9SLJ/1rXTPGfuMGFRPA
ZPdaAS0urTRzw8coUv8BXEyF8SkONzRVpG4YqG9UXAkJntuX/pgKrCL47h/Cb5SBmwCpQo9+T5kb
u+pY+zyw7HsBvyxMMk08PPxEfN2FnjyalFHcxkFppCjPW1sb8/PMo5a6szs43pzyLtxZ2UYcNkps
H5bgxAmoooSl2y+LeVXJGLHpaymNBiPO562X7KZ0gWE9FsVDHnuLCjsjKiyUsgl8S8BVLpqndG6b
HgDnnVAByE4+exBl/JiK7ww7SFPCYMFsYKCLRK//Ew3TyA2Rj+GHSdSbFda3LiSc4L90ZtUYCpPY
//omopd9J3q92dcMzo+JcqYhF+ifHbwz/MO17lGhmjKK6OVW1anZtrJAWPs+i6BoF12EGxD/edVv
Zi7LfDbAkNeSm8/wg2G1onp+J/5HQExxcFFbOpX6L+dlFghEnhl8BN8tJDuFnx+MEoZzqFT6DsMN
sPozE0+PZYRthyTFe9+xjWXgJM5G1RISwwpK3sZaIhB4HRFJBw==
`pragma protect end_protected
