`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
jVJg63YmByem+Wtav7SIzpprDGz7RSQNCQW+mkwDAosg+0Y7FU4xCDv7RWEvxYhMYQr1HZr2lL7S
i0IkxYlOsh3HZqCo7A3z5JYrJMHbEOMiHrIdzFZsmr4mvtERA01sK7gQW1xPpzI2zbvRRHC1MRWb
/5RqkEK3pvELDji3CdV1cPvWCJtpfsbVDAtCGPeYYovWil0FhUcW9oxP8+ZGf6swemamMi2Q3rt9
hFYZfo0gMqNG6gfxNcS+gSdEfvZML8du01++B6Amuj+QPoJEbF+ycwOnBPLIOL8Vvt6ix1nYT2dg
Irlq+psEfvD3cJsucF0ToG46chac24xCzLPdeg==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
YQR/N30d/3MzvaBdgjszzavwRagI5XJnhYadI3iOIjLfepvadFGyqn6pQ8KEKP6oDYDHvP8ov5SE
jM0EN78KCtaV0CyEHgqUOJqhrZFZYnaozptycdOClzyIkuGto5JziYsErITFmFPD9pdCu/g4AW3J
PL6rAb6ahF2urtNw3Pw=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
M6MwtpD2/ATABecZRVPX9/3/r2PowGsag3NhQB7zm9v+XAkpRB3x1zq3SWJE5exX0j9YfcGdijqb
GgUIt0ulGTm4P1LG0T2NeD8k6c39Zf8qUQD/oBoQodRRpbg0SL9oShHwQ9/s4fNTqzsoPgg6kZ/n
ad4O+lI2O8iMVJZNXhY=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1600)
`pragma protect data_block
vgcrQN1YIdXyKxjvZeCtUVT6ZE7yGMtgRRHrCcEFfDTkKutsNKiXsai44ZeoQuLLO+qrsVoO5VdP
XLY2q+PSmXie7jsbIWg0X6VrEVWuNdmpntN3DtXA94f6aqF0jQuMZe5cHsIad7jNBu/Gsz05+/jY
T5sbuhLeLe9TJ7+WZ57fX+KME5BgICextqOeziKYgJXBMzHoNSi3sEpcvk1Ut2+YaxzS4EIzGCWO
u0/TFMHYn8GSK1UDfVDt+RYJUilYzIifBqdjfH9qBzB5fk2KMW5oCMs3yJEn4rOJJYz3jdkabHm0
3VTRJxkCe46rkfT/0ItKKtL6C6Sd4nvFoYew0tNKUL0wBMoM0+maXY9RZkvmtYTuE+1ivIlUQS4Q
AE2PlAxzPGBSiz4BKK1ziWUdQquqg9eRiAVmd+j8tB5mTgFUFBSObyfWmFDlX9XMTCzY9MXHXBZt
15znrhaqS/A37azNE+33xiYxmTRgQw4LOiFyEPNzboVdL6GLxfViwNGGt0Z5ctf9E4UGGS2D7H0e
0Bf9FihRPAvcZ0QBssJ2LkHwpEGkrhUSXa0PDTB4FtZDFHIt20FCHB0BUReFGdD5kw2yOK9Olmpd
1NakrcJvTdUp5MfftILGuJWgs33ULuY+GSjXAmRbu1eRVRCMmMULwdIo+DfbR7S36Rhx5LqLAj9m
lgJSoY0rGQMoBGngvnBoIU9mdUHIEHlLJiI8SdFl8xTKqFYvCnJXyzyT5CUEngxiaoecjbtqEjsq
DCpMrWrYeddLZNnnKp/8RlsFta9H7K3rQUKrsGEARUHCdtw49or2yiXvBR/fJrhu4/lhC46JdMU2
8MDTuVHSuYQHVDE/28XGvdIRrI7LeS60VHDJycUhPFlhO0z5RlRBe+jdDN4256HH7cH5XJY16QGg
znGq7RXNyJVNZFwOzreDycGvnJQt4tGqAPcapp41AdsL6SS477k51CcsDhUhNdThb84jt3qN8j+s
z5ZqAHjUpNg1OK972wGPi+06ouP6pHigd/2UkOjSTvGoQFZIYTO4tWuz1+d0oaJEtoR+5ogxPHxM
+gOiTfmCKzWKTYjWGXf6R2Umz3Na8YWKACQ888suhSaYeh2NVC5/M0DobvtjHZjF6kvjDVPMjCQU
AW2kaB/TVya9cfnszfP7Bte/ipE7KY2iIwYWQACV0OU1wcTQFCBI6yjkcOyJIxN79bgtdbpvTL1f
VvsFq2LRMpKOo15wJRcXKTaP8rzp2qTnD+gOGkEXU5tvULbKGTZEiuIVkzQjWWp1CTwPEM5aysyc
ThwpDlRpF5qGdup+o+S+7lSDkDn9/iEcU1HttrUqbGM1cf35m9rX2AeieDVZTAMkZOLlKB6K+UMR
RUMDBBHfxoNeB/HrcfX2iCaQts/inzQQohDmR8fKUj2Mcxm/mgLaxOarsgYPwRRUUURp+sQ9ymvN
dHSGlDHVbqETEhrfWvNzUmHlFNtHOsPIvj7kRAe+91XGuQ0h2k+wx9gpxYveIwl4i5sdt+oo2ZaN
CE5DSqGXCLe9vvOBPytZfKw7SsKiE6X3H9UPCmq1rDAi7+D5ZzRNZ76aRV3eGCh/+0CBtjUp56wx
4jEy+i8zjL7YyytqLaCWXC1xS8b0mGmEBCL4ukoAOe6b7j4pSH9ZXKwYB+4SsK57gRi8OeD1Cwdq
rS7wt8Jl244BikWKFdgkNf1rNGS4Gpl/0tv3fqIuJ8FXtvM/PS5wgZ+s0Dq3mi1in9xtr8YYR4Yb
1OaNWdemaHIR7hREZk/qRohEJJW0zOUCkpz8Vw9VUK8stJrdjKVZ3Ot+gN6LRsivzFs5LTBlXxd8
v3gHxn55JxpG4XV5bmMCk3jAOSk5gwrHIrqL84maEUHSRCWkEYfOfNW6DHNo8YyIybyOGRSDJqfF
TSOU44IoSchHw5MW3s2ozYVrSX7jI4RT3Ua5/24bUo+2WyTN5QVb7TSe2t1oy/+9EFZq04z1+3Q7
yxmCx0kcTwYgXQcp/6hvpzbrA7MXhKODSEvc+lOuJFBHm/5RSetDEiJEUjUa3xtRIxtsMMMQL7h/
Nsg0x/9uL3OunxgVRI21mqVWO2bSUsCYVWw9LXcuzUOlYkUwo5gt4mwoo9gXISeYlV1siLvcOcmR
z3niog==
`pragma protect end_protected
