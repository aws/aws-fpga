// =============================================================================
// Copyright 2016 Amazon.com, Inc. or its affiliates.
// All Rights Reserved Worldwide.
// Amazon Confidential information
// Restricted NDA Material
// =============================================================================

module cl_dma_pcis_slv #(parameter SCRB_MAX_ADDR = 64'h3FFFFFFFF, parameter SCRB_BURST_LEN_MINUS1 = 15, parameter NO_SCRB_INST = 1)

(
    input aclk,
    input aresetn,

    cfg_bus_t ddr0_tst_cfg_bus,
    cfg_bus_t ddr1_tst_cfg_bus,
    cfg_bus_t ddr2_tst_cfg_bus,
    cfg_bus_t ddr3_tst_cfg_bus,

    scrb_bus_t ddr0_scrb_bus,
    scrb_bus_t ddr1_scrb_bus,
    scrb_bus_t ddr2_scrb_bus,
    scrb_bus_t ddr3_scrb_bus,

    input [5:0] sh_cl_dma_pcis_awid,
    input [63:0] sh_cl_dma_pcis_awaddr,
    input [7:0] sh_cl_dma_pcis_awlen,
    input [2:0] sh_cl_dma_pcis_awsize,
    input sh_cl_dma_pcis_awvalid,
    output logic cl_sh_dma_pcis_awready,
    
    input [511:0] sh_cl_dma_pcis_wdata,
    input [63:0] sh_cl_dma_pcis_wstrb,
    input sh_cl_dma_pcis_wlast,
    input sh_cl_dma_pcis_wvalid,
    output logic cl_sh_dma_pcis_wready,
    
    output logic [5:0] cl_sh_dma_pcis_bid,
    output logic [1:0] cl_sh_dma_pcis_bresp,
    output logic cl_sh_dma_pcis_bvalid,
    input sh_cl_dma_pcis_bready,
    
    input [5:0] sh_cl_dma_pcis_arid,
    input [63:0] sh_cl_dma_pcis_araddr,
    input [7:0] sh_cl_dma_pcis_arlen,
    input [2:0] sh_cl_dma_pcis_arsize,
    input sh_cl_dma_pcis_arvalid,
    output logic cl_sh_dma_pcis_arready,
    
    output logic [5:0] cl_sh_dma_pcis_rid,
    output logic [511:0] cl_sh_dma_pcis_rdata,
    output logic [1:0] cl_sh_dma_pcis_rresp,
    output logic cl_sh_dma_pcis_rlast,
    output logic cl_sh_dma_pcis_rvalid,
    input sh_cl_dma_pcis_rready,

    axi_bus_t lcl_cl_sh_ddr0,
    axi_bus_t lcl_cl_sh_ddr1,
    axi_bus_t lcl_cl_sh_ddr2,

    axi_bus_t sh_cl_dma_pcis_q,

    output [15:0] cl_sh_ddr_awid,
    output [63:0] cl_sh_ddr_awaddr,
    output [7:0] cl_sh_ddr_awlen,
    output [2:0] cl_sh_ddr_awsize,
    output  cl_sh_ddr_awvalid,
    input sh_cl_ddr_awready,
       
    output [15:0] cl_sh_ddr_wid,
    output [511:0] cl_sh_ddr_wdata,
    output [63:0] cl_sh_ddr_wstrb,
    output  cl_sh_ddr_wlast,
    output  cl_sh_ddr_wvalid,
    input sh_cl_ddr_wready,
       
    input[15:0] sh_cl_ddr_bid,
    input[1:0] sh_cl_ddr_bresp,
    input sh_cl_ddr_bvalid,
    output  cl_sh_ddr_bready,
       
    output [15:0] cl_sh_ddr_arid,
    output [63:0] cl_sh_ddr_araddr,
    output [7:0] cl_sh_ddr_arlen,
    output [2:0] cl_sh_ddr_arsize,
    output  cl_sh_ddr_arvalid,
    input sh_cl_ddr_arready,
       
    input[15:0] sh_cl_ddr_rid,
    input[511:0] sh_cl_ddr_rdata,
    input[1:0] sh_cl_ddr_rresp,
    input sh_cl_ddr_rlast,
    input sh_cl_ddr_rvalid,
    output  cl_sh_ddr_rready

 
);

//---------------------------- 
// Internal signals
//---------------------------- 
axi_bus_t lcl_cl_sh_ddr0_q();
axi_bus_t lcl_cl_sh_ddr1_q();
axi_bus_t lcl_cl_sh_ddr2_q();
axi_bus_t lcl_cl_sh_ddr0_q2();
axi_bus_t lcl_cl_sh_ddr1_q2();
axi_bus_t lcl_cl_sh_ddr2_q2();
axi_bus_t lcl_cl_sh_ddr0_q3();
axi_bus_t lcl_cl_sh_ddr1_q3();
axi_bus_t lcl_cl_sh_ddr2_q3();
axi_bus_t cl_sh_ddr_q();
axi_bus_t cl_sh_ddr_q2();
axi_bus_t cl_sh_ddr_q3();
axi_bus_t sh_cl_pcis();


//---------------------------- 
// End Internal signals
//---------------------------- 


   // AXI4 Register Slice for dma_pcis interface
   axi4_flop_fifo #(.IN_FIFO(1), .ADDR_WIDTH(64), .DATA_WIDTH(512), .ID_WIDTH(6), .A_USER_WIDTH(1), .FIFO_DEPTH(3)) PCI_AXL_REG_SLC (
       .aclk          (aclk),
       .aresetn       (aresetn),
       .sync_rst_n    (1'b1),
       .s_axi_awid    (sh_cl_dma_pcis_awid),
       .s_axi_awaddr  (sh_cl_dma_pcis_awaddr),
       .s_axi_awlen   (sh_cl_dma_pcis_awlen),                                            
       .s_axi_awvalid (sh_cl_dma_pcis_awvalid),
       .s_axi_awuser  (),
       .s_axi_awready (cl_sh_dma_pcis_awready),
       .s_axi_wdata   (sh_cl_dma_pcis_wdata),
       .s_axi_wstrb   (sh_cl_dma_pcis_wstrb),
       .s_axi_wlast   (sh_cl_dma_pcis_wlast),
       .s_axi_wuser   (),
       .s_axi_wvalid  (sh_cl_dma_pcis_wvalid),
       .s_axi_wready  (cl_sh_dma_pcis_wready),
       .s_axi_bid     (cl_sh_dma_pcis_bid),
       .s_axi_bresp   (cl_sh_dma_pcis_bresp),
       .s_axi_bvalid  (cl_sh_dma_pcis_bvalid),
       .s_axi_buser   (),
       .s_axi_bready  (sh_cl_dma_pcis_bready),
       .s_axi_arid    (sh_cl_dma_pcis_arid),
       .s_axi_araddr  (sh_cl_dma_pcis_araddr),
       .s_axi_arlen   (sh_cl_dma_pcis_arlen), 
       .s_axi_arvalid (sh_cl_dma_pcis_arvalid),
       .s_axi_aruser  (1'd0),
       .s_axi_arready (cl_sh_dma_pcis_arready),
       .s_axi_rid     (cl_sh_dma_pcis_rid),
       .s_axi_rdata   (cl_sh_dma_pcis_rdata),
       .s_axi_rresp   (cl_sh_dma_pcis_rresp),
       .s_axi_rlast   (cl_sh_dma_pcis_rlast),
       .s_axi_ruser   (),
       .s_axi_rvalid  (cl_sh_dma_pcis_rvalid),
       .s_axi_rready  (sh_cl_dma_pcis_rready), 
       .m_axi_awid    (sh_cl_dma_pcis_q.awid),
       .m_axi_awaddr  (sh_cl_dma_pcis_q.awaddr), 
       .m_axi_awlen   (sh_cl_dma_pcis_q.awlen),
       .m_axi_awvalid (sh_cl_dma_pcis_q.awvalid),
       .m_axi_awuser  (),
       .m_axi_awready (sh_cl_dma_pcis_q.awready),
       .m_axi_wdata   (sh_cl_dma_pcis_q.wdata),  
       .m_axi_wstrb   (sh_cl_dma_pcis_q.wstrb),
       .m_axi_wvalid  (sh_cl_dma_pcis_q.wvalid), 
       .m_axi_wlast   (sh_cl_dma_pcis_q.wlast),
       .m_axi_wuser   (),
       .m_axi_wready  (sh_cl_dma_pcis_q.wready), 
       .m_axi_bresp   (sh_cl_dma_pcis_q.bresp),  
       .m_axi_bvalid  (sh_cl_dma_pcis_q.bvalid), 
       .m_axi_bid     (sh_cl_dma_pcis_q.bid),
       .m_axi_buser   (),
       .m_axi_bready  (sh_cl_dma_pcis_q.bready), 
       .m_axi_arid    (sh_cl_dma_pcis_q.arid), 
       .m_axi_araddr  (sh_cl_dma_pcis_q.araddr), 
       .m_axi_arlen   (sh_cl_dma_pcis_q.arlen), 
       .m_axi_aruser  (), 
       .m_axi_arvalid (sh_cl_dma_pcis_q.arvalid),
       .m_axi_arready (sh_cl_dma_pcis_q.arready),
       .m_axi_rid     (sh_cl_dma_pcis_q.rid),  
       .m_axi_rdata   (sh_cl_dma_pcis_q.rdata),  
       .m_axi_rresp   (sh_cl_dma_pcis_q.rresp),  
       .m_axi_rlast   (sh_cl_dma_pcis_q.rlast),  
       .m_axi_ruser   (1'b0),
       .m_axi_rvalid  (sh_cl_dma_pcis_q.rvalid), 
       .m_axi_rready  (sh_cl_dma_pcis_q.rready)
   );


   axi_crossbar_0 AXI_CROSSBAR (
       .aclk(aclk),
       .aresetn(aresetn),

       .s_axi_awid(sh_cl_dma_pcis_q.awid),
       .s_axi_awaddr({sh_cl_dma_pcis_q.awaddr[63:37], 1'b0, sh_cl_dma_pcis_q.awaddr[35:0]}),
       .s_axi_awlen(sh_cl_dma_pcis_q.awlen),
       .s_axi_awsize(sh_cl_dma_pcis_q.awsize),
       .s_axi_awburst(2'b1),
       .s_axi_awlock(1'b0),
       .s_axi_awcache(4'b11),
       .s_axi_awprot(3'b10),
       .s_axi_awqos(4'b0),
       .s_axi_awvalid(sh_cl_dma_pcis_q.awvalid),
       .s_axi_awready(sh_cl_dma_pcis_q.awready),

       .s_axi_wdata(sh_cl_dma_pcis_q.wdata),
       .s_axi_wstrb(sh_cl_dma_pcis_q.wstrb),
       .s_axi_wlast(sh_cl_dma_pcis_q.wlast),
       .s_axi_wvalid(sh_cl_dma_pcis_q.wvalid),
       .s_axi_wready(sh_cl_dma_pcis_q.wready),

       .s_axi_bid(sh_cl_dma_pcis_q.bid),
       .s_axi_bresp(sh_cl_dma_pcis_q.bresp),
       .s_axi_bvalid(sh_cl_dma_pcis_q.bvalid),
       .s_axi_bready(sh_cl_dma_pcis_q.bready),

       .s_axi_arid(sh_cl_dma_pcis_q.arid),
       .s_axi_araddr({sh_cl_dma_pcis_q.araddr[63:37], 1'b0, sh_cl_dma_pcis_q.araddr[35:0]}),
       .s_axi_arlen(sh_cl_dma_pcis_q.arlen),
       .s_axi_arsize(sh_cl_dma_pcis_q.arsize),
       .s_axi_arburst(2'b1),
       .s_axi_arlock(1'b0),
       .s_axi_arcache(4'b11),
       .s_axi_arprot(3'b10),
       .s_axi_arqos(4'b0),
       .s_axi_arvalid(sh_cl_dma_pcis_q.arvalid),
       .s_axi_arready(sh_cl_dma_pcis_q.arready),

       .s_axi_rid(sh_cl_dma_pcis_q.rid),
       .s_axi_rdata(sh_cl_dma_pcis_q.rdata),
       .s_axi_rresp(sh_cl_dma_pcis_q.rresp),
       .s_axi_rlast(sh_cl_dma_pcis_q.rlast),
       .s_axi_rvalid(sh_cl_dma_pcis_q.rvalid),
       .s_axi_rready(sh_cl_dma_pcis_q.rready), 

       .m_axi_awid({sh_cl_pcis.awid, lcl_cl_sh_ddr2_q.awid[5:0], cl_sh_ddr_q.awid[5:0], lcl_cl_sh_ddr1_q.awid[5:0], lcl_cl_sh_ddr0_q.awid[5:0]}),
       .m_axi_awaddr({sh_cl_pcis.awaddr, lcl_cl_sh_ddr2_q.awaddr, cl_sh_ddr_q.awaddr, lcl_cl_sh_ddr1_q.awaddr, lcl_cl_sh_ddr0_q.awaddr}),
       .m_axi_awlen({sh_cl_pcis.awlen, lcl_cl_sh_ddr2_q.awlen, cl_sh_ddr_q.awlen, lcl_cl_sh_ddr1_q.awlen, lcl_cl_sh_ddr0_q.awlen}),
       .m_axi_awsize(),
       .m_axi_awburst(),
       .m_axi_awlock(),
       .m_axi_awcache(),
       .m_axi_awprot(),
       .m_axi_awregion(),
       .m_axi_awqos(),
       .m_axi_awvalid({sh_cl_pcis.awvalid, lcl_cl_sh_ddr2_q.awvalid, cl_sh_ddr_q.awvalid, lcl_cl_sh_ddr1_q.awvalid, lcl_cl_sh_ddr0_q.awvalid}),
       .m_axi_awready({1'b0, lcl_cl_sh_ddr2_q.awready, cl_sh_ddr_q.awready, lcl_cl_sh_ddr1_q.awready, lcl_cl_sh_ddr0_q.awready}),
  
       .m_axi_wdata({sh_cl_pcis.wdata, lcl_cl_sh_ddr2_q.wdata, cl_sh_ddr_q.wdata, lcl_cl_sh_ddr1_q.wdata, lcl_cl_sh_ddr0_q.wdata}),
       .m_axi_wstrb({sh_cl_pcis.wstrb, lcl_cl_sh_ddr2_q.wstrb, cl_sh_ddr_q.wstrb, lcl_cl_sh_ddr1_q.wstrb, lcl_cl_sh_ddr0_q.wstrb}),
       .m_axi_wlast({sh_cl_pcis.wlast, lcl_cl_sh_ddr2_q.wlast, cl_sh_ddr_q.wlast, lcl_cl_sh_ddr1_q.wlast, lcl_cl_sh_ddr0_q.wlast}),
       .m_axi_wvalid({sh_cl_pcis.wvalid, lcl_cl_sh_ddr2_q.wvalid, cl_sh_ddr_q.wvalid, lcl_cl_sh_ddr1_q.wvalid, lcl_cl_sh_ddr0_q.wvalid}),
       .m_axi_wready({1'b0, lcl_cl_sh_ddr2_q.wready, cl_sh_ddr_q.wready, lcl_cl_sh_ddr1_q.wready, lcl_cl_sh_ddr0_q.wready}),
    
       .m_axi_bid({sh_cl_pcis.bid, lcl_cl_sh_ddr2_q.bid[5:0], cl_sh_ddr_q.bid[5:0], lcl_cl_sh_ddr1_q.bid[5:0], lcl_cl_sh_ddr0_q.bid[5:0]}),
       .m_axi_bresp({sh_cl_pcis.bresp, lcl_cl_sh_ddr2_q.bresp, cl_sh_ddr_q.bresp, lcl_cl_sh_ddr1_q.bresp, lcl_cl_sh_ddr0_q.bresp}),
       .m_axi_bvalid({1'b0, lcl_cl_sh_ddr2_q.bvalid, cl_sh_ddr_q.bvalid, lcl_cl_sh_ddr1_q.bvalid, lcl_cl_sh_ddr0_q.bvalid}),
       .m_axi_bready({sh_cl_pcis.bready, lcl_cl_sh_ddr2_q.bready, cl_sh_ddr_q.bready, lcl_cl_sh_ddr1_q.bready, lcl_cl_sh_ddr0_q.bready}),
  
       .m_axi_arid({sh_cl_pcis.arid, lcl_cl_sh_ddr2_q.arid[5:0], cl_sh_ddr_q.arid[5:0], lcl_cl_sh_ddr1_q.arid[5:0], lcl_cl_sh_ddr0_q.arid[5:0]}),
       .m_axi_araddr({sh_cl_pcis.araddr, lcl_cl_sh_ddr2_q.araddr, cl_sh_ddr_q.araddr, lcl_cl_sh_ddr1_q.araddr, lcl_cl_sh_ddr0_q.araddr}),
       .m_axi_arlen({sh_cl_pcis.arlen, lcl_cl_sh_ddr2_q.arlen, cl_sh_ddr_q.arlen, lcl_cl_sh_ddr1_q.arlen, lcl_cl_sh_ddr0_q.arlen}),
       .m_axi_arsize(),
       .m_axi_arburst(),
       .m_axi_arlock(),
       .m_axi_arcache(),
       .m_axi_arprot(),
       .m_axi_arregion(),
       .m_axi_arqos(),
       .m_axi_arvalid({sh_cl_pcis.arvalid, lcl_cl_sh_ddr2_q.arvalid, cl_sh_ddr_q.arvalid, lcl_cl_sh_ddr1_q.arvalid, lcl_cl_sh_ddr0_q.arvalid}),
       .m_axi_arready({1'b0, lcl_cl_sh_ddr2_q.arready, cl_sh_ddr_q.arready, lcl_cl_sh_ddr1_q.arready, lcl_cl_sh_ddr0_q.arready}),

       .m_axi_rid({sh_cl_pcis.rid, lcl_cl_sh_ddr2_q.rid[5:0], cl_sh_ddr_q.rid[5:0], lcl_cl_sh_ddr1_q.rid[5:0], lcl_cl_sh_ddr0_q.rid[5:0]}),
       .m_axi_rdata({sh_cl_pcis.rdata, lcl_cl_sh_ddr2_q.rdata, cl_sh_ddr_q.rdata, lcl_cl_sh_ddr1_q.rdata, lcl_cl_sh_ddr0_q.rdata}),
       .m_axi_rresp({sh_cl_pcis.rresp, lcl_cl_sh_ddr2_q.rresp, cl_sh_ddr_q.rresp, lcl_cl_sh_ddr1_q.rresp, lcl_cl_sh_ddr0_q.rresp}),
       .m_axi_rlast({sh_cl_pcis.rlast, lcl_cl_sh_ddr2_q.rlast, cl_sh_ddr_q.rlast, lcl_cl_sh_ddr1_q.rlast, lcl_cl_sh_ddr0_q.rlast}),
       .m_axi_rvalid({1'b0, lcl_cl_sh_ddr2_q.rvalid, cl_sh_ddr_q.rvalid, lcl_cl_sh_ddr1_q.rvalid, lcl_cl_sh_ddr0_q.rvalid}),
       .m_axi_rready({sh_cl_pcis.rready, lcl_cl_sh_ddr2_q.rready, cl_sh_ddr_q.rready, lcl_cl_sh_ddr1_q.rready, lcl_cl_sh_ddr0_q.rready})
   );


   axi4_flop_fifo #(.ADDR_WIDTH(64), .DATA_WIDTH(512), .ID_WIDTH(6), .A_USER_WIDTH(1), .FIFO_DEPTH(3)) DDR_TST_3_AXI4_REG_SLC (
       .aclk           (aclk),
       .aresetn        (aresetn),
       .sync_rst_n     (1'b1),
                                                                                                                                  
       .s_axi_awid     (cl_sh_ddr_q.awid),
       .s_axi_awaddr   ({cl_sh_ddr_q.awaddr[63:32], 2'b0, cl_sh_ddr_q.awaddr[29:0]}),
       .s_axi_awlen    (cl_sh_ddr_q.awlen),
       .s_axi_awuser   (1'b0),
       .s_axi_awvalid  (cl_sh_ddr_q.awvalid),
       .s_axi_awready  (cl_sh_ddr_q.awready),
       .s_axi_wdata    (cl_sh_ddr_q.wdata),
       .s_axi_wstrb    (cl_sh_ddr_q.wstrb),
       .s_axi_wlast    (cl_sh_ddr_q.wlast),
       .s_axi_wvalid   (cl_sh_ddr_q.wvalid),
       .s_axi_wuser    (),
       .s_axi_wready   (cl_sh_ddr_q.wready),
       .s_axi_bid      (cl_sh_ddr_q.bid),
       .s_axi_bresp    (cl_sh_ddr_q.bresp),
       .s_axi_bvalid   (cl_sh_ddr_q.bvalid),
       .s_axi_buser    (),
       .s_axi_bready   (cl_sh_ddr_q.bready),
       .s_axi_arid     (cl_sh_ddr_q.arid),
       .s_axi_araddr   ({cl_sh_ddr_q.araddr[63:32], 2'b0, cl_sh_ddr_q.araddr[29:0]}),
       .s_axi_arlen    (cl_sh_ddr_q.arlen),
       .s_axi_aruser   (1'b0),
       .s_axi_arvalid  (cl_sh_ddr_q.arvalid),
       .s_axi_arready  (cl_sh_ddr_q.arready),
       .s_axi_rid      (cl_sh_ddr_q.rid),
       .s_axi_rdata    (cl_sh_ddr_q.rdata),
       .s_axi_rresp    (cl_sh_ddr_q.rresp),
       .s_axi_rlast    (cl_sh_ddr_q.rlast),
       .s_axi_ruser    (),
       .s_axi_rvalid   (cl_sh_ddr_q.rvalid),
       .s_axi_rready   (cl_sh_ddr_q.rready),  
       .m_axi_awid     (cl_sh_ddr_q2.awid),   
       .m_axi_awaddr   (cl_sh_ddr_q2.awaddr), 
       .m_axi_awlen    (cl_sh_ddr_q2.awlen),  
       .m_axi_awuser   (),
       .m_axi_awvalid  (cl_sh_ddr_q2.awvalid),
       .m_axi_awready  (cl_sh_ddr_q2.awready),
       .m_axi_wdata    (cl_sh_ddr_q2.wdata),  
       .m_axi_wstrb    (cl_sh_ddr_q2.wstrb),  
       .m_axi_wuser    (),
       .m_axi_wlast    (cl_sh_ddr_q2.wlast),  
       .m_axi_wvalid   (cl_sh_ddr_q2.wvalid), 
       .m_axi_wready   (cl_sh_ddr_q2.wready), 
       .m_axi_bid      (cl_sh_ddr_q2.bid),    
       .m_axi_bresp    (cl_sh_ddr_q2.bresp),  
       .m_axi_buser    (),
       .m_axi_bvalid   (cl_sh_ddr_q2.bvalid), 
       .m_axi_bready   (cl_sh_ddr_q2.bready), 
       .m_axi_arid     (cl_sh_ddr_q2.arid),   
       .m_axi_araddr   (cl_sh_ddr_q2.araddr), 
       .m_axi_arlen    (cl_sh_ddr_q2.arlen),  
       .m_axi_aruser   (),
       .m_axi_arvalid  (cl_sh_ddr_q2.arvalid),
       .m_axi_arready  (cl_sh_ddr_q2.arready),
       .m_axi_rid      (cl_sh_ddr_q2.rid),    
       .m_axi_rdata    (cl_sh_ddr_q2.rdata),  
       .m_axi_rresp    (cl_sh_ddr_q2.rresp),  
       .m_axi_ruser    (),
       .m_axi_rlast    (cl_sh_ddr_q2.rlast),  
       .m_axi_rvalid   (cl_sh_ddr_q2.rvalid), 
       .m_axi_rready   (cl_sh_ddr_q2.rready)
   );



   cl_tst_scrb #(.DATA_WIDTH(512),
                    .SCRB_BURST_LEN_MINUS1(SCRB_BURST_LEN_MINUS1),
                    .SCRB_MAX_ADDR(SCRB_MAX_ADDR),
                    .NO_SCRB_INST(NO_SCRB_INST)) CL_TST_DDR_3 (
   
         .clk(aclk),
         .rst_n(aresetn),

         .cfg_addr(ddr2_tst_cfg_bus.addr),
         .cfg_wdata(ddr2_tst_cfg_bus.wdata),
         .cfg_wr(ddr2_tst_cfg_bus.wr),
         .cfg_rd(ddr2_tst_cfg_bus.rd),
         .tst_cfg_ack(ddr2_tst_cfg_bus.ack),
         .tst_cfg_rdata(ddr2_tst_cfg_bus.rdata), 

         .slv_awid(cl_sh_ddr_q2.awid[5:0]),
         .slv_awaddr(cl_sh_ddr_q2.awaddr), 
         .slv_awlen(cl_sh_ddr_q2.awlen),
         .slv_awvalid(cl_sh_ddr_q2.awvalid),
         .slv_awuser(11'b0),
         .slv_awready(cl_sh_ddr_q2.awready),

         .slv_wid(6'b0),
         .slv_wdata(cl_sh_ddr_q2.wdata),
         .slv_wstrb(cl_sh_ddr_q2.wstrb),
         .slv_wlast(cl_sh_ddr_q2.wlast),
         .slv_wvalid(cl_sh_ddr_q2.wvalid),
         .slv_wready(cl_sh_ddr_q2.wready),

         .slv_bid(cl_sh_ddr_q2.bid[5:0]),
         .slv_bresp(cl_sh_ddr_q2.bresp),
         .slv_buser(),
         .slv_bvalid(cl_sh_ddr_q2.bvalid),
         .slv_bready(cl_sh_ddr_q2.bready),

         .slv_arid(cl_sh_ddr_q2.arid[5:0]),
         .slv_araddr(cl_sh_ddr_q2.araddr), 
         .slv_arlen(cl_sh_ddr_q2.arlen),
         .slv_arvalid(cl_sh_ddr_q2.arvalid),
         .slv_aruser(11'b0),
         .slv_arready(cl_sh_ddr_q2.arready),        

         .slv_rid(cl_sh_ddr_q2.rid[5:0]),
         .slv_rdata(cl_sh_ddr_q2.rdata),
         .slv_rresp(cl_sh_ddr_q2.rresp),
         .slv_rlast(cl_sh_ddr_q2.rlast),
         .slv_ruser(),
         .slv_rvalid(cl_sh_ddr_q2.rvalid),
         .slv_rready(cl_sh_ddr_q2.rready),

                                               
         .awid(cl_sh_ddr_q3.awid),
         .awaddr(cl_sh_ddr_q3.awaddr), 
         .awlen(cl_sh_ddr_q3.awlen),
         .awvalid(cl_sh_ddr_q3.awvalid),
         .awuser(),
         .awready(cl_sh_ddr_q3.awready),

         //.wid(cl_sh_ddr_q3.wid),
         .wid(),
         .wdata(cl_sh_ddr_q3.wdata),
         .wstrb(cl_sh_ddr_q3.wstrb),
         .wlast(cl_sh_ddr_q3.wlast),
         .wvalid(cl_sh_ddr_q3.wvalid),
         .wready(cl_sh_ddr_q3.wready),

         .bid(cl_sh_ddr_q3.bid),
         .bresp(cl_sh_ddr_q3.bresp),
         .buser(18'h0),
         .bvalid(cl_sh_ddr_q3.bvalid),
         .bready(cl_sh_ddr_q3.bready),

         .arid(cl_sh_ddr_q3.arid),
         .araddr(cl_sh_ddr_q3.araddr),
         .arlen(cl_sh_ddr_q3.arlen),
         .arvalid(cl_sh_ddr_q3.arvalid),
         .aruser(),
         .arready(cl_sh_ddr_q3.arready),

         .rid(cl_sh_ddr_q3.rid),
         .rdata(cl_sh_ddr_q3.rdata),
         .rresp(cl_sh_ddr_q3.rresp),
         .rlast(cl_sh_ddr_q3.rlast),
         .ruser(18'h0),
         .rvalid(cl_sh_ddr_q3.rvalid),
         .rready(cl_sh_ddr_q3.rready),

         .scrb_enable(ddr2_scrb_bus.enable),
         .scrb_done  (ddr2_scrb_bus.done),

         .scrb_dbg_state(ddr2_scrb_bus.state),
         .scrb_dbg_addr (ddr2_scrb_bus.addr)
   );

   axi4_flop_fifo #(.ADDR_WIDTH(64), .DATA_WIDTH(512), .ID_WIDTH(16), .A_USER_WIDTH(1), .FIFO_DEPTH(3)) DDR_TST_3_AXI4_REG_SLC_1 (
     .aclk           (aclk),
     .aresetn        (aresetn),
     .sync_rst_n     (1'b1),
                                                                                                                                
     .s_axi_awid     ({10'b0, cl_sh_ddr_q3.awid}),
     .s_axi_awaddr   ({cl_sh_ddr_q3.awaddr}),
     .s_axi_awlen    (cl_sh_ddr_q3.awlen),
     .s_axi_awuser   (1'b0),
     .s_axi_awvalid  (cl_sh_ddr_q3.awvalid),
     .s_axi_awready  (cl_sh_ddr_q3.awready),
     .s_axi_wdata    (cl_sh_ddr_q3.wdata),
     .s_axi_wstrb    (cl_sh_ddr_q3.wstrb),
     .s_axi_wlast    (cl_sh_ddr_q3.wlast),
     .s_axi_wvalid   (cl_sh_ddr_q3.wvalid),
     .s_axi_wuser    (),
     .s_axi_wready   (cl_sh_ddr_q3.wready),
     .s_axi_bid      (cl_sh_ddr_q3.bid),
     .s_axi_bresp    (cl_sh_ddr_q3.bresp),
     .s_axi_bvalid   (cl_sh_ddr_q3.bvalid),
     .s_axi_buser    (),
     .s_axi_bready   (cl_sh_ddr_q3.bready),
     .s_axi_arid     ({10'b0, cl_sh_ddr_q3.arid}),
     .s_axi_araddr   (cl_sh_ddr_q3.araddr),
     .s_axi_arlen    (cl_sh_ddr_q3.arlen),
     .s_axi_aruser   (1'b0),
     .s_axi_arvalid  (cl_sh_ddr_q3.arvalid),
     .s_axi_arready  (cl_sh_ddr_q3.arready),
     .s_axi_rid      (cl_sh_ddr_q3.rid),
     .s_axi_rdata    (cl_sh_ddr_q3.rdata),
     .s_axi_rresp    (cl_sh_ddr_q3.rresp),
     .s_axi_rlast    (cl_sh_ddr_q3.rlast),
     .s_axi_ruser    (),
     .s_axi_rvalid   (cl_sh_ddr_q3.rvalid),
     .s_axi_rready   (cl_sh_ddr_q3.rready),  
     .m_axi_awid     (cl_sh_ddr_awid),   
     .m_axi_awaddr   (cl_sh_ddr_awaddr), 
     .m_axi_awlen    (cl_sh_ddr_awlen),  
     .m_axi_awuser   (),
     .m_axi_awvalid  (cl_sh_ddr_awvalid),
     .m_axi_awready  (sh_cl_ddr_awready),
     .m_axi_wdata    (cl_sh_ddr_wdata),  
     .m_axi_wstrb    (cl_sh_ddr_wstrb),  
     .m_axi_wuser    (),
     .m_axi_wlast    (cl_sh_ddr_wlast),  
     .m_axi_wvalid   (cl_sh_ddr_wvalid), 
     .m_axi_wready   (sh_cl_ddr_wready), 
     .m_axi_bid      (sh_cl_ddr_bid),    
     .m_axi_bresp    (sh_cl_ddr_bresp),  
     .m_axi_buser    (),
     .m_axi_bvalid   (sh_cl_ddr_bvalid), 
     .m_axi_bready   (cl_sh_ddr_bready), 
     .m_axi_arid     (cl_sh_ddr_arid),   
     .m_axi_araddr   (cl_sh_ddr_araddr), 
     .m_axi_arlen    (cl_sh_ddr_arlen),  
     .m_axi_aruser   (),
     .m_axi_arvalid  (cl_sh_ddr_arvalid),
     .m_axi_arready  (sh_cl_ddr_arready),
     .m_axi_rid      (sh_cl_ddr_rid),    
     .m_axi_rdata    (sh_cl_ddr_rdata),  
     .m_axi_rresp    (sh_cl_ddr_rresp),  
     .m_axi_ruser    (),
     .m_axi_rlast    (sh_cl_ddr_rlast),  
     .m_axi_rvalid   (sh_cl_ddr_rvalid), 
     .m_axi_rready   (cl_sh_ddr_rready)
   );


   //back to back register slices for SLR crossing
   src_register_slice DDR0_TST_AXI4_REG_SLC_1 (
       .aclk           (aclk),
       .aresetn        (aresetn),
       .s_axi_awid     (lcl_cl_sh_ddr0_q.awid[5:0]),
       .s_axi_awaddr   ({lcl_cl_sh_ddr0_q.awaddr[63:32], 2'b0, lcl_cl_sh_ddr0_q.awaddr[29:0]}),
       .s_axi_awlen    (lcl_cl_sh_ddr0_q.awlen),
       .s_axi_awsize   (3'b110),
       .s_axi_awburst  (2'b1),
       .s_axi_awlock   (1'b0),
       .s_axi_awcache  (4'b11),
       .s_axi_awprot   (3'b10),
       .s_axi_awregion (4'b0),
       .s_axi_awqos    (4'b0),
       .s_axi_awvalid  (lcl_cl_sh_ddr0_q.awvalid),
       .s_axi_awready  (lcl_cl_sh_ddr0_q.awready),
       .s_axi_wdata    (lcl_cl_sh_ddr0_q.wdata),
       .s_axi_wstrb    (lcl_cl_sh_ddr0_q.wstrb),
       .s_axi_wlast    (lcl_cl_sh_ddr0_q.wlast),
       .s_axi_wvalid   (lcl_cl_sh_ddr0_q.wvalid),
       .s_axi_wready   (lcl_cl_sh_ddr0_q.wready),
       .s_axi_bid      (lcl_cl_sh_ddr0_q.bid[5:0]),
       .s_axi_bresp    (lcl_cl_sh_ddr0_q.bresp),
       .s_axi_bvalid   (lcl_cl_sh_ddr0_q.bvalid),
       .s_axi_bready   (lcl_cl_sh_ddr0_q.bready),
       .s_axi_arid     (lcl_cl_sh_ddr0_q.arid[5:0]),
       .s_axi_araddr   ({lcl_cl_sh_ddr0_q.araddr[63:32], 2'b0, lcl_cl_sh_ddr0_q.araddr[29:0]}),
       .s_axi_arlen    (lcl_cl_sh_ddr0_q.arlen),
       .s_axi_arsize   (3'b110),
       .s_axi_arburst  (2'b1),
       .s_axi_arlock   (1'b0),
       .s_axi_arcache  (4'b11),
       .s_axi_arprot   (3'b10),
       .s_axi_arregion (4'b0),
       .s_axi_arqos    (4'b0),
       .s_axi_arvalid  (lcl_cl_sh_ddr0_q.arvalid),
       .s_axi_arready  (lcl_cl_sh_ddr0_q.arready),
       .s_axi_rid      (lcl_cl_sh_ddr0_q.rid[5:0]),
       .s_axi_rdata    (lcl_cl_sh_ddr0_q.rdata),
       .s_axi_rresp    (lcl_cl_sh_ddr0_q.rresp),
       .s_axi_rlast    (lcl_cl_sh_ddr0_q.rlast),
       .s_axi_rvalid   (lcl_cl_sh_ddr0_q.rvalid),
       .s_axi_rready   (lcl_cl_sh_ddr0_q.rready),  
       .m_axi_awid     (lcl_cl_sh_ddr0_q2.awid[5:0]),   
       .m_axi_awaddr   (lcl_cl_sh_ddr0_q2.awaddr), 
       .m_axi_awlen    (lcl_cl_sh_ddr0_q2.awlen),  
       .m_axi_awvalid  (lcl_cl_sh_ddr0_q2.awvalid),
       .m_axi_awready  (lcl_cl_sh_ddr0_q2.awready),
       .m_axi_wdata    (lcl_cl_sh_ddr0_q2.wdata),  
       .m_axi_wstrb    (lcl_cl_sh_ddr0_q2.wstrb),  
       .m_axi_wlast    (lcl_cl_sh_ddr0_q2.wlast),  
       .m_axi_wvalid   (lcl_cl_sh_ddr0_q2.wvalid), 
       .m_axi_wready   (lcl_cl_sh_ddr0_q2.wready), 
       .m_axi_bid      (lcl_cl_sh_ddr0_q2.bid[5:0]),    
       .m_axi_bresp    (lcl_cl_sh_ddr0_q2.bresp),  
       .m_axi_bvalid   (lcl_cl_sh_ddr0_q2.bvalid), 
       .m_axi_bready   (lcl_cl_sh_ddr0_q2.bready), 
       .m_axi_arid     (lcl_cl_sh_ddr0_q2.arid[5:0]),   
       .m_axi_araddr   (lcl_cl_sh_ddr0_q2.araddr), 
       .m_axi_arlen    (lcl_cl_sh_ddr0_q2.arlen),  
       .m_axi_arvalid  (lcl_cl_sh_ddr0_q2.arvalid),
       .m_axi_arready  (lcl_cl_sh_ddr0_q2.arready),
       .m_axi_rid      (lcl_cl_sh_ddr0_q2.rid[5:0]),    
       .m_axi_rdata    (lcl_cl_sh_ddr0_q2.rdata),  
       .m_axi_rresp    (lcl_cl_sh_ddr0_q2.rresp),  
       .m_axi_rlast    (lcl_cl_sh_ddr0_q2.rlast),  
       .m_axi_rvalid   (lcl_cl_sh_ddr0_q2.rvalid), 
       .m_axi_rready   (lcl_cl_sh_ddr0_q2.rready)
       );
   dest_register_slice DDR0_TST_AXI4_REG_SLC_2 (
       .aclk           (aclk),
       .aresetn        (aresetn),
       .s_axi_awid     (lcl_cl_sh_ddr0_q2.awid),
       .s_axi_awaddr   (lcl_cl_sh_ddr0_q2.awaddr),
       .s_axi_awlen    (lcl_cl_sh_ddr0_q2.awlen),
       .s_axi_awsize   (3'b110),
       .s_axi_awburst  (2'b1),
       .s_axi_awlock   (1'b0),
       .s_axi_awcache  (4'b11),
       .s_axi_awprot   (3'b10),
       .s_axi_awregion (4'b0),
       .s_axi_awqos    (4'b0),
       .s_axi_awvalid  (lcl_cl_sh_ddr0_q2.awvalid),
       .s_axi_awready  (lcl_cl_sh_ddr0_q2.awready),
       .s_axi_wdata    (lcl_cl_sh_ddr0_q2.wdata),
       .s_axi_wstrb    (lcl_cl_sh_ddr0_q2.wstrb),
       .s_axi_wlast    (lcl_cl_sh_ddr0_q2.wlast),
       .s_axi_wvalid   (lcl_cl_sh_ddr0_q2.wvalid),
       .s_axi_wready   (lcl_cl_sh_ddr0_q2.wready),
       .s_axi_bid      (lcl_cl_sh_ddr0_q2.bid),
       .s_axi_bresp    (lcl_cl_sh_ddr0_q2.bresp),
       .s_axi_bvalid   (lcl_cl_sh_ddr0_q2.bvalid),
       .s_axi_bready   (lcl_cl_sh_ddr0_q2.bready),
       .s_axi_arid     (lcl_cl_sh_ddr0_q2.arid),
       .s_axi_araddr   (lcl_cl_sh_ddr0_q2.araddr),
       .s_axi_arlen    (lcl_cl_sh_ddr0_q2.arlen),
       .s_axi_arsize   (3'b110),
       .s_axi_arburst  (2'b1),
       .s_axi_arlock   (1'b0),
       .s_axi_arcache  (4'b11),
       .s_axi_arprot   (3'b10),
       .s_axi_arregion (4'b0),
       .s_axi_arqos    (4'b0),
       .s_axi_arvalid  (lcl_cl_sh_ddr0_q2.arvalid),
       .s_axi_arready  (lcl_cl_sh_ddr0_q2.arready),
       .s_axi_rid      (lcl_cl_sh_ddr0_q2.rid),
       .s_axi_rdata    (lcl_cl_sh_ddr0_q2.rdata),
       .s_axi_rresp    (lcl_cl_sh_ddr0_q2.rresp),
       .s_axi_rlast    (lcl_cl_sh_ddr0_q2.rlast),
       .s_axi_rvalid   (lcl_cl_sh_ddr0_q2.rvalid),
       .s_axi_rready   (lcl_cl_sh_ddr0_q2.rready),  
       .m_axi_awid     (lcl_cl_sh_ddr0_q3.awid),   
       .m_axi_awaddr   (lcl_cl_sh_ddr0_q3.awaddr), 
       .m_axi_awlen    (lcl_cl_sh_ddr0_q3.awlen),  
       .m_axi_awvalid  (lcl_cl_sh_ddr0_q3.awvalid),
       .m_axi_awready  (lcl_cl_sh_ddr0_q3.awready),
       .m_axi_wdata    (lcl_cl_sh_ddr0_q3.wdata),  
       .m_axi_wstrb    (lcl_cl_sh_ddr0_q3.wstrb),  
       .m_axi_wlast    (lcl_cl_sh_ddr0_q3.wlast),  
       .m_axi_wvalid   (lcl_cl_sh_ddr0_q3.wvalid), 
       .m_axi_wready   (lcl_cl_sh_ddr0_q3.wready), 
       .m_axi_bid      ({10'b0, lcl_cl_sh_ddr0_q3.bid[5:0]}),    
       .m_axi_bresp    (lcl_cl_sh_ddr0_q3.bresp),  
       .m_axi_bvalid   (lcl_cl_sh_ddr0_q3.bvalid), 
       .m_axi_bready   (lcl_cl_sh_ddr0_q3.bready), 
       .m_axi_arid     (lcl_cl_sh_ddr0_q3.arid),   
       .m_axi_araddr   (lcl_cl_sh_ddr0_q3.araddr), 
       .m_axi_arlen    (lcl_cl_sh_ddr0_q3.arlen),  
       .m_axi_arvalid  (lcl_cl_sh_ddr0_q3.arvalid),
       .m_axi_arready  (lcl_cl_sh_ddr0_q3.arready),
       .m_axi_rid      ({10'b0, lcl_cl_sh_ddr0_q3.rid[5:0]}),    
       .m_axi_rdata    (lcl_cl_sh_ddr0_q3.rdata),  
       .m_axi_rresp    (lcl_cl_sh_ddr0_q3.rresp),  
       .m_axi_rlast    (lcl_cl_sh_ddr0_q3.rlast),  
       .m_axi_rvalid   (lcl_cl_sh_ddr0_q3.rvalid), 
       .m_axi_rready   (lcl_cl_sh_ddr0_q3.rready)
       );

   cl_tst_scrb #(.DATA_WIDTH(512),
                    .SCRB_BURST_LEN_MINUS1(SCRB_BURST_LEN_MINUS1),
                    .SCRB_MAX_ADDR(SCRB_MAX_ADDR),
                    .NO_SCRB_INST(NO_SCRB_INST)) CL_TST_DDR0 (
   
         .clk(aclk),
         .rst_n(aresetn),

         .cfg_addr(ddr0_tst_cfg_bus.addr),
         .cfg_wdata(ddr0_tst_cfg_bus.wdata),
         .cfg_wr(ddr0_tst_cfg_bus.wr),
         .cfg_rd(ddr0_tst_cfg_bus.rd),
         .tst_cfg_ack(ddr0_tst_cfg_bus.ack),
         .tst_cfg_rdata(ddr0_tst_cfg_bus.rdata),

         .slv_awid(lcl_cl_sh_ddr0_q3.awid[5:0]),
         .slv_awaddr(lcl_cl_sh_ddr0_q3.awaddr), 
         .slv_awlen(lcl_cl_sh_ddr0_q3.awlen),
         .slv_awvalid(lcl_cl_sh_ddr0_q3.awvalid),
         .slv_awuser(11'b0),
         .slv_awready(lcl_cl_sh_ddr0_q3.awready),

         .slv_wid(6'b0),
         .slv_wdata(lcl_cl_sh_ddr0_q3.wdata),
         .slv_wstrb(lcl_cl_sh_ddr0_q3.wstrb),
         .slv_wlast(lcl_cl_sh_ddr0_q3.wlast),
         .slv_wvalid(lcl_cl_sh_ddr0_q3.wvalid),
         .slv_wready(lcl_cl_sh_ddr0_q3.wready),

         .slv_bid(lcl_cl_sh_ddr0_q3.bid[5:0]),
         .slv_bresp(lcl_cl_sh_ddr0_q3.bresp),
         .slv_buser(),
         .slv_bvalid(lcl_cl_sh_ddr0_q3.bvalid),
         .slv_bready(lcl_cl_sh_ddr0_q3.bready),

         .slv_arid(lcl_cl_sh_ddr0_q3.arid[5:0]),
         .slv_araddr(lcl_cl_sh_ddr0_q3.araddr), 
         .slv_arlen(lcl_cl_sh_ddr0_q3.arlen),
         .slv_arvalid(lcl_cl_sh_ddr0_q3.arvalid),
         .slv_aruser(11'b0),
         .slv_arready(lcl_cl_sh_ddr0_q3.arready),        

         .slv_rid(lcl_cl_sh_ddr0_q3.rid[5:0]),
         .slv_rdata(lcl_cl_sh_ddr0_q3.rdata),
         .slv_rresp(lcl_cl_sh_ddr0_q3.rresp),
         .slv_rlast(lcl_cl_sh_ddr0_q3.rlast),
         .slv_ruser(),
         .slv_rvalid(lcl_cl_sh_ddr0_q3.rvalid),
         .slv_rready(lcl_cl_sh_ddr0_q3.rready),

   
         .awid(lcl_cl_sh_ddr0.awid[5:0]),
         .awaddr(lcl_cl_sh_ddr0.awaddr), 
         .awlen(lcl_cl_sh_ddr0.awlen),
         .awvalid(lcl_cl_sh_ddr0.awvalid),
         .awuser(),
         .awready(lcl_cl_sh_ddr0.awready),

         .wid(lcl_cl_sh_ddr0.wid[5:0]),
         .wdata(lcl_cl_sh_ddr0.wdata),
         .wstrb(lcl_cl_sh_ddr0.wstrb),
         .wlast(lcl_cl_sh_ddr0.wlast),
         .wvalid(lcl_cl_sh_ddr0.wvalid),
         .wready(lcl_cl_sh_ddr0.wready),

         .bid(lcl_cl_sh_ddr0.bid[5:0]),
         .bresp(lcl_cl_sh_ddr0.bresp),
         .buser(18'h0),
         .bvalid(lcl_cl_sh_ddr0.bvalid),
         .bready(lcl_cl_sh_ddr0.bready),

         .arid(lcl_cl_sh_ddr0.arid[5:0]),
         .araddr(lcl_cl_sh_ddr0.araddr),
         .arlen(lcl_cl_sh_ddr0.arlen),
         .arvalid(lcl_cl_sh_ddr0.arvalid),
         .aruser(),
         .arready(lcl_cl_sh_ddr0.arready),

         .rid(lcl_cl_sh_ddr0.rid[5:0]),
         .rdata(lcl_cl_sh_ddr0.rdata),
         .rresp(lcl_cl_sh_ddr0.rresp),
         .rlast(lcl_cl_sh_ddr0.rlast),
         .ruser(18'h0),
         .rvalid(lcl_cl_sh_ddr0.rvalid),
         .rready(lcl_cl_sh_ddr0.rready),

         .scrb_enable(ddr0_scrb_bus.enable),
         .scrb_done  (ddr0_scrb_bus.done),

         .scrb_dbg_state(ddr0_scrb_bus.state),
         .scrb_dbg_addr (ddr0_scrb_bus.addr)
      );
      assign lcl_cl_sh_ddr0.awid[15:6] = 10'b0;
      assign lcl_cl_sh_ddr0.wid[15:6] = 10'b0;
      assign lcl_cl_sh_ddr0.arid[15:6] = 10'b0;


  //back to back register slices for SLR crossing
   src_register_slice DDR1_TST_AXI4_REG_SLC_1 (
       .aclk           (aclk),
       .aresetn        (aresetn),
       .s_axi_awid     (lcl_cl_sh_ddr1_q.awid[5:0]),
       .s_axi_awaddr   ({lcl_cl_sh_ddr1_q.awaddr[63:32], 2'b0, lcl_cl_sh_ddr1_q.awaddr[29:0]}),
       .s_axi_awlen    (lcl_cl_sh_ddr1_q.awlen),
       .s_axi_awsize   (3'b110),
       .s_axi_awburst  (2'b1),
       .s_axi_awlock   (1'b0),
       .s_axi_awcache  (4'b11),
       .s_axi_awprot   (3'b10),
       .s_axi_awregion (4'b0),
       .s_axi_awqos    (4'b0),
       .s_axi_awvalid  (lcl_cl_sh_ddr1_q.awvalid),
       .s_axi_awready  (lcl_cl_sh_ddr1_q.awready),
       .s_axi_wdata    (lcl_cl_sh_ddr1_q.wdata),
       .s_axi_wstrb    (lcl_cl_sh_ddr1_q.wstrb),
       .s_axi_wlast    (lcl_cl_sh_ddr1_q.wlast),
       .s_axi_wvalid   (lcl_cl_sh_ddr1_q.wvalid),
       .s_axi_wready   (lcl_cl_sh_ddr1_q.wready),
       .s_axi_bid      (lcl_cl_sh_ddr1_q.bid[5:0]),
       .s_axi_bresp    (lcl_cl_sh_ddr1_q.bresp),
       .s_axi_bvalid   (lcl_cl_sh_ddr1_q.bvalid),
       .s_axi_bready   (lcl_cl_sh_ddr1_q.bready),
       .s_axi_arid     (lcl_cl_sh_ddr1_q.arid[5:0]),
       .s_axi_araddr   ({lcl_cl_sh_ddr1_q.araddr[63:32], 2'b0, lcl_cl_sh_ddr1_q.araddr[29:0]}),
       .s_axi_arlen    (lcl_cl_sh_ddr1_q.arlen),
       .s_axi_arsize   (3'b110),
       .s_axi_arburst  (2'b1),
       .s_axi_arlock   (1'b0),
       .s_axi_arcache  (4'b11),
       .s_axi_arprot   (3'b10),
       .s_axi_arregion (4'b0),
       .s_axi_arqos    (4'b0),
       .s_axi_arvalid  (lcl_cl_sh_ddr1_q.arvalid),
       .s_axi_arready  (lcl_cl_sh_ddr1_q.arready),
       .s_axi_rid      (lcl_cl_sh_ddr1_q.rid[5:0]),
       .s_axi_rdata    (lcl_cl_sh_ddr1_q.rdata),
       .s_axi_rresp    (lcl_cl_sh_ddr1_q.rresp),
       .s_axi_rlast    (lcl_cl_sh_ddr1_q.rlast),
       .s_axi_rvalid   (lcl_cl_sh_ddr1_q.rvalid),
       .s_axi_rready   (lcl_cl_sh_ddr1_q.rready),  
       .m_axi_awid     (lcl_cl_sh_ddr1_q2.awid[5:0]),   
       .m_axi_awaddr   (lcl_cl_sh_ddr1_q2.awaddr), 
       .m_axi_awlen    (lcl_cl_sh_ddr1_q2.awlen),  
       .m_axi_awvalid  (lcl_cl_sh_ddr1_q2.awvalid),
       .m_axi_awready  (lcl_cl_sh_ddr1_q2.awready),
       .m_axi_wdata    (lcl_cl_sh_ddr1_q2.wdata),  
       .m_axi_wstrb    (lcl_cl_sh_ddr1_q2.wstrb),  
       .m_axi_wlast    (lcl_cl_sh_ddr1_q2.wlast),  
       .m_axi_wvalid   (lcl_cl_sh_ddr1_q2.wvalid), 
       .m_axi_wready   (lcl_cl_sh_ddr1_q2.wready), 
       .m_axi_bid      (lcl_cl_sh_ddr1_q2.bid[5:0]),    
       .m_axi_bresp    (lcl_cl_sh_ddr1_q2.bresp),  
       .m_axi_bvalid   (lcl_cl_sh_ddr1_q2.bvalid), 
       .m_axi_bready   (lcl_cl_sh_ddr1_q2.bready), 
       .m_axi_arid     (lcl_cl_sh_ddr1_q2.arid[5:0]),   
       .m_axi_araddr   (lcl_cl_sh_ddr1_q2.araddr), 
       .m_axi_arlen    (lcl_cl_sh_ddr1_q2.arlen),  
       .m_axi_arvalid  (lcl_cl_sh_ddr1_q2.arvalid),
       .m_axi_arready  (lcl_cl_sh_ddr1_q2.arready),
       .m_axi_rid      (lcl_cl_sh_ddr1_q2.rid[5:0]),    
       .m_axi_rdata    (lcl_cl_sh_ddr1_q2.rdata),  
       .m_axi_rresp    (lcl_cl_sh_ddr1_q2.rresp),  
       .m_axi_rlast    (lcl_cl_sh_ddr1_q2.rlast),  
       .m_axi_rvalid   (lcl_cl_sh_ddr1_q2.rvalid), 
       .m_axi_rready   (lcl_cl_sh_ddr1_q2.rready)
       );
   dest_register_slice DDR1_TST_AXI4_REG_SLC_2 (
       .aclk           (aclk),
       .aresetn        (aresetn),
       .s_axi_awid     (lcl_cl_sh_ddr1_q2.awid),
       .s_axi_awaddr   (lcl_cl_sh_ddr1_q2.awaddr),
       .s_axi_awlen    (lcl_cl_sh_ddr1_q2.awlen),
       .s_axi_awsize   (3'b110),
       .s_axi_awburst  (2'b1),
       .s_axi_awlock   (1'b0),
       .s_axi_awcache  (4'b11),
       .s_axi_awprot   (3'b10),
       .s_axi_awregion (4'b0),
       .s_axi_awqos    (4'b0),
       .s_axi_awvalid  (lcl_cl_sh_ddr1_q2.awvalid),
       .s_axi_awready  (lcl_cl_sh_ddr1_q2.awready),
       .s_axi_wdata    (lcl_cl_sh_ddr1_q2.wdata),
       .s_axi_wstrb    (lcl_cl_sh_ddr1_q2.wstrb),
       .s_axi_wlast    (lcl_cl_sh_ddr1_q2.wlast),
       .s_axi_wvalid   (lcl_cl_sh_ddr1_q2.wvalid),
       .s_axi_wready   (lcl_cl_sh_ddr1_q2.wready),
       .s_axi_bid      (lcl_cl_sh_ddr1_q2.bid),
       .s_axi_bresp    (lcl_cl_sh_ddr1_q2.bresp),
       .s_axi_bvalid   (lcl_cl_sh_ddr1_q2.bvalid),
       .s_axi_bready   (lcl_cl_sh_ddr1_q2.bready),
       .s_axi_arid     (lcl_cl_sh_ddr1_q2.arid),
       .s_axi_araddr   (lcl_cl_sh_ddr1_q2.araddr),
       .s_axi_arlen    (lcl_cl_sh_ddr1_q2.arlen),
       .s_axi_arsize   (3'b110),
       .s_axi_arburst  (2'b1),
       .s_axi_arlock   (1'b0),
       .s_axi_arcache  (4'b11),
       .s_axi_arprot   (3'b10),
       .s_axi_arregion (4'b0),
       .s_axi_arqos    (4'b0),
       .s_axi_arvalid  (lcl_cl_sh_ddr1_q2.arvalid),
       .s_axi_arready  (lcl_cl_sh_ddr1_q2.arready),
       .s_axi_rid      (lcl_cl_sh_ddr1_q2.rid),
       .s_axi_rdata    (lcl_cl_sh_ddr1_q2.rdata),
       .s_axi_rresp    (lcl_cl_sh_ddr1_q2.rresp),
       .s_axi_rlast    (lcl_cl_sh_ddr1_q2.rlast),
       .s_axi_rvalid   (lcl_cl_sh_ddr1_q2.rvalid),
       .s_axi_rready   (lcl_cl_sh_ddr1_q2.rready),  
       .m_axi_awid     (lcl_cl_sh_ddr1_q3.awid),   
       .m_axi_awaddr   (lcl_cl_sh_ddr1_q3.awaddr), 
       .m_axi_awlen    (lcl_cl_sh_ddr1_q3.awlen),  
       .m_axi_awvalid  (lcl_cl_sh_ddr1_q3.awvalid),
       .m_axi_awready  (lcl_cl_sh_ddr1_q3.awready),
       .m_axi_wdata    (lcl_cl_sh_ddr1_q3.wdata),  
       .m_axi_wstrb    (lcl_cl_sh_ddr1_q3.wstrb),  
       .m_axi_wlast    (lcl_cl_sh_ddr1_q3.wlast),  
       .m_axi_wvalid   (lcl_cl_sh_ddr1_q3.wvalid), 
       .m_axi_wready   (lcl_cl_sh_ddr1_q3.wready), 
       .m_axi_bid      ({10'b0, lcl_cl_sh_ddr1_q3.bid[5:0]}),    
       .m_axi_bresp    (lcl_cl_sh_ddr1_q3.bresp),  
       .m_axi_bvalid   (lcl_cl_sh_ddr1_q3.bvalid), 
       .m_axi_bready   (lcl_cl_sh_ddr1_q3.bready), 
       .m_axi_arid     (lcl_cl_sh_ddr1_q3.arid),   
       .m_axi_araddr   (lcl_cl_sh_ddr1_q3.araddr), 
       .m_axi_arlen    (lcl_cl_sh_ddr1_q3.arlen),  
       .m_axi_arvalid  (lcl_cl_sh_ddr1_q3.arvalid),
       .m_axi_arready  (lcl_cl_sh_ddr1_q3.arready),
       .m_axi_rid      ({10'b0, lcl_cl_sh_ddr1_q3.rid[5:0]}),    
       .m_axi_rdata    (lcl_cl_sh_ddr1_q3.rdata),  
       .m_axi_rresp    (lcl_cl_sh_ddr1_q3.rresp),  
       .m_axi_rlast    (lcl_cl_sh_ddr1_q3.rlast),  
       .m_axi_rvalid   (lcl_cl_sh_ddr1_q3.rvalid), 
       .m_axi_rready   (lcl_cl_sh_ddr1_q3.rready)
       );

   cl_tst_scrb #(.DATA_WIDTH(512),
                    .SCRB_BURST_LEN_MINUS1(SCRB_BURST_LEN_MINUS1),
                    .SCRB_MAX_ADDR(SCRB_MAX_ADDR),
                    .NO_SCRB_INST(NO_SCRB_INST)) CL_TST_DDR1 (
   
         .clk(aclk),
         .rst_n(aresetn),

         .cfg_addr(ddr1_tst_cfg_bus.addr),
         .cfg_wdata(ddr1_tst_cfg_bus.wdata),
         .cfg_wr(ddr1_tst_cfg_bus.wr),
         .cfg_rd(ddr1_tst_cfg_bus.rd),
         .tst_cfg_ack(ddr1_tst_cfg_bus.ack),
         .tst_cfg_rdata(ddr1_tst_cfg_bus.rdata),

         .slv_awid(lcl_cl_sh_ddr1_q3.awid[5:0]),
         .slv_awaddr(lcl_cl_sh_ddr1_q3.awaddr), 
         .slv_awlen(lcl_cl_sh_ddr1_q3.awlen),
         .slv_awvalid(lcl_cl_sh_ddr1_q3.awvalid),
         .slv_awuser(11'b0),
         .slv_awready(lcl_cl_sh_ddr1_q3.awready),

         .slv_wid(6'b0),
         .slv_wdata(lcl_cl_sh_ddr1_q3.wdata),
         .slv_wstrb(lcl_cl_sh_ddr1_q3.wstrb),
         .slv_wlast(lcl_cl_sh_ddr1_q3.wlast),
         .slv_wvalid(lcl_cl_sh_ddr1_q3.wvalid),
         .slv_wready(lcl_cl_sh_ddr1_q3.wready),

         .slv_bid(lcl_cl_sh_ddr1_q3.bid[5:0]),
         .slv_bresp(lcl_cl_sh_ddr1_q3.bresp),
         .slv_buser(),
         .slv_bvalid(lcl_cl_sh_ddr1_q3.bvalid),
         .slv_bready(lcl_cl_sh_ddr1_q3.bready),

         .slv_arid(lcl_cl_sh_ddr1_q3.arid[5:0]),
         .slv_araddr(lcl_cl_sh_ddr1_q3.araddr), 
         .slv_arlen(lcl_cl_sh_ddr1_q3.arlen),
         .slv_arvalid(lcl_cl_sh_ddr1_q3.arvalid),
         .slv_aruser(11'b0),
         .slv_arready(lcl_cl_sh_ddr1_q3.arready),        

         .slv_rid(lcl_cl_sh_ddr1_q3.rid[5:0]),
         .slv_rdata(lcl_cl_sh_ddr1_q3.rdata),
         .slv_rresp(lcl_cl_sh_ddr1_q3.rresp),
         .slv_rlast(lcl_cl_sh_ddr1_q3.rlast),
         .slv_ruser(),
         .slv_rvalid(lcl_cl_sh_ddr1_q3.rvalid),
         .slv_rready(lcl_cl_sh_ddr1_q3.rready),

   
         .awid(lcl_cl_sh_ddr1.awid[5:0]),
         .awaddr(lcl_cl_sh_ddr1.awaddr), 
         .awlen(lcl_cl_sh_ddr1.awlen),
         .awvalid(lcl_cl_sh_ddr1.awvalid),
         .awuser(),
         .awready(lcl_cl_sh_ddr1.awready),

         .wid(lcl_cl_sh_ddr1.wid[5:0]),
         .wdata(lcl_cl_sh_ddr1.wdata),
         .wstrb(lcl_cl_sh_ddr1.wstrb),
         .wlast(lcl_cl_sh_ddr1.wlast),
         .wvalid(lcl_cl_sh_ddr1.wvalid),
         .wready(lcl_cl_sh_ddr1.wready),

         .bid(lcl_cl_sh_ddr1.bid[5:0]),
         .bresp(lcl_cl_sh_ddr1.bresp),
         .buser(18'h0),
         .bvalid(lcl_cl_sh_ddr1.bvalid),
         .bready(lcl_cl_sh_ddr1.bready),

         .arid(lcl_cl_sh_ddr1.arid[5:0]),
         .araddr(lcl_cl_sh_ddr1.araddr),
         .arlen(lcl_cl_sh_ddr1.arlen),
         .arvalid(lcl_cl_sh_ddr1.arvalid),
         .aruser(),
         .arready(lcl_cl_sh_ddr1.arready),

         .rid(lcl_cl_sh_ddr1.rid[5:0]),
         .rdata(lcl_cl_sh_ddr1.rdata),
         .rresp(lcl_cl_sh_ddr1.rresp),
         .rlast(lcl_cl_sh_ddr1.rlast),
         .ruser(18'h0),
         .rvalid(lcl_cl_sh_ddr1.rvalid),
         .rready(lcl_cl_sh_ddr1.rready),

         .scrb_enable(ddr1_scrb_bus.enable),
         .scrb_done  (ddr1_scrb_bus.done),

         .scrb_dbg_state(ddr1_scrb_bus.state),
         .scrb_dbg_addr (ddr1_scrb_bus.addr)
      );
      assign lcl_cl_sh_ddr1.awid[15:6] = 10'b0;
      assign lcl_cl_sh_ddr1.wid[15:6] = 10'b0;
      assign lcl_cl_sh_ddr1.arid[15:6] = 10'b0;



  //back to back register slices for SLR crossing
   src_register_slice DDR2_TST_AXI4_REG_SLC_1 (
       .aclk           (aclk),
       .aresetn        (aresetn),
       .s_axi_awid     (lcl_cl_sh_ddr2_q.awid[5:0]),
       .s_axi_awaddr   ({lcl_cl_sh_ddr2_q.awaddr[63:32], 2'b0, lcl_cl_sh_ddr2_q.awaddr[29:0]}),
       .s_axi_awlen    (lcl_cl_sh_ddr2_q.awlen),
       .s_axi_awsize   (3'b110),
       .s_axi_awburst  (2'b1),
       .s_axi_awlock   (1'b0),
       .s_axi_awcache  (4'b11),
       .s_axi_awprot   (3'b10),
       .s_axi_awregion (4'b0),
       .s_axi_awqos    (4'b0),
       .s_axi_awvalid  (lcl_cl_sh_ddr2_q.awvalid),
       .s_axi_awready  (lcl_cl_sh_ddr2_q.awready),
       .s_axi_wdata    (lcl_cl_sh_ddr2_q.wdata),
       .s_axi_wstrb    (lcl_cl_sh_ddr2_q.wstrb),
       .s_axi_wlast    (lcl_cl_sh_ddr2_q.wlast),
       .s_axi_wvalid   (lcl_cl_sh_ddr2_q.wvalid),
       .s_axi_wready   (lcl_cl_sh_ddr2_q.wready),
       .s_axi_bid      (lcl_cl_sh_ddr2_q.bid[5:0]),
       .s_axi_bresp    (lcl_cl_sh_ddr2_q.bresp),
       .s_axi_bvalid   (lcl_cl_sh_ddr2_q.bvalid),
       .s_axi_bready   (lcl_cl_sh_ddr2_q.bready),
       .s_axi_arid     (lcl_cl_sh_ddr2_q.arid[5:0]),
       .s_axi_araddr   ({lcl_cl_sh_ddr2_q.araddr[63:32], 2'b0, lcl_cl_sh_ddr2_q.araddr[29:0]}),
       .s_axi_arlen    (lcl_cl_sh_ddr2_q.arlen),
       .s_axi_arsize   (3'b110),
       .s_axi_arburst  (2'b1),
       .s_axi_arlock   (1'b0),
       .s_axi_arcache  (4'b11),
       .s_axi_arprot   (3'b10),
       .s_axi_arregion (4'b0),
       .s_axi_arqos    (4'b0),
       .s_axi_arvalid  (lcl_cl_sh_ddr2_q.arvalid),
       .s_axi_arready  (lcl_cl_sh_ddr2_q.arready),
       .s_axi_rid      (lcl_cl_sh_ddr2_q.rid[5:0]),
       .s_axi_rdata    (lcl_cl_sh_ddr2_q.rdata),
       .s_axi_rresp    (lcl_cl_sh_ddr2_q.rresp),
       .s_axi_rlast    (lcl_cl_sh_ddr2_q.rlast),
       .s_axi_rvalid   (lcl_cl_sh_ddr2_q.rvalid),
       .s_axi_rready   (lcl_cl_sh_ddr2_q.rready),  
       .m_axi_awid     (lcl_cl_sh_ddr2_q2.awid[5:0]),   
       .m_axi_awaddr   (lcl_cl_sh_ddr2_q2.awaddr), 
       .m_axi_awlen    (lcl_cl_sh_ddr2_q2.awlen),  
       .m_axi_awvalid  (lcl_cl_sh_ddr2_q2.awvalid),
       .m_axi_awready  (lcl_cl_sh_ddr2_q2.awready),
       .m_axi_wdata    (lcl_cl_sh_ddr2_q2.wdata),  
       .m_axi_wstrb    (lcl_cl_sh_ddr2_q2.wstrb),  
       .m_axi_wlast    (lcl_cl_sh_ddr2_q2.wlast),  
       .m_axi_wvalid   (lcl_cl_sh_ddr2_q2.wvalid), 
       .m_axi_wready   (lcl_cl_sh_ddr2_q2.wready), 
       .m_axi_bid      (lcl_cl_sh_ddr2_q2.bid[5:0]),    
       .m_axi_bresp    (lcl_cl_sh_ddr2_q2.bresp),  
       .m_axi_bvalid   (lcl_cl_sh_ddr2_q2.bvalid), 
       .m_axi_bready   (lcl_cl_sh_ddr2_q2.bready), 
       .m_axi_arid     (lcl_cl_sh_ddr2_q2.arid[5:0]),   
       .m_axi_araddr   (lcl_cl_sh_ddr2_q2.araddr), 
       .m_axi_arlen    (lcl_cl_sh_ddr2_q2.arlen),  
       .m_axi_arvalid  (lcl_cl_sh_ddr2_q2.arvalid),
       .m_axi_arready  (lcl_cl_sh_ddr2_q2.arready),
       .m_axi_rid      (lcl_cl_sh_ddr2_q2.rid[5:0]),    
       .m_axi_rdata    (lcl_cl_sh_ddr2_q2.rdata),  
       .m_axi_rresp    (lcl_cl_sh_ddr2_q2.rresp),  
       .m_axi_rlast    (lcl_cl_sh_ddr2_q2.rlast),  
       .m_axi_rvalid   (lcl_cl_sh_ddr2_q2.rvalid), 
       .m_axi_rready   (lcl_cl_sh_ddr2_q2.rready)
       );
   dest_register_slice DDR2_TST_AXI4_REG_SLC_2 (
       .aclk           (aclk),
       .aresetn        (aresetn),
       .s_axi_awid     (lcl_cl_sh_ddr2_q2.awid),
       .s_axi_awaddr   (lcl_cl_sh_ddr2_q2.awaddr),
       .s_axi_awlen    (lcl_cl_sh_ddr2_q2.awlen),
       .s_axi_awsize   (3'b110),
       .s_axi_awburst  (2'b1),
       .s_axi_awlock   (1'b0),
       .s_axi_awcache  (4'b11),
       .s_axi_awprot   (3'b10),
       .s_axi_awregion (4'b0),
       .s_axi_awqos    (4'b0),
       .s_axi_awvalid  (lcl_cl_sh_ddr2_q2.awvalid),
       .s_axi_awready  (lcl_cl_sh_ddr2_q2.awready),
       .s_axi_wdata    (lcl_cl_sh_ddr2_q2.wdata),
       .s_axi_wstrb    (lcl_cl_sh_ddr2_q2.wstrb),
       .s_axi_wlast    (lcl_cl_sh_ddr2_q2.wlast),
       .s_axi_wvalid   (lcl_cl_sh_ddr2_q2.wvalid),
       .s_axi_wready   (lcl_cl_sh_ddr2_q2.wready),
       .s_axi_bid      (lcl_cl_sh_ddr2_q2.bid),
       .s_axi_bresp    (lcl_cl_sh_ddr2_q2.bresp),
       .s_axi_bvalid   (lcl_cl_sh_ddr2_q2.bvalid),
       .s_axi_bready   (lcl_cl_sh_ddr2_q2.bready),
       .s_axi_arid     (lcl_cl_sh_ddr2_q2.arid),
       .s_axi_araddr   (lcl_cl_sh_ddr2_q2.araddr),
       .s_axi_arlen    (lcl_cl_sh_ddr2_q2.arlen),
       .s_axi_arsize   (3'b110),
       .s_axi_arburst  (2'b1),
       .s_axi_arlock   (1'b0),
       .s_axi_arcache  (4'b11),
       .s_axi_arprot   (3'b10),
       .s_axi_arregion (4'b0),
       .s_axi_arqos    (4'b0),
       .s_axi_arvalid  (lcl_cl_sh_ddr2_q2.arvalid),
       .s_axi_arready  (lcl_cl_sh_ddr2_q2.arready),
       .s_axi_rid      (lcl_cl_sh_ddr2_q2.rid),
       .s_axi_rdata    (lcl_cl_sh_ddr2_q2.rdata),
       .s_axi_rresp    (lcl_cl_sh_ddr2_q2.rresp),
       .s_axi_rlast    (lcl_cl_sh_ddr2_q2.rlast),
       .s_axi_rvalid   (lcl_cl_sh_ddr2_q2.rvalid),
       .s_axi_rready   (lcl_cl_sh_ddr2_q2.rready),  
       .m_axi_awid     (lcl_cl_sh_ddr2_q3.awid),   
       .m_axi_awaddr   (lcl_cl_sh_ddr2_q3.awaddr), 
       .m_axi_awlen    (lcl_cl_sh_ddr2_q3.awlen),  
       .m_axi_awvalid  (lcl_cl_sh_ddr2_q3.awvalid),
       .m_axi_awready  (lcl_cl_sh_ddr2_q3.awready),
       .m_axi_wdata    (lcl_cl_sh_ddr2_q3.wdata),  
       .m_axi_wstrb    (lcl_cl_sh_ddr2_q3.wstrb),  
       .m_axi_wlast    (lcl_cl_sh_ddr2_q3.wlast),  
       .m_axi_wvalid   (lcl_cl_sh_ddr2_q3.wvalid), 
       .m_axi_wready   (lcl_cl_sh_ddr2_q3.wready), 
       .m_axi_bid      ({10'b0, lcl_cl_sh_ddr2_q3.bid[5:0]}),    
       .m_axi_bresp    (lcl_cl_sh_ddr2_q3.bresp),  
       .m_axi_bvalid   (lcl_cl_sh_ddr2_q3.bvalid), 
       .m_axi_bready   (lcl_cl_sh_ddr2_q3.bready), 
       .m_axi_arid     (lcl_cl_sh_ddr2_q3.arid),   
       .m_axi_araddr   (lcl_cl_sh_ddr2_q3.araddr), 
       .m_axi_arlen    (lcl_cl_sh_ddr2_q3.arlen),  
       .m_axi_arvalid  (lcl_cl_sh_ddr2_q3.arvalid),
       .m_axi_arready  (lcl_cl_sh_ddr2_q3.arready),
       .m_axi_rid      ({10'b0, lcl_cl_sh_ddr2_q3.rid[5:0]}),    
       .m_axi_rdata    (lcl_cl_sh_ddr2_q3.rdata),  
       .m_axi_rresp    (lcl_cl_sh_ddr2_q3.rresp),  
       .m_axi_rlast    (lcl_cl_sh_ddr2_q3.rlast),  
       .m_axi_rvalid   (lcl_cl_sh_ddr2_q3.rvalid), 
       .m_axi_rready   (lcl_cl_sh_ddr2_q3.rready)
       );

   cl_tst_scrb #(.DATA_WIDTH(512),
                    .SCRB_BURST_LEN_MINUS1(SCRB_BURST_LEN_MINUS1),
                    .SCRB_MAX_ADDR(SCRB_MAX_ADDR),
                    .NO_SCRB_INST(NO_SCRB_INST)) CL_TST_DDR2 (
   
         .clk(aclk),
         .rst_n(aresetn),

         .cfg_addr(ddr3_tst_cfg_bus.addr),
         .cfg_wdata(ddr3_tst_cfg_bus.wdata),
         .cfg_wr(ddr3_tst_cfg_bus.wr),
         .cfg_rd(ddr3_tst_cfg_bus.rd),
         .tst_cfg_ack(ddr3_tst_cfg_bus.ack),
         .tst_cfg_rdata(ddr3_tst_cfg_bus.rdata),

         .slv_awid(lcl_cl_sh_ddr2_q3.awid[5:0]),
         .slv_awaddr(lcl_cl_sh_ddr2_q3.awaddr), 
         .slv_awlen(lcl_cl_sh_ddr2_q3.awlen),
         .slv_awvalid(lcl_cl_sh_ddr2_q3.awvalid),
         .slv_awuser(11'b0),
         .slv_awready(lcl_cl_sh_ddr2_q3.awready),

         .slv_wid(6'b0),
         .slv_wdata(lcl_cl_sh_ddr2_q3.wdata),
         .slv_wstrb(lcl_cl_sh_ddr2_q3.wstrb),
         .slv_wlast(lcl_cl_sh_ddr2_q3.wlast),
         .slv_wvalid(lcl_cl_sh_ddr2_q3.wvalid),
         .slv_wready(lcl_cl_sh_ddr2_q3.wready),

         .slv_bid(lcl_cl_sh_ddr2_q3.bid[5:0]),
         .slv_bresp(lcl_cl_sh_ddr2_q3.bresp),
         .slv_buser(),
         .slv_bvalid(lcl_cl_sh_ddr2_q3.bvalid),
         .slv_bready(lcl_cl_sh_ddr2_q3.bready),

         .slv_arid(lcl_cl_sh_ddr2_q3.arid[5:0]),
         .slv_araddr(lcl_cl_sh_ddr2_q3.araddr), 
         .slv_arlen(lcl_cl_sh_ddr2_q3.arlen),
         .slv_arvalid(lcl_cl_sh_ddr2_q3.arvalid),
         .slv_aruser(11'b0),
         .slv_arready(lcl_cl_sh_ddr2_q3.arready),        

         .slv_rid(lcl_cl_sh_ddr2_q3.rid[5:0]),
         .slv_rdata(lcl_cl_sh_ddr2_q3.rdata),
         .slv_rresp(lcl_cl_sh_ddr2_q3.rresp),
         .slv_rlast(lcl_cl_sh_ddr2_q3.rlast),
         .slv_ruser(),
         .slv_rvalid(lcl_cl_sh_ddr2_q3.rvalid),
         .slv_rready(lcl_cl_sh_ddr2_q3.rready),

   
         .awid(lcl_cl_sh_ddr2.awid[5:0]),
         .awaddr(lcl_cl_sh_ddr2.awaddr), 
         .awlen(lcl_cl_sh_ddr2.awlen),
         .awvalid(lcl_cl_sh_ddr2.awvalid),
         .awuser(),
         .awready(lcl_cl_sh_ddr2.awready),

         .wid(lcl_cl_sh_ddr2.wid[5:0]),
         .wdata(lcl_cl_sh_ddr2.wdata),
         .wstrb(lcl_cl_sh_ddr2.wstrb),
         .wlast(lcl_cl_sh_ddr2.wlast),
         .wvalid(lcl_cl_sh_ddr2.wvalid),
         .wready(lcl_cl_sh_ddr2.wready),

         .bid(lcl_cl_sh_ddr2.bid[5:0]),
         .bresp(lcl_cl_sh_ddr2.bresp),
         .buser(18'h0),
         .bvalid(lcl_cl_sh_ddr2.bvalid),
         .bready(lcl_cl_sh_ddr2.bready),

         .arid(lcl_cl_sh_ddr2.arid[5:0]),
         .araddr(lcl_cl_sh_ddr2.araddr),
         .arlen(lcl_cl_sh_ddr2.arlen),
         .arvalid(lcl_cl_sh_ddr2.arvalid),
         .aruser(),
         .arready(lcl_cl_sh_ddr2.arready),

         .rid(lcl_cl_sh_ddr2.rid[5:0]),
         .rdata(lcl_cl_sh_ddr2.rdata),
         .rresp(lcl_cl_sh_ddr2.rresp),
         .rlast(lcl_cl_sh_ddr2.rlast),
         .ruser(18'h0),
         .rvalid(lcl_cl_sh_ddr2.rvalid),
         .rready(lcl_cl_sh_ddr2.rready),

         .scrb_enable(ddr3_scrb_bus.enable),
         .scrb_done  (ddr3_scrb_bus.done),

         .scrb_dbg_state(ddr3_scrb_bus.state),
         .scrb_dbg_addr (ddr3_scrb_bus.addr)
      );
      assign lcl_cl_sh_ddr2.awid[15:6] = 10'b0;
      assign lcl_cl_sh_ddr2.wid[15:6] = 10'b0;
      assign lcl_cl_sh_ddr2.arid[15:6] = 10'b0;


endmodule

