`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
ha1tMYw+ceIaAaE/e/beNYUiddD/aqwf8lYMP3p88/D0lWcuJesqIP/692OUSJKb4QyENY/p2llD
+oBBIVPomLp1/jrlbLchOvp/BbYuritBPZ82XIOLMRobOr87ZKx7e0JKXFjTqk9T703J0Pw0z8IO
ZwwYaHt7ZhnruYXudmuhOrPM9AJ8tRCDYMoU0DZxwtPhs51QYegupV1bW5jntdpadbu2e2iGLwCE
BIScvw8qwhmYxALxE/6kGCnyHdhvSKa0wxSF+u30EANFL/TiKQ+CacTdDdOj804Mqu6QCBUQ6ypE
7sSH1IvfWvsJc9j3fKWmR9tJuskwkmCQYr/2Yw==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
hZlP1AvojUOk4uzW2R5Y1fRAzLNBWOkVZ0BEEnNXMkkNT+kXU1lh0LJqNec7SgrLeBYfgeOkGtiU
ojx99vyPT6x+rVWlKSVbXi98/yZtSYIlUYiccNpG2HKB1bWm966cm/2T6OcnD1mTXkNrWxABpZeW
WjUEQ8KoPlH6EbTtXWs=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
D78YQBUWw89jvnnAYC7uc2hI4ogEXAdRCYJktkjyQ6iMULCrMU0tJuBchUAWfDj98kHLA0sj0W/F
S0CCyzGLNvjFyBTtbFTShUCofUvNEwbpXr3R8aZeIAelI5pUoXTTM3y9YC5YRFxjyNw0tatjuEOJ
/EfcxVlHqFGmV2V+FWY=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2688)
`pragma protect data_block
vBqXsBG7U2RW2eNvrfnuHIhck/wcmGHm1TblkRjQLuuIC4rVGKFACn/WWnSV9mn15huHNYxr/Jxt
lTAsAZPJ7j29/PWn0oyD9Uxx8IkaqSnNbFyMbygZt7We8Fuk9MHz+mWfJHPC6ySqrvLiy9VZ4aZe
+6r6nMM84a5nKZsa/Y8SA8AWoB3GIJBByuO5cpxaV62KVlLC1uto5RfKSHXDudGEWMfFt86fH4pu
UeNNhORGFIy/SKongRN+g7H3Ce9D9dX5KYHz/PnlfjOzxvklf09+WxuY2oqJUUgqZQNC8iFvhP3k
AiOm95kdl1dWjuxMvpyPge/3rnKdAUThC/LIHMJFSQkROxXfpkLt+Zz8Ligij+69xPzmYyWh5B6B
hRsnBW7PZ6JQ1wO5ZNKnMOm5yJOvyUDzcEPQ8yALlUvli7h89xZ8Qtvo1DZj8VO16X608J119KVq
BheGM0yecbDCbEJ9L/aY/XRHSkWetJ8uCzP1MTH+f24GEnHg00VqD7YIzfRqBBPTT6jACMbCiRgB
ITZtrmotGRa0jEHffj+hEpKMbJ1d165gm0FP4WxoGDFjiwAQUmnk2XzLUJfILu8mmbfBzRhvpGuR
6KBWhxh5z6W9H8y05F6WOfUzaXLxWescerAUxUupR5IjBK30rZbCn5JBCi7lbEpyM2ihaEwB+K9i
JEO0hBrOiT6ZOBd02gIPONyCtb5owfJLECutJUYR904q/dOF5iUFrsdybBNG491I/TWbll4O3VoB
IwlSAocdE24eZdDrebu3xQzOZbzgXGRopYlRx/SEvj7N1/vZ18hkwXn8vjUy33pPh1y9NSr0Yb5j
EuAJgYrhG3M9MvGttCcEYTlerj2r3OT7gNatGimwfgsI1GFl08uNAlRy+UQNu3pQpSat84bmg4Zb
BIsjx56AxLt1QvZrs8tWO+mCr9JPeoy0r2f/Vaak2J+gSAnPCmQiuDiBCrSlU6Em3tbIQiv+Qyg8
wXHuvFuDkPJXoVYi1mdiWGflhiRGw9xE5jkp/yryZK9pgGPFWxn0lBZ2Wm6Fw/n/2LSEeiUehP9Q
RhfgEAjIKUgpFu1QOYyto3A89wMs2ykL4fiD/iutdSMTW8k7/v1M/m1rZlrhbY74TxktWuq+M3KS
QxHijZ9dD/JnMeH1k5QnTX4aNMTS9VDzDGU/aOAJpCwd6PvelLU7rXzyJN4Iliv+2O1s6hUGGwTN
2AaKJ+sc8jK83QBkCD5WgyYln0Rk01mpoit2rPFB02iKiFNPWKbVFSZSAcL4LE3Ssof4dOcNjj5J
rbrhsHsq7EkZ9rIch6VweABgo22aXW0qUBVe0i+4jm/hsOIVuhEoqQz/CyrMcIpJiXIKmMVJw9hj
cYf+ojGcdGIzDV2Jwg/6YrYphTSuqNc/LC3SLk5KaZ6rClfs3+miy7kRBdBb+52MYbE9gkPyvWrS
exSLwwNoMAT+6YqyUzsG4DrS2nVApWzlWGrQM18p2DDv8Bcc9GNPotfofoy69W42QMKGPeKFalt8
IBEGtsGZWzYX14bw0bg87sY6KkOSUe+2FjJ8/N3tMqjhLHeSp91+WHAkYwOe7GHGCCg465RyCCyC
C3BHZtM8WCMtrjbmbVJKWOQqBA0CoOTrmdtSaTxkfnpNQ2HFCXV9No+yQCFh13Q+tW7V/LLThdVp
RVchYo+RQvHj9DZSZtCjOhpcRBCQGu5jm3g4M41ahCHyD6/6xZaoXJX0Y0fNsGoqVYQzs3W84r50
Sc41pll2liUNJ0CWvKz+tjwvCnJ2sY8UntRmqb5adcuvsCRE17Y9T+OO7q7pDmgMuVKvWsv44+i5
S1IV5AMHJSOZzFgNxrydiqQyR4DUlX8j0MeBwHhzfO/NZiGciviQarfUq2SzsjHVVW0MTnzyM8ZB
QatuZv5+AOrI6Lbvky8/xF7ytQ/XzAmXUQJ5QgskmEJRxJ02VlpnmRoX+iFzYF2VPSR9CHKcauTu
EdSnzDMCRSHtXc0qSrD3fLyqF6zOavE4VPC2HI2Gl4tct/JwKMpU5NayVz53SX7/0PZj53CdHCGH
Ay7WfdMeJgD0V6RHraMIzc11n3ynczs8ccg0lpE42uqXygnN8GQYptDw1d1VDln0IeTwnqsLGM/S
ewQZCx1urLAUujhdcM0d4TnmeDpP+uYv2DgRaabDYp4ZFjYCa0Y1ewBdZ/nD2YJX53iJcLqvNFQy
PzOZYSRTYCuExpoChauVyhV6fDGHJNLESlz8Yy0qG8Ei/5eyqXiW4XNEN+ab5I76QtzulV4Hz3Fx
iBio/LCl1yZKQj6bC0Aaf/en5NIjb67LjRLC4SbGdRLscgu1z0qsiYTZM+joxsdjwJ5OVY3bQ/5O
sFMfrBv+NZ9Lc1SBU7bvlCKlAIXwAoHVHKBUQ9QtRn70RVwyv6hf0Q54kQtEGA+1dnYGrQEBqe9j
cmo1qy4z7rKrG1ObgMj3Vn0Fv+ry0ZPW8H4xOzqzeaxJ+52il65TO4Ib9ZAi69c1aFhdhAw5FrUg
hO6Aa+kWSNysq7MN3lqcbFSGWnZHQPEvkURFliFahsqj30/Pktk6Wrt0MF6wOJmOJzxb4ywidlfW
v+bYriv0eCZqNFf/xpOBMrBvEasF0NENqE8c6N/p34apGG+ftQcMGe+dDhfbWSPYRINJuRInR+It
cge0lufiT7htL2RPdZOBJlWxYEZdJh411CyHtIDgp9meVQv+pfrm2LoObVOCL6hNAZa6qf1WnLHO
EvB6Or5kUKnb2dlkk32l0aeqReR5D+2FXTBHffTkTbzzSbBOZo1ZHvWUelsXnrrLbB5xZvOTfugt
DJ58YHpKAXVb4K4+5NvoQWV1MZ+SdiY23hxx+7c2Mc+P/blUmHHk7wWbHYewDlrxmx/1xbWtn5v6
wsM0hg0MuKC4733Nahaw3NC0INXdWf5ds6Nxal54QOiQ2KFbl7LbOeupLczaIr+46o3ZDf+ZwxoE
X6uRoSU3lWFjWEYtsYoKp8jV7CW+LgVoWKSdJQrlTkTw6iz+7d5+rzyR7z6Lq74A1BbNfeN+WMJh
wZCiKY3wz1pPQLjMosfQpxJcYWrG4A/KqIoAkq7N4pyZFGkD5kPY+7+S/nAuuShImTPyWBnONnGu
Lb2rZIEA3MAi9sTs22FHBHRajk9e9ccxRdzcREhnWP/kzZ0HduuDlko4cSuPME1REFYDjPnts1tL
X9VruY/xpnmW9XBd0zq9bN3bBbQuBVogjrvSLfQQ6M76493C+cKY8TbENNc8dI7DFx4s446jSNk6
Mq4z48uM3L3TFpoIRaGgSre9ulxmAX5ilpJLPP7uP2C5G/h0dHrn37HAk27hsyO2M4Zy4CQXwdgt
On8UMVYpugAhICdHICmAiERP6oAsSRBb9Dlz5uC2VyjhGEWHkDFi5cTJn0xjlrHY0K7DsI9PsaIm
OJc8gHxBN/2iXAaNyk2rrPu6ZAhvtjWeSPqs9JeWdP3KsiWTIRPTf/47YxNPuC6HIfozzMzwdr8v
NAt5MMb7s8UF9h/aur8GFhJc8rOPzOkPduDZjF+ujEwS8bXT299Ehryyn1f/q7MAkMyuE9y1w8Rd
CbtSdjIUQJoY
`pragma protect end_protected
