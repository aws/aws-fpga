// Amazon FPGA Hardware Development Kit
//
// Copyright 2016 Amazon.com, Inc. or its affiliates. All Rights Reserved.
//
// Licensed under the Amazon Software License (the "License"). You may not use
// this file except in compliance with the License. A copy of the License is
// located at
//
//    http://aws.amazon.com/asl/
//
// or in the "license" file accompanying this file. This file is distributed on
// an "AS IS" BASIS, WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, express or
// implied. See the License for the specific language governing permissions and
// limitations under the License.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Gx87JJBq2wxinn9UItpQzN93HPLB8MXXRKbK2CAcry5T6/hygofNhn0nTz8ku1A9Smgpz1ZBqqh8
d5fTq8q5EbV+vCYF4XbOLJbkKwPvlPti6G/rSq39Yv7ihbn29rWoxt1ugG2RQPORLjS//jSBcw69
GlUGKbBv5thTKKp/aQI5oU4JFnHfdFXhS0JED0VtsXlsn0Ivr1+Fu9Yur3VR485qe+AqSA/BD4Ew
f1YuTokSI/H8lzu0Iq127Yr4jHecngdKDO5t8OwJKINWE5avC68LIu8vJc591iGVE2Ml+PaOU2F+
QG5G9QAwPHOY5ZjAEmv+DrzkOFs8r+RX45TTfA==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
AwmKLh7GAjEZj+X1S2vn1XsMx45y0UlPh25jZ4rrLl+ekbxc887qrj6zFFFnRXPJ0+f+v0yGLECx
0DjZCLhX64zRnxOihgh60D9CGb6FEcdaDpZQRi2X1x3l2TAklS67VequDiyt9s9zvXQKOtVKzt3L
zg0GGaerc68UEwdtnAc=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
arLDZk59TdmVAXn3Mr8ipwpe/j8p5isVfGTKmR9YJHIXzHsrbJleL2ddqfYo1nQJfNuwskCujTop
/swyavGJNNAbTU6gBMHlvzFIFKwm6UCQ/rDAsbf44iSoyKG0Vq+Il6/TAWb4kneCjay91czYorhR
zMLZl4cYdnA3tx3vD3E=

`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
j4iKvHFemFVbUFisf4iaF7vWn2BBUxfe1lj1KXguyRwvwHfhGUZM4nFjgzJeAbgOo9ZkuXNAX277
Sml3zdNWCQ==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3504)
`pragma protect data_block
FJ67Mmr3HmhMIddkBsTH00xBnJrbTASh9PQTiFaeP+Mr9KpYnJIhHFWctxvXhYWo6YP35Tu52jvc
BeSJKC23ZVvDEmsNvStPAd10WFJLihjiYW7G73CByArb/ZIbMr3K/zBs2dmPVvE+RW0EOCj4WLZK
5933+hWLuhtKJ78PiMH3otDfBc3rf8V9/MWZPnoM/Alb+07uVh+0f9q+qVIWTteVJ6viHghPOzw/
lA36CR+KSDWCMN4OCxYoRD1fsWq+8VvTZJ+6vZsAiYiuFCoT1b62f7yrsb8etUhNxKlTQ3D5jxdT
k2rVDeoUl18q5ub/Obo6iO1wOJRQZcf68vjdO57QzudIqWFyEQNIy5vWroRXkyCX1otbkMlQF9vt
Vehno5psrDWvJVu4lgt38ORl2ixBUav/8gCp62/HY21nfq5bTR23JVU28ogaVBF4d1U+aErNfbVM
sbX1QAsDhBGhD0rs7Eak368EKn6WsqqM9AP8M1/laBhdk4oIDunEjfMKwm8ywtAKNaaXL/+cWAmn
zMsE24BUDx4Zo/swJIV5DafJf+t8wqrlMV2G1tidYSMSrleUfaNBz3NsKgJ4UdF8j1HHwloejiQv
Fs21MuevSYAQUz8PhkQtxpHecTgWhMvV3LDAM1BAAii4JXQOEamH0KLVSK8DLwewBlm4ybk1EvwZ
kHlYcyoaIz3fg0dCI0BahMj6gzC0O7QN6Ox/pkAGY/95URZ+kZlrVg0xG2KZHbC6BMbTYKFOEotq
NbKP+on4yI0pUt2T7wAmYfmBltJYm69gHTKQK7m+tOwkgtzzOymdJCSSq33+xC4PRkDXmQlbTPh0
URyU+dyDiVIddTL3n/6mtMEJH9rXas9TxYeY7TIQg/6ONhHCGnWwKwYffNXG5d2Weu4WZ2ESf5zx
k0uhmI4pLmJJk88gkaC0Opv2M4b5OjpSKr/WoD2tholPQe7lPfrMEBb4ETb+yuT7JHDh2oafpHRq
05pBEYK7Vo3Q1uOg4CRi4BPD4QLeMRx/pzxRIQqLKktl9iAoRoWN2DoUKe885zZkvaLLEJxYU1KC
oZg4eGm9uOHwQrgBkaqg+6tpypXxOE5/xw1O0MiUHt2JgBnr5/RKLLMjaNbwjz1LLD8y3NtkkJXc
Iz3U0H/3iFFDx5aLy90O7B96+QNkhGU0JbBZimjHKECEPKuVimykASmJvWHPWytc9AGx7BNUIVHT
rabXhvBi5MzSTYd2hnmWSvTs1lhHozlC/tqWrnZZ+cdEdhhoQf3vnytE0CgQ0bKwp0bap+HyGS8W
wQXMkRWHMs89hCJk4DfscldpvgoQfOe0A/kLkgimRIRPL8N0KnOrtMCOdrT+Udu9D9b6BMMneK+D
6ZEba4LJ+dyTIsOw9wBbxE+Q9EynvvmhMeBAWvPfyqjNNEur0DaTvyM5ZsXnaPFHTQQ9Dh209UGG
eULGseNthcdxo96Gg8JrtUsStJgBpDR+wHSDwnfzU/LUKBAPtjz+Yr6qIDW69Cas5kPNdL+iefsO
xqRkl4OtxejziTWiZ9NL2E25qxc+L+9nnRlqbv2zVrKyzf1jC5ZaXvuxJSYapjLjL/tAJIy4zyo0
Riwn6Xmgc19cI6JlynIErAgRjvD7S0n1cfJCI7c9yW+V1gtSvYP5tZu9pat+70hsom8ZS+Dnndkp
/Pfktuo5IEvgsTzHo1EUujs3X0KRtY1RRe20pOq5fU0ALEB9Jpl0diBSZa2mqskbuqIktaCDY+b0
xaYcH/W+ZLaoBEvdJTVWOkOonlxkrIXVVTd60PkKsVTwSE1uBdppPxXfXiQfXYMvTfa4kLZGsiYb
sGb3RynkyLUEH42dwFSOAN+EE6uGN7auYpm3GO9xF2P/0CWmizOXwlUWl46vkSX5Ip8Y/U0BA8wT
7KgAG7/8q8MtRCi+KjmxXs8nrlN8WcxPbbnbcvGkAji1giCM6pbwO73KcdnouqF9pxbjLdENYPMO
uwQ5iWSrBbsqO7OCXEpu0wN8tUPmnL48DPNj5PfqmnU/skaeJJvVVkKHEucO7Ui77/J4N77yvAba
sQzhaSmXYOwZwtp5tg4mYNds7+/NLorQX2VkbHoNrM4+mYP9bxbPq/mFNsRFASmz5axzQ0Us7W0l
fvpWHAC1rbuATPFOqCpTVGDsj0mZUJSJKyLmoLT3rlq01esoPrChI++2MzPjGI487fCN6GobxuiM
mrI1CxBXOq5AR2aRX5jmu5mq/mHEiu3RXGGRLDCsihr4W+Ci6RUK2yp4G7wL/BoGgWBdpAPHGVfb
0O6KFkKTAZAfnozEdWNi/y3rNtCHnkxf3HgkI26VpwVvRbrEwZE+UxWqMZ09tqQoNc2rJHTgPRMt
Xb5op09CYJjUSufXNNqK1vgjEkAud1WW4ZitcoxGBD8qonYcn9OmH9w1RMQIpmVNcyv3vOKBPqcT
mc8mDUm5CAljnIG2P68C+d/TSW09lDiyuJg2ltfvstfXJxLGjnwB+uK7ffWsNU4USbskdZ8DCk10
Ncp26r7oeT+e39aaSiyXEUooPwpcQvc747NTwjwQ+u4UHzPycXqvf9uEqt5Z61C+HoT+UaZMRSPC
kyS8ALkp08C/ZAkO66NbHfm6ZsP+zAqg0gvZIFssJqrUNTDgUEzgD38qW5/EDgO/3rfkCfrtqetu
FXvjuwWggNclm/slRdo/Vgc/43aMEGzdQOArn1rsiXZYXKfDQppCDN+ZbWFmbdupfVZ8Bfyi80Yq
nUt8EkWXlIKZve3JBeWsjxX8/Cg8oWVnoCQFk1gwjEgtCFyGGQbNYXz4dqlEEn/7bm3ZbxtFhvLK
5QyTW8c1fpQnKOktpsxeM7WDAy3HwGCUU+pnvUYoy3nMjtdJDyFt7gQmwFl6rbG3M0oZLl//nxzM
jC70+glMQfg7UTYn4Q5nwwd/qQsNsBZvdNnY50+ROeUqrN5x1Pq1mSEfhuaGIUO5M8EbHaJQemfz
PLgGq/uhYOMJj1a7mpgl8A6nN6thqg4CaQ0xLsnUeG1vFt/zXOESlSSmmuyc8T2wNb09Y056VEF/
1eqHCEtoowtc0w+PE0xJDnhuUYTQX9jNw8cg1LKcYjFSbW38g9YpbuFQIsAfDlOkJlx0ghk4oxiH
HY/Mj9vp8+D8UwBPiYSX2vXhsYHHnlILHsmoq/D8iYluwvAZXYl3E2kkDy3u+lcYDwbMEbUI3t+n
kamqF4DwZCOGV8EOudEEapoxy0RWwKkAqA7Z6NkWbQeLCH4cWlQeVwohf2NYwPAB2BD+yT15V1yp
Xkp1lWWFkyPYPrAasx8+y9yWiYzDttYDy9JQVup1CAtfF1WUZEqkvCASvaUlzUo3YPHPeb8RaOLb
gYHaKKEa4msrAnqZFVRU/lMQt812K+AZeduVegT2ZAimYb0I0y5NJdH4dmjdK2M/DMpKz5r1zu2W
93JQh2WD9olnqulI8iCGY4gvPYGFXoDBMkMzhS+WLdYzi7sdcmATZNpCFETZ3fRE134oJ073NBU1
BwpKU/T2vWAYc8/B03IPJ7ZEYu/Cu+d21AS5guiBC1Tl69yiZMpmGpwuS3QvVFjccYcMloEwHBOv
1WbTXGfPLoBL/2dXk1KttTJ54esf659KbV/qtRxWJe+bCG3SEqwp9MCfAc+fwRBNTC7zXAeKhi7j
G25EWYOeA260x98i2c6dMq61if6CYcm2wM/wwMviczqTJ9yPZu6fmQOxMHFsak1lAhR1W/Yv+4SJ
1CKh1KjZXybK1gdKyl1lEgxuT/2Dj36gqQsz0hk3vff4KZUElPqxf3b/ZLtMy43ecEjce/ANkhlt
T+XD8JjJs3LeBgds4MFT2H6NW4iXAF/jKiF3unt0y78wveqLlAO3/DhTA+6RgSJw0AWwQ8SRBE/2
y9Gx8Jp0RkEsYtMXYi6xqLJGhnEZ2XuXrYpQgtiEGKWvTt3ozkTjdSSvzv9KSPNOi3841SOHM9mb
4CHNGC1slIWFqLhWSkQ+Bu5lz1S2tMKPg+r/zB1wxeZp/agwBKRVjnjivRSuVjhkVIO4lvzyqWQn
iNuWtGxUY1XZ9XdczHcgV4q0EBqQqrKl5fnKDiygjpkSydd/FgOXpfTP6/K8/T0/LaGbXMruaFU8
FZsSvbTlO8VVTWKvjRCFYzarfudR8ZLl//PjVY338Bws2tn7y/ON2i66PCXJYN/cAFZeiUd2ruav
w2y4rBoOdgCY1zdEa8DAZhbZQqRVV/d6VAaENKOQgng3R0lapThjGdDSs0Ul55//+MnHvcEvMkNl
RF8Bqah3ihm6ZjmiTjf1+3cpBX5BGPNuNXxumgvpbP8UCD+siEXDSx9N3eTiV9001FOoHGumhD4n
yBIVhSdCHQHTVUvZP0Kl4HUpsrDklGGpgxD/mYsOXkoaa6WQ7evcpy+BjPVdlnjfVywmhB560qzC
RCuwvISfZdlMZDmXQwC3d84GKcr3e3KfDn1Zb6CEe24Si2d/ajXovoyTw7SorXlc+HldFC8CMBEE
gNdoOfydLgStzTSbF4WaOqs8MY+nJ0JKNX90D2ExqTnOtRc446mLS0xffKtvkeQ/1JFSIUygcoyA
Jx/JKaQ1oPzM8FDQHRjvBpI20HyLN4MECCCH+pZJS1vjHRpTX2nzOj8IXkJFhu0iNkghe7FhILtl
xnj6yYfW8s60p2phlylD6Evbtabmhhi17V2S
`pragma protect end_protected
