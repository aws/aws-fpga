`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2024.1"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2023_11", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Am9rhBVZgqXuSn3VtP/vHsucTnLQLX3tApa1HTyU2Kt3CxUir7kYqlQosmj6cZWTG2CFJu5lCVYB
YA9eeU/U2ja7Ddi/rA6F0qh61AUzpaRazp+HGu6UWeSuzv/93fv+BnUyTpzADkDjF0atbQkPXvNR
daddEOIQqAcEo6JALAoFbXJXUbJ3ttnYPPTZmH1czLuhmz9UWyJ2Q1/HuBJtZBSFOcbi6Uoi9A9L
tPoaeD9RKP1cXcjAVnt56HTZQ27wLeEsGN/XAWOzRr+KNruaOACamakzxjSwtNjC3e2TWPFUBG2p
kttnBcfXsXBIWmZJm0dIcteP0yOSOyoxEXWxrA==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
TA2WoPkGU4Fh2DbqfNsgxJcC12nf2yKLPHY5peFN4aHIOsUjcMcna032BUQLlfHAFqIq4pnqPv1E
AkLdw5K8s8qidT3SABWp/MPN2UH6mbf87v287hKV/PHLTp2hzqwDulDkTID0q5WMEQPSYdQoACkQ
6KUkooFn+Wk7mEC/YnQ=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
V3f4JhoTzMuwekOOff8o+Bj4uFV4xQ1ih3Wa7sr76JXPbDSGwsnDhUGcG/ugKrv+Xi1aLwok7GWS
mvm43+En2SuSyFC73b4ys90tYKxrPziuu4i+PePurScv7PgqRvJT8Bank2vWM5VS8sWDiYLihZi2
uTNP8BdK4fYua+lvdis=

`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
AW/hkFGSX0rHy4lvzgFWn9XaHRSZAWB6a4gjj6/0v59J84ijQ8fPa9uy5xZdrTQcxb048GpXbGqW
2WKuG3GBlA==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3136)
`pragma protect data_block
X9NfS9NXcPiXMvyBkhWD18kcwGxAlijOewWYTzq4OE4pFfIwJRMr84yKOg7gNlcsXIId182rcq/H
8jmexZ9Rww3sG2GrxuzQUm4EArbeXpsI8Vb0diae0KGFHe3+bT2uQw7eHnSivxHZdBzP33D7/KCj
tiINIjazaJ/JXGQDaKnYrDTVAwL2Rs2YOQdV73QJCbscIhbjePUbQl0ctPMoJd53+z7j5Tv/d/rm
iezoNVROURTfyn/iaxZtdaFmbXn1Phb39auVJvROgs8MY2LKP373V+Gz6o2OMDNPEofvqD13lLhn
YiUEQjgGKOS9CxjRlkRv4xRm2pDSwpIiXg75iBOZLUM8yC3PxflcIxVatafCws3wM5zCS18ZF0ub
XUdVo93Q6vaFjV2NTTHyLBvkgQFV5wC4GmzjB7A5lB0yymfcfhtBBhhi4PVkKWD1NuzVP1fcmpD+
TeT3kcH9yvXkGmE40FXvNWRdky52eFEQg1U+FXbOu/VFR/fU3vm3aC1sGJZhjbKoX6gIGnjrBbvr
tBYP57SQPW/zWRoy+BZtbucKrXpP1qv48B/1ZYClzGw0OHDrb9SHN7CKdC0BgFa407XnVnqMOxCY
RzBEGBARM2bxvQBNcJYWXdASVE1UwWIBwbYLvaD1/erSzwbsOzfA/3i+hSYJQNXMPdM+DkurMaw2
JbkHZPduGKkPyYQ6lgYWON4MOeiKHoEpFjmpsZHjIpcE6QR3c3fueu7jtEGrLrUayngLDaNDPyEB
GqZdb7Sj6xv3tkR9EFFA0R2Q6SqLqIJCxvSSbOZSzBMyjLbbpH6KywRzz2nr6HZiIuv5NdBwUMTc
tYKY0yvTGg3yQz45g2kOeer6p7NFD43oKiUaO8PhvIOyMR2t+VztlTWyJqSAXyYYsF9DPTsL3ks6
cAgnXC+uoxMrt3Yrs1nEKz4FxJlv4JzsUFhfnb2j4yjoZc1rPYg8M1arKTS1HaQsMKciSuY0g8/c
La/j2ZLAUtjYhY4HqHCmBVjiyKBp4QjlWeqpisaaECuamHlHWOzQHjf+6WG4IJUxFokbNN9qazda
auLwDlQNbE7roZAuo6yJJwDK2AgX3giOcuLIUSdfuNDH9ZnXObySs9ZifxpWwAxwfHbvDoOEiHsf
U8afyFLLi63opmSOH2bgyrPuiVrYYXxS6apNCnQapTMqdB8JKC+lEAebFk+Ya3VLxBjA6/0+sDrd
9nr91zYBS25GkWHYG3cEC9OyKoiIcnJLUSY1d14S8tIzvLmPWycAB93xLabmZxXKLRM/JPjdcv9y
Pjpd1Eg1O/W3/YD1UcExr/dYexdOQEBpFbVzzny8g49HE7D58+o127g1Oz9stzgOvQFSTmRbvQMt
sFcAiKisZJKyLcwyf29/BX/myMrA83OJy9TSRI6hoKKeDGwhgAjoHyP/JMBFVc2m+tg7eDBEddsr
6cjovHUaaovvJytOT5UOtF7u1lVp1TkTIRaBC2ek4bwq2bTantdH+slakZ4oh4RVQ5udMQSTq216
NviPVx7zYycgrU/UP3L03YgQWtbKIuadAZGVcJfp+KEvlVDYawhF1912dcd0kdfS1K7ZwSc+5whH
0eM0rTlS0JufUppWcScEfyHtZn4e2aCguFmCk1QsrIoZayeCRsFHUL0W5nIa3Goq36bX9cHPwGWf
PBaCOSx1kMNMCUoWSfF7lCuL44DjOfVllTCSsxMZVAs+zvmHuw8MNJdVBNUHf+0tsZmDsKJtYOhe
NcwS+vVOotsIwopa4y1uV5J+46LMFuoPh7mu4Q4i0a+z6Oo4Epe3Cdqz8YB0+6RPdy2oTWU4w3K/
MTgHuUHfLk55gA3cWrLKjRyigt7RZP7S4dZUzK5lD/croin1ENnMWIHlo3pGsDgC+s9znhPGg0uU
woSXBc1L28rOM3QX7qYDt9vgFbul5Cq7hxCsr2X9T2r+7uQ+6m4AIaLT05e4dgGs7Mstj7qq7/NR
H3t4oLsV7tFyy6ttlV+myLrg/zIU+VM5+lH9+qC10KgFhSH2+OuaY1VNsW9gRm1dyoaJ+aJrSYrv
5PGCscnr2b33Ta+WUmrvEk96UggFML3/UkKQuwQGx2Thg3r19sl8bStwCu245lJ+/4Ktu738H+Vk
Xx2eMDydueoNoXXwJlcEdYut9MyH6pi9cfwraPEBt2mfXn2WrZaxLalCiVqYzELd9VW16uaABUCX
0xED4KVCg7WzfxmfN2dJw5pyWBo5qdp4EXisRF9odvFvhgh36GnC9cRFlGa6CrnFBlfZwiZjybF/
x9u8PYLB3xSJoCaQTvVJPEImAfGuAGHEV9lcpvOVujhpF3u+Fqgo8zd4Qou/IhIcF86uYxkUaqxC
wlsFYClFJVXksqa6UHXrQJf+VmrGHlYI/Nb9Q9L8kSDReUwCKBO2Coc+slAUVeTLG4Pkm+sRbvVc
Z5+uRmeiDEFUtG6x/ZYQ4d+TusRPMYRZl5xIN3TLvki8KNxazbW7zpIhSwHC59KJo6faDwdu5pzb
mXAwEM7ttlIoIA+YTNjqxsO+ow6Lunzocr32ly0+ZCIoGlSjMrv1cSDzkrbnwj/ij83cEbE4iXSv
1tTh+1zmD8HIo9446iBkhRvmyjzY7D6FXo4GWTR7K/pMsmKe2l0W9tj7S9UmeivqYyDXOOiEmMCH
nleWU1Fz9gyPmFY30zNEq4ASdvyjb+elHGMzzJdQnDulQUU5QKCbJ3mCDa8Ts9DUP11+GgBGFBvK
wB4CI6IN0jbfm2sk63TsNTgiZ6Ob3EUNijIMjMwrkDpy2Uhm5vr/wJHH/FN5BS7n3Cf6Rix1xJ06
vn+wnCq/jLRGKt+Iy/pZ7w2r4lePI3iVkSdhtqXfZSntJXkdh+jkPCOo2QE7wA58ih2ZVVCoafdA
5ZkElMlGiOQwmcr7ZdSVuBwlSTV7eV7uX4YAo800dCZSULRxcydPWJuD7kk5vi00YiVbNtvhtoFb
hnH0TyjgLRDtEn7C13JziUWKWDw8vt6zvIJoL0ZjWWGP/NfdDgUQGtZt79o56SGvuHuARHa3ZNZe
604wXs0aPYzQ4qBKz5p4NkxGFukWAPnKdXKNbK9ojBcdm6w31FT8Da6Cf2CptjQk6kpXaWRTGJfk
nsLF2MJMi2AbJbg9wTe64EWe8j5jVxorxRNpwx5xU4PQn45LArZ4vADe5UTvddRc2anHA8S/zS3t
xCkwgtUNTXeJ2DrLkYiQ/I4t2Uog5jERrcQj/1p1FWBJf+ThqmV6gwEI0R9tslDaPwtFfkzflJEC
b5nRzYlGNKhWfKaZJ7+KjrbRnnurJlVwtEwIkeBKqFvrWNlAWYpJrhOZPW796tIf2RGuqdVxOKoH
OvMs6sJt59Tcvt9Wv/kcI9zNacVNLtwT1UrlkeSwTIc2TWkLn2AvmvFw1DlkiRQXzIGdDh9HO5BI
d/kjKshkTwOBCzz4ccXJca5LWLoWyriXvVtWjSgfodyWIAa6H5j+Gn9r00pWeb8/c4xg/DGFesw+
b32qJEIqD/ctaoGk8JV8duwQ/1t+OmnQq5uxIfBl7MfPtDpaHu8V78BNJvscgMnjpU1jbw4YtZ7m
ta568wI5vCg3C7adkYn9et2jbcWz1dkC8C26xWP9PfVGvn721aZJL2C2eXBLnB+nfvEyDCy7X3+0
CLPLmi4QyACxlB24tPmGKZgIcwLUDcgwHM5rH5VUhaX6/KspGk0C95burWQjw1MEFY3HnxnS2qi2
l0Q9PxJE/Vk+jgy7qV1SxcRI+ZwRFmUVrZaWv8+E2eXpOdmNQWEBg6ExmP01iPqyXKKc9rWcFN4L
SItjaf4h0qDSDV7wSsxvF3hEKqMGjPiLLdutknR8qF9K9/H3CTNvhXhi+5RaZyLXyNyS9kwXaP4q
B2si/pgMJj4pQlVcwdldzkWyHB0vd/tm8HECVqPrteMAiKqrLQYY8dYZweIqsYHdVvh29oSRPXSm
orLQk3T1feD1Ri644TKxYbgF3IqCipr7AdXsMtbOZFN4nf38CHhZYQi68NnRFp8u/pcrviOjhnsn
vvbWVROYt3p3H4ZIdH9wKZTgnlH3yJ2gP7vGrCuFUCloHjCpVRLyjG+7+HD0ylxBJZPgm8ydOmw1
L0oRnNYKBrjyd3zjuFDcx30EIvBqkDD9kYYb8FRP0uC18b2CUfJBe/DdfH4W70iK1165VLMexTQ9
gQ==
`pragma protect end_protected
