`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
FYnCCFndqLVMJSdcrUmQ66AJ1xE23M8L1wvNGDmQMmE4eISPC/Of52KlKEZhvnBsxtF4gd+lWWdP
XnTu0OjbYoPq5u1grQnAK56xr7vZahBlyn9V23uOkFRmcH7LseeBIZVFE8wBxpfpvopuf9SH/Sbw
AExjvHHrQpe4orlnRMEWsIIi1Ykj9bl9Dh2W5vHxsyURyM1uEmGFTUAG79zQTce0H6EvL2h2se3u
XCwjRO/WrZ1X8WsSvFX5wNBrX2sb1PbIapfHdFQk3/gn8XmveaOPI0l//qHad1P/Dmx7F0c1vZ6K
0yVctSo78c9ClByIMoI6IJAkM5vkDil9qu9iyg==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
f9HwkPKPnBzsoVBGiwwHEYwhlbW7Zqpa11YhzGmhI1snChFZfrVy+OCbK3Qlv6LIbCNb1HEux2ZG
FtXMgzJ/zqNc/wkSi8b6PMv21lXUnnr0eLFghXXTRMrmuxHOO7aG0el37vRSGVw3v4oY/Gog9CA1
B0146rwUu5TxN8/fsVg=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
V8+R6/XL+sLF3xEkOvlG9T1/sIn1dG88kMPDgSqblhCCvoO6Vz6X6jqeEhegPj9yNOIqKEAmYpKq
bIBRr145XUYtsGt/fLsrC8W/34LZq35mn0AH+6UXRDghKPmecIGmeSrJP4TYjewFxGUrnbs9Jnk/
CRJu+/KIBRVSJUiqyUI=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5008)
`pragma protect data_block
a3CcWJ5Fb/oZzZdNcJgtdxSmi3ko1Ks2IrWS5JwW6z92iXR3n2e8x3P/mqytcdQx1lWiGWLi1S4G
TwprXCAeKhr1vgpkxH+OcEeo4pFVStIOOo5QZ2TeCoLg5YaNYiFtAPptsr891q0lfhVkDMdzZ62p
uO8J0mRp22oczjOy4baz/h7TP1uOpHN+SSqE2tvVoLdcv362ns4IiqNUSb0npu9vojr8WbOJjxcS
LP0t7Bc7upTB1J3QH3PAWlx1XtK3kaXRGgNqX8JCm1ot0xJEV80Yy/prlee9iR0qS/v+yD7tzOIK
YLXYCEcQRZ/DeGC6WxAAIfBl5U1JyJepIc1YXuk/+iCqdJLwF81tbIx99C+FYIuUiPe2IrNxyzMj
gMCvDwikd0jEIMx1n3QjCuFMtUFFLbI+2AAxSSlRNO4wzfK8DDoapaKprbCW1xVakyQTBVsJM5nB
YcSiI0p2ALw6oPjAHSaASVu3m9IK2v2W0C4INhrRphxv2feyDDYtD/gzwtHU6C9Dn8I9ggXnpi6J
U3VbpSNSWhkV69BW7yg/mdfh1EVzuux++wuSVnLBCSG2SkNG+sn+/0ZXFVPy0VCfAmDmh6oJNqmi
dwuDJ0AOJMIxBDOhFDrnWN4CzfH2+urLyAWX/cwQa1aH1j9qTrpMtKyb5vnMWpR8pBoaanqzs0Ap
w/4D7s0mAAA2tuJAUdVGWIsSh+XODztfuZNjGP37Kx0ykEm8bzAeB2fbn5KW2f/QwHde35YIZGE3
QJwIIO4uPBV4tW6PSCmDug/maREacmRaMXd2d2Cmm3iRT7kj98PHoEpdrJfD4U/f7o4B22LwQAa5
Z0OzBYWcEJ7+1/2ya/UXulSEJBQKEpLjSE0MxSNANZknqMjv4hm6wAZRNMWx6Kvri1xZ69QQMyRW
3xGeL3VLxxq+JXw/YfecSC+ZaisvuBaC5ntFHjz1QA9h449F/MAVQL26PIs/jm6RvbqbUlqplSSg
443OzCn+KifAgeEzw7xKiZHwwx0rYdaH2cFGe5pW84DJ6VHanOttDDsYAsy93VSlhZz9eQ+5hXjn
gwLuS4Rei4j9hLwK/bsIdimtKarF0Q3L+7TaT9ZqQT1Mx0txInb6iOgIpc7dGAnz0zyREaWrC/+1
5ezpnIk9iVN33G/9ZnXzJwKXe1dxxe7oqCsD+3L07NSY/Ll1W6RFezMxvv3C1jRxzxZlF6oGsZjB
fXCRsrynaWKhdQaMbIpdNGgF8iD4m+fPQJkZ3ikdONwywS683NeSs5oIXSyPfRyJ/M0p7/HdwReG
48eeEpxefSct08LB41fdNOIZUIzrWFzK9gsc89zMCY6Ra2hq1clKegrAAyHAuXXGfWaajBEQrgB2
wESYwbpQXxqw3qTMBeI898k+iHwUytkErQG1CVWfOXtKCT3Z+HgKTvjwIE7CmW7rrei39PCQsKoV
Vh00usJziRsGFXzdRrhdKkr+dG8Mtz7/Yu0XjNQiBvChsnhIeBHbkLXDpRoKnpcnZdgsmszxCsjw
qN8eDEkaoTBYwGBZX2Udu/+cHhpfrrsPBXW/E5DWMZN+QNecBiEWGEpxJWtq2dW3AK3M2eAzk2nD
QRLZJcA4lllmaqhQYsu7Q3MNBp8cBJTctETV0KGi9RpmyuUMIDxuMj+auiRLDLN7HJ8qVK9q8NUc
8uQ5JhuW/SPre/AObqc7y3Qtj9So+HGrJJdkp0pSOhAOKVzLU+XvRaLaOWmoNCeFHpUYeSHi7Vmg
AQpL+85KkvzTcC9e1dq5ynQLA8mPf3omCSrwCu9sRxFMCy/8IkrVwetfJubsKJLiYlPguhBHgv/5
vAsyKzLuH0S/3TSO1U2YleZkQyRYSKhyawabPSlc0I2mLQkoW3906oc6lfdxL27YgXalC1crhmX4
l5BMVaaolVX9k/N5DsVs3MfHmN7jSv1OnK/C+U9FHpRhlqfh7xcnkiwMZXb0quB8z8Ye1LGvY1v/
dXcgwWNC9Sq7TCyVwKF/WeSDdbxnEi2tAlbgQE2wYZtsKufNpuLR9whl+GdkJ9ag9Q0XWacxZLMc
KnqC7PC12yjuwaxW6zH1vu+5ZEsOLYR/nz47BAB7kVO3SCtK4GX+1JZdnM1SohTpI2e0ogqAFH/C
CflTUoWD0MOz0rXd71u126qSbd25+0kU0hmNpnWToVOdbYEBCEUNJ+K0FNy+gERLny6cqi3WsDZB
uRbvcYOmDCnQuCmpHFJYxTRmoPv7WJduxJweLtPufPxZGDCzGFdagub1n1a7D313nxfn9BGEF2qh
UinkF/IMcPpG/h9xrgT5807c94mafJD2CXORlB6KPzHZEhJH64SDGl5tZziSBqgbi6vOq44y4Avv
cKXxALafErgjtCmgWjU6YJ1BuynZ76Gl05tlRp+zVIhoLUDLUWUSb4BPWEKfmuduDg/XPJGmNz9t
YwpmsgNzjqtBZO6ggPAhU+boiNifvPdmj9+l4Tu/7jvyKKJllF2nQGNs5jKaKq67FgE1w2QyZA2y
0LMZ6TJNEeKbqCUclu7vhmtkNKVJHifcYAS6QCaWpVFM4FZAzmDRph3ytWp2s3rPRWkpCN7c/XAw
I7vEv0Zgdc9MJqDa5YLzUSXz4QDPjYDONjM1LmtsBx7cGZWA9MRJYEpsY2KCuKg49IokbbXvGoud
GW8r+XF4lKXq0jthbDALXvUqVhjvdktwIqo7QSbotYs8/TA01jwMpYn8gB2QWfQWXQbAMTGCMEfo
gYdhM8SC27C7d4BNx+u1BjhDxRGQrQF79AccetHoHgbsXGSaoRq+wx/ROKVQeeDI/LNpBTe7AsA+
hAUG0m4aY4OLkaLs+b1bJhkQsDCLjyqan3fLHTjQwCSwlIGY0Ns027L4BKcnrupMs4vRFzTy33CN
pzyhJiT85IFNndvce5T95ht7x/VYGoi0N2zLbCBpdNBXjxoI3RPDUVcQ7WJQ/Csa7sR3dEcgGdFS
IVQ+sX6NIkNX+7Auco4eZgX6G9ttZPoHQhi+qMyg5kIvs0pCGhpAmjmqPB6Q2G8S0UwwbG4cgIJl
TvtKiL6R9vF/t4kCI+5LboS6gPnZ4WzUTjNQs3tDBo07q6shhYjd+pxiUqhTiDDqsWlGYMJmYiW+
f6wVjNjHn5l7KdMlwTXwW4W1aHzgRd2Egs03UUTf5xTrOeXuWMoO+XeAX/qqzdcQsNl4XZlStaDn
2kEqif3ujC0yZmvN4nfV+O41TduQov5USyqVPDwQ0hZNNshAd7FeuOTU4jPcHhVezUPvD++6NhOU
f7VeEqsVOnaRw+qgKL64dQVQioq/jMr9xomhBmjuLsQfa7G3yUyTu3m0fDsVo7goPs8bMK+yF207
ZaUyfdEvtWQI7b+m40RoBGr4zUyoZthpVg05YirwcAyUCFZtkk6S0CTocnD5scavdDoqgncqAxgR
dwx2umCo2FVKbfcaqpq+IaOnPVBwFKpH3DKdZMnNWaapCaZKc6G0QZG4NoTsOzV5Ceg2GCjnLDeg
O3psqH/YDmtvVBaabVUqZfEFHZ+xjyXbrW/DPHzE6ZFv3S9EL0sAGZXt8aqWmVRPdSkn6wbFRKqR
pYuXzNMB/+JaViIXXl9f4sNCcujlYvqeIDeGSk4+HIGJGXPoW3J2brkdj/iWE30Y1z2ENrurrZfL
7ReEC1zNvHde7uTz2lrupF/RZjiWW8ndm1XSV4s7oyiSrfyUYuQNB/vwEDj2VWB/2qtQKY2ril3K
BWWbBbYUrEgAUscMpxHhH6/V7X4fkwyXq52va2ALVKZNDYlkl/TeaFZadRwpujgazaxl0fezeRiL
MC4wkLHx/ksbUFCozul/kJOG2nFPrIoUtvaQaQXkJT90LAs90XTYTBPZ5LC35IAf74/P3FryvOze
Wvsjg9/fmhN/h/rlB+0wMWSv10dCxHYzie6EP8m4ALi3Ypse38DnSOP2hD9Mj7ZdZFwodqnMXDpv
eiF0U6vZP5xoE7PFUKYTd7D9QDIX4PRT2KNUH6b4pmdsQ+nlc/cXYSA1u3HktP/tg7wpg4Np/qbJ
nxY2uckux0I0fCHS18EI7d1lUEutCC+b6SDnqjpS78pMFFMoggOb4xDuM+yr+XL71FouvvJSroxk
xtD/lTlatDIx8UFUmZq2kj4xnm+C3Mvb6tzUHV5c3XJaZYIMm2inX1PuCkKxQhef0796aAXkbZuN
5VXSHbY8vqXknXPt+8+aBERuiGx8lCR/FS1LNNetewnjcDsJKH2MZsGCkWLqqXvGlGg7mq8Ez9pi
yCC7UVIeyu22gvli6gsXW9BuTPi0MLRIWCVXEYoRkbFRq/+I9mRvfF9EUZdfFvr0XxKR3IWKcQJY
nVwoglRfxr/WWGEHr9HBlIC2gLTzGHXPhQgEvwEv5wwRG6le4VOiQgTyYbwSp/EBr++fWpWC+b1v
yd0jTils3ilS00bEw4WHH5dCkvREi/CHd/KJwLD/veq37+ecCBO+v1ouxVA8AqoVNDdJUyCbCAsn
jevmJzFhKHfUFQEwxEBymBw5bB/bmrQelvjis6EqClVs6hRW1wuCWW0tPvdHqiRZGmLsDVBMrvFN
Cd7Fu5x8wJ4y3vCzKTFqpPBXPP6LQdnOQEx7b7HT2OvPBCbg19o7DuEj4YEPLJZ7w1MxRhLvGBTQ
Vkad5DJ9Fc8TbQo5SuSYGcQR31B2ROua/50BB6fbRme9kOmQmzbqCXURhzLowQRqYQy/4dLK065l
FYd/E5IXTVC9yR19cRwz2fhA8Z7s3Bdg14kYkOPUtp4VCPR5MIYdTTRFKf8lA7G/p+7WOG1b56VG
ZC2yE4ThMrYVp4pg5ESGGZpGfO2RH3lLXLH1/r1a+Rb0qDOCAFOo+RQ5hDTD45ts9tjMptPW0Gpx
hTS58hQHMvoQZDFgw7bZh/y3GAp3aEAtrv/LUqdQYM/pBdC+l2wCXqWmeSGHnlEpr0EjtASkiqD0
Idm2dV1G7tbUrj2d+kkZTJDa2i7t/txnn7a1nLJ/ffJcTmpfE1JFTfnN5lfhB0oRUn28oQFxud9X
KgSA/IS+GuYePECnUvsbV5FcxdMz6x328d5/z5wNRYK9lXVaackTc6z8VrGnX0lIc1cgAZLnOzZq
ulwCuCMrsC2pr6nuI+mDQyqhCK/k5DEWaEyTvzz3fE6ZhMMi1I+2Px8RBb3Hju1wV19RpICShGO7
GdS3d1QP5CNblxd6Eud9dyoJwoWygCls5LUPseQf4WO6p7VkHv3UIPZRqAlIUgWh9q9rId/biVlU
nFqFChPeafotb2rfvbf2Jo0IcBVmE5s3WTeBNUMUgNVgRmm84X4r4tZIGITA+HeogFBlxmFxbto4
woAqqVFAyR9+eb/Jq00VKLbDJoOuf+rAFckJRY1z/FjgZgQm5fXfzBKgk6/qWMh75SNU5/wAl6d1
QAXueAe0VxgVYl9HPI3hoFCrQzQOSqhzdspkMz9UaFnKfsJWxKgjEiRYSQM+EEbmMuw/SKw+od+A
uY5bcoWvyKOcqnDKVgDAX5p+kmiCDfrxul/vJ74Dm/5kjroJ1kXKsL+mho0JMBgAfg+1/76yhqPl
gm80hyGwprQpYotviUxnZi4mW0Iv1ihlQ75R3TPnowrEX3IRydz7Y4z6v/0i/tuoA0OQNQMhHlA+
9WEuR0COYJ0C99gQzEyLn5uVDzhaGGJuGkVSV92DDk1rMvs59s3mO10HMN/c3rJU3pfb/ocSy2zl
3+8OOxn5ycgLugWqqlB7H17VRrPOFxKYgeeqb3Kw73sPAq/z6+Kp+KLIHF0K1FKGJosepOTkxpBz
dcA6VZKBPZFyBt7okxTNq96bITb/qmjTCdV+gxbDWVV705p269zFrJjZd75lDn+flmGyt3OagB9c
ZjkB1Wmd0G4ihP5ro27Sz914epEaT5DnAQe9x36gM1Ue+FJQrCGq2pAB/R4JOOML2oMFJk+mOb7g
UAaP7mUHsMAmIelDLWvZaETIXqHrHnkpzJGAFr751H9naK8jaCoGmPnjv+RygtU0h4s1uqqDanLc
ZJFxkTg6aGx7xMUDwBkxnwxYDIXabyWtYYvbrMZulx8TJMB4xKsbUEft+1mVckMTZfM+md5F1n+7
Aa5Bo/pCfrZR7Ovz3UaUsxOb7ivu+dHHu3Af9A9SjLxVjRHz1FlLRUe19xQ3IOftMqxqbVdSYl39
Zy+fw+/Tl1pzPA5MB0QfNzbIF8xY1AXbGs4nhH+xj6piL+diNgZH/gBgFRTCTt4w3xbZzzZAhJ+p
/FOmQzTbNJEfBtOIkdsavbuZPBnFlubLM9mTuopZLU0/wjwM19gs5G7lg4SePyaVSVPLBG4KOEbv
/liNL9aJFG+wuBmjAqGFgoqvY+CiydTHECEh/U36Dnx+Go4b9PRuZ0yXltcc911JklvhD8X/OSYR
ZpOvzeqP1tEt1hux7czE/Tz2wZgLo+khgrRiAXwBXaSuiCytstVcDDwXkFqpba6fhJZ2pIr1r1De
7OuJk4hbBHBPBlqmX57voSU+STD6vDrhigD2HCl8OzF327JmYpQdYt/0ME+uiQtcvwJ/pBm0Ffui
ia0+eYIcDZc7U/0CpgVHo4ftSw33DeQjhfkWkEVx6GJqACSdd/JjJQHNcQR2gqakJ2mGZtaPuXuv
iWqF5t/RG08fwf+LbE3ZGf+Gu/BgiUkfPmKHbl0iX++Ownv2ZDXKlqCuPOvqVPBnIg==
`pragma protect end_protected
