// Amazon FPGA Hardware Development Kit
//
// Copyright 2016 Amazon.com, Inc. or its affiliates. All Rights Reserved.
//
// Licensed under the Amazon Software License (the "License"). You may not use
// this file except in compliance with the License. A copy of the License is
// located at
//
//    http://aws.amazon.com/asl/
//
// or in the "license" file accompanying this file. This file is distributed on
// an "AS IS" BASIS, WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, express or
// implied. See the License for the specific language governing permissions and
// limitations under the License.

// SHA: bddf8457046b3a64e63d28d7e334020b6f1d09ee
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
J4FOGjMXPu/gn7ghXA5CacY2v31ZubI7gOi7zscw1iInvlhnE28bHjS+1lwYpPT4rPrFGjapFszI
BF4nKRaC6F2fgaEheRMy2r1j44nhGpyhy6SZ7Gf+cpH9j1miKydHHaEK89/Fbi6i/RFJX3uyo0e7
0UPyMHvwvc6gKcaLJ6G4iDXzhUTVv5UE1elt/yFhYrbUe3nRucnPvRcW6kfJloUIV3naUb9004SY
cpYrrOeM8PVnHCOS+0ij9O2Ff8xnUkl8kQb3mEejgJYzveJf4n65OmwLpUfuuTugcM/eKByQRcbC
C188BnNEuewi8fWRpe43YiOJaM9BT+mgynZI6g==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
EZ5/HbFQdgP+fn1FVkd9FrTqwjf7/NAE48ZfHD8Nqd5YDG/EX1g0huC5qpts17jLFa18CuomLPUm
sAdvmxD6P3ghNUK8UC8V/vTNqNlmBSJSfKlLDdNtTea3AtaOuFP0j3usX4vs93v/8AoeEu3vC3Hn
AKamrYys7mKOkN8JNL0=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
WYYVBZ3O2JvW1Jpc1cWWWpCIjxm8oY5N0On8n6LEy1KCmUzNsFt5v/VTF7y/Dx3yZfECvx0vCZ/q
6rG6iAn+chPuHv4q0+Znq7wI1Inl/pkm4+BvwWrA9ufNClcKb3M00COGbJ4z3IsFF890Um9E00/4
ZIaVypMT1EUMOjX0Wcw=

`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
SEQKzb2DEoUIhLf45OawB5dCSSTJm2uEIbuG2yJpFskGqu7fw8mUpn+Rlr5mUwXcZUQhJXRpC5cq
10/ZxLe18w==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6304)
`pragma protect data_block
B44B3o3bdrC+g9L/BHxop54K5aS+lBJXr2WrvFfgrcGHBNIzpQESQA86vLBumSDtyRtBwY1874pV
yMSAcL9Yw2/svKLMNcErPQufgBGGEQxwNDT9C5oerPxXToJcRTUGihvHtN9FpRbGQXlQk/HBQ04s
UdrmtG6VRPNfQ1t4i76WXnL4wPUkwVDGidbwxKHWSbztrNsVg/DkcUfCXyV36I3ypJgys1mIZkSC
1PB98Z9u0jdOoxhc4s+7zj5cDPl4qHvGTtlhgwYp0OnasrYO+z/0mF3ABAFB0Ce/j30PjimqR8VW
eLQHRYTpwmCsYmcJEJ9/6eRdvfRLD5uNaszRTakWF8glDWp+sXylFFcl0et03ct+24RAywFUUO81
ixNL70lnEYI7JO139MVyJ/liwu4+iNT+96r+vEUrQpKkrlabiwmR6tin3SlzwxO8o8vNb4OMHr7s
y/NwRPQpCNrMMFlN/0WbqWvqbcLD5zOFp/0dvON6oN3LS/0iy3RPbkMMPx3yGG/4gyBcOf7w8S3t
5tgK5LMV7Sj1MiC4oKBNfQ1riTTZTKxZ8I3BvVrPKU/WqsgqjYOK0XR3+qp0H3Ms5uiZsOwUMhPf
BT2gtmFzH0JsynD+4P3+of7ax9kHDZanbUspPEVVemwIT+r4fKJwu0YhL5nYRw/o+dmammCn8XPQ
I/or8RjlsOqhXxGvgu3wKx7iyUi15y00dOqZIjZ+ykfUCoK33RPrDhXL21MMnvRmuJplVjpVXIot
82tx+0isOCNYROO1VRftIbjzfPPbUw08l+quYlSkAMepUCzNrYyrj/C96RtK1HBpyshMO58qbabN
djHjW0cG5WizqROHfRHTjUZJsgY2mFpcBRnCz/mt7qNbr5p3O1TJck6r6wvlSFX3QvKDZgeE839W
Dw0sTIWG1F8F9BrdKg7q4atE1dKLZzNgHjEI7s6z8jVvyJ2lLz+13iG8ndljEHNoQufGqxnmhKuv
nbR4nge6HWdRYDysUECTo6ktCgr/rgRiJokoh3/MGuNaEGg/R1nSjG0w/+cnWJuqKGQvobLnanIp
hkeCEKlHwUo/IsRD8+NszM1jVC+MHKPyikZ9hYSw/DWL981WXDQfvOBhPFJsa3zOG7sL5gUNO7al
T3Bb6wQSEdMLuQuKfz5AwQBi3jTwaloEJ8/fBacJ6mNv2e9JMyc9/Ag+j6x1VSnXDMcFowOIAyep
Wc97enSUmFEYeFZnIRIz9Qg+8QaNxRmZN0XnkqrZQQrmUMjbIvQFYwgbFXxydOTCtteL1GXZ9oDl
80q7z9RJr+jbN5C7NbH+3z38cS29SzFq0RglDkUF+KCLuoFh0qgnNn0nxtccj/Aq9blEfm5vsMFZ
vcboGwXxRc0wObmFpaX/Bwt3KwCyzLMQu9/D1fqOZFZf01gxkR4TZDsMSIsMlgyO9dH59bJPcgze
sHEaXh0unm/iyQleftj1x3XNB+mj1L3KBhDgSJibUclOYmMOJiTQ7g6iPvIkpkPj6ZOi6pVfJWTW
kScdNXmUQW4f2bWUg+7ali3HW00Rv60v6wDtT/JyxSqEZU5Yz4Tw6iYS2oGW/ZRf7Tdxbht5pxwQ
eGcT+KYaTO7b4aoHvVlyArXyqVdCy2h90n2UOZxojSkrwIOv4jkhUCnQTBNV2iN5MtOmv0LJDu9t
+3p/KKOvnOyN44Yuavu+KvvXvh13H5KHX/3UoGMWSkqlRK1CB3kp9+OxxDgBh0KIgUEyxkciF0ly
vXbsvhJUGl4PzeWqf0nIl25MFgzvXIX393MTyFcWgMBl/cjKPN5Gdt+wXf3hD0tWW2k7P/P2OayZ
NTbaieai5KPLpoxX0+HQCbdAIOZ6wJIxCF7XcMUXoTT4B2W7UQDRhp+o0eHK2W3XP1s0xONe4ZNh
dzrxdaNr1wnYvZfm2vG7xgY4mRl/4p34EjROSHSXoO3DI0MUkg+k/tegc0wGmeILpCm4//Kh6vKm
qrG14P9wLvmcYOw+sg4heKfXWDoTc1P7/NJKrUhj8GzPwDyNqTnngO0dpqklCg8NDUV4bMgjXGDN
RoMphgvGkiU7nGfUE4Sjm5fDUWodth4uOpEWSOhN3miFdfUe29YoYV1nhTXqbhjOSnn19zRofADG
RPjBBp1omDdWT19+SPdYYVMqOrPKqtbvjBBN4M6b38dT7Bgj9YyksM7/Xe0W8hI5k1dh9Xhh1z94
qBtFkFFnnOYqD7KHTcNqMcKC8+9+SOZk2TAnoMF7+KF04TqPVCOihErpTPVUF/nQblz9mqgeZn2j
CFcs+dX7nuIcoWEvLP81w8NqhlLQn45CbQygVikSefoSjTuFQYxt9I7D+6kosEpUVw2uaRJhHfXe
FmyrCfy3BxQzXPFQtqlmP+116hWMADqB0Bv0E7FKTYeiQXYsLzE0tJWatcNye5YjhZfJAwqEFTkZ
1R+xV6hdjCoQMhXmWqtJi8dkKCRY6mH/FRKZqQqiGuUaWOLzIOG9g+U05us1UQdZ1Q4+rOx23mRx
SVX9hZhUTJiEBzW+Iz5GWpMnZLgZLn+FS8kHJtdkVp1hbvQGXqJSrpKaqJV7+YAIWmqYyLmyu4Nb
lg15JpVVTeecImkCPpYnMz68RtFvepaD7oQi7AetEun2XO3FbAotiMyMXATpgUFaVfZwxh0/XD+1
J3vJ2Af3fAm5KeVr+i2O0I9nlNOHuRne2iA5Sb18Yysgau6X6JeKECALwx+cBv0jfdy/NlG1kBen
dU5pZpCraaW00Cacu8qGmJrQfNa1y9/+kc6AGNrnnjbYs7jgsTtsLV9TVbPKb9U0q5dnDWI7Tu9I
m8VkwjrN0fmv7e7WewtpRnexfWY6qFSF9F87QjWmVI7u19NgZcUJjJdHYkfNiXdXiE1kUCU3yn8G
1bI73G0g6CcYwWH9UW5szTQ91qrFjElRQcoTSR0b9SB01OElOjFntEhwNp61Q8SRdwED9paTaQKb
W9P6EjoJiZP8l/PJHL+yGYvxmAJnexroDE+NQSUAVeAU1UFfAgzSwtokhBLgt5qZe3brbYJ/1cSG
tt+P8Y32pzKeV4NSUgyBakfxDkiIEChsQZdy6nmf5X0jg81MCbxoWYXUAquTuMENri+R6J7gr3XT
ClbbJzzuRRUb3ccvlCngOAP4B4iHRjd3z3QLeAKaaz2n5WwVaemlDwfi1O2PE4WvvYSmf+yrtJZ9
lYaO9x7Pa2Nz5CXhpDOzRfKPGQ6XxXZ0HWLINgy1p4N3unS1N+hiDkCuWwR2Ecm5wVthmYEFO8/d
FsrUaydk4wdbkgxASKy96OIDHOXc9VZgsD+bal+6EsDuvjAjKsjJedoPLByj4EGRSCprHglnjVyr
1NBRdw0DBIFVtSROxKeKnniKFDKlRUfFT6wCbbdPWvjehH1rU6tCmVLv3J3uA1ddpvVICwgHCWqx
CDl0jDEmNVvWe99Q0HLYsssDky+VTAOTry/rd2aT/aSyurhvTyTf1xHAXsD2syl4m/w5MriNYFix
67zquupmssejx4atRtrtekJAXsCeYVovEGi054ity6iui/TlUMzs3YIWFeH/AQjPp0GSKenYOzOc
mRPCatWg4z9PP5AXzLEBhhO3YzmpLVc5P7B9hLF/ZSRI3qe0QCVf9skkJMwp5qGnx1aypyDLtMIi
G51aLqBByhC5x6VxsbvAKXveQr/ympp2Odsx2wD5xWRbOEGhrKn5Fl7ocdLbaKt3cGeurgUBmpSs
Q5FecvfvrxmhJPmdlP3ANf1hZlOTxDSVIBwnQsgLdpMuHsYVN2vFPOdj0vh0/7guI6QUPsC0Fm+9
i/f6gs+YDRw2UM1y8qV8HJ81Us9QjPujUtwreXUnBqWPso6Ql4dlhXAgjgANq+rvZR/Gej/NGbJX
cCMQUHTjoKiWNVJhbgkeGapSjpbRoXvKXa6kU0lRw9/YxaS/rdCVs+U0eij3dvUm1jRStAvT0IMv
Ulh4h0vXmJmYGUwo3GVwU6xFkmRZffImXkxYXc5fM9Stm2j840cPhz/0j931KU3fcgNiUjv1dRfM
wFyHhA48rN9sUYuxC4MzeNW4Ubod01mMe3fLEOp0suIPzuXE+OaQe8J7AjZpNStDkdG3TyzEr5dg
7TlA+ne5+4F+W92rRgqzTTnWdklOllA5QKX2TzkGQnFWJtI/Z42KUia6zcchlxlv219Vwe9XiG8L
74LT9lzsX9fXmawjNp811Q2GmTN5oePKpeRZOZX/eXcech18nVP4n5emftl+9/0ao5peDABb6ROd
YHxjv62+QPBjOL9cw9uPE5PfVRHOVT6+JnUxOgFMSnrm3wq786vYQf7VaBwX+4JUJ5xSGDutZRTy
Ya9ehidwomGE6+1rbcWRGynxMYKVP+Y6UxqdIHgYe7E/JW3XIKl9HXLm5rXrQ5WLk6QeZF6/nXlS
kMj/ZNc1luaZZ2SsDCUanxkIn2D2EF7HMG4A+0+BDTip5FgW/W3vOOh1UonmJv/wxMu1v5rzaDfZ
niSPrSvSRx2OVOt4rfv1CM7Z9D5qOKSbKxBeZtkCmAhTu1XOuJAYlp1bm5yHG6GmMdezaIIGeZ73
NgJR/S0sYEvDzeDesqQNWNpn/XSaYz7nuvg5tgsVOr6QIGxxp4DAJc1Lttxs02Hi1VWPuh2M7eSG
WQc46GUEcf2x7r8VnB6UROdUJdT1jS4issSjxQEpqMg0NynSvXjuuZVOhploOlNp34AGuOhcVGwS
QxDIGV5LOkDno58HngE7ereDB7kGPHSho1spN90MSeu10ti0gX5hyV2JcuDGczJA2UohCZ9tbNAx
40FD6w5xZCxaQGyJ9QbtXqpe/Od9pSgg2Q5tFgk4EoA0CYB25tkPrNtwQo7dfEcUE+t3+L6uWWOX
XNMExSHf4Mau5Pg3VFdgoI8KAo26i2rXp1UrI+6iuky9iJu+3VXbAcnqn16n4IkMQyx+SJkeYCYC
c4FOvRtHk7XjVu5PEh076wKMcPy4hGi/tOEJxxOlzq4TsyydYgAjsSNR1idFxXBiHQZbCS4SEjeh
fKw0Afd5fdXNcG6ZcwrTiPjJ8eHIAjIdHeTpbQCtkauGLgQuyfiGRUN1SuAaQqVZEDGb79OZgnrv
ijw1aVZrOrs4KT1p4T2jNljBBO1nD3Lzlk3Cxni2kapv5XW1dLQgvngkO0JmSE4XsSWTbYgzbwfm
KFdUDqbZDiFV81DIvU8+Lnj+glOaLGj01UyXGF7DHmfFGTIko+HlFbLYJl8QLiAhiWKNPsKqmQ1Z
uorAtHcqg20J4ES3pOS/BUD/rAQ8qUpYotDZc5d/Br6mHCZkYB2fMHoT6mksfKe8nFc495Puk2sf
xGqGD2OVv1pYcw1PczkFOPEHqVSj/5BLgwydGZr50r5Cm8LajXuGfHAnVlzQFwPyM+22k37TYAOA
U6UkmoGY4v9cgVry9SFGByN30kzosu7/cph/0V2h9Quj0wlmh18AfueMXUEsDEPXEMZb5IKnzU9U
3CjTsOGePdiPN13/prVNpNtAY81SCl8j8IKOjacthX5JSZLUC14ICH+83nBaaQTiUeNbHnMRTfpH
Wtp60Zeq2hb7IWVRWDe0mO7EM8dXh3GA7Bs3M716gYP3hI/u+UWkXaqG9CR+v3Oq5I0NIATi8h36
DubGxNP2RMSGmE4epo1FQ7DCbibGH8zmcqWg3YOn637QKtM1fSZNO+W1SIp34XKOxqyQFvGfN43W
brxk0F5jOmemTWp4nVBlwFEe+NwmBS4rH8cqa4buC+x74huF5IH8zC+xo9g21KWFhHwdKx3Q75cf
Nr99AKxlWRcyyNgS0zFHTscg1n13f1bD8juwEqgL43GWu0Y5KBLPN/MsaTK12baarv6/dmanB8PA
Dsy3h+9lc8MmhptHsiZk7lINoWGusQ5yGDsUN3wVw8Ym2W/tybPXF51U+evf13xG8xG4ATEB2cMk
46lX5QtAn0W4O1ZEl43DL/RElbJn3jmVeyu0mdD1vYkqzuL0tm5QmRWUpIvevWMXOlerrn1Kd2IG
f/+vbPRnjz4Dk/zsmg2ips0TxSGO99I5cc51STinL7sikBgKrvp1xgb54QSIf5LJoTS7tj5yDg5y
4bQH8U9FheGIpfSCON0zfF6N/8dmbbNu0d5CTf4gZtVpbZv7gAWvN0OqJcTgZEC5yTSyVjF7uEiO
jyQ+esh1I4tk75kR1/Xl5u5IjnPVuFWqr6nEOBxnvjfF3di4QsiJmNfQD9vbRM9toB8ByIJBZ2Pb
hwG+r4ZphaMFZKEksyhxdCY0OyPNsIead4+WbKYR+bz5XwKEXJKRCl0I86GlrIqat3mJ0x9sENdO
MD50gs3CaTWN1ggGj55jwdu+GFPw3XRuLSYTs7XFBnNOeB7uAkzvjnam9insc2XrUIqEBxPez3uT
MrtI0HwaeYjC7I0bMkAHfUbmo47/FesazzP9IkypWcGad0UtCfc9rA4/Xgo8Ag0S1zX+LcnJQiRT
GpT9yzaIvXtAWOIy8INj4IU9DD0kbdxbIiFlarLPfZVW1tHZlEUNIzwF40zAq1gQO5RxInF+U5iK
isJYoQJzDfqN4xTfXzdzM3VO00Cm4/uCq5Ia5hFhMyQdiwL6/2eoajShnWugkEkkwS9K8y+SnOOL
O24sgICeGwFCrMeiaS6Z409fq2mDjqYEsBnnUDLqGJLrtoEisOI4WkuPNsYJp3KEMRXX60mwrl7e
eUq0T8za+A8+H7nGp7Ao6ER2SPpSi5ssvv2zaWWeWq4NkwxUbQ5F5xi+zYMm4dGw31BDAaUqgrdQ
vdVjZpgO5YlEbZxDYRmWpb8rA4zaPq/VoRCdxmwhd8O/dywHmkFnJAeIwj5VpkfcB83JkA3BnWCj
8hAnFbtvPnpHBRWCn62h9qCJpML6FBin39Tkpu7lHw1EJXq5qDTHmb+IBWVv8N4Gnq18bs+zWRl2
nuH5pD+/cB4BPi00sHkaPc1u98SROKasgmhu3B2TP8w0JW7B1U0g/f0MQr/UnKPXIKlbccBr3VtD
f504QT8QhXLVyy+Qs8MDtLvfAaC7pJMOglWMwtuw1VKWOOiG/hZEb9+YSasdhMckUNVUheMS0YyL
s26PoA2nnB483eSv2s6d7sPtBRoLKlyhGk1XrmmIiZEF+Y/fwQGUqFWF/q/HrMxQ3ZY49+SF2N01
At+97/vwgBzbLAxcj6GhcQKCZzgCdnLG52EjszB+v7weCHE+dIK4P6gFNACUR2VobGxWOw474bWV
F5/mCWgL3zi0UOv6OWmi2wFtN8IaqOaCsiN1tIWrfbJ3Qeu9lrXzfPqZmtvlXUFySOBZZtXb8ufr
2BVQO6sz+4aMoebDABPmyIStHyynblo6jdbzOg96CqW4mw7dAWnL2z2+55pjV8aqS1Kw8v79uhPs
75EU7LFQhZ0JVPIfZ3GEbLHv5qXIejeh8RxLdR1W2Uv70aGmzTmE+E/ObAOMsk4UJxHNvc9BHWkR
YclEMtGS8ybmAJMuSLlGokgr4YtwjIbe/XtKAumiE2mGcGVgN//KY8TbHCkPkkehxyK6VGlpy/LW
nGiNzP8uX1lKtH9ktqygBct6gfmDpkWqjxd92FVn0gZVGioSj1gwuteRyuaxNpyQhFPh1ftpkaqB
6crNf4dzfcG3ljfwUdvB4CzB4eCQCjQHYjTE5+5W9C5EcZvNMp8bhE59ctqWsqFDkpO+/lWTUFhb
1bY//uYPJ/api0VHFUaIPA33TWlfpv3bREr/PMJhgG+W/5TlQm+eU6ti0Pm/qZ5kFGOIuxt5ts7b
QsJX3HZO+j94h13lTBQabK41kAhi7+LE7lQj0jKEkryC1rf5Gv8yuETAtRkrDvHnjsQ2IxqBgXvD
TBqIaQneeMJOpPpRPlE7Qi/MJDN4OAIPZ4u5eH/0nu6ufp0MYuS+ndWRksJzjpnlaLW9WTJXsEKV
QgIv4YMgejgoxYNs5+ZiLvCwasmmP6HJEIXVNDJE3XgmDMnPf39HWc5LMaskDY8mU/w7weqA4WI1
fw4BProg6HtIlFW8qko/UHf2Yc8JmLMzkAjy8W/XTRet7UFjGXungDOuWFpEOrfJz0ZdY7AFHTX2
5Jiv6BQdnyasNiq+5jM8bWqGEKdof3+G8+EEsLTMPZZYCYJaER9HbMzMzk9UH6N5Q6ZDJGib1wFI
Ii4p7APA36J7dCaUpt2BkTYLUCBEINAVrLNzJiu/3GrBUkgoSZveeLxlnYRQke9KgCRAPIg/1FL4
CxMBHKyzyKEeVv2IJwW/MP0ER9aaHNDmWr/5Lv8Ng4Z/tWLngtDnJxUnw9lEGn23hDEafgbG9D1n
xLdCahYMQf0PQyfK0jsaeqP9K07mV6yBNW4BkOsit55KMQ9azuxSVkG/sxgeQ0elGyvhKX8vQquS
rN2L3sijk+Dr9I/q5WQ4PsQfy5kpdwTPS7kC1sW112L1lQ==
`pragma protect end_protected
