`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
A+43fno5xQumKGU/iTEfiUyc9UbKjC9g60Ecei8aES21FioEUlpKxcmh+6hBy7YeiO6/eTkdgWt9
kIk3tC29eEr8BKG0eZQk78uzPXS0/KxXP31jWVnCSkG2JDcyzxm1QbP5RnomflyCjySyxPFR+Bp2
p8Ji1PWIPzwWBBYZOesjhjcHHjN8jx8gZgBUjBsO7Yrdm6C4+L/tIzV22Q6HQBTDjds0hmxrdQ9R
X2hPfQ1K5MioWHNiCEvWEW8Cb0W8BykuTplKYKM7Ty9mp3nUY65/yayZKvolOVilW9iyBQOJtuuD
/iriAKOxpC1FxfdHauEKUsCx42RctSLIWMZftQ==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
cqrICfhHQoRBkvY1M/JgEESiWRgP1HCwF/2JaV9PeMkf6WqwmjhYUYCo3hnazXf4eyoSLJxawbuA
aMqJnH+ol/4OSLNelFc17XKKHiGvD5G5E+7bZOaqPVM75RekbnOzzKSJNMDbDX8yyCJu/aezB5AT
jO8F5yLwD8AlwQ1/QG8=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
YLTcOhqwMjgVd/Hf2XlYfCoVK3UG8edBZZmT7Gq4Q4vVUwapJ211M7UWrpWxLfAJl1DZicond3lO
r/00bsfLgYxp+/C3kSPJjNyjWCqBAOIWUhFzotP4n+Hh1Y/ikRMZjW5KFvgexeJZQ0v80Y40pGzy
fz3L5MBxHSNMLYKD4h0=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6048)
`pragma protect data_block
2dwtM0fES03ueJs6vuEQjayl6iAH2uGo9GsfthOH5YcLxlD2R58H6K1/3NMx5wn4+rh84kiwE00y
2LH704qsM/1ZqQ7r1iX3+bcLnHgj95gRApW4Qh2Upqwp7qCKyH1Jj6N4EBIUgAGCfpWMProgIJQN
zZWEyhkMcvE0JbId3XrqLuNKJKnkOBPeS/hWC4P6efEdoNQbHBcZo14VjBZw3s5UnSm6FBMtnPFz
HEZwAJJvOHWq5DKcQadfmIqakptSA35W+I5QXjoIvzGEYlAUXNH1Fft/rjwC6L+pgC9g8i4cVPjG
xIwUZwjr0tnggQPXL/xIl28HNa3i4xy8Wt51JHn60Q8z8o50sA/jxrN4r8vgKvoDlKrpzeSbxEXR
sbgN05IRkGrUyCnwJa4BdH1EniUE7yRsvJ+KNAlL/AbpgQDRJG2FS5UROCHRWVK9iQiqW5ZcHA8O
NzcRAZR6qtFGPtBWcGYtAboazlaZduQCu46WGud3AfnqQb7DBqAG5pkbcyp0NGUJZrnMDgiIZqXt
mRVMb3AGOIz2wbLOT1rNHg1MFZFe4z6SMAzh1hnUHXqCI9wxgwzdZVjvu1rlUFMtLJbUAi8OFtyn
c3X0w7e7onox07Y1koGshLyUE1LGy/8lgFqwJ4DmwQL4N3tzGvHLFZ6oRhsw3wqed325ijFi7h0b
CsuJDV9skPM2IYDj34SdQf0UXCnxKdpOEGMO/gqQuT4V2IV2jYMd2kN4XeAPIQzWLapxYcaPL5YX
WP8uVxCQNl8chiTFXlLlKGc87+NoQHPrXpbGpj9dEE4WxayqcmRDwj5z6HSZULz+HA1V+OkdnilN
mgFlzcylsPeotEjpXzLODP7d50u4pdQGzVkH6HbqKdHHfSpoiwwfBewVuXASA2TXFjCKjkyxOgyr
JtmQ6VeA5AerXuBIPjb5wwmArn2gRN0RwGcONXK5AHXt7Ikhtm0/JKMLMdaFCXgPW98Jpuw6HQdZ
a9N6GPbaDngkA12qD1ktgsLNuBw38WzwhZ8vaUiaHyXGUndaLTg9kr8nnIjrXhpaw4mRIVyYj9qc
deKwYX+0oRG0cHM7P9QbOyM1e/pv12WXaPE2Q3zK/+cnqKrK+vE3r6PLtUeB04RT8heQeiFpBVWX
xXf/CMTWcpEpUzqWpIavj6l4nV6AyN/ZHa9M1U5TCsC9JZOuY6NtUAs3yZuEYnE+P4qW5OJPs4PP
oCTi4sM+8i8x/c8b85un8JMvXpDeAYnk6MnAYqq/mjnkoD/pjaJLrzERYKxvXuMZogONR8CdvSQK
vvEbPom6hpc+L8q6uGmnNfsmM2Y4HlddRr42MmYV8vaTjGXqvyRikVG3uu0CPwWvwvye6WOCFt7V
OBnKlaNOJO0SNJputBJFdQ/ym4SDTXcWXsqOCGX6qaSRXoZsPLke1biD01Bwt+IFKiiJMJMgJzNN
9qOKwS7NrTxF6QdfnAok+eYBHLwaKqj39sMP6SotNf2rfB3X7asCVXLcWyceqBaX04INoUwgjrpJ
mrtciykpdsv8Y4cwcv3/Cs2W7K1zkufFjP+axa2ZarhSSWHHbpmDvbpeL4A6s52T2pt3SHy0LIhR
aEn0RHzvbHLLFO7YPvwYVebsstf7xtJSbVEJexHSAx5fjsnn6zlybo0dBEImHAsngZDP9B996WDq
gx4D9+TlfBG+KViCHykvFMs0VGZnIYkdjB+TbJ7JUSSC3YkIDLNAMlu3W/adCn+ydDiRrCkA5qtx
AjEo7TrFq/dUGhc8dLOrkh2VtoZiB+FY2x/I1xGFA+jiOS0Yf9mSCU3LCVbxyWO/HKdJ8naEROJL
N/CyJ5IjT7xjh06pguR/dCltFk08j1ior13be/WRHFHbNW4wmuT8hlTVavk+ZXRamrylAMVrnkHA
/EJHx4rN59VqUB568xsuaq/a4P8aHKDaCpNhu0xSJHA+H8ZOzsVl6AbIG52ZWylpfHRxj1MUMIt7
929zqTvfCAv0gLMeT8XJ0WAMruTLqE2Sri3IUqlX7brH+FApZDCFaxBFJeHNK8pM2mXsWHCqz+lQ
mvU3MEQUKnYpJPxKEV7qaSb7ykVZKM1oso4gkmKJ293QeIWH4we0liF6WDscK9H8MDXrvmfh2Lnd
sYjX03bjjHiTgst9nQRzCgdunyMNo5Qqn57FTJOR0qH51pkEsaDGXirW6GDT5EZ67D1bzAB7gMNb
A/hr7zpoM9WgshLDvAOQ22JWT79FGTEndvwhVdOGgYaP6StfBoMVY2KjenwBrgnULBhg0Z8BD6LS
nxvWkxqiWt3LzYj4Z/WgR3h0nanGzk3Xe360HQTs3cyv3hbUri4JrsM3OzeK6hzxJVP33zdX/2rt
Ugi96lcqVtMg8C1Jf0Ic/TZOHrzOoPghf2Qa3aY5+hI6ylPSInh7OrPsoPfyZ41iwE9aLHKcYeLS
vcsosPv+I+BJb5FmhKJ3RkdUveLcBwvtLII4/qDXq8eC85jUNnU5Bc3TGScR1Azfmy+x6hy82g1S
FV2a6zf3PeradwUkW0ymyOkaZXc7440qsknvG1A1ztmNbbdfBXs77D5XfRCzjkZpndMWZOjnZAr6
YMk69chTW9vCu+jiCc5ltF12myLIRKnwzznk1IjSham0iRn/wjeL8cy4KfuHu9Go+q25gzXf37gA
TLGOFtyWqTCKlk9pLtKhqs3S13PVCTtpsT6CcSQhOt/qX/VCWTILu7TWEHUTczoqkdiydQC/wSmz
PPXcHh2K7/3JzCxKf5jF9+axz/bOv6kIX9se6p8ODrKlNj8u7SFqjvWOzSTCWvOvH+YXUz9xJ4Gf
n74CBEuprIrROQEQT6oll0zA5T8NUFEv07jaonZZRGXa8qC0+7z4XM4AC/IMcq40qXtqIXb6dfD2
EOevnsV91g/Lf/5Sl7XxTxnO6YiRgPaViEsuCIphD2/Y1MAaqMZ20hv1iZz+MklJSs33tXi9FvBh
BQZ3RMUfRL3npT4aOl+AEUv92qFlOpTJjSR70xGS4IwlLfQjYQdgU71D+0roQ6Etz0EHVaGKOorE
Hyjv5jRP/zvFx+3c2qRVZ8Ox0bn3uUtHHeTBp+Se1VFTszMxp/a+G/2g5oSgBweomVqysQ0YHatO
j6n3zQWPofTARjnZu2Z8LJVDgHL4r5xm5LnRUIcrARPrthB1RAIBQOjbnx+LCzM4HwB/vgn1fVh3
jyTEFWRQIjHgrTmkA3vk64nZEXtJVYz5xzSPaaWmeHCctAfJmnu4gSEbRuv3czW9P0Pk4TQCwybK
TEiZqgbGkk76qXGS8PzO3oVpYWN5oUc/yb5oFSnhESJkT7EJK53k8R1di8Yxe0BQLSsxtphk7z5l
olGUEGFKMJFAwqcFsY1Y2Tu6qOlRUVtHckwJ8kaVCHqz5WBiAhyGKI6Qg5i3SUy9+wyUyzOo7Bnd
6MMwwMyUbowcu19E2OWLzAIDmk/fE6HwSwORA6sdeLbL3bqsPllL7uKv1C9lBj2QmL6e1IROU3D2
IlSw8WMB7CvOAj3Of0NzW2uJ/wVXWQLqmRSNh7PVfozEazK7uQSckQDJQW4Ic1o9dvh7GMgaDh2p
184EUqZ2dsiiUyST1UTu9+jMHWGiXgq26TJAIOJqWzGxJf8gB4ty/bEYlHfDOHfBiXeKx49LJmbL
E88b8omNkdxjw5KN/PEZSe5Ej6kZHoxPbUMZaLGDaeJpBqzCsPg9qZ51QcW4gzDSKmzcpwqABcf2
B+eBZHaqB4N+5KmRNdYeMl7BxOa/HyIxR1N+3PKI4OckhdDu3J1oT28iWGtNpV3SSd4xXJ9OFEZj
fV+omppa1EwWoTXBlqaIZvoFr5XHrN0Bde3adxvEzpub7PCheu9h3XXe5HFYol6YXOYnVtVrC8dG
XkyBJ+UqS0ILUapC7wXHXeAefFHWwNLPYEgReKjpeOQq05NBQwtcAufOBrnX4iLXlUQjEMx7rT2o
Ac2TFEIuzPvyiPH9l9iVS+Vi5eGzwvzJV/qH8TpN68zd7004BizRY+3p/lirBQe7uBQFLv73TzPm
dLyaa9uHQHFEOaixrq/N4j43FrzVuiMExTllPa8DzqST/hp20tFPqiMH2aDTFjLCjyUnLjgHJ7vU
cMCcEahMrBgYYJ0TFlkpFkNa/8f5s1pp370ErteShqfQ0o7ivokeCtwXoYJih5/Ydn0qqVFRO2XX
aJxChvmnoVhx2L0OUG3tvU0ua+T49P+PUy96D5I+IXBNQMJ8hYIOeWtcq9r4i7GIlgUwWxB2bELR
WJ7MYGOvE7sTwEg0CFugI+pd/7WvepP+kWJyZrApbm/rVRDkpteidZ2q/j8GAWt+2cAiLWF/0mkf
ohyJiIWByAX8ST0QlANddhSqtwsITnpjVD6Kn8+yIg/mfRbrjcT4vPGaBGgKWrgyCi/3w4bOYNZ5
QGyETvN/BuhC1qKgU3BlmUiVWqAp77G2PAZItqZr44rcg20bOzZFaug1liRfyM1K0NNRm+gvNouU
ZQqlXf3a1NmjNIU9ETNjiB/fDrE3CuwGlSbtXoR1OobCXaTxV3flXy3qTYqVCq9STX8emIUMRJHs
/IWxblLvgShKoKAao+/otXtZpinjMP6b+bPQwLkntOsfr7ZWxLkLWe2byAq4e/aXNvJYGXIuFVqS
mejN3Pv38smdL/uHbF/h6Jd2wrKW3sN7z+akBgTBYtL/iZ1gST50mrTqbu1wmCrRMvE0ttBGFxuJ
XhQihdIw+4qHnd5u6BG3SQcolQtuo2mUkiDy6QzujTCeyAeEzViqzxC5WedUkALvNUPs0Htm8c/b
wDa4ssTBvXNjZI0uEZOAFKxdN5AjuwOhBM4JSD13JZLfFyKM7xCoEG7PYa1Vim4RrxhH1VziLK1y
GcTKSYntfRr0uk2ZZ/NqL+BbfqPyQcijB3UQX6JCkeZdbAcR8yc5brIV9UiFWVFv45Unlk65m+cp
1MfMwewYIBxCcwagjJrv20IxglQQw8b5UNkG56AhOn/c50WkKJerqNzccXEDfq5CdJpKsOo6Nm0l
l0ToWIMsr+L+Dk4mlPCog51mLEHJRVc60yHZ4ReQ/m2bD5iO5f6TFfUpb08KFVwizp9N4pdo6jmZ
lsTB0PRopO2rixcr4nopE8P9HpuZdlTMbsdCtn4YVWtRq5YVpF30E9HCNNOudLaaoLSUzpfUnxWN
PC/YnDXQva+r0qdaydCi29WmWCo8a7nfoF6X7a686lwT3lC61EJ+xB4KJpSBpyw3TSm07b/ICQhs
7zn/Pgmq/rTyThtwwjDRJjkA5UDgfVYlJOk1sBR2cr362mRPgt34HDEbKfwVe4xlbUAyX3yHlZTe
SFvXrimDya4no0kvafLFHz5V4cl5wBWF546TK0MUSTmBjBKiU2vyLUlvsb5399J4p2dLLvwYNaQ+
T4bgqwGlAtt8Sl7Rhf5ezG2ja5tPSTqc144Kvw9/pnvgsdnZCujPiyXQfEdSElqYyj92jPlWtzXc
CIoCUrezLrMYKzTg2X6gx0UWaCM6hgXxqU2qL0nwr1wm+Yweq4bgdoDhWf79Oj90b6mx/yD1cUV2
wztxPfaBi3F+WBKjn0pYU1jP4+X4jUiGp/Zn344kU//4IYYYEHW/77pODc3SOZV2VchT50kv8m0F
qrMgZM1SyRJ7l2IryShLMDhz7RPVG6WkAoLW5FRzl2sDB0wQM2ewtLULxtkT1nHEplT7lAx7g3jq
89HNkhNlYg23BWFKiTtuhG70osz8nU4RpvwJITMGfeKgFXXUjzwDIbEqgymKkDI3N+JQwAqXTYve
RU4kaJ/WPf5+hhkRBrzojYNBKR+g52yl8h00qAz9h1SMqItsRO36vcXUGJpAGH6vBgeHRNWgxxu/
V7WBsv3UtDcdrNoHhc3G51o6wbrk7TbDfuISR+JpJ1CdMAPKRYj1c/Livp9VOAGW3kNs8iIqWZOa
0i/CN7h4rkK6YMnVwF179xEsBCQUBuBfDnIuZd2ILATf1mzCitAMoQPjeWU4VNDhXSOKShxlcqOm
pfdLtVQi0nfGkN4tTCf68esi8Y+QeD6JdzA7G9W67Lwt831SEBzW2TLEVXGiq2RTcPVpwiO6uHj/
fFRKqsdg99wJkX1H6/raX5534sG2nBEIJJxAF8065hjsI0mdVSjZnLESAkAZsuimkBPJdM0KBFmB
nq31IEbBtr2YtfpLN9Ika8UK0BNiR7DioC2cs4MIms0Of7WWzkHMz/3aJq/yLwRwRuuYfZZ60FpI
3XUu5SY99uoqKSfw5+Ud2QyXtqIdAok8emUQQgzgRmrJfXMufPEaZaKxDIbVq9FcRV43h9ipg48L
kdA2iinqgfVr0RUJtdsR+bx4JnlqLnphxeEq+8MxfYzcHPBGuwDv8R6Dr8GRikqUw+318wp4yasU
0/YYLZIZP/N2M98j5h4iQrI7o2RV1MY3CtLjxVQQVSyrhmHBc2KKlG9bC/3BxHtVLFnbV91peXrP
WfjDM4EqaJkGeE1zQI0wzPx40aCSycbhLk58+ThvWoWFt2Z5S5yqrXadUzBpWvGZKXUU7xrQs58c
szDX3N0dczrNxobdClD7x9FIbopf3suAlcfFMZsL1vv2/MnT4L4IH86KsxAiTh9A4w7W6kXw+YRj
LR/CQLxIKPzikj7pdiZE2QynuC8x2Yfx7j0hATQAxFbYb6mlpxlvCj/7NJOrm8mriVlTgD0aBBqI
gexo6ufztmvs5oUuoImCO4ncKiPWLsx6sV7tg6ILsnk5QVIuUz9EN6UfOx2T03ngsM3gyi/z95yL
rwxcmoItj8sJkBmY6peUVD2dj5Cu/wY7i+xEbWTb+cBrO2kanfNQnM1HMjjIY1g9ydIwkKiiwLXx
9v/rqBnCTXCxnsgIz+M23Un7w7m3gMg49EWq3bv9eH+qAnIWna+oVZ68Wo270wEoZTQaGJDfO/l5
yToCdBZ8KQjBj2UsYLIhYHORae/p67Vop1S3LUrPL5u7CDvlj5xqgHtM29kB//Brq8dyTcv3cqP6
L0bQvdelJYHZXgtSlfwaikQ6GiQeD1R21IUQEnfXRnsKD4ooBI9LV39/kUAsoHE9D4IJa4X5aV9w
xhFwncLhEpy6t6bEkv0UHyoWYLQVRg8OomsbdUY6R95yj7hI/Wznh/ROU+gU+fTREVlaAPHrgRIB
sAGdBL5CBoJeBtTrJmlECDiZ/yx2yFlD7bFm+hSve4yTdeU+f9OO+O6Rwm2fpqctUaFdJNEU0GFj
51JZ/EWIOGRGw6aCDJgqvy/sHOr2TAdSdAit0HEtcUxn11DIqqxmMwsQxINCOa5MBg3JVQob0E13
EIU5UHrtoz0J2ozyzjpVoJYRtJL4vD+rSW+SyotkeNhboYdzcyBsOV1UKvFSZJnjVOF8wJAT7Y6L
jYHms9hoc6tqgKoeAHnRajEHULa6HX1j9hdV53uDZw5raWGGmzn9j3WWIgEQfcXVUiF4Rb1x0Mw2
UWpFScTpQhaHq+2NHxouZzGSk1kuUHUP3ltqmXqkhH2uMbYHeAOlmf9ISkS/9KtI4z7cNUCvV+Bj
KCluvGCRbyHnzXOdWXrd1XvB/CKPFerxFeiIwe0NjHGUqsUCE7YDS2jaegGZgh3qq1bzkDq+USM1
M39GshHnZXJnQy77S8fFe0D8EtwqVBfbxlsYHp1pLVdahyTrGMrtI37nuktANuVsDhmmn1gWOur+
N5jc3CCF7TNO0cKWvzHXbklR2fclcRkSLjpecR5Y+6ZN8wfH9T60sgvwVsJ4uliHqlTlt6L2QpnL
EdafYW9iYirit+cT07pWwkr+GKjR0F9Cx9hbfdAS0qzXkyW+PxgcytrDh9JAXFvS9lboktCdeSbM
30+JjPZebF2mfgIbwMwBMP0mZHusjn7eR04ToqeFW+o4pJi5OPfXkNYUrRb2RSklB3pt2vJ6CkNc
K7vp8QWdNckino67Jk+43YK0yy91VJ3ClusfYcZgsc4OjubmNuCqDJqqtm00gsSucxJVe/4Qdlup
hkipTPbdkdUKwx9MgjYnt8C9aRzS8wMDXmAWqMSuRZ2phtfoTk2j6+kiGKblWJghH69YtEDX8IJm
m4dwbnW+
`pragma protect end_protected
