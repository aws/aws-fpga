`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
V13KFaLxe50OHgLWJNXCv7VHz4b3k/ZRhHEQlP+puWHeesFcSX5GAMq6FezLjBWwRQm2BdBnoazB
afKzHSXRINVPOjMtLmeUvfEOMy4ghTdpA5KaaZ8Km8kH3Uvhz6db054GwRqp+tJZjBR2Ycz8Gq6H
Eg7ismN3KCX3jAjAQLjbqj3j/tFRm945M/OdPONIeIjrgHPWsoPipxMybKkzNzZ61zhKWDZMe1Of
LdgrMbFrqnG6MBVGFcb9rLVyutjPB2YGcQRiWzNLuxAtkLUs9MJ8EvScRfsXhQTul0ihy+KFR06F
uvjnV1qB6WhEO2cexfV4lh6sQ7mv9PaUh/UQlA==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
MDT2EDN0xoCyoiu0SE1LW/EhJMz974VM1wgdYqZ25aGbq2JxJRz9l+6jDIhN2Q47I65DT6GJYWGt
XK61cV8tHPPKRKJfnadBEXFHHmOvJq/qiR9gcYb0XQbeFabXFZxcasoD1J6I40dmMiPZ1R0KtfXo
mA3GNSwNZpZaKDoXSUo=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
FIo1IFkNUC1rfiO14qqDFO1LdIIQD2DPW5VtLTHBT0CThytFsjiUS2Owi9PRqwUve4EzGlx0kOp3
sR3pgK1ND4Osv13nNXQhj1py3Vw/zZeBeS1WKlEYMNvQPl7FqfZXN1TnoaGz6mu8wINu1s3oalG6
CHi/nnpC1q48leig2Gk=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2160)
`pragma protect data_block
zZvz7ea0c0hbs6M9hfAZADODuWNKY8xiMphrRjCni2cpz/Tibl2ShXHYQ3NNnrz6nHcT97gg5WdV
T+ccXhiQiOH/8qS2jEdns/X6ikUHiZVv5j7jG0qHDM9iTyeEfb37SlDxJ5EfKmxrNTQ7LcREinMN
e8QXd7/dzrXhMRhg4CJYIetaPHKOy8qjKK3/iHFv7a5OCGLFZTn3i9JGnh3CLPK6iMyzQlZAgiXe
vDe8TF1copxh4uwthHBr5SYqrudep3+DluYNDvoK2mitE+72RqPms9Zwy1h3JDghVOyeghs/jtEU
bdvPsI5zj7u1xiQaLN4s5+9Zx9IDGV+ACjmO87ZnmTWl/Rm0GURW8u2tEak3QFPCo4yiF9aZP/2c
zJEBCPLS4NQSO4Ecvmle2IUK82eXx1pj/oPlk6rgqnJIAIEI8YnHBUrX3FdO6OwYXzZSd1LtLRqY
ii3IQjLap4fGqjo6Wu7ai7mFR3ZbHX74kIOIHjYnGrxHr/MtxxyJo18h9axFyLPj3d1W7zvlV06f
JEZphd3z4I0kXtMX6OZ6TRdPkl3Zi8BvBadUAQTj5Q11NOvUkNOvoDdZTTZjABnTweae9x/3bp87
wyQsf9i/B/HhsB38rbj4gHNBscZLAGxaRBo4FEBcaU3QAK8agrRLBraWkIoFMeKL/FPISnuh+TLm
b2rQNwxvtpjxh8UP+pLLQ7nd0zGVQA6ikVEH+BCGHJLit4E8RHJKgVG1lqDTH8+HGwvDtiaNwVMk
DnLEb9Vf00MbYBsiyb9V0xWsjg97d3JTvgU4+lxVZNqQl11hWCtPkl1H2Dlb0w9NAlk2qIZbmimC
xktZ0mElIDPJWHhXSaUBVugRbnueAGdEx5RxKxEO2s3xqRsnOsIr1JSYT/XN9b04/tDtGWEKpxPp
4g8x84I64CYcBe5/fkQZ6Hb78LvB/KMhmudPzlR5tMR5WoGXOvZ0+RQi3YQIRYG9Hw0Vx6xIBC57
An5Fd4ukUt1m3eoMtFoMe2OIpXKBndxWsWH9OPEHIPHmgf2RbbPqdgW+H2rAChwo+g+SSe1ukWZW
dlQo9RXxduIN4fBjwqC2gfwcJ5yXIgcfNAZOkHgy6pI9MmUmKWTutVHgIGZmgRX+C+CDqHWTUUQk
uCDVdRRnMt5Te9AGu8tBUCq9rzBWYKVWl580ubkWrhSjEYIr8IoHs1T+jAmd8gG5VYWUL+c+Jt+s
ttOfKZunYyU19Et2Fkr7v21ChpYMPA/3cJVEPd+JR1YOnXgX9Tt24H/0B9rVdtw82YmMVomLSr3B
NXiJ9PZVr3cCXs7JRTqcmFVXSU417lACuUVbLh2l19qMZx2ev9WXisOElpYp9DXoQr5tfBforSed
PcT6gjtahkjhH45IAJMESP30TmW923rk8W7/Nyvprm6lJknS7Uo8X76TkxT6Eq1Nhym5uVtIZz6d
BLyw8N4Ul0xtJVhi94nLH+XQ2I3/SODIVhOUtsalzY9sIq7CH+P8kqLwD6EN/oaocCs5aafZy6rC
/7Q3vgoB0O8OeTqI59ZJn0I6gf4JNy1eUkiYpVtBacHt0sXLZOZahZd3Rx4WELs6FJBWI3cZ6s/8
+cp4F3cNmg1Hqre0Wo9lGXmoTSgPnBpONrwxdQ/FqjZw6YRfUwWYou9mcgYoChUv+kVFUpq7vtX7
czIw9TkgqUW+RDyBcosFemcI9XIZzHuASknpy3aXTbibHcQxOWXLGNG58DT806St8hZSON6k5pQO
BIJGUj1Rjhycojs22VKbrkwkSp2wzfCS7P0SJiGyyzTJP06j1UvWc2np+qdU3RtZdWAIOslH0lxv
CtTgZE9W/5J9s0gwk6GeWd6bh3Ff8joJRwQrnYsziF2PBUR1ll2Ds0KblMQO0yfDs3fDSGPJ+G2Z
D/HC2Vdf5BA9xAm6B3hFGlXczt8TPN9Cwg855YgCm3c1fsmpV14AbinD/HkgOcowbYaxi1t02jyH
q6RQ91Bet0YqPf4nqAamBc88RqyneZD8rTkpBGnbQW03AHDkA/dTeF+1NM00PAq8ctwa3CNq9a8X
1/lygWa/ab61RMgOk8W+i7xyl3JF2iu0Ii6/hcnKMmFWLLfLpEGCaBOMclw6s2/7H/2eqL9bSfdO
xXyjlJXnBf0B8ka4pOZXuFp9FE0oRqKWx5zuG25Wg2DZ5au7gOJvvcTzbs85cgDEjIksFOO9qORy
rF+ia6vs+DRxeav0ze50gqxnE4MTKeqchzvXcHVE5DZFEAFwXoq7K7YeoJFJVCdaDDIcXvKbbFu5
kCIEplEUPT9n51ZJ252TNdcitC0gAKxHdDrTqIfSzVgsozJ+CLpfl3BpWpVV1rDIaWi3h4WrUPsR
dMFUK+La5DI8Zh54j1w2aJomusX62Vy9EamhVlDrDClarEKM6MhlWhU7J0kyZyYxuu7gwZPucYZd
d1lhZhlMU5GKNVTmBVoAwvXpHz8+yrojHDMJOr07IuoPOSDJSMi8eOaVxWrKCGJlA+zQGR92aTbJ
DZb/bU3UHYZrmk+lgBtgl9aaqB9ASwdY8xSvc/KZex+fvxkfjFtMS+KMUpQaTc7OCMfJO4drWMyy
NEdgjgoRigo/sltnpHmATB/2mtpmrWlE+as//z5uGh2Gini0V8ufU6KDRMX4siyap/WXVuyDE42h
BzHK3dHPMXq5LLCNr/liYxOa8PIRQYdSwN+I34sjn+gnuT3sqrszSyukd/M83Yg7JiYmyj3TWEes
aPjZ0u25OgsY6UumqB4SFsAOottarDJ2muYfm61C/qu9GWPyuDKRDbukpTdWwqU4SjFGT1co9209
eHgOr7vbj+UMl2YaTHT2Vy/y3ERT01Fa1EjlibwvIL71Gu8/YrXKyXKWn5kxiWatYY19
`pragma protect end_protected
