// Amazon FPGA Hardware Development Kit
//
// Copyright 2016 Amazon.com, Inc. or its affiliates. All Rights Reserved.
//
// Licensed under the Amazon Software License (the "License"). You may not use
// this file except in compliance with the License. A copy of the License is
// located at
//
//    http://aws.amazon.com/asl/
//
// or in the "license" file accompanying this file. This file is distributed on
// an "AS IS" BASIS, WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, express or
// implied. See the License for the specific language governing permissions and
// limitations under the License.


//--------------------------------------------------------------------------------
// Stats interface registers
//Register MAP
// 0x00 - GPIO 0 - read/write scratchpad
// 0x04 - GPIO 1 - read/write scratchpad
// 0x08 - DDR is ready status (bit 0)
// 0x0c - DDR reset (bit 0).  Set to drive reset to the DDR core.
// 0x10 - AXI Address - AXI Address for accessing DDR core (refer to Xilinx DDR specification - pg150)
// 0x14 - AXI Data - AXI Data access for accessing DDR core.  Read or write this register
//                   to read or write the Xilinx DDR controller registers.
// 0x20 - Write Words Low - Stats, number of words written (512-bit words).  Write to clear.  note is 64-bit counter
// 0x24 - Write Words High - Note can write either register to clear entire 64-bits
// 0x28 - Read Words Low - Stats, number of read words writen (512-bit words).  Write to clear
// 0x2c - Read Words High
// 0x30 - Self Refresh Request - Request self refresh to the core
// 0x34 - Self Refresh Ack (read only) - Self refresh ack from the core
// 0x38 - Restore/Skip - Drive these signals to the core
//          0 - Restore
//          1 - Skip Mem Init
//          2 - Restore Complete
// 0x3c - DBG Out - Save/restore debug out (??not sure what is on this)
// 0x4c - XSDB Select - Drive select to the core for save/restore operation
// 0x50 - XSDB Addr - Drive  address to core for save/restore operation
// 0x54 - XSDB Data  - Drive data to core for save/restore operation.  Read/write to this register triggers
//                   a save/restore access to the core (with XSDB Addr setup at offset 0x50).
//
// Interrupt Status0 - bit0: AXI-Lite interrupt from DDR core (refer to Xilinx DDR specification - pg150)


//--------------------------------------------------------------------------------

module sh_ddr #( parameter DDR_A_PRESENT = 1,
                 parameter DDR_B_PRESENT = 1,
                 parameter DDR_D_PRESENT = 1,
                 parameter DDR_A_IO = 1,           //When not Present to include IO buffers
                 parameter DDR_D_IO = 1)           //When not Present to include IO buffers
   (

   //---------------------------
   // Main clock/reset
   //---------------------------
   input clk,
   input rst_n,

   input stat_clk,                           //Stats interface clock
   input stat_rst_n,

   //--------------------------
   // DDR Physical Interface
   //--------------------------

// ------------------- DDR4 x72 RDIMM 2100 Interface A ----------------------------------
    input                CLK_300M_DIMM0_DP,
    input                CLK_300M_DIMM0_DN,
    output logic         M_A_ACT_N,
    output logic[16:0]   M_A_MA,
    output logic[1:0]    M_A_BA,
    output logic[1:0]    M_A_BG,
    output logic[0:0]    M_A_CKE,
    output logic[0:0]    M_A_ODT,
    output logic[0:0]    M_A_CS_N,
    output logic[0:0]    M_A_CLK_DN,
    output logic[0:0]    M_A_CLK_DP,
    output logic         RST_DIMM_A_N,
    output logic         M_A_PAR,
    inout  [63:0]        M_A_DQ,
    inout  [7:0]         M_A_ECC,
    inout  [17:0]        M_A_DQS_DP,
    inout  [17:0]        M_A_DQS_DN,
    output logic cl_RST_DIMM_A_N,

// ------------------- DDR4 x72 RDIMM 2100 Interface B ----------------------------------
    input                CLK_300M_DIMM1_DP,
    input                CLK_300M_DIMM1_DN,
    output logic         M_B_ACT_N,
    output logic[16:0]   M_B_MA,
    output logic[1:0]    M_B_BA,
    output logic[1:0]    M_B_BG,
    output logic[0:0]    M_B_CKE,
    output logic[0:0]    M_B_ODT,
    output logic[0:0]    M_B_CS_N,
    output logic[0:0]    M_B_CLK_DN,
    output logic[0:0]    M_B_CLK_DP,
    output logic         RST_DIMM_B_N,
    output logic         M_B_PAR,
    inout  [63:0]        M_B_DQ,
    inout  [7:0]         M_B_ECC,
    inout  [17:0]        M_B_DQS_DP,
    inout  [17:0]        M_B_DQS_DN,
    output logic cl_RST_DIMM_B_N,

// ------------------- DDR4 x72 RDIMM 2100 Interface D ----------------------------------
    input                CLK_300M_DIMM3_DP,
    input                CLK_300M_DIMM3_DN,
    output logic         M_D_ACT_N,
    output logic[16:0]   M_D_MA,
    output logic[1:0]    M_D_BA,
    output logic[1:0]    M_D_BG,
    output logic[0:0]    M_D_CKE,
    output logic[0:0]    M_D_ODT,
    output logic[0:0]    M_D_CS_N,
    output logic[0:0]    M_D_CLK_DN,
    output logic[0:0]    M_D_CLK_DP,
    output logic         RST_DIMM_D_N,
    output logic         M_D_PAR,
    inout  [63:0]        M_D_DQ,
    inout  [7:0]         M_D_ECC,
    inout  [17:0]        M_D_DQS_DP,
    inout  [17:0]        M_D_DQS_DN,
    output logic cl_RST_DIMM_D_N,


   //------------------------------------------------------
   // DDR-4 Interface from CL (AXI-4)
   //------------------------------------------------------
   input[15:0] cl_sh_ddr_awid[2:0],
   input[63:0] cl_sh_ddr_awaddr[2:0],
   input[7:0] cl_sh_ddr_awlen[2:0],
   input[2:0] cl_sh_ddr_awsize[2:0],
   //input[10:0] cl_sh_ddr_awuser[2:0],
   input cl_sh_ddr_awvalid[2:0],
   output logic[2:0] sh_cl_ddr_awready,

   input[15:0] cl_sh_ddr_wid[2:0],
   input[511:0] cl_sh_ddr_wdata[2:0],
   input[63:0] cl_sh_ddr_wstrb[2:0],
   input[2:0] cl_sh_ddr_wlast,
   input[2:0] cl_sh_ddr_wvalid,
   output logic[2:0] sh_cl_ddr_wready,

   output logic[15:0] sh_cl_ddr_bid[2:0],
   output logic[1:0] sh_cl_ddr_bresp[2:0],
   output logic[2:0] sh_cl_ddr_bvalid,
   input[2:0] cl_sh_ddr_bready,

   input[15:0] cl_sh_ddr_arid[2:0],
   input[63:0] cl_sh_ddr_araddr[2:0],
   input[7:0] cl_sh_ddr_arlen[2:0],
   input[2:0] cl_sh_ddr_arsize[2:0],
   //input[10:0] cl_sh_ddr_aruser[2:0],
   input[2:0] cl_sh_ddr_arvalid,
   output logic[2:0] sh_cl_ddr_arready,

   output logic[15:0] sh_cl_ddr_rid[2:0],
   output logic[511:0] sh_cl_ddr_rdata[2:0],
   output logic[1:0] sh_cl_ddr_rresp[2:0],
   output logic[2:0] sh_cl_ddr_rlast,
   output logic[2:0] sh_cl_ddr_rvalid,
   input[2:0] cl_sh_ddr_rready,

   output logic[2:0] sh_cl_ddr_is_ready,

   input[7:0] sh_ddr_stat_addr0,
   input sh_ddr_stat_wr0,
   input sh_ddr_stat_rd0,
   input[31:0] sh_ddr_stat_wdata0,

   output logic ddr_sh_stat_ack0,
   output logic[31:0] ddr_sh_stat_rdata0,
   output logic[7:0] ddr_sh_stat_int0,

   input[7:0] sh_ddr_stat_addr1,
   input sh_ddr_stat_wr1,
   input sh_ddr_stat_rd1,
   input[31:0] sh_ddr_stat_wdata1,

   output logic ddr_sh_stat_ack1,
   output logic[31:0] ddr_sh_stat_rdata1,
   output logic[7:0] ddr_sh_stat_int1,

   input[7:0] sh_ddr_stat_addr2,
   input sh_ddr_stat_wr2,
   input sh_ddr_stat_rd2,
   input[31:0] sh_ddr_stat_wdata2,

   output logic ddr_sh_stat_ack2,
   output logic[31:0] ddr_sh_stat_rdata2,
   output logic[7:0] ddr_sh_stat_int2



   );


`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
dVzUBpXWl3SUrlDYkqUC6kTUPggnVQv6M+Jzp/+EkbdBgAmKfHHYByoimM3IhVaueD7mScU2/IN1
uPpzbxyNpy8F3aFizTrX/0qFWbWHdX5DRoK5v+VxU65W5q3CsPFfRfx5YeuIrjf0+Z5pIYR+9yS0
XRYM4QCJcJBUAGJJIt7O4L58wATrLrEBEqljbxkR9c0Zyo759EX8ZaULH2w478K3EUgFVly0r1MS
P3qIm4n6bSHIPPfkunc2bs1EQH6rrFvEGdjl2UXOjpALTEzwrJkNtpcwEeK1NQQCxk2Ylj49bcw5
8mqVO3zK0F49rCdVFfh5HsmKBTbqp2RjsrxVQA==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
NncSUCW1DM7EMZUeWYWUx4KltzZtnRg3f/OpMvc4EFwmSoVN4ypQ0Wtz75vyNxsmd2EJaxbasL3F
FPsNNuRuhOmHW4ZM6mdZJkAjyLdhwDJmVv/iU0Q+PQfM75zIw2LK7/jPlWb1AhswM+WO3O20T1/S
Nl/PKmSjpY2xTrGhjbc=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
UylrRK/EGsc2eOTbxbOznPJUEaazRda3lFgUmEvUYwy5q2hv2PdTCGCwKmAbKlbjUwg2muv6eOLf
GUvLQzUf8dad4FtYdWwgWbPcfAgs7SJvORAn0hot54mw18FZU7A8brcsGT4GBA01h2BOXkA4u9MA
7fGEntenAqcVEQwu8j0=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 56192)
`pragma protect data_block
ohUsUkBNAyweAYY4Nb4R9dTq1+g1ebUEiwR1xZS6SKeOpKj/IXuoboYLNaQ4BkEDVDx2gDQgW/Op
zY/WoGJOFnV++7xUGMyah7I3CuImkJj7amoPaVPnMcVh5PG9HxkRGPQqNTpZ3phpWGT3EMCvtO7e
G1ShQ+j8o0rxbweNxheJh7FrNmY8UaVS56gP0nHmkoSJJRZ7nhuG8Z1JA+Zltgxm1BPE4a9y7NhX
kSJV70Sy9srsn61PGwLHZoo29lyK96QLFikEwGjQduKyi+zlUHEDtC2hAR11uFKvh5LQwkit5CJ+
aYuCADx8S2NiljjJmQgfJN0epMwUk0zaoMF1eYTEyWBtAYpw5AedZTMk2RVffnsVvP3DDE1jLwu5
N1PhvQ2XZtt4+KZ9K0ZeUYozbyav1gk3ggsBi1vzRcu1J8LXNtjwtzYBUdv9ClqwCjHy0JCCHzSC
HsNiLLVC9dksb5niA/RAAXNSEOTAQ9xnhcJqkEUm0BZoXb2j7IpjWxeLiNevRLG5pGg/MtgtGCpn
AucbYpGHKH+o1WMr9ql7tdQ2weL9/XAHsguHbmuExMbshe2UeJnGYvAu8TGu2sQTKIQuWvDXtTjv
Covqx85aLhPm0t/uC8fh7WcwBuLB6Nky4kasQqajloSXu+0ZFwHpIpoa1utyFc76aB1yiL/s5j7P
+SMCnL0uqYrOsE+QOuE9DP0yL0WAVgkMYyuVtqEMkbBCxWb1sqlhnJxA727awIeksop3TD52ylQ+
UPtJrwliJNLT/kIXlS+rfxu83bIMliMVyb1hVdk37E+FIaWJt9ZLH36TPj4qEepUudvyiHxT2wnD
MjK7XW5ZigzlO7KcKPQTBnS2TBk8JmBeBgR4VXj5R7cmJSzjJRE3zL4QlR1hYoZ7YZLEGOdmZURR
V1mIsmWzPVFdLsf81jaVE49X05G9VOoy0AYelW/EmdR1EziPMurH3IowATKyNwpcYWKxrWfiDXlL
qUq6MwnkWa99mpshyppddBqpTqF1xEqot1xX8V9pDJNYNjA17470BXJJ0QB2s4+yHG25T5NLRz+T
EccXVjKVsQQsI9IiHEf/p+imNDT/9d7BQC3LR6I3JfPPGzl6XOiEe/eWlx7852GZJF2Ouh8pE5ok
PL/VPui/o0QQ9mePxkaV9ysJIgs1skqJjBwUwKLDLt8ehJSNSBnSU3ksxhU8sPIa2grqR+Q/UY8Y
7sQppmI1EzDfUiCj66+eCV4aYtYn4fvuyi/TygwSct4SfGTZorWODw/f925Vo2SV14VwkFnkGQre
ujrr7mxZrvb5GMh6dvF7mOq6lTeqXbNVlMweiiBhWnEXxOdC3Ie2wcZmTvGH4Y/Glvpz+LiU9FTb
rvd8trTVmwJXveb7lipMkbKaUsIfaLS28fgNUJ6nI3Epca9roekkqOpcx/6+Y+P25yJONsrTmyZR
lEQt6mJhOBFT1jYRDw49Ny8eOhVVmsZg7YA41JduVjRxvaooCiaK/Y1m7KMFz7h8e2j4zp7rPh9S
5cOxM1OtYApE1RpQaEDPhLvF9BILcpmD5lSDF81TA3W2vygRA3LbMwmvR7dtdWoHlJuHWLFK+b9l
bi9ngMdtcBxH/FHbkWJRLIGmsDfX/PffdQ3KYzlX+r8ixZ04scMZkvKeIl3MsOI2W4XvmeOjqET2
8vh8hHhKso8X/zZh9XZ5JPw1MCUFYkfXKGKsOzpjcNeMvj3IAuP+PrWYjR/sZt1aNvevT/KzxThl
fdJkcvGl0LNdCEiNVYcTI0UTewoqeZxcF6RrQuoyJ03lnxhRO5Gi+Olrp7exch9rKxD+cavyMsVM
jK9Cee76qahSep0l1+dt2yZU6z612y273fp4PFb1AoFIDWOx0psYZeP51GJ4Bh3qQMLQk8ONSa+U
7gDKyz0MzlA3nSfg0lRAIFrDSyRxid/K3mzWi2S5mwXT8OW51NSHPqh3RI4ae3Y/kh4Wa6l0WIKD
iSqQr29tyQmExZ+J+eM9naoKAdXuiWMRplmLxeEICKWxxVR2CM+5j+m6JX3qs5Uz7Z/SK9Uo8Ycr
TAoIIQV2nxw0YhuIzyApU9UyjDDN40zl04vR/1Rpye3A4qebKuDKmfJkYpoVVP9gky0ERXwtT9ZC
2qa9pKlZSgd/V3gYKv7pVTNsnJYIvrXw9waaMJnbYpseeW3FTFKRngZOwrZ915VyqIYoCLPmhPyk
cRm3Zxub4A+xy7map6Zfgjv6fHhoxTe8A49d4qmbpP/08yuoj13wtZTvwjI5C3mPO+opk1JjD0qf
F6+qnzfoLhAxzlrLZEUG+vBp8VN4JJpl3rBRlSdAb+yCa/64Hhvup/tsB2s5HWoZgBl+20JiK5R5
Ff0AxRAQ5W1qMgV+BiGC1xQAZfRWaCUQhQ/DExA/fx19hwHwLOn7eSoRRnJfmTmuGK3d5ijE9bmh
rY7USJD5zmwfHljYp9y2eB3GC/NOwhubWISeDc7QZCT7afP8ZSaf8zLhgWZ5IR71QvOBA7L539XM
/o7wfPIf7cZUVsl9mkz09hAWGZ4Tzx2E/rnYDkBOMD9BeucqeN4j9z6lDu/lQOSeRpI4EBrh2TTK
w8+Uv5J5zX93csuuoKH5+Fg/Wnl07OmPldbt5RVabw7HjGrKy2X5IYVJWx4r8CRCXfpXdv5n7GLI
oATTyqCKqnFpGjfpT8CZtcas0ZVK8eAqD/Or4gtfyY91Q6zayOsqwHBB8ZZI89ykUFDlLnGAUV8w
shnR7xuXEBJw00JP33OopAtmFrqDn2wkKdie7LALy8WKoiENHvQ3ek2DxBOB+qf+yABMKXmUTzHa
LU3qMtlzHly8uNJ7aWlWHbsNBZ4hRiO2edDc+w7kXxGWgKNi6UOHkpJRU315gWxfCEnCpbxo2ba0
Qn8jF3ByUAZPU9fEEKejMgvh8IUKDWlI9HnneTF5zDPrJHqt2nIbNGq5UzMH98RxWwFf4+b7NnOg
ZsrvrH8HVBGDlqdYLx1UM6dfYZBDJ1ZbrM2uGmqJRRRw1Y6K2YE/YDblLP4Ld2LjmxDQxwEOm726
KxP3h3BhUxpHatKWg28Q8fj/FwNn0INg8QRI94va+RME8xv0EJ/FlVzL71q/yPbFFeFFOqSfAbDc
zmPaQOKspdYrvr3r0Cl6+JU/rhDJ6oAE3Ll+VzNFW95bhEaSf10g8Z8WXAOBs0Fh27gKBGP/bv2S
IJjf/CQX877iB9A6ES5Kzc1q+I+bCJLHbBlEsFAAgYTJeyE+AWNVJVWdanDuoaS6Cu9lgwfjxw0z
iSjwqK/99DwUkxmudlaR2RK/aZp0eMjh4jPmLcfjLZRiKokpvsaPfXUgJoAdTGqENXkABG8RSABz
S6UUuEVlh1NxQVXKWBqV9j78h1IhhjUVd+fwHjZl2h/WlrNfHGRd+dNRvsbxIjkMhcLst2aCR/3N
yoV9oOyBlcp2yGzoFlrRAol3B4GLJlKv770BuDWJFbvYfEwi+WlG/AX72ojEpsmm0HIRiDe5rd19
ReBXQ9BD9UALDSVcshpfxUA2cJRYAFc60klrvXj+sRP8TER9FzRNk/3663UHLtIAUD1MZybmit4t
PhVhz5mhuceuad7BMcTdFzxSY8QrL7fztEKVIQRAiZP4WQH2NNO5aw95W8YoiYi/ectM7UHpO80W
oeNuotpV/Q2paon6oQA2P9+OwsTuaW30LwXy4e8IBLRJPB4IOZOe2pdXcIbN/sdLsE/5N6ZdOBvR
WJdNDlK4gVpdn8fnTgEgqdy34wk3rizkR6SQHKFgK5NSPxTpXi3/JAb4I35dMjvtuotU5Mm07Qi4
YMZqFMCnHPYU1Kz6UMCvQj0c9AKxYD/EYqv1MyUUityg4i+122B02lJSdXLoBilkr8EnkfWcg5cT
mq3eP7wOPQ9fBdBm8QFz7Z9YuhhOyhOjCa2lbPCt/sMrI6mbJE2ha5/9y3wyVXUiyHH5U1kvPphI
ZqKKWxoqCXS/+QwTsyygES6BKVhjBVlwKzgk5is4d3dh/xX+EmVMisKWDF6QxXCN4dhSsGQ7wriY
pMxSQJLayoE/k4SgDc3iwlqlIWZSdIXRf8kSa1fwA7iXtzVOyDHwvHq6jfzuwHl5/8Yt/SKNj6dW
f238OvtGZn3ddO6R6oInmIeYH8fnmOcZIC1USdObBo8wIUay1JIXh9WGqh3Ba3iNuavPGcPUNoE8
dmqTJz5Fu+n2yhXwqhxUipEkoylERVvmsYyY+YsN0RCnGJ4H62Y2/EAliV6UtuqZQUc/ANTj0K4g
lODFKbIvd3lZXLU7moZOpRXJByFq6a2fYx6td+2Axr2pdBnadNvUtnhWPEQjYMhYjCVVnzHKLSxs
XAWORdS9I+hAshrzLsiTBTqbyOIZzOsbv1HEkTfvi/eACckL2X7x1GRvRNGL0tpoBKCXGRDjxkHg
MhOyl3zJkkkJLY5KDy4ybNWSik8DdamvN0Q3YLoqL9t/vsLVFYp0nOx2UTk3N0tZqiV7HYwvJwG7
Yg+l8L+QWsbif76gVss0s0D7Nip68cPDcrfxQvZje8PG2CHgaf4H6oas9ZR67ABFOBeaBxpgXC3+
+NkTDJJsc0dqnqavUST9Pci2xDzsNN1+JdNioHuxVAtK3tUH5iHsbKPpaxdgEFa6vwS1mBPKGXRb
BWA7JnLoHEkF3xW6gJClB1jYS25u4ca9SYjahNyN/JLHW5MFDZbhvSOg2qVplk3c+XA08tRS/7lG
PUHshjYolL5Ur//QHgvDEh2OJaXITvZZroMtSxSqg39Nbg3+nlA16V0caFjjf2RXPNvK2hyIhRgL
IFAk6LDSJDfAu7juv5Canje7T10RmoGQC/CLKQOicsuQM8TpggyYeKorz9G6aIkThUx7h3XNqKIH
42fAqYBf0iWVEtXq2Pjz74eNi9U1v8O/lc5XSDmofIxULW/j2ipcVLOXmtB+GZBnS/b5QbD4A81q
+7Or5j7mryjUonzcnSKVR2eTbIQI3ZD3xFh35MpnMkw5b44/vR5KfoBhkR31B8dMAsipvrHD3+P7
M4hYOKiUXHEyWnUnLbSi80Ve0X6RwXbnDSWvRJa4fGIyuSIPoF1QfJ+c+5BE2gZvhOpwUo0j2hbE
W0eZZQufC1pX7J0fnVo7KYdrqthsr7SWNVOGj+eX18FDK4RZImN0u5DmIpSnAVPJcnN2aXXwE8nv
FFjLAUcldkJXBxTTrBs1rNoOGYyi8uuqeM8j+virXvQKluLbDKQWAla0I6DXWsIj7uTfMYXymlSw
eSfPguiSQqG4sejMA+BTX/vaBi/TJkbbW1RpOFJsbRQt5ANQzNeU1xC0eBuXFXdYgXak4RMpCwOb
YT/gUpBRJLj/W5/fQQ2CUbiIQ/tQCXF4fy9+KeEJM9+qMF/CDlqyDejK2x4iF9EybomiGx1VE2Mn
IftMcR320pONI3Ta2/1ZBa+dn+HpDj7goB5p3FD9O4JFEV1LeU+aNM9vkhvo8EB2kD1++p5ML4EI
rGi9BkyxxIIvDHKwd6fKqzLrfPtDWh9DGw06kXGRPPLwPIQx9feR5lNCCjI0XEoU4HbT01/XV/Ms
GfmRpz8+rAF1kKqbm1U2QcqHxpTVxZl+X94/iVQcnlhuZNwiTyuw/tA34K7a/HGDN24FEQIp4uKx
TFK1IL8wfj+Gqv7u2rgPWSxzrfqxEoJr7aCi+3ZYZ70jwQ2xjrOtjgODiHT5oZfwzO2D/YC4K9dH
2a3/2n3HAGV8QMd6WTbTA2XIlqJpWvncNsL9FgBQe3BL+BFV1QDj5Lnkx0YjHLce3euOGVnXNNEw
GfVyiQsKpJLlhzHWuV1rVtAPJfP8Iz3TobittlBWX++8FU/N5SGG4OS8ARPnULkZFr6cQHSto6FK
4q5ISMB80vPIlUWFQ3AEU9QPpD8sBNEKiem/cMpbqMwUV4q/MGG/6FHVXIWx8AmzaQD/zZT98oKs
72CfH/MLvUKovf65xoi6DfqRSzthrmUGuHv2fJpfO+S+BLFzM5hSfhmwKiUS9PxAX6E8Ipe/mjhv
gOaqa/kwQm2dNeKqtoGNbDJsbG9R3vuOI22q5ML6jPLSCwWYhYA44dCPwqwQJx8mvdHxyVFl234+
8bY9UWLbOeDNVxOqqMvbDosT2z+6+swjj5Gp+nbDTRjAk/DrU/AHDcAwx4ejpXKFP2JU4BMvhjtY
fZlE5I0LrE+QIVj+QMj/AnrUhbKl72yO/uT+1qm7i6WSMalFBo9ZKnHDKsKO8XefSyLA6HIzY4XT
TYNFMYCHP/KDvJNaN8tGtmZ/wyGxoUXk3eRukfPWI9oV9L/Cwy0/GiO7bBoGZDAASuAq6x8saCmJ
To1e9rKQbJ5PBgfwP7MhzUGqqV26T5uc/JRKSK2fs9Gyzh/p0mAY3Fg7jSdYK8cMzw2JjRNb86wj
YDVZVzy5raVn/w/PFKMQ0kVGCzookBociWhIY9mtAgd2TReOqQAf1lybx3b18klGp5ChJ9g5D2nT
Pt28vnjpCIpeZKojcpQlyzuD+VQo4DQD/Jc/eTeLiM7nHWsPQnNcEfNIQpRl+GVb8B8ze5XBESWz
nWDksjg9Ipnn2R5voXtS6njEogaP0aHxV616oDv/xZ3PiF/f4Fvw6npSp9oCOizTAK0jo1E4wynP
xi9boXJP8lIlFR7yxEwFozg0w0lO6v8Gbu3am+pHnMxWXx+wNQ0QmpNeb+Dg9L325xhF9kGOMBL1
JPdyXcRpcQKlWhVw0cyKlokz7XUCPv5tvJCUd3O1XQwaZGdw/CJTBF5qYnLAzByqWRyk5QhGWswD
x/ZhamY/Z8Bksq+A48I3nu1DU7YdB5nAg5B5qF/Excmzuh1Lhe2mQExUZ1jGuXJAXSHsrUvQKPhH
EhWB040pxVggjL741oPp7YuuGu7MmoQ/8p4kpE+XfTMUlK7uNubsHeHfGKbKubOJenUvVMgp7D9L
vA+wG9z+Ix+Fbyjg9eykC+04xr3LYoHjbuMiA0/mqgEecWgfr8H90gnpGdJbAaChWJ1Lta4gHNuD
2mcepzhVfiZNE50Ouxh1Ysr/g6scNK1oZ3/GbRbpoBoI2TsEuugMgVwUrHJVWIorpVFwDdyNe/XN
QdmltP+YBwYlLsq/X7r70ez6MDZoKzJ8iqjTLSPPo7otKbB60SXr/IxPLh9GAdpsU7/62DBGpNaQ
3/qEz+PMjFYtFvWxmqCfc3TxaWUWeQE0uKXUWiPMpLGhSWo2ZdjBCFnKP9OoyBBBqOyjqVMlq7JE
7+r0D+e+coYedv29c43sDWkwjLcRNpdk30VqLfTgPOV0QvDSrGZHzHQfShH10AB3gLEXK0Uj82wt
OT8ywoN8x/cNVfFgedsvy6OuPThHeBnjNzpMmSu2N5gKkpd9WAoi3bvBgBWlQESgV/pX3kqi3ZUe
WPaG8EqCH6NKKpkXVFp62QTjRjK3t2DKntTjsC1wgpLjCHYlYX7m0FdWeLCA4Z/voIIsLvmcc1XQ
t3xXlT6zNYaLq84QudH+qoKHLL8yJoNTrF91GNaXkC1zZ4bIt4Yb4DUyFZY86V1s2Ark1v3BCDAT
6jiSdYN7iSTpjCpLUwLQ1tSh0cjMVA3uL0qxTAEivnKLBaeX+u2Soe1vK36+pPD4OdBxACXVlUps
t/N9X/K4uoTCG6D8/ebRt7mHjP++/+vw+nNyHLGgUYaDDt5agt14U/mDKU+jVLu4iRKPtkP6xE/0
i0FTdx7CFHQyKj41m+hSeh7FHcC/NAiLg1ZT2Ye9rBLcvUoNvB2At33CXYJSyEv1UbnyDQQw1s83
Qh5L12wczRxfH5dzkKi0rWMwpIKMojtRcGKdAJFPd7h+E3k8BHOiUQRoP0r33ophF8NlJgwlcMxU
brfAeJcGGPtTZief0LoTr+dRFd+s/JWd4qoUVwSGvVMEoNofY3eGjSirwh9D9GrsAb5HQXAUcLgn
hp9PH2IuNNWfab65056tSqk620m+H0eze+kfPLj5ajea8c2atAlIdMR1Xlf9mGFLuNuJWvDw673/
xgd8RnyJGGR3a7m5PBHPjn5+VXyMtIOjwEW3kDqXaEc8wWcxhYARytvzOdAZCb4vVYDE+6bx2AGD
p9XpLgtuL803K8nLsJXMUDnm6nIuh1v2JneDfI8mhqdsJL7vtl48++8Pjqbx+mrZNhm7zWAxLF1v
QliE1N+pu6ltY/LTFn+u7FFmcIR+TOsXpFl6SgV9G00rsxy9EwpLif1UHXumWD9JX9ciPrYklz2c
0HuBELdFiix5wIZ4i1hETxYQaykKEtXfeeEaCAKUuQXRvQxELd0yhEGhVVk8kL0LdceAeF1OJy60
YRBwNn+cj1enP/PmBLZV3pF6n2gtpPVXskSzWV0UJsVV4uW/dYAGDYOOcVehdwpzlfhx6kCoK8VY
cYaNT3FxmommsfEaT/JHBJHCgWBapoEx0Mwahm0DbJTqeRj9lqMZVDu1w5Zm2rPinQ5valgQ+wyC
/zFZ7HLLNmuIyoCzbmPD93qmDa87l5QEPCHWpdaUQFTmnFWTh8pl94GgngaiUXoAiCTPiuolacid
fhJ1gTR3NZ6dgB7Z/DaQk2DsX5C4bm+QvyhFJs7QLN4h/GZc+uvFB/aIbxnYVuVwbI0Lw1C0UUpV
1rv4RldKES2lSZ7HHaHTAkRijmyX747kkciMOKGYktjWE3iwlsAmpwoMsFot1efC+j5aOHFvaiPU
9eRP2PMzMjL8xzWno/Y6bz5ZdOu/XBaMDtzsflynlFYvqUtZbLu19TA5UFAg9MzDkEymlICY+ZAG
MM10eaJv6O/0+Ji8n8F+hJdltcHw01Q05Mxzv5RicKRELz2o+3ZNBtO8fClG26VCA20GTa58G5AV
IT/5pSbp65bWvmRdsxPgHMdAwSvfY2wclFSRRMv5GgKAK90U7oE25L93LxZszaGogssOtUfxddMr
WjdKbzIxJw0fsm1bQT6fIU8eh9lpQdnWC14u/SR0Dub4gWmDL/D3er3kTxEDJzktbhMT/HXId0a8
OMXB9xQba9F3eB7q1dGRnqTN5ZIf4shyBPNaIc98/a+K25LV2oBQFXI8U/1BneByOHWtmlr2NOeZ
O45JO3irD9iY/uo+ntBjsXOss6q09KScQSuoXJMSWhekH+v8Uw1uFqO+4sfxG3+P63q/YCjZC5X9
mW4nF2dG+urKjwSO2iC+lAJw6xJCg4SGfHoBDtjEkrceBZj1xziQu8G2TWylvtlslkd2aMFzpxWI
O/8wH9QwHeetuY8rakrA/+YY0ihtET52B+XA8mp1xlgpTQEXDN3ycBL2tzyB2aIgL7qh0Ybumqzf
BMdgql9o1zmOnk5k9h1f1s6m/QbOvBeqhPq2tNfR5SHiDOzVOyCwXgK2iyBCNMJvFOT0rkdfGe7l
BGHHcBR6Wbf4DxRd5Gh3eLTrqShVJl1vfPfisgG24qbbYjFWWm3djdEbWGtJ0PusB+K0s+NUk5n0
YwY7Lm+ZfH44W6cYPRzEyRl2l32/wWosnXlVj2Y18KiWl5sHLMBVL1i+7gKzS1q74IVG2kpQABp9
8taJ6ZlBB6UdUnjF/IUEXD6TwsDQCJsvjynJf1KfcwzA0bFUOYZ38H/NFYGffrnOqmecC06HIG+3
CMjBJZVJO2unjgt37gN/u9+ypy5XwN0epn++x756HwaPVKMPkTJBueihBh5rhG7NY9RZzcEzt9AZ
RvVpTCa/76jOzQ60S/unUKS321RiZq4JsNHrKaJhlMrWtAADdg7BSkXoZCZcUSC5XagpHdA7myC4
kAmHNTx6Mp0wOXxakZCpwXUb9s8axB90SE2dhdyXdOLmeGp76L7jfIT1oEhc8V0NfuQWQFWZLGHG
im1GzNpYsSpDxExCQjFpRQ/LMVgX+x45gywUqyX+SH6sYgHLElYtKw1Swn7wymE/ptl1QE38c1UH
dGLDenOrzbRJ5T0RUgasB3SyZGPEZNuseZgCKp5X7Sm4HHTUGNlK0iB151/fpQ32egwKXOneNXVM
Au88rnbePr4RERbVfk3RqXEcmEXwyChJVKrfpoNbK8VEY2lMZVXWFKGuAAKsCYmnE5nhMe3DgEQ2
dTeKatcFvlq8wmrnUSK7oKqjaAo3PwxbQtGra8K5nwQ62pkymn7HeaMtKsdMf8oWRm5M2Et5t+W9
Tb1d8Nf7lcwwJ2n3ZyiCu0/mzG+tEB1KX4xwlopbdl6JHTvz7unWZ6HoOHIBTqvbXyQOuLt95DvK
KXiZ5XSNRY9YTLgVj56fteAdI1/CLPkDiJ8JQKQi9C2/E4xFwXk1qTB7jiYGDemLLyoQ25VBCd6J
U8HuuyzLro6L4wjxSDuTL0ZzJCOM9REjIvZfaZFGlUu4rBPo1TcKvfPtze+98UnkZfBSBu6Kdbr2
Oe7dzbkGKfGR5vsEeEeQvp0ZeomiSB3KxgyJt1LQsiYXhyb1MwERScgxYRp5GQkXxJcsWjAvpnWT
faGehNqbpQGVj6xJSPOVWC00m1hy1NwExOM9zCedJ06U6tmLmWLUBkZc/awOrMUdKA1IGR6FK9UY
3Cz9Fe9C3ZDgwgWhGaAoTLCqJNNBuYcPjSFR9xRIDYU8CUw7YFKam0nMHre5mH5MlhIEFth+V7fP
7aU1qiG+GekUBHYR9UQ1vy6lsziZzAzb7xhzjmitUOMyrslPEE6yzmZxwaEog6UvIKXxvZNcVylo
kK70Xuc50lPoPu39w8BtB/OL12kaCVkemFAyU+qxgVyhctkmJ26KlwV3/hFSnFU47+HOk/KwBR2R
vh1De8NJr3G9P8jrJLNW1ckILn07lVWs3GGpvXf4qvOuUJbS3Th/iMdcJoW/z405aZTWTwdVTU2W
CLH1fE08FZ5MAajfxWnOQu0fxecgIAURHOhZZvzP1RTkERv/O2ynhP+q4fTRexCoYBTajDTblYr5
fsnHRcRoKacL4ozyG6g+0m9o2J4X8XKmTDiTYp38nxJh2HnQPV+HAZnvhxDaiBDp5MGAM2N6gnqB
0V6+70FLzfj75dR42wPjucR5XSv7g1oUVtXnJAmdjWqrQOud4eTPbqoHny6axsY+5KjeQoO8mtn7
00T7LB9aSL+ebHYWEZ+jkssc+Iu6nY8QwxCCGT9QcOA5yi3aUAt+wgZ2Qg9Jyya1GqpADSjSqfLF
AD/aP/DmdrUY3yXt9CMyZWB9wfHeRTAWouAm+Xah3aYLLozlT/R3Ap12UKXfdRtrLqdG8TbSa8Uo
1paq/B6+xH8zYhb1se27KRKhMtgsIv/NwG6rC9IsU7d8vqV/+YvRqOXA1WzhrVKuXTQ12GNx3bZJ
qYyakvUDVy3MTIKbpE6/ZKBFQPlyw/7EgECEHRB+GvM5JtUon2rieoGFTtW9C0pLuX9F7/9tH50J
uQyVPd8nuu2bGI2kYVd7wOBm75icwuUy8a8MAIqOxKEQb6JmI8MHgppJfrXtIta/iaC7AcAcgP48
h3Lh2/SiE1i1+7N7k3FToQSI5E/l9Z/CGGMvKWbPb2+060ZSr8pNA+wJ3V57oeeBzyJNnkfjuAec
zfXDovvp91wfIgK0OlJdYhrV/5ht6+EPSGHjYzsx9Ecpi3x6sjPYFrOir4NNNfI6TdiqBvDjNIjQ
lRoTb8MmNpuC+ZNcS7VPr5LJ+t+dXtF/K7ZkeHsHR89FZEQ9hlgR2XZhJRPLnWEf9gK9hnDjpUuO
KNZPHGLz7hy/B0xLoWo+SwgloxbrsgKEuPc0GKhSOqZMiMh03tM4tMq0RB1tQHeYHVNpKdtZhJdG
bLHotVH7zRTmnZMufJs+QTlvAijZ+045vq2cFuZK1+dXdttGZFD9Lny1k9SGHR4GRNkukXSRTz3m
vWiqAKTQgwm1fSK6mRmtYpOPhxSGsyrng/I+olDnrj97m1Tf2PkOPGPp6JSPeVbUVKfaNct6TUB/
Oe2HNEpgDUbs8XNy2uW+sE74Usz7b1n/VhCTwDqaTCIJx5WLNxQ0VRYX6dmpn8qV5FE8r/93Hx5x
rW8/gF9i3qpOUYV4DCH8XeOe420UxgBoYhcWbpPy9dA8qJqF9MWQIwrpueSF0+5+ArXJwbjXboN6
oKl5HVBtFu8eHY3cSKWw/9ACNO+UO5rZADx4+g1vhufG4/VE7jx1oxqdT7a7BP2q7P4kaJ2kbaZd
oFNDEVV3UskCakq+CA1e76dPlha6BckcKH/G78WoEyA8NvivzTX9wAy4aQIzUmr9aHaLreiHPjcF
4wSZfc7VxEUNaY6NdOBa+1Emsfj9eI92aDTBrYtIBWkn5D7lUnuS3alQ7FX9gH/ESWV7zODVx4MP
AHe4uFte6AK2gOUvb1tJkMdoJtWf9Giwpsl90+Cwb6T2dsu7lSX2c7io4Nrn2wjHCSrdxLjlibhO
mJgkaExUR/Ozv/t8IDjnmBwc1vnTN1ElHfrV1ALQtuPH7rZWc94oKl/qgE2aUA91Y4lo4PM4g+rf
r8DqK+SjtFpw/ecxBeBzG5HzXD1cXxVquGFIfbqfBbsCkY25yIybVXU5ABB8WrAlRYDusZviTH+J
Pkxuufp9EDJfKb4UVDoPt/1Quupq8AI9Rn8EVEBLIh6SInvgRG+qPNdcV8p0R6QJ4WQFGKTgLU7x
2RI7vfO8H3QSDzrftNJL+UX88VklN9jQlSnpwkeMgN7fbdHDub15mZpX0yUcjb/RCNbovdM36byR
8k6voSS4rTbLOPcWm20k+PlKVhLDl+tArwL4nXRCxdeXYtN+8+aXt/ZgTcTyEWEDjpenJVO0J9FU
M7C7mzIvzIPAlARqiRaIgy8t/mvVeJz2HZs/Vupd3iI0c4CDtBYYO59D7cFIR44g6F5dgwBLc96R
+sCXOkZzEDi0tsKcvMiDvUok1xH5rHMsHvnTg3YXUX79UxLbelU5oa13XKfhwCE8KkllOTS5XDhO
ZI8W/64OPO6Rc3of1uQ2sRq/PHVGjWPaMtweJhiEyKPhyTq8zwEJTqSmVKs+Gx1AIdZXpELJR7LB
x37+IfWfE4sKmbXGevUfoeA7LBBu21hRkC6bzDgmHd3TqYlB6cnCl03AhLRzljMbMdh5ysaO5y9N
8c9KWBRE3rQeKRa9RnmtJLiOxxIIDRFIHyi4YubwJM8hjZTAI1nX5xq9GYei6XyQyUjaTYkU7oWA
2dzxt0Vx5DGXzntn8bcwHyjDeApHRNwf4vsNGWHo0GOix7MEAxuNvzD/zydJzgkNkUkKFVEOyzn4
BtsrvNO525i5T+wbVoqKH3+wEsIbSjc13y/JFqhT8zDZhjm9yZvReJ+aZUiUkKwNaF69CNcm66LK
g47ssA9KJ5bmDVyTiDzsCiEPyRE1yU12iSf2bJXjWKIhcQ37xq0kngCPZ1rUmMGHa4TUWMn5OQAG
FhrVS7NFrzSCbPnG7TyciVnmBxRfX9ZH8EC9abNPcp0/K7FRmY0NukrqbrlcprkDfGKhpT09r/d6
HSW9a8WXpUGgwOwUoWZZmVEckvXWk5JFS8W0ZwuCZAnEFukthLOG7yTjYr5uC2Q4LhfNW+mveJCA
4roeyTtYTxUevL/rSklkL4diGkXfj991ZRwwe/0AUpVMVhXidsaWUEB7bJR2laReXPdLK6snrkB4
PCi33wQiPIE0C0bwH+N07GNDzUEHQxHOt5n8QRuNGPE5Yp7fbyct7e/U2U41sQ6G365HjjpJlWsT
sjtr+iFyAKbD+e2Nbbw8k+XZdmaXJ2Gk+Y4aRrwg2KcclPnLvDwQje1kUvUttILFYFJ4s0Ap3kyo
DjV16y18RUCHWcQMFJN/INm0PdQfG4U20KacDe6UapHrbflfJEyd2Ip9j+1q88byNW2dLmdSGk/E
0d9sJJz5xqX7GCbyRgv2nABOMb1UWcqzGlmPT2Em1igu3NxOs7eDoSe5qkPn0lWi3SkJi9DVC0hM
88WobZkhc/r3azC/Gml7AJR1sxmbxWZ+0c/2c35f3nOJ+edRAvhM4knhzZ7A59tIkyEdGhP93rM6
PpV5VltKdxy5au5NMKb7Jib+EcknxK5GUtSdNL5Nurai7ryf/7Pqrq8OdbzdH4bfqD1q5jE9bZ+E
W29FSib5zM/O1Gn5SpP2NO9D97V/LBvCC595Q3+hnLXMZwcbsOYlwWzuz3+fjIGE61A769TsptN1
xCXbglwhDiffRKyAOm1YOSML9Pg3iKX2lzI5Ap9RWxav8KGxVxg/nhGeXR4pXK876HqIuIAaWtKR
GwQqDIN5cN0J4l6SzBbkDnJleL1+9TTUont9Zbqo7psgqCGR46MLTleQWM/pQED69OBBfQFkDhQZ
t3O6uhBLN0gjQsGsh+SldOV1wSZyB755Nk7P9CbE8C5fQMYTSJHCTU9AxXUvAJK9i7h3LtxPXJv6
3UvmszQpnfwC5bX9vFhCs7TDfa08yHgmpZI8trdZuv6KwZ74VxHR89OH0cbjV8f8D8FTam9JGhOt
C39ik1wFJX+WleoPh06/2fMd8MDZJo5g+WHyv6AeVUuiSdU7cNhPPjNS72Fu0K6mDX7g1cxgay5d
eimfeFMU3+9DIGnuF4C1d0CZGhWTP1cNQ5VIDrNMLnVld9PweWQ27gz4Z6MVpUbgH9weWFWCnVwc
P80twui08yXS68W13sn3ZC5CwwQGUJRQZm2uBrJj7nK+Lku2x51jaE0L3qqbHLAo1+B5SLmt3ifc
LT/abO9rNHgno9bsPsOzJTKJQV9aTSgd93bC2nP/8+l4thB2VV+LHL22Cpt+pqTvIQW74Co8Td60
V6N/r0B4j4DUv13dNbe5qRXAl7YU8SBZ8yA4Lbiv7jjPs2gxe6uMhzvTsK+RLwYFOtY+GBI8DOcT
QwSWNb2qRIzyIHjx+HWG2BBN3rc6eaBV5x35aWEmoKNLFkL5EtdTypf15W93SiMobrKSJXUAPIF5
1SuCJI8fLYXR5gzn+AYznMGo5Fu4k1JSC+RiEpfNoTOX7DICZeEMwn0UQHQTRyMGcH/FVV6pfzS3
6vdGTg49a3IBs7v5cVPVyoOGUxqfDNMNGQPmo3Z/Lt0LoCK/gAsv05RbxY2/xqcqnHKNHqyTO8zF
7QacMbRleiyXUqYlFsbO1YUYbyOISb2o3NF4rYS5JrI2NUwEn/CM7mH8m9XBCIbugB+sHzh2fxrK
EQy13EqhhFH9UKLfYkNSyWjVvkkah8NiwrHo7pS+7MiTAwT+7yi0DWsx8XLK4NzFmKhda70401cj
r+4ePmLSXCHPZ00OQcfx/MEA/Gm7k4mefp/OfItyvYlKwrHHGhjltaGXEH7679M3k0YGRmciHMa/
Dz7cubDDhy3Hm1vMcXCYyUbhllKpOlYtkEceKdvC7/HTSEes9aQH5QxJNupHaCf1hctx4+ZJvx03
c6h5bcdz+NNVgsTDmHRaG7YgBfKIfTO1jVpSY3xERUVar3G9DTOk1RNcxtPd+2tXnBa93tghw/oN
XMb5+804i4l+LPxgFwOCyaKxMdM5WaoDJI2keAXBq9GHWYqQkIYTxgQbOIdUSGozxsjuuy2+k0su
JICM5UYAxgC5IBW+9bbcib6Rw5bz+22C7jzu8RXjBSAC8p2WL81q3ghJrMZFBjPbJeZfelTQJFav
mch1RFDze3ab5a/ivZ7HC1kCxQQZeHbiaOYiJ6tVnEEageCz7AJEvscsS3aft0+zq3W1rqoTRkJg
NLQnhfGKTqDq8QPhXlOZ0x1V/eiCgNwacqKi4MQYpVoX93e32Rtty4pz7UcN9KHp2imlyO/WgPca
CH6zR+NwasfdHg8l4wL+4C3jovNO250UAWFeHhuPlEY+wiXa0ebQAfmaKGRjrGHPXkaCVEV7NWfY
BcXLCi640AwZLBo28WHOWYfoxfLreAZ4tkag2mKL5xYKEG+ffF2YbbZYM2X4rL6T/vwDGnVJBVY+
BcQ4Qz49PtO2KLkpIJj2UBWnopLU8/G/PSClmxW+jNytEqZFrSpQLWajrBKlMUBzeS7mWyuxNDF0
bxrLled7sx4zLYmLYI7eA04JzYcf4Xvecvl5uYkf+dlAqu+uZGFnM4XQVkmvoF7tNzRIhmFc4HKN
vnU76b3VXAcCnE0sfSLtt3qmIE1R9XKdtX7E23epx2J7LhsvYBC5w38Ig27Vofa0vK6AbRr7KtC3
mWC7ERcTlXzP+CLDbn4iorq2R4E6//TcVxJ3RzkCrIeUWXtDwIoySa6WLKm/6/uMVLHEzMP61u9Y
D3RimwzUihhBTrLcb8Zxxy8y+xtHuctcmZcQrBI+GAqaW6lOSxc8R+gsllqhtS60NyIGemrjWw7K
MAglK05ITHRMkaCkrGsGIrxg/VOyGkkv09qJPMsrKKas6xbdHJiUlO8bqFVaQdL9YF9DSODhdnII
GEfomYralkWntrYUP02RXv+MWK/fagsmYsilz6aiQoZTC8fnsD67D/I9ww9MKEAocgO2OUR5Il4P
S/aBcrPBrxtEgUg3CKccOLXgdh6GT+ihkR6jSj9I6WLWopLAA3nEnn1i8ruxeFM5pV/5Xv7JcpLT
Xm3BWh2Ptospg5gzEYemmX47VbfQUq4u+2TIHJ2w/6Erqnk1dkNzbwbIXElxLGR4DJM1ayx5cu6v
q2BPVdGvzMeE+W+g9BUZl+0aBTMGdreiTl5HONa0d++9wjfdH3oTOXDqz8NnyKXXV4KD2AibPXhA
OpU7kgdSKq74+sk+roWTyvnx3d/YzAt8KchzR+RNcDXINMX4TQaoSaTq6fcAhwK1TFa1nj5jlcs9
9VAAvdNkJz0CFA1Rcf2QJ/xBbPJfhFPDDWwIZuh4WQMI+3qMbd/EgwyNgzS31dCC4l8g4kT7L+/L
dK6Upc6YlpEePp07dLfgJAh5jw9YIDgxYKVgTCaezAqS++Yv2npdtSdC2s0wImV/DVfIB1P9yUH8
delX7182evfAkgVsltrVb/aTmSbIqkZZXW+EPUwetgrcbTnfJAvLT7y57aO72PV2vjq8QhBRU5FI
7oGrQy76c18RofS1BqYxbAjPXQjY9zdtPNP/cds6VB5w7flcuBktKed5ssuIrQLht5RhsJUiFGVj
jjitQMmhRNYhRYHZmGe2DYUFLOdCj2e2AH0d9Tpv9DJ51zQnrSqbIysxrFA8XA/+gDX2S4r0xjI/
H1DG+18RKI3gHaXdhX08nPXrXgbD2qUjenjl3n+Zhg4l2U6vm0UQxvbqRmhK7wCnCIRYUWYEW9NH
7P2SnyriSMsXppZxn+KCIiMYs+RhcBH1dfFMMmSentXZXBAeigQBKlkegWnCwHGa+uUxRCRdiQKL
OGcS9x0OSjO6ZXG+L266lDvitYCttkOoEss2ukpfZ5PRaZJIcimCJT6Fu1nCce7JMz71d8m6ya7L
+U74CTmjEH27vWYPy0i+8FAEyA/mQHp8s2OSFdY5qMhdtSRlU94aB7WV/tyT4oabndMbQ0Sa/f3e
ErECGHEe2RUB5BJlhR771fmPZ41XesoyE3DPIjMJb0mYhoZ0H3gUDG2+8tJSSUaAvecUV0cPdTH+
/bkGcehVeXxP2qLl5YT+lTVvFtp9gD/c3eiujcukoGKgMpPMkVxuzH+x1+1JDWfkfEnuSlF/0mWT
pELw4Ibc6PCO0dfMW4hKNOCzrO0p3EgRFdj0oPHKU9XbBFNRGgaeUDwT5Wj3dAWSVX0rltRikxjN
ViFHJW3LQQKILMk2UsOTjDerZby50+32dXet/fcwEkCS9gykEOoMD+9I2Gz5KmdS/O8rWcyWd8Jh
9vIAO7azR0y/5XO0hC0IC3PEvPiniBgvSdoERWDy0ucXQpJI3hy+LP3Y+68mjzW01IL69Kz14uVP
mhAnmiD0LJw0ewPAZGPN4bl/WeTek9Trnt9PiLPnL5+LXcqHUqIwQtXQQIyOUt8nSPvK8NN7A0IV
lncA1N9O6Gz5S7xzJbMN3OSINYHQYN62oZiKId9TKwjlRWLRm2XLnOAIwKwvmj3lGUdMDrVc4Mfi
4Kfl6ahRnU45JFe2zFEm4WA8MycDg14iseZmXj/WclWgMNQxKoYfD8nJfPsledsxKk3770vc71wE
XEm0i6FSaFdbZp9XwD8VqShZHdrJRauGuA2maYyAWpyaSpY2Tlv65g68X4R4v3ziWpFM+IC6FInK
L4v0dIOEgik12Z4DkKTkNUmYO23z8a5197Al4/Lh5+0T6d/bGGjUXLu66UL6bxeqbArTzOhe4EfH
TmwXgiiJK6odLhHGeIh84YvzrqmCPqryG0Q+aINbs3AZonbVVB6GTBOz03mLTnLyBJUkmfiX2tQR
sONKzso3AkhNUyoOaTf2kDNbeQhobsx5so6WSytiTKqhfwojXi3GKP6HurKhAGWtusIpACTcaLJq
T3Ibj6rVmNGdvfZdQsCZYZ4Vtjur7ReLaRxny5LsNlnphWbheT6Lhwc3z+vpcXuzvh5dlaU/+rD7
/PNtOqv79qABiclsA0JvECWeP4YuF4V6pMzNTbvs/7JVGlH7ucE1fsNUxIoYhpjOPnpD6oQqlz0/
BpGb0suLMbbg/bTtguBE7EHXDvkB07BSyrOgyHZ/zwy+/nJNfPPt2JTeqRBkMzrHC3mCETMQUwrm
gp/pKxsw2MouA8roLbnhLdh0zpN3ZHywhZVxh2Cg6yd2p7VYiT4GG77QXSxg801ikZ3jZbBcgYFp
j0l32WHmoiIROIFdVhyA7yOvkaS+RWKs0Dlbg6/+oV16VDXUrN1EYGSztrZX+u7XcFowMqTLBJXm
SqEtAgol1HuFPpP+cC7LGFWm2Jv7iWOwR1i11r5tZFAEDZP58hnX2/XGqxPa7BLtXmL124/SUoQp
q6NJHTgKYztJRWCTSfA2CHR6mOit8ZXqNIQJq/KX3PaKG/OiTNboe6IsHpoHcJ6ZgGpgh4ntYAJZ
MhotiGRbaFZOkiYmquOMmoidwE6YTW331g4jUkNxhYFIaYqhhfaREfFpqS8toGjJTZkMsKKiCuqD
E0vwUv7GxGK2h491ALFdOimZE4cnUEKVc+thZJ+hAfVAFFe5skjZVCvFi1ECYPd3O4K2XcyIRwN5
zfOnEPxoU31hllSozbkkb7b25ZBuj+nTB07RaYVitFnfPPFwXRXmN9IEyH4r5FrJAbhpdMKdCavw
Bp/nrqjRleD40T9nx0Ylhkd9nCPveXPUPg/d2eByJcU2w/USob/eu9xCcgbRflDoPYiIRxURpwWD
6dk1JcqXYvdsjTa2ccRwjp5XRTXRWNTiNlWfDLv7YJhSguzRxuqK8oNJnxeM0R1M0DkgoVj+/lC1
nQpd3j7Wh+VgLI5r5413rfgSZ+Yo9lRcGAg3t3mWMExmBglOIe4C10cY3MWaaHyT4knR/MF+xy/O
2tdc8m9AEYnyBMuFM0qHiF6H8vdFQZdpOPCA2ALcWpHKyPA2oHOspLHNATSy9m8oL7f2pRthIbx1
MViqMtckOUmtoxlkH81fN6UdPYLgMKWKEJDiHLKHO9snVmeBXALJFDvlFBI3kEoKibkzgSSpK3hJ
UIjF61gq5kZHNbvexJp4efndfobLO2JLLbx3oyN/ZqOqOwIxI9IDUxlDZ+UNVICVb/O7BIKeFsBj
+98YMoJmurPZAnoX2ZF8IBHQdutU5J+5C1NPEjiJG1zFN3G81LkbPNLaBe9qwZFPWKERt9rZtvTE
KtT6Php8EH54MwaZcBVeYZvR6iR8vBf+jkhXr8uScnrpWUn9caeKZAfCC9wWx5vr2eUD30HneXTM
/kGZJhX22csr5Qgn6voMh8m4MfjmVHpBoRbKvjT+LyVQkv94pvhRCgessXVb3iXWv67wQouUy7Uh
xhs+nbR9hqB5EzbqyStip6dy6oq5xAQbfssuzM8mID1yPvXP1rJb1VWtN9z60ue70mb+8SEb0+BC
MHX6eJZnyGEsFsV5QivUHw6M0gYJqoMEUF5lAwPZ3cfL+5yZF1SlSR1uhe4ef0iXY6fKH3kOVy7Q
7kbPbOo8TtyOta6HG91lqR9FB4UhEAgAQBPAG4XbOo3du1WgI6ZnG9yBQQbdg6HipPS58fASMNmR
Oobkv2y0a+ANt+XPn1H2mnf5CSO0KLUm3knz/cLw2wQVE9+nBqASn3bnMoFasnirUlHzWhlvxml9
g5iWQiX1FBQGi4RH/GDzF0PumUv39rTwqQF7+d2tNTyhN60XHog2pbRach0IKnvggah3uaXNkMKg
hpHnM0vCnA36G7yzaQzUcrtdQV9j2wawWy936H+2nPV80UampoCR5W1nNKkkSYKyy8mDNfhf6WDj
Z3MFfl6dqHzHWbskBxykTwq2JaYG+9Jsd1eST3QRCjhchuWCNgad/bAciKZZJpRDQdjhhNqAyQff
sGdNErYs9XO6GGYYQE74MHm68Kbvhmm7yjfif8dS08ydAjVoZ8/0JH70/+63trkRePXg3M6uLdoQ
aOyBxt02TcHvSTCpMu0A3iLjUh7HrSrOJpn6b6/zrb83Gzdz4vJnasBJ3AWJVINj8IrsVcOfO7w3
QH3M/4lar6rYqob5mp0nTcrH94tXJqZXvDcksJeBoCedw1VV5lGUVl+Cd4oBnnTk2Me3VR/c8UQz
Vnd4ySUbJG11jWjRO9eo/7f5lxCZm8w97ic4OedI9SkSjSBXkOc58ahWvm/WB4lOXsUQtZzxYLwb
7B3qQdKAKuClxJy91T3w/3tlHUI8Xt1Gej+iZl5tWGHnUj3ifpcnvdOr0kYGiVwyQyzouCI6mJiW
gfDtrUv1Ae33Xzgi7cekZXr82iQDD00jc8fyQdvxDfQTMH1kE3bDjtnIl1BgTjshtHUf3eHeTXN3
rUxK0nTC6vIWXjJGRzXxA8f9R+xeZC06E/tK0HPyGfy2qdFbspRv2IZMrd7bAw0R9kHKBd29KhmN
k9pG33juL9Qft4tr3Yzjvd3FZH+aJH61rq2ZuOZ67w7h5itpyfRi1pIHbKgjwQjx9+rgdrWwOS5B
WW5AHDj/DH0FW6xtFOOJja6VnAo88u46MtObCB7dVtmREqw9lyBV2tXu8lEVeNczrhsSGnnZl0Vm
ABWKqeO38zQxzK7CmXVJ7nEjiAjnLwdiFEbYUfvupN+1P59iEOm6uEc9rw21LXWpsQ5w/zH/wgW1
g4TDXic2ArrbxBI2SKjp1ncd+B8kWFITt8wOsslX0y2YQXV/G3Og7uONU+O6/aDoWYppPY9n8elR
1ctkdCoZQO+0a+2KTjQQfsgMaj0VClltlZPFfaMgKCD4bG23zujCrwOzJR5Ehf4JDGkMwjIdR+jA
8zI5rL+oGbHbC1UhpX9cqzgMygQPiDxm8me3L/dMIE2o6f0Tmxculeq6P4ME0IeO8zrzIjzWbz5T
6bAzbQBsRlAGIkWr+9C/7zuH7D3NxlLZGe4ikHT9UB0tBMdezYct8h9B495/U909eeBI9vjAU1pE
qk3zLINEvYTOOcwxCjXOQswvBkzthRRXd2q0oHiW9ndPKUF3tr1/v53oyHQJJIa1GY6xniDrVia7
ODjJQ3nloYLhmGoX/BqTS7my69QHo4NYTOLuVNRZgJQvIlmsXjyr7QN7nYHKoGXkVYi/cd38rXaU
GNqj6ReLRibTCg+CVqCx2jmKXrs2puhU+SdpF614wr800Bx1/diKrNsMYccJPOUweiOZCJ1UScg8
9kvp7vZgz59HuKJFJtEgAAeCKOnfOWmChoAsfDIcs+2sXVAbbstkVR9AivGWpMUZKqZcZ7hBTTaA
FwFk4M0Cq3M+LIq7jVCYk97scMDVJH7PAJdPXyIge+67oXv56BgfgKD0ruGr27xKOw9e1Ojtajrv
fzLq5CYTFuRW4KnTPGL0BM7qEf566QVAsCsCNi62+VvdPy/xT4K5izWsAUWQkCLifi2uVXKrx2zi
0aA0ZprQeMlmkG3Ig+dI6V4HMcvxrZ4J98Ho2ZQc1y4Y3oP/s9p4fTEzY8dNmUpIILXOdZhKcaen
n5lfB0+UfDDGErLUkhnc/A0dfhGBjLxo7Xx9UD7eOtwP62xw1vSWz/k819sL9xyNGfsTQirV80BF
0y8L9njcOQKdzlJdJB+uligVVGriEf9drEXCjdFPzPxZeDsDwXkgtBIVwifN2bIkDGRiGJBU6MHX
KQmUxxWpIRAnMLody30XiwNsj7wnehazPiZ9D6Mp9503G2mW/3+jhG11NVop1frZ1bELhjrQ+99i
Y7c6diSMwkOk8GghKu5O08GvE60oT8kUESsIfsuJpmoC8QEE4lf/NDT+qQGrzfcNJod1iaNMzNT4
tQdPkaMnFiPiE6GFiQiPpFo86BX8s8ORQfjbrQHOBzIM1uKAJTQIzS2We9wkJ693nyhi0b0OIUuY
rUHgP6lFUOGbdysSDwiqL0zcZ64QQsBA+ru7Rx39ntYIqWYvkHFL/NWTzydyMU0YZB0LN1E7HGug
vERLRmeh1AyJwNs4jZ9R+ymIOCDwk+Ftfj2ZEP+Ss55jZdg0UL665NEO9N4CT4DcJxgurt43iaZE
FDz5JYoKJm6ijU47yzIHuKEBaQCgqYM7tk//Ed0DUQ7NcdTNBx8mStjmYJUywhhMANGAg8dfNqqV
jSaBvRwCChUTdZ18+bguYc3M8ZkxQPWM4TXf56Ho17+15W4cV3llDT6FIlLIRLpZl9eLs/UNNXUs
DSSC0pZlv2KKINP69xydpyzQpy09xmLplJxShglydFj18cGnsY1AghwB7zOljsXF4uzjlPcLKJxH
g8sZlePhuXkLTaTb5h3Z01/KDooKUM7aHgLOSJ7auNh1zSKjth73AV+pr9IFznqajtkowWnG3QgY
WPUGwFY2KrZB8QsW5lSOVrle8In/kdip0cxR+g1DsVxfE3fWy02WMnO0C+EF8D6UkYgD+rR8Cp5P
TpEga2+evjTzHX+jzI6cLAka9tL0YN+Xmjs+2KItWJXHqIkiPMZNIb16nEx7xuJCB9PFFdln7xlX
io+c4uayEA0noM8jAAYsmskq4pU/O+LCptzj4MmbWy23Bhz+1rhp4uqT+h+WpullI4FGosmlxhZA
4cwxQwidtWLEbNllBvXwOuRC6PlLgthWbGcDr8AHRJmpWqb8YteKIRw3roOP7lUtzw9IVbdhB6b7
wYuyKPXmayQ/QoNmzTxPqRwOyINfWLZb/chURNjWluFanYEoMyVs+5XYXyTqRfZnS5TscOzG+Ruj
HwWaqY3GylqxjVSYEHT7Bh9/Oy/bE38XBY1CgtRs8eCA1RiH6zhF0sN40rKPacTyITAJneiyPDrS
+LHkTsuYJX0Zn4ePeRAAiDWuxM3kHQrnqkJYBIQ3VGxiBxQNqANuFJuts1ifz8+eo6SPA7oiqM/R
vAVVIyJcm04ibstayZl6JrbaypqLKibrS991z6N52l9iJhLBnxp7Rih+9LzyGUeP2ologqulEyPH
y6UvNFCi2cXaSkkB0+XxpVUKGzwP4D34FIo5knyczGtm+xiyTGzEzXw6WHwhSyJ0kpHzUp4kGb+F
iXH97QKK0Ez42Tt6E4GWmrtvs7z2PTShDo2P3ASPczVeh8y/rpOyEBMk20D9KBO/wmRJBIzVFYgX
/XK860O38Dofp8VT5XgKSOhE7kv0wfpHEE7zVhwq5wcGBTgEpYnNTVAVLm2VOy3FpmRKJGak7xAD
bl9p2TCQMhpI+EEwF/rFOLQXVMbFq+w4JyxzrhmiDlOtzUbyTsBY1EAZfa1CNUB6xUIf1vJyLyyw
BNpba4fBy270EDgZMFOWI/Tk/ol6oVp8YkTDmPQVstm2rC2BywYZeKWlNMHXD52GGb9y6MOiGs0U
j+YyWQtov8lF5jxYdfwM7f8IdI82e3h10icgUVwXgnsQ7O0ZGF3S4Myoc+CmQAkJC9eUJnhALWeO
Ev/6kvykijcaC8+d4xXct62iT5chVmv+u/3OESurFDSo17b2PNbKzMmDvmwZP2iGcuOSsUr0NS9k
c3I+R2QyHpUTd0QQCApwhi3x/XEQRXFRUnOyD5TlIgHfKDsEb+w5oNKGCAmGKAVnZHtdxb23hK8U
Lqb1kNxivc5ECPVffyUhhWmDyRCeROSMLhx7K6S2YXCHT4Z5YNHtUZ1OB4spMB/WWvPcW+DescHi
ukXl99X3e3lFelQtoW84fXY4zopRsR5g86cDgDPZwdlUVFvyjSBq+Z5/HDnKFwKVHTTWb11HBLSN
hogRAI4YQEIzTomTkTQzZWwYawXb6eojuzqDAk84wPMZ67lB50hErY3zOUVwMHn7KvtbI07FL3ln
R4n5etRsjGMBRxPd2lbstaYC0AUBFvvN9MCF3d9/CkIP4X5dYJu0TJEKWPobJRNhbbuQGyn1sR5a
SnPH+Jd3bUQyXZwM7S3SDsq3eOP26t4IMUn9xZZiYALO2Soukc4iERTY/5B4F8Kia95DrA11AfHd
3UFNktUMMjWMSrb9IIjzeg/6oVrMPfazwJCF6aCZY8KT9xYMrKV1Viqq26PmL/4RdBPFxUI4vQEg
SpSbJHJflShc9twBpMSFA6CrHoyL8WBZAK6F5zg5Y2rhpf8Rh2VjqzcNFbEmeA2gjqiZ/i4sO0e9
DpciARNzMQV4Rh7jNext9AWWcldNSB1VWNBdomWgz+2Q2iDU8QOU799ht2Xpmku0meLWkZc68fdB
mJ8mqcfGRteRuCKF2R5g0xEl32WOumGTdizNSFQYPwMMNUxzBtjwlfrAwN2qjtZlkrFfl6DlK1CX
UU5Yel9GsziHOKAeneOPTCU+srCX8oOG53LMLxiaKPoLeMV1BYBotZ6vtU2USO+v+p0JEXWIdnDu
QPKcwOdGEHXExFZuTf96qRri2C+QefAsu7TLroK+b38tHkDDFu2wNU7aLuVkBsOLgsrNXh4EYHE3
XrjK161XMUJAncLrYaGJrku8534htpvvJwPXuGtdBuRv5SGzqaT7UWXgOIJmXnHVUrmGSbgzS9Ic
7eDA0umFMvK8jRL+KwkfZpLmOV4Ft5MnV2VDY5SyGIlcv0jo0B4qLwMNHAGuKARcl7Dt53hzCbBa
a76m7aKrJaE4pmu0PArxbw/KNgNHj1D6WgSNZIhDwW865M8VkYw70QnQLx99FMV6NTK5tOpUs+rj
+EHOC2F6zEb29I9VUiF/x7Gu3oOB1LjR/fWK0UHvgc7iq61meY8I/0VBWNniUOcAQNQCQIKa1sw5
aCMTiKMqU2K7eC5f2fD8468rdZ1zuSB4UAbxuPpsRpU7SEksLz0mBNANPMQ+N0dJdmpWLOVQibup
7NuI786v09BCRCxYS/69dI2muTbhTAcQ8m/qzLRCSUemxp0MjHxHPiy53A9ppPJ6/Gj1PMPq5ZRt
M2VSNds/6kbK8De70Ll/ENXyN5U9sojo+5cFmz8KfrYf2i+XikWJmr39EMKNb7mr4la1S9tNvx7j
/Vve0Pccy5V5Fjx98qf8MfHSUNvrCBdEebzpGx5T1G4zQcy9t+h8QA2ICvA1OU2i+8Lun3KY61gR
pjv8ItHrX23wX33hfbpjpE7NDpDMkwcLYwkebngAJxdMRUvartW7/O/BuGpARY+mVYv8ltGcik9N
sILbGG2JMCY6A1WYIOF8GlJgJYHaQSonoV4zAuH9AUbpYIUQbWWdoZ6XbKJmJ0wUlUhbLu/tkZzC
50UaCpGaFWARKs9pvnTmpctUDeywusD+WvFBetZEy7q+iTirj1wbp/0AJUwzPe+OCvbf366Ti1v1
uQt+R72uYIdR68BnawPMioo9F864Ypwu3M+8dueJnNs3HhcqMYZ3bj/W4Ywq3JV7o3yQMC8i784E
QcuYBDUpG/iH/Io5XLRG/5/I+4JKr8sLYzoT/cCILazxT1PIT+Dlhfxw6MK43a/5hRyGjtDKsHnw
YFEkRlZ3V7FBug4Fdvic7d4kBhKUqpxyR2UhbX3KH+4J68IGeP7c4JqsSIRIhkfIunSnXbY0kNcu
guFU2j0qgqZpcdnmFWuD9r35dOR7Q5s3RTu1utBb4ypcpMHVJOVQ+vizzwgcbYsvEbG1a/rCG2QC
CD99x7GloijFTBDffYkGwNYlelmG8wOzubcilN+dZyIRcFpWBl+QtXHe3Jw5TXGkogHsEyrVUGaD
lp5XdWlnm1nT6JH1a7G/4hGEUQtau10gee7LvIgBlrC6gYBR4ddmP22syg9EpiVZYDJok5LgGzLj
dtJ0auspAoUHNaUbB+x0rON/eNkaDrcT05OLtp69Jr9qEBpKF05wRX/qGuUgrw5d5jxz14yOgVwS
9njKj+ijosjpfWLbLHxFXtojMJYYfYDZb/soiROsi1GGO7CV5WxHCFpwJ9AwSWTQL3HpC8vgKxSO
Q3WbTmMywBIzcH6VGI9Vh22nH8nxLhgGkBddZU3iJYB38i/qZtyEjLkkvcGUc307CB/dSCnFRkKM
9Qo04lRAdSEZQV4yrQLDifLCDmos9qwgP0IX3hSuAAhStR+OPSxMx0Zk/VGC6B1lrW28PQeS4RYf
WgHK/Br9pu1LlMfOHAt1Uim62pufV9EaE6LVCxDDcGYTRs4Q/4CkNAt6ndCtTvp3eci1jDAsORsr
f+31WXi7Kq6QXca8v2Xy/KWSVN8pINZAUsDjDIF8I5ne+TotGIuy+I1EFjREjzS7MhvHrdKJ6k1b
iiX987oqoWc7YRHCxcmmXtAZI0x+9Bc3S/2aIukifCzZ2Bzr6HPxU5E+ued9BoW8r66nV2C48lZk
rXAIOLFlvyTSMxNAW6sE8zlVJ7g2hapXhz6K51xINBDOKD3YITurYVcZ6dEkDYcxqcTJwUc6ep7d
d53j3Ud3yp6arPftk4f2185Ft4Xes0ddRnpAy2GL4lglWTd0n6z0gMY89WUnDpbgNF7ov72qgSdQ
wYZcTJpL3xdfdcQF0b/z7cU3PbvMGUosvNODAmCPF+XAPdI7Uf4YZ9sEuASj7RiK2LKupkfV5Es1
ApBb+ApV4XLN1Ta5l21MkBIY/2FJEW4RPUdb4yYfaR8u/d/odSQWy1M2j6s5VA+E+oun0tbcYc2F
D/cTEhV8x0BDvfTqLz2DTJIuTPdseAdC1My9hN9Ly8cQpd1YhPA5QrYs+0qokeWQWZVr276Hoj+0
zRFE1Ee5BFNWvrorIlSngPucU+Uc/DxyURqVHMXlO3r20bJs9joTwjxfHzs7vYAJRRH09UWw32Vo
w6HiotL38VJ1ybOAlk5j7dyW82b1Ya02XWAJUWzl+HvdWXcJ3PKVcSBiRMospAF96asKDb8Jv5fT
iI7baOpPipyqfyhzHLLsdEVjfNkLls+s7zcKC0GEPlo2V8VxSDTZ3dQyh+eeM7nsg+JJvDMXeJGy
ZyKZs6jJT99zytlHMAYkKk+5morAOX79CWd45A62oBZSjuLNd06Bb47lve6pCifAyu33j5EbXjxU
x5nC23kyF0ERTRlW9oNipls9ONNhRF9Ul87IEb9dvcmNecG2rVCSp4bT7+tQkZDn2VZ3SqbPNEpI
INECKG02ZGkYiwztvPVj/TPuNXsVt2qtdtuXrGc3WVfG7gCSxRgbUlJaTgUpIr8ISyJhVyn9FP71
h7DA21/jNHbAPElKGc/1hiYPrfGFCSWMeU+t34sIZCZTPQTe0wenHTny6+dBXiW/gnDBoUQJsH7s
pm4n73X3oEP/Lpb7h7zvfOHYf4pSthL54nRZTKB2dkUVuI7SQV+XD+1SlJOpl0rOfRI8N9Sdhpg6
/ohGdEWDmP6lhAODWKCuv1FeagSEufPzZ1tB0ih64R7bt5DzJhf1VDOv4QX8RaR6XWzae5E7SaVg
DMvUNQxVH9IM6lc5cCMGzeD7uLM0bmGOn2r8PzA77PSEaGFwNmkQ3oEIpildbkTSoFvvJZLOCeiD
QcpnKeht+56eiDocp4DR61qUHl/LxJRNExx2b/QbTGnxcj3lAT/VsxVaIQkcV8m2jWQ2vF7wmWPH
NN+QqlLDxW+vktfgFb+g7WmQofR64ny1hp4seCuGm6ViGWRT0HjDz1erAS9hxyT2LxrjdGVlcriC
ZW2/nShzQvu+CdQCRxnEggVj+ad70rPQylIV/sq9V6M/2LtS3RkDSYhRPIAskayaEsKwqCnDdlP2
K/7t28gdLPhP2SEKXotxqWfIjAhkgXLmSvo2rEwVi0wEzvsn3QbVYfZ+fSe+4ZHfQn3P7MxwS6hH
mddUp0Z1+r1Z6yqFXua5JpZiJc/GpZJifXm62Sg2RWGTyxAXJh2b5wdNuc0G0JdrWynfZywIIuuf
Y53gHks3PdhJcJnuAUj1JE/z1rNZ4wvIwNDVZWzvIO6B9Zt+LALVh3rux92TNyi7DBs0vF/j4MFm
93ZpPVdCLEurXX0EkVcpGFDIf5Z4+U9boPMLN2+rNLdimSWabrV8lGgzTQ0GiwgItj5MjfQqRg1v
/K82SuH8/T+wQ4kJnd5ILp7u5WryBrItRUThj+RsG9cv+DUMBeguq8MKcPZCy5eU8lP+XuJjV7kP
ClHbrehlcqZcPwTjYA6X5xI+fVVxRs+wMFLg3IAgZbmk7zTjFMcNjjIzuB9YUPh7Hl6VGLqUOND+
eJEZ4n3qnMb/Z45/H2eJ/HzuTTDOKkIb0jmOGEX+ZihLck9TOdW0A5bG+uxowZV5PYsXM1qkz8ba
xdOX8JBNOTXfUytYfrvU8YXCcNqumTatQY/alZgAkicxYZOllMaimwOfY+3A2EaEdhzB7UTcO6E8
houEUrCbYjRiV9sjzfykJIceyLIVGP+zHu1dAv6y+6c6NtpnAu/e5PJRQKRCox28uwLuKg7Xh6kg
L2+4YR2+gknu8c6Vckx52dDICGkdkkfMyZBgiAyUBH2jA9xKVl8aOewzChJ6c5ZVmviIFTsZWJBE
l/5+ZmRrNfPOF+1h/GbwrC9p7c8eO7wypxy6tCMWco8xwZRhjfUsGXJmO35ELCpj3oVYQATQZECK
5JNv0utnWAXdEKE2wbCRLrXeyZ6fSLpaPvIS555e+UIvTBii9xr1Hn/VyQul0HKqlwjgQmIsyLBO
ZuOz/Fci5jzuHPSf6k21VkeYmQ5zm04qvjzMHOtstaKkk7rnHsuduu4chBZD7XEjOcKj27t6Cf5m
nT8+UYdnQVAzFTYQUGcGbvugciHF5MkE0laV1kcgfQKqDGWKPsKcDoI3C8GOzfDDVrFvVmfZ2Z+R
pCXT/XkDKlVwSstgfAZcDE6ledHSi46y96DhFCesuKQs+l2MfKurCHdE3Prq75Gez8v7XRdSM10p
nMTy8pzNRCMT3suxU3EMjD0HfeQIwrU7KbnYICPdOvMvCTF04KKi5FZo7EOvibHIZYqNV5bH27l5
V3TXwv0fPGOhkxHGH5BRqaDA/N2LvrffH/t86T+cjdeFsif24I8NEUnK2d/N4Az/t8UHZhXTl6Vt
aToqGTgHl05uBiqszwy0+Me1ZL8/1IYcZl+AN3jIOZtNL4bmQ+zHV+7vTiG8CaMWYETmW8zs6+gj
Oee4YEbT9uzmd/s8eH1O4+h15hogxcVFhGsuQWLrJm95btzVvuezoXYM/i2XOO7OU9eP5rKf6QNo
cy0NsfLs+v5khiYvH8tXoLxOr55i9j6/9uUXCLVvjEsvwCWuKJeEgA44NnhHV9D1L2ZJijrUdvI2
C7u7nAMDJ5VNEMpWCfdBcv+fSLy+KPJsDvB0Lhz02PYhW+JZlcUyqe2FjhOHKbVlipnZrET6XOPn
WaXe10GCc22vUOXn9Q3lPBPx5acaFpiQFoAemL872qhXx158qGahf0elr5codnuZ4n5OWEa93ZWJ
rUdm8yGjXQ4wHy2+WasZ1jSplP+rODg7OZoPOCEdf2e5WxIhzr267aGEWjy9rTY+eclu6kImxrCW
+5UKdN6zyxEMvgimyy/c7mu8Jh/FdQwgyBOwBuiIP314dbzxhq7y89/i25bOdWUrn60l48n3uZB3
E71AXhHxfrn/iFo8K+q4QET90W5IyqTCZWaFodh6HpPjD5qePMULmYXIE9nNVConNkLn/aTVwxN5
JHS/SRkxQN4DMPyFy/bVrqM9o0ZA3q40bOSj6Q7iuvVUXuKkuPLDGZJHd94fSuiaKbKzzhHDfrIk
cieMYiSLMsuOYInAbh1wtcGvLs3Tl0Sv6imNH/Ic+g8j52JJrAlwOjtychIlhgGNKPkSPBnfLHx+
6ewhFnNeYvg33cim2a9ylY4Yk5Y8hgyRzdnckYqx0/o79VvLrlLg2j5tXFg96sA1brlTVGvMYSz7
WaTQobTpd65Q9CaM5QxDRKu0KY/C5LfQQ8khQfj9F1nRlpx5orxqJeTdoMZz6S2OgiuFVcH1Bop3
d5nP5zSzKb+CUwuIXFwKHiknQBjAHCkzclVl5lUdGhOrAYyCMMpvWBH2JlR24I2iF8xEYu/ZODkU
PgPGdI3Gv37igQ4D3gg/wtda8TLsIMpAgrjgBhIuL4CC76wJ7JnA4x6LXhi2tQ5Hb6aCp+wpmI0E
22CATDKlLmZYjN+sCxCTUj9BV9KTBm7FtRpSbtKYKapmKem5ke/q2NPkFYifUVxea5u2QJItSdRi
6PEyJgTAfSavDOO67er47hRzopRSLWiUjSluavLXA433oip7Fk4GjPNJKpUMUIiJQpEtx4Ij2Lqm
IKC+Y3ZJ4hm4UKp87lyxR7MlaV3vyeOhhJvxYzRmNLefN0bOndznKTM2JhPy0oH4YT0YtMa6lIYl
2k8Nm9xxQ0UUszp1EftcZbFy34pdVXlN+9zDRoAzQ4zMtdiszhjuYiMSSQDZJ1+F0cqDtpfSxiMU
Wn8GT1Lyg98Lb76thHsmE823ZCAZ2E6NHOpRisrjPi5VX/v2zJQ8RYnBVfsSEwWPHvFtJA7IIEBW
mzGh4UzHgqq2xJO4tdDM9lo2o+CzC1U8hik6WD5D2D49dCatZLE7dW8Xg/B/R14SpX9eBY25gvo8
G7fq6uljFHGt9TfP/ZACO0K6qKIFXK/2aSC4rm/aGVzyMLgT7pmtZpQZF6nBRjv27PDRMUwidx5f
vW1M1TnLR9Cy6a6l1/gcnaS6uzWu3yzobDBPpgUya2Znf81adT6Qr0/YhvvnWwaNFM5Iioai8gW7
TqKOEa3JAiVg2CByF5dqgpjTq0qIEqxph6EiIhpg4UFiCZZ+hIxoxV275izK7ILEI+4GnfubJLFP
FsPbXa2DhmgOC6qEDQfq0/YJ5Y7Y/u+1HepZArzDGRGyeWmPQTih52705nBMcUncbY0GBbYha+l+
WLYDpe8LAdOWAKu+d4FsEX6YqKzY011n2Y4P0+/6hvuyqvM5esop7iaG01ZxqMrHPYxk1LzEbrIW
L8eC5L4q34mWLIsoItGuZtxcY1vNOLZeTdnfcxURAkCrB98Zd1QsjUlS5rRII25Q8jvc4EJ+fVf4
wqSFg3kb5OKZYwj3D+LgRwZnk0oh+1+Jwqg8sLmAp2gXftC+UVKIBv1g8iHPSRlvcmy/qO7ex0vf
gDuJagND7T1VyxGRNoI+ENM3mvhRpsWp/E5NX3hhwbvihgbKzce+T97VLlaw1mxV11dn203ljN3/
TXoIkYuEhGsnARtsCQEG8c0ThSk49ic7U8DR0KP/cVKulUNmYQQJmWRq90A0bAJnEiYlwFS2vfXz
bT//O50E6iklKRGPg7IhMB+v7BO38+6DeupHJ60URhLuxDimlLiMVfskrAhdhwFIsBA6Fe+dLs/e
4Rl9j9g9lhmjojORWXGA7XzuecH79c73k0uzb2pCIeKm2owKZSC/M/w3XM3WRBuJCqd56zcRf+ID
tAsozdNvTZ2Ib/YKc6Mr1mqj2lkx65HLROmEdKc1WlMp6wxGoZObycXhOazkA+53HUL9glsOqFii
7fuN/pLV7g9nQ8hYlOfUE1qarwiJyWA2J40++ai1+KjUijcaXSEmmh28OEPba8fVw4WZEqnyzDRW
M3VxYAIoIZZVBJLPjoEVC1kpSE1NjWpIf8B+SFgbEDvthN5M4AiHYn49W7/MspEff9fwOve+IcOr
Y1zcZyC3fGYYbFX4HyM/vpDZ/pWEZ9x7d0PfI6OoQGEaj5HaGSX9IPzxl60n/eF60AvL7RIRzaq3
qP6ySK6R3XOuf/5eRguImUux0xQpBmDHFO/6CYQ/g4kSuKct034uRIBJSRKuxovyV07y5veqz5zY
BpRlXdCC5uese0OpgWjAm5U67QtMeLiGEhzHsPV1K0evp6YyVO5t+mVtFbmSftmA+bEcyIIMp+wB
wIR1sk7uL7FSGdSKbQgrxvp0ihIRhHr+7Nr5wJfHHNWSbApamw5jN9QLZicoVZ4rbwJP/jvRxtzp
pjXD2V6XcMO9vdi03GUtinyQ7t4pMEHFsQIJxRymjX4f/DMAwQFOcKaYJDOW7FHxYwryHzpccPX6
RnkbY0a1osU0C+bwN+YjyrvmEiJXSCbcnTegBD5XKiRz2vLFBZzcdy/EuOp9UJ8hm8WJRZq3q6MK
gagPBb8WiwP42APA5sqSmcbqQRDlY4eO6UmxPYBx1S5bu+ROc2mEeXZYLnpemDtfs33u7bBkSb8s
6YaXk1Wf2tAnwbeDmsuKQLBSwqYJV2NMDF6gSqcVrEXUcjCUrUZjJCJv/CguNwhrWVInxmIxH0VD
1aiN2wMFZBlvNbKo+nXZWxyyC5kp2qeM6h+lAwwrV4fvYIHMspHItH3ygjK1K7KPWeRQCP1aKLM7
wVv0eL6TX9HOL2Bhrs5E5E1HjAdqEwudJqbF6Pi+K3OS05bt3pWdlSZRGG7Fni6pT+DInmihQJMw
liy4xwksdiOUe7y97XMDhNJuHPodrStKD1jxAaatgwGtrlLql8nlvByi0SQ5ckamuQHOO1AVEx32
aoHtlxM2YZv2NnCXMqj0tk0WOVI74pVZZoJCF3Qm8DgVQgjrRJ/J3Qvz7ncAm2hEMZHDdnH3g0KT
x8FQAuBoHVx9rjSW/Vf6coa0qTitv3JttXwsQBOM81cbVcSLOzOL1zw08T6aAcQrv1OJlGaxGpYK
2eu1j4Fpw2hDorMZ+KHNAElsY7G5Mw2iQ9RKuOWLHRFn8I7L7wja9MIYfnMusRUp8yj6wjYZtV2P
qKIYaRzskwwLMLQfVhMZoP9+j3pgTRUTZTxbIpq5vIKyfcq8Sah5upylBvqywENKAstTwgNTYIv6
qbaRK4KLOVmlBO68KS+hLw2RUVArx/1FKOGMLi06+e55+yCXXMsi8wfAw6xAOEIrl9wPC9dkiojd
u49E1sSlIsDi4q8uFNVWBtC3FMrK5cExkHjN6sPaSftdfYcvqaPX0MysjeQuQi4KEZxDWF/rfDD0
GAcOjtddKPutyGrx8BdlHaycb2pWwkemtqn7Ehb4fncOGJwSSw/tYjcNlS/5+tHSAFTcVHGtRW/s
MD1EQe1IbCn/J/jdAmGsmEd6pqWtZTH6JYMH+YZr8GkTOb9v+QOEPAxyhxf5bEVXwVutZa0KVjPZ
ntP2T/bipZY9cdb8X5WJVvTywq4hEGm8UH1jFA1LXvR8tP5Ose6yNYzh04/a+idKwN/jNTP3eBZ1
7EbJm9XQ9UYOzNiQoH+AJ0mukgydvp0CtkaMpEy/7rKI7Toz+hW1GBg5s3OZmTpxs8fMMO1KMkvq
t61dmww+LCuySlzJxtUFuwzHMQbi93wJJUtW045MGWp56vZDm2PFueqxKV+5xMV8V7hCPNQZFwy5
U94orGk2t4QYH5t4BUvm9wjO0vAOCzFUwlY+c1M/ygnbgptncwAp8kHltj31eIbBo1NF2t2aWB+z
SmncYF8GScrqpEEoNgMm6DFOktYOfWy6zf8lb2HDq6A/VrZWQD/0iySgcTA0HE4e9OdvXitj/Dde
aRocThToYElJyBfi87qtr61l2wKLswVZXXQG5nTv5Xo2EgIEH/Bgv04EUrLwqZdczcS/YnDQyLCX
TdrcIs/6h1WLsYlXHA1GytzHlJuXwAFQsDS4HqiupGa8cR2PSEsItwT4ZmyHrjGlZF/5DgR4uwtR
3XMs7osmSqmwAfAWAFzvYgsUKDwukZsBG3vkFHkGSNLB2yEhlQvqTXcJHEzBgAe8ncqF8j6Sse6o
3kw2qkh4uKsdnIiYAspIcy4gdtikiXA/t0Jp/bvYo/9e+1grc0bBDZ5UDcUOZUywJ5aWdp3i8NQG
kImzjbVnoYfnWfC2iQmNxaZ7OXhIPdSn76DX5PHEG96FR3BGCaQqAwKmovco878Evl0tzSKPW8Bo
0aR/bh1ufvZuBGWO5hRF10Fu2apFjFkTV5hR8WSngvEpA9cC4F+z6mPVJASusW8/AdWNE2xQ1jPi
ObPDI1cC/sQWgeGIwbi0lEliLjwtExvrBYNKxqmoNe1ONHvmHEe0xDj7PkNgQl6FJUOL2gHvo9ga
NtF/j8B6Wh1dtreRTg2uJjqx16nH7BkeV7Gt31Fgfq8gSttmf6ULmw0s0LhO1MZolVoAm0ntdNld
Zb0UCVaWqb+4i+fR3NJKl4b1sh+6ag+wNYgQVtuUJ2M27c6F9Y5ytPntgLmK/zWXzHX9m90TBoqW
0LPGvGde4crOX3zP6F4+d9xMHPjVYHhg+V9yPYx1qPRx1ytfJplUrUci5ACI4GiF7ak0lUy/HwRf
cPEcw02Vx/7Wf0IKV9t++NYXVfBMEdU4U9TX+/ZxdIqrOkTZrt5vmx45/ypHscMReE5609/8UbfM
pesRmWsoi6bps0MQpVYMDAj/CAH7yfQ1tzE3k2UXcs53cuCQrMOtfOiVafzzs4X9RVyt1YTvsyhJ
dlT3ZsIroYayJtBxxuWlTyPD+Jw/YcJLmsT8Bi3gjWm8MOzGVQ2IoCJFZZ4LHcSlmfDyO9fjYf2S
VPPBcAqX0NxhYd+fQvI/XluOdRo6WqVLcDRNalnj7O+8LHIormrREpv/O8iJtDlZlHNUYa85oCRJ
DyIF381E5ghWMVQrmHeGRCSkIFE0Vihfu3Yzm7F+Xj0aCGxPixgoGBOQcN+vBfOuP9Dmo63rwjsR
ioyS+TCJZwsRPE4Qkia99WBBHn7y8U37BfW0be/SK3kqYO+afZ9P1EJqP/HFFqv53XkUStQRygIC
zYxYApkgQM+WkFhrwtpgf2f1GFOPITa4Y7HvK7ukwtJCiKPBxgyxj7aiatX5OXt7Mg4Z3EhIIoEW
uaopM0L2gRmozUfEKP5Ac9Tj7xhepqEBr1NJBMbb11jaxD+7r4CbXQNWLGdjwUyOXFIVg1ZRS5ie
hlSiB7Wi2c5fMKFg09oDAiyobD92KNtfBqIuPhVb5dVIVO9JhWomf8yM3YSgapg3Nw6izuF9PIOA
64sQ4+bkXoLRc7NeiVrY3BtOtGxYe1v3utyRE7Y2hQ+ePI0VZlCp/uNWi5aCQijPe44ETq+OQV/Z
02o3o0zHzyWbOk9MksHXc49EFe5Iv14GqcBTMbPlzBArpzgLgPYap1Tp5wDO1xhbT+7cDmlfzcdf
UZZ67+k9pNcqNtJmd+QjT/z9V9ZF7hN3bq9z4lHkBiIzj7EIsDul8j6uQq/nAMfjLBKDVAoxUnB+
gsM8yBbaUiMazua6PgjGYPwVY6cow5givRHCW1iSbe4OeTSZ66QlxpSZLFw5nheTrm0cud5jkdlZ
Urg8QjGUXDV0wjeuMeLTNIaT9qfv0BPvofUq4UJDrYIN9ZNWq0/YNGaVP9Oo9hGs+HmW9ldHgwB3
7wiBRa0JE0EMrPtIARnmiZPzLoFediEmMtnjsU6Ydn48mIF/5ieY3hC3mdljrwvSR9TuqvEaOxQX
icKoBn9jX3G6c7p79iCeR8HwV46FZvSkoFtrvohGHyEjCnaYmxxWvBWXueZUaURxA0v+4umRXl4w
bl9zynZc59wvM2dBlVIyIsOfSLSnGI5QdDTwTKn8+iITEcAU1AcRi004BYgbGB2z8f2DOXJQHAnD
yU3zIFEpw0yXjIHcwp8sHBORCdozpLKFjeJ/bEz8tmQLN3UAWOgQIiA+I+II5WHfR7Gu8tEcjYXZ
qU4E7QvXwoBDeRyLmidQaJKiRtMDIE+fKiKLSJYHd6Y81ddhObesairiK8oGnXSDukC+utWqpy7k
nnWpkkBQSEkpyE3kYZkmcJZoyGkOqT574PtmRRLSBl4o9kSQ8Ybltnef/kcUi6blakaHAbpxbKSA
DCk9t5eU1+IiEg9sb2PIltxDVWS2R/1K2UkI0PSEnHZPQFfKOz2OKAF7GHqQRfFbxEgds4L/xKA3
K4k2Zl9ClX7nWglg2sFK6702kdatuwmQkoCtqP0pILoorOQBvQG9yJm4tDrkfLnZVobrS43s+XSm
JF2k7O/gkQI/2ev30ImYbYwjrg48ILEbu4Cgi8F/F/XmzNVNIkbcuX6zmDmXwZ2KM2q+x+o6f/dJ
fODDGH41tMeAJWi5NgXCbanq5zyCx2Cy+gtmA90N+3poqjaTt3Y/h6SiyQoT1YUmLwJsiHB2tMZK
YhdC7dQ1yjxBYCA4CtjSWriDJr2Kr3Ac9HL19mtmFT1zUhdVnCwIM+79P96rtNg0JOwmhrX4+vxr
SN08W+QoCypTpR80ogibNFKLMqoaxDc+XRUpJwpMQ0TNCOaiY+bcQ0FzmgOfb58zbGgfeG01vCI+
A1ui0XO+d7c3Vdm8VrrUa28Sbi+zpu5G927XEY4BFEpg2TI57Y8yVMXrD2s6w/5t4fjBkV8zwx14
k+jEDROFZQd8k6kVIXo6HjQdVbtL4hHPXXklgYppZ9b5vUKX6hvukq7QBY/TXW80Ehrd3lwkXbDF
lDt7w26W6IE86/+hepa/l9VOc1xtnBz2xuQLUPBmb7OvL6KGpcLJrI7Id95OO3Fk5ilB5aL28VkL
HS06+v3Rqgn4u6SX20iFh1KpXecWa9W6izlx7jHd9x3xXwsPPJYXE0SnlAllA/03Zyc8UF3d6CEu
7OH+L3uLpJM7n8aXVhYGrcxJPKC1WKKgcszHIDAp4PpeJTmZszhohU66/fvpzQZAQlTQW0wJNvpT
EqgXEP95tZSiQjJOx6PsYXJDlUWV+fm9qt3XeBLcCrF6rn3FvV9C5WfeXYpu2pcovzyVKbZgnkqf
Sn3Pa1+4czmMjVvRT3RDslCIOpj2bAZFI/TIbp1SML3kr+eukYOOWvW884JjP4Ha5Zk6habmnry+
GfH9rHG/J6Y9IPYug3bXNvsiz0BlI41SCj6uwBeZqeW8NATTkb39zb7fxmcPU4s1km1QzP37Eiq3
O2558j8dpXbu69YzP/ctSpl7PUAZfs2ip9vxjTEj7PhXP0yLXdK+c2sO5og7I9oReadKflskrpR4
oisfvFZbl12bGRiFPT/8sBOtjASOlZeYbdjV/ukbgDzZjgO/0OrURHYnwU5Hs/39oRY2eq/UodBt
hn5GHLJVF7q/kbEmolxpHTVapf1g9GmZHyRCOMAXVmnpbXOnBCVb4SjPka3jyzYzit81jVgJYsu9
AjjsfeiBVhvAU9Lth0whDY/2/Ui76aC68GqwiLXOhqB/mLDYnScW918XXApkLfXiy9h8llPWh0NA
4eqBGKwyHYJvJZXcona8qArj8bWqTKghkXYAmsBgGu9aKNG4GteXcxlBwCwwdez53RsXv0ux3KhO
ZlfmUWf6pa2PEop8wKjXYyzpooL0i2MbfMeNRUxv9iosnQuw5Cxzty4tGovQWkKXzyMxEXNlAQjA
5pN4eZ1Y1Wab8FBKCUGF5WO3ySrSmjaskbiWmFa8uQ1NVNbeLR9xsf08zmikw7IstwEKUdJwpDm+
tfGSMkS1cwOv/lNPEkq8CrfzzHdJfPtalpRZuBQA7jP61KWidYT7+E0yrNW3+N9bEPU30uODcRnR
GUe0S3vQASXkp5J5aBh1Fbhps1vwN31AJrzqDwsXgLGZfuO5ynt/sJksZHJuuOZXnxVpgjAnDdmI
15ky7iptEwM6KUmDxGLxNVNEeGORelMe3ydCnzyRqz1iE6wJv8/RJN1ebXa+yaYFiX2pdB9w//OJ
tPtIdQjB/gNqSb3nlKhSt3bZ+MNq/tPTuk9u1YmO5VF2htViRnp7ML6ePx1rlurEWSFQrwpV3Z+x
URGzn4jNRnHezDE9u76eW9wmMXBxWIxuSqwJ+wiy1yrf13LLhAGscAb1yBorFpkh1jEzkfolPwvw
Yw/OjxyLRv0J8W1c4GnYqlc2jp5QoG1QlwmsqxhUx4epyMsabQBRCSI+SDYbua/IbVdptfS1I6GJ
zTOZGrWYVJB2cGyL8cWwMGTIJZxTVH6Aub6Fydge7uyMP7xgkUvWakqklk/795sM5VyB77MZdmUS
VVihkv9tuW5LlIIfLlAieMsucNDaGERDLvIkj9VP0KGgGRnX89q1VeGpPxT9p8ReBWcnfph1x6g4
VF4vWH9MGlpzTpRJVN8+mYZcJtgG99P1z0AuiD6gvBs8FRKdk1c+sywBH51075UCUG2OAuB64o9H
0YGVmgTd7ACUICRS7mXVSmrjp/igkV7MuaawVpw52e/o9k3Xwb5iar8EfRwEmC8+JKS+1d5lqAhv
Hyh+/FQdwvr/vvPLJC6OB34MQk4DtnbTG2izlTSnjgpJGFjVH29RxmnMHkNM4q+nV4AJTn1hbXp8
/E+pDjJW3oPKoMSv7iLOmt8aAnxcy8rVpUr5w6mq427mV0SDfzBGXseQdfEQ4Znc8OW+yzRTsoVI
SEfZ8VU1QDjoWhrVFXz/+olb8Sh3jHWaHowodrTlFa4Nejg5kCJBAo1NqGDLQR+DAcy4Fgo4OjZZ
ePFQ2br8TMHPQIZsRoPrpkGpNyifDwq2+xtFvxoJaLEFfdCRKDpkdcOTcZpa4O+pBMT8OvDwe+ki
F8W8AU4emOu77z/07TRERRNF+S5ZsFivXs6wh08cu22h0dhj1xqD6Dns7qWIubZv6IDoPvYhTvrV
ldn2PEtRLCLD8NsUcbIacs02KLMekbFccHVHA13IdbjeT5p0GHXcH4EO3G/YinkcHyLWQiWLPQi9
bW7NChZzfPHWWwuYD3wbZ3xlP4KJudTlz10Nvs7rWOPCj/5Rt1oIQ11+vXm5xSSxllXCxb3clv4S
QHASCK9NPT5GpFeRMyXoFasWUcUpi/zxmFxvpZLNfS3/QfjwMGte/Xbgv42e+UY2yoymAm9L4CC+
mPhBViCbptIKkDc4gPofPoPLYqGGEX8YgmtWa43+lkPjNFA2HHPWUJR/TZWoCabDaxbFlfve7GGq
6o94EvRS/M3N0duka4oRk8ecBGSEcBQYb1EMrAz2xchqclibAoE1U9fyHpvzipJV7ghSBxobGYah
XwR8r2hh9/yx1KL++tGsMhJZgPSGa9jXTaASuaQ17ZN0IX3JdWDrcxt9hKDD+raveTzGI5HXL6Dy
iTg+WSxcA0JcijHfUtZFcHADD0gU532ZvpvBs8cNug/j4mg7Yg0u7P/2YeifCLElY9B4BZsNxb3H
6okEnnzO6b8k+I0XfqgHSCJPTZA8kPV4CTv1GT3eyTlF4VoVaEIXAiMmUYVWUNSnOdYu1L64K2ao
RsOnhHWbAEb9i1ADeV16ywwMv4zhh42ZnD+5vfd/uB74cTFyq1jdvdkdLjFnmyZXxkYjwUhMkmns
erNeB+7voe3ipVUHC5vmUp/txGf9+s/dGGRz9eM78a3267nif629OFp3NlOzc8aRD4KKwQ527yFa
XZlsMeb943xxVH16tzxsITe1TGF6V84ryxroZ9PtxRj8neE0yoIYAHqWdsBAJbNlLPcoOCZ2OVVQ
PsTDsxJ0pTLR2xTY+XHYkKLsGLm3pKH0LrbNtPLPtbiY+uSTiI/F66ygVcyjsGRwMj5fDi5IXxCl
PRGLuOUtchBRGaVuJZL1McX2iMLRJvB1iQqybaS+2cZpCdxaMY5SuUcJ2e9qDJJ6gdAjUaL6b0fi
rXLcce0oaHE0/eIAr19G+QYXub9qz8mNa2oxN7cPO+QB72O4xFq86AfPp9Zj6HUd2SVQxHNRYUQC
UBN+QyMcFpPOcfGZU0ScobR8dK5eGAG1EtOkG5TSYdpShBotbX3tOj7qSAorN8egeQGzkfFZuNmh
wScaNvljLBHyrocu91b1qVNrilGxUbVKK5wRncBUJYEIh4lVose2Ptg3LV6biO8krG9uGdH4LF2T
I24SUpS1L0+bOpUo2iYkcUW0zTRnhI5nEpOJwOd9a/6kcUWnTilGtL9vrk+0IluyLG2L0NleFNjo
YwgzSE8vyhltMeiTaVQKbuKgw5f4BylpjXpVoW0CLi41qVPrTYIYm3FYqLDyaORctzt7a+zTXeOi
RbpNqEkJ88qBEqOQtg3WsZV3lv45XxWIZge75MAIWAdreZTULozAJ8mGxhcmpqT5y/aVleLkll29
U7TqdBs1VlRKEPJhFspwbvVzlr7w4C49MRdbZE8FJIdUkGnrQSNnIoFW6YTytOnxx7DC1RFqppRd
juLsP+1VQhsClQZJq7ST7az32B4sx2Ht/mglOxjB9UQYrbYJPQf5JLRiRQkhBpHyANgxCqaAeCCW
3ZnappwINzaxDZCzRNtJQiSQkdYHabcTK4nUtsZln+V5pUBShqqD866ujH3XSV97s7eDXxcypD9Z
VNB+vEWQXVetmyP6P/T4yvWe68UvJVphM8EoknFq0P75p2AfYlR65olh1HitZKWiXb/o40/VPjCP
eBb72gx/U9kWzZ0jeWGZf9ZHU6s6+NzpZxL+2Fv2n3X99iXRwPeGfsFkKsgVuH6NgWT6lHdKBDkU
G4Mbc6HQXe7F3GBNsNOsosCwkzdlo1c9CZdnLjoXISmthAta9KQbM1b+rcV1KEgZMJiA9mkMCeMu
NB2cdjRvf90X1cSh40E+mil+y3b5+zPvhyXnStMX6UOnJyEU9MmexiHRk42OSbpqr3O+eONgzm0p
OQdZkambWqQ5Pc/MuxTQOYMvSmGK/IN9oHU7IvaPbG/YcwaXhSXERSRgqMzHU7DF4zkwQC5VLYDO
tOXmRQ21UJSZBxVEYhGGOw6HSgYzdbevdXU9UUhay5FhFN0oNQOvdTVaZQygKXPWmGVqoDswnwgW
BOxuL+4PvbfClteGeTC+vuWyKH2IW0ZNQaqvQYYPWZWWQ0P+EegGoVZ/Nq+YW4c3uUVLel94O5GQ
yp449xWzFV+MVG/whHAZSrt0tu8sDPNVvXXOMSLqP0HC0J2Vpod/i0NDnNmkOlG2zWO9OxWhaXjG
fIDihPV31HWiHfPulEEqyOrVq/F1mQDrCfCAbKaFtjKcGHDhOCzS9bqTfP5rM4em0Ve0K9Bzzu8I
gzKlbRu+u/25GEKU38ypR5IDl6ad0TxlsSV+FkvhfMIpw77Fbp0zpSc7huhgKnNgIoibUXrqeE3Z
hHqB+hzUvL70STK7avQoX51U3cCEKAecSpl93Jx3n2dsY5ghB+jhHwS71JweWlMcwx8oVhN5OGJS
wegm1FqQsO+GBI+gneV+riKMj65x3kvd0xlUYqHzhPynB14aVfOjLOw2GbMsJrAKnwNu4oZAinOW
P62MOjVwQG98/WgqmDxxAtkwyv/TPI0ZzoZ0VwGtDPsdTe+jM+Nda3WA/KBF8vIhKJMcq7rIOz2m
RXV8nBU2igj9op2vqPum7zqM4q6d7KNoqKwqo9SCWqzUxQ6fYSsQTaGhaJc74R8oC5Hv/Z90u/sI
jMd+THicDM/XimMiD/LXI34jfCBnMt+rBotwYQVWawYGOL8v+p58dOex3ZyBLyJq9xphmdkTDYcu
izf/9+U0+wwQeyh7hipIFLJ9B1S2DrsaSMmf7y6xYaBWgMYASeFA+038UyNkntpv4cdqG6ULajS5
PfcTl1ppBScnxLYvwqfk2ATkOOlDax4vksI4YHXInqS3ba7mJvld6LJsUg9E5aF197/V1LOyyXpr
QdiQmBTc6ls92/HcvBBDRkgfQif/FaTpQyT5+7NxEoJVry6UTFt69h6SnoWBbQUMvClBADsKoRbT
qw/c+vXGyqUTt3jOpMTkDPzVaeoEZBEQ3Ge28GFgkrvQRiqDajyVNx21xC+ii/V9AZboXIGZ6ct3
rTK/Wn9nyo8il/aESkMqpyusJwPh5C2DQxOz8scpKL2h6jx5a8nhAZeijebUJpcugSCx8T9nrLz2
SSw9NFv2j8B8ggGjzJYtCbpoeI+bPJ0m2UtCZ23XAQ8K03hAFP9Btas3+MZ8QzKZZg0BKXJIKRgo
3EvwqaH3ssM2R9wST7n1gD1/u4eI50+gy3YRweXDtg7bq1PJOJku9apvJcajnjqrUUbv6lI/wn57
eKVV7vsXgDYfS4FO5/O7dl3mLxhzWnk5v6Bpgax+YUEZdPc7U8vtrvl3MRuvx3IP7lf4R1prX0Wj
XZ9TSeIlVZjtHZ92+RQSjzO7gcdoY/lHqNmrOAZwjkjmcknd+E+mvA8NO+FPIGp3Dkc3HJ4dZPfO
OmUFodMRfjX5Q+LXNIWcCD3YeLNfVTlq1ZNC8RNPTL8a3xaJa2anTMtcY+sTnOG5dgbI98jEX4JT
y83l3CzgBGKofLSL91jqkjgck5Nj1G2d9K4UGooM6WG3duarjq9VXYsSOqJTuVmlKw8feqoQTdq3
7c21c4K/79UFOzWPql2z2zTtOurJQh6H21+nL1i3U3eGCFGHSegART/m2YG6MUMMKQa/XYCOtz53
PjZWSxWTw8LaQHp6/c5owMwwMLg+1/2/1a51Mmzrt1suwDUjLAHhipTaEym1pppdM7H9AOvsTe8m
wCaLS9KBrJaHbQQqJVKSBSA1bKJt0ukkCyG6wNVhd6NjxD3uOcZmB0fOE8/YlPMMRHXnZT6CPqdU
/gmCSFDJXRqfnv753R/nx+uKrEXMwi4OB2UTugcj19FJGQZwyZmWSzpeaZgRsaOLmc3zSwFr5wV9
zfGGPe9DSxwdv7IAdRbYegHVN/3V4V1Nwm/0fN3sxpWSxQJ8wv/WxirEx5YCQq7gUxpq3E5HS4+o
u6umqURBXPGN94VjEcTIyuIx9eJnlfX+l6RjJQ+fmpVDW5sh60LgNXyMsz/xWriWYroF0hbYPsJY
jKaH2qwR5VGcPd+HvIyQG0/Q3jIJDahRDG+s3j2GI8Cu3qHQM/z0p63L8SjGADDZ7J8QPlmIHCHy
R+G1wbgSSJ9i+2EEEPeB/o0VFdcqw8dF07clVolk5NWFgO9JVzX3rAqsur+KdKKEWJFCfdylhUZN
xe05IY9orDTCvdZ0D9gbrU0g3zozEfvyC7ZJes89TkbkCTaiSNWtYCUgEkGGD7O+kRSTYUDnaQMd
c4z8pPXC428c/gfoOQWIMV21SBuzO4klvNFTiL/YHwXlr3+f/I8CF9gDwp4gx299jOyDeJWoXLV8
XWK8Khiau0XKMrJkf9yB0R7W1U+8Q5lkYtV+N7VcURulnu5HkjvlZC42pZMfUmb5HMRQQX+3XMgB
sVJURUPTpNuhoIlFOlKfuZvw4z0KOSIsVnZYdrCnt4BLiPwfCV8gyKYna4JVN7Q8mrywHlAJPYZm
JXVoNH5WKf3JrzTYLZKYzyN0NhN01nOIjvd+UBSz73oVuZaMOq+/1KQS41cKbM56PNGfvRz9XLfb
FIniTtYjeC78eOKzynIXVi5dNVFoCe+uHM18/3Oonm+ixD7sjH2JAxNHLve/ZV7M6QBu0megqTiz
JpcBwty4ocqYHhpPR26tEqvv8KJ43dvS0/MqIK2Hm83j/Zz199/Uiw4f1B9ntznhcmJZxdE/4W5l
fS/J/Bv2mcKVAMS9xrKeW2JPJsvKw5RvzJ/NukrDBLH9pOrwvo1O91A78N3rtNhtYdaHHWgeSK1I
u1Kg+4gWZxgZ/G9Vk9v7WQl+8nFKNPeX1CdoiBu8GpbPW9yrkbkYx6Rbxti1lw8fskYjvVd1XGms
X3aSGrGRzNJuFOAZc+MG84/Mu+7aZM1K+6jNJ/J5ClcH0rxoF4spYk5mZUa9UjdYQbbMM3agFTDi
pxROqvwFT2Rsl+9BkcBhncqcolvpK0PRJj/Zhz+wwe+pSlFv8o/0fQ8sn96L3LG3D1LYTjWB564+
Y3e4QddhOfuU+fzKMnWi00hL0Ol42gLOAXwHVwwrbuT4ZOsg9XBUBkzmbyY90F9DJ5vLnw1cg5Sv
QBtwCRJgRPM5fW/m+a38ZUr2W8uT6A7LZaGLU2gw90RRZTDGfoopCL6g0SYDmbntZlYhVyxlAcEI
r07rPZotLa0eGSRJDtvXJqqM/rZ+mCA1SkObvSWUtpRpfA+l+5yQhfS1kDhrGvPzSZW7z8ZkDNG9
TRQrhuqC9id3IysJSBPJDd29eyZE+qqCYRPk77V+FAI45y8AmsFHl9vaJ45h0kMnI6GOX/wwRX2I
gNzxkAeTOtC4CcYMl295IEK5PkUFaItuNztJI/+dKKGJR/bqUvlAT+W9HkN4TzjdE2/smIHrIPVR
C+4rGHEjn0ZptPfrMJiiEuhFiS/rgSv5Gy2MPLFD7liSr2OjbIpz/RWId6Y3qvdvkJeodxfiZtgj
NhUqRNZtyOyJQ4uNL83ll3ZM4YackR/Tuo32D7YASRvKCq7ljNMkHyVQ58Cmi64ZwbqvyWfcjjao
S22RkYvB3dc65LiQMregHsWMNcMewfUiX2rjuxChT890aCHJ/Z/rVUi5kZl1fLCQMsblrDyJpyjS
jqIw9WyIUrW4mmYX6ZDkFyoO3PN9tgvq+VRxXLa3QZRHiIZiXxM6viGJZZmIdG7ntv9HfYc6TPoO
+LroVZCCi69Fh8LnrmheFVzmYlIKcC0qxS++rZLW/DYu4iOItiy7WuKgC+vYKLufSVMDjV7mPueH
U/t1qNuKDPsm/MU0/LM++9r/CRoJr5AEZRPChrVLE4XogHoJpe8Gq5apqYjVF+6V0z352Od1KJC0
mXx4Bbow73AgBekWxRRsCDi9+z7qnktvl7fepvKq5JUAbDJL6kBH10x6dA5Wa/mpTYpDuSkvr70Y
d5g9Br/CQB1UpyLqLWLkOqBzJ3BpbCpkq9rMUkMXpCurtxJeTkSJCQsNfansxuQQAqUc3FM5ZrBP
Om5PT49iSq81i2/bWtMewRE0KwNxz40jgrZ4gqimX4kMKXkl2ARtjQ/i1+O1jU0EKKZsmlivfdj8
e7dycVvPD2jnWqphgsou/ILzF1I8q+5mLMhKIE10KB49iP+PyLsSJGWOg5OP6waK4if0qYDu9ITj
y1J1AJtdZGfLHQxmRlepNhMxbTv6MYcY8dgxXqtaMm+lyEBSg7PJRpX9W0OIXJbZAAFtFXv8iMBN
eYofoMkzB9bcxY1R6i8YqieZ0nPuLH6+o3gLTWX/zQ17u1ykrT0oCminv1PfGlaynxYO17kebuBs
ZGkoA6R+1qhL4n3UAMmKltkH5FlgxoNjE6DR0cBPcVC4e4gdIeePs4vv6eG8/YUH33Vgx8BkUUDf
pWXfCWM2LOFdKqvPZyjDPTz8b2/Avlf65FfgC4xwPLEYhdJBAheQifOQhkxp+JkJ19qIUN1ok7kN
scK3R2EMcH+GRObQRmzKVJVGPk7xLdWEsNTQQXff+oPckM+s+1CSGGjFnWNy3fiFqBR5JzplXL8S
aGETN/QQbp7mWa4H9FOPlhn0R7GQjxmdUUPexhsQd1WZw1WZ1Pksze9TYsEXRmF5CdF0/JD5rZ+z
bZUdKed2Y1YglZyjxg21enNUV0ZBXpcxCuPrR3PE7WovMk90q6v+CypA4tjsHDdVfUH+uq3UTzwn
COCmRqlhyiFLa42/BfwSJ+v5wTRnmGTSiPaN+muCAntXLY7oFXEXVTCx2LDwgMGwPquPG9PEJCQn
CccgDyLqERt2HME9TqPUFS41GbB4RQy/1lYNvDYxwjdWtGHloho2TWgu3OF2mOVUUdCMbDPQrffy
m+NQZ6mMor2pzVfAsIh/xGIgprNmb1SheimopyNt0Rs4xEuwYDycLEp3JrNUOzBl0FnUSIcNlLo1
16S5RyuGjYVwSrHWK31naRR9wv8wyfU9VvKAt5GNsIVL2NoKjoRwlYGOfTJEFokA9KXBDUruukPx
C3YRMB3NZdmnu26wF6y/rVuRctMnXhaZmGWBi9BlixJXm1lxC659Lg9R4LzRzWbzPG3RZwCuMdF4
jciC+OFhgH7YuY9ZUtP+OQ9ylkyBLH+cTVGrWrB8IzxGj8lZknprSXqSshyrIjPln+LXZ0dbikNe
kFVbxnsCZ3W6VS5ZzEcOXDStfNn7aCwK96LQIzFbTiUznhrDu07tIDgTTF6UuieCZeVeUFgFnug5
DIDN0TD2utGXdPUEyEmUb0tsjHksECoXbfb/Cu3K1GGMChidhwWif+l7s3G0GbnzK8nX6RgO1Caz
7tnmcLHx48cioUZsRxX2THYf8LGtEjd64T745QPl4SlZcKLp/RwCIKoLBeSARf5VBp/g5lKw8Rvf
khZCM5VqwKtTWhKvQdVSHJGzqqD+0wq1irGzvpli5cG58zBHseWSDT/ZhfZBUromBUN7BY5ONVAz
ZJ9v7hsk7S1xwN4bJZ+aNPC+3w9e0ADD91PIrwnDjmQNMLw+8YtQWSFIuLBC8wH700AdWifx0t3W
mpjULXXvxvRfgGLasla5IKvFkrS4b/3hy5aamOGlHrSlqOva6uSLH0s2GlWVgUiZLSqSSL0WVFZv
Xa6Toz09jIWHcpNbToa5jqnRZxM+Wef30+jbSuSAM+oZISfupD8GuBrqWpxR8SRmhQZamm1BLHRG
/DAxoNUGX+ZljXf/3HOQOcICL4ptPYGRRxwGD15/40PttB2UDRRCTZOEXRJ7bsv0YteOA9+hGati
fzHB+ufkXlLIHaQIinNnEAAO0zncq7XU6/wtfTK4KqVeFmQEz69o/PCpbqroHq02jHqCuwy3mtCq
QRf9J2tfAH41XZivJbH/nHmKB+kkzbOOk/tbOldBZgEg+7ar1Xdq4cVI+2Zo39ZpLBIWh2l04vmf
tlpWUArJHHCDHhEt3iA2T1EIQAMIhrX404ZsDC91Vxxbgbc0KCt1jw/qUN/rlkaBgSTcmhPSkwZO
DFFErc5N7h976IRZeOmkTyMHDDgPubU9aKccv6cslmoufSvEp4cERbpbiB8BBUJ2vvjiyiTNBFos
dLeU0bRu9LwGlSomJAasCQgM/ITVUQS0KBLpfD11bH9jRBYGuITdxL0b5XfhbIWFENU6TgiIPblF
7dvq4ZsI5EMg6+ssIxP6J9hK6rpb1fmDL0hnfFqnO148a8N2IVo3l8qBprXWdIqbgTRYdGSeRDz+
hZGsRss1H7XH1au2rcZ2oLMnvkKF9miVrCWpr9aOqYH849MNRPFCpH3ba29GvLRG7M6k7AuUh/Fq
c0Z1uP8KdZ//8az5XWc/O1s6hT8Zmk2GLWUsWaAeVtqUt4vHjrSUr2SHslDjvmvoPoeyN98IIzt6
RkkqnuvfnBdI+S1FNYUd7rJOGV/RKXBOSCM4xlnf42gZjhkJJrQB3WMw8psbqW+uWVW6+Gw2CQhC
OW8neSZGsCcR+/D4wxpUG102qmO731cCGS6WkRwXVpyglDJJXvnrvQjN5Hy25So7xz/j/kq+FKYC
ioZwhMopnNvU2BVJzmTWfA1rRBThhfP+XD8u3+g+GAqqb8P/o6Him3GOUr0O55d4eFBNgSnKCHEN
RWHMM37rrgVHEO8vvkF3KEkVSLPvU5vypqIL1Vm/D7QRVvw7SVROfTNAd+EbEBNFmiyF0K0sU4QV
Qtr3yIGC/1e95XcF2GY4YwBTSm0qxJEThzxgmSdzFCiHEiq/FHFkqy+0kEpKXIamkM8itMkB4pra
7cHiZC/TyfiapH3VX0tKeYr7VB92l+Hq+p9lVMD6n5cRVWIjjrD+F+itqhA8q4XEvhAVLTabzib9
hYFRs69SK2uSOPcNnMK1yXLCTRd2ZTx1XvPEZ6pROIhga037/nUyH0lSRE6Yivzvj88J4KQI+tgI
ZCC5D8F5cnm2YXLhph9qLD7bXMMSJF7emWmy9I9ATgNpEgCrbKLh3Z0fDSMfNXAdTuOnu7u5FeIH
Nxf3ctKdrzhAmbaaWQyZ7OOCI+JnEnvKw4pmxUn8ILj1YhQkhtKEY19wkVMm1peF51x8dc17LkIZ
ZaRK1289KA1b2bWHQs7DJF4oFPHb2Ay/p3YzQfN2JakkG3foeKx10zKdt0bwvso55K/NiWYWdhqT
Rsw9RBi7dhfZFfv/0wl8/WqjxRHZvcHofroeRTckqY4I35Oeu+UxLIN4fzeWYFV47W5qDCJdjftV
yCik4HvQEEB/9XiTj5AvHBkQpouCT1DM5rIQ60X3h7xqTwKuRcP4ZEgslmuIKyunxxTLJ2iyfMkh
v/zC7C4JMYYCnByZH5mPpLBK3y9vDTGGSIlUBMG9Bm2czKm3zecAOK4y5xL6BolGgLW/+ZkV9yRg
lCiShZUfU4mDSMjuJOc4vYxCQz8MMaireMHaBKazOpt9e9Gj0+sPgzYeizef2J6/Qe95gU9FekRj
eVggeBD4B4widGjA0bH9w+duVbtgC3kAaQ0/h5LlQK6U7F5BzF55809i1vFgNNFTvHhLwU3UDnWe
h8NifSQqz41vJqIAB3S0s2Xlt4BXOPM/7Kcud2VJ7vYjzRthWDhq8r422V2oomrKtMH6oAJkhIhi
pUiHbs2/+cxu8Z4BGUtWkz42l7+38ukN8R2/v9awIBKP8dphtdyTuZayxN5G8iHdei33H+q1xQDs
D9h0Uiv1+kuJBlLErpyowZqysP+TAdIOEnCAjU8l6DXWaNMkEzXkMk73qt04RPVieIIhktlNVoV8
+P1IekeEtMEN5fwxthAvCCuPOxHWqAQbNvbegM9uLoyfclQg9fwk2LGMcJCnKjiQQQCDqPm1Kwq1
zSiF8xTNTVcUo7YXoUBsGVoMnXesM/ERv8KK7PwXBK3Id+ERyzvD3cfa9gueiMfzbiLxoXQ6OPNM
0qNmIklrDZIMZZcrAKzsWR4nBo2qOLMEGh51NZKj63e6BEYGR9csEoPP8ZKeHokoD5/IiBxoZ5Wa
jmKFiSP8IYmajbfAXXw/8WE+NlGjJFIbxYu9Kx8DoLmFThMghTM+55AbqmQcvNZyEzH6MtlDVtm7
qVl5KPWuOipn15DhLa4UyAyYOqU7BXE9nHQ+xLL9MukT9j3B5dPC+RZo6q4MlT3xUahfCPjN6WI4
jMw5h9WqHtb3ae0aRUURovRFbhrxKLOc+hcNEphb0HlEgDqYpqCu1POoVwtcN3sX77ADuwNqHr3W
YR6ymaeOmBG4j/9inHBkSODkujc5XwX++cI8zEF+4LfpMyl9/Z5vQ8VWH138QxROrFbT7wNDyaH/
RrotCgqsMa/BWn+FS9C1tqRv36EZuKI+sZfb3ghvAuIHvnr4SffSKNi2MGVVTknS7DcSfPyoTp4u
KP3qDM+LHrHdTF5yxWAVjG+VrA7/GB8KYZhHJPf8ppW3vL4jqpJnfTVXS/hbADW8ktpc3NJ5H08I
BMxMZ1ybysQuRMgXjLg/H0SEkKzENTSCY/75CWv4JULsE26oH/8B7Ca80qbsO9Od947d/aUjfFF/
OL6bqGmfN05UNRr3L05oSSLuhp21v+zPl3gkQ4zD7TlDJtNPJiP5nDA6E9Ynjyqk0yvO1seChIKN
Ln/+EZQttq0qY1ZMxrKktTbo041G5iBGKg7OISCdaEhvMCzYy5aw6xAcwZqYTMxuH0i+4jfPS4IP
dO6kNGMPViitxyKM9z1ZrM4crDTzJ7bTCumPyey19dfgkGdgekTXPeFLSJKEpeph+hLoV+aj7bHU
5ywrLrzDcEsJETCHoGx5tPxKwa29dXMe1GmMZQEz4E5MU0IoRZAvlDG/7+NhIGgF3aL6xg2svscG
qWQ+0phnpYI9OYOf5LKaFee6LmD5z96fCfszNq0gDoOKY23WAo08lR/zbPwJ1pPJQ6t5cQwdDm3k
jGoPAHKYvpMxBaNSD9QsvF/rvRsJ4esmge3xOBcT8Lj+v7wLbcU2CJuZAJcuXnT3md25aQ4dFYrl
21/LkHx6inyiTtmWSlp0U+Xo5XEnBjLPXP78y5gw/fybJlzR5TI4BPXR4L0i4FwS69uWGShIPKsT
hbj936FsnHoryh9WAVcBMbbT3vVV54/DeBzEq5xc7RsPeDgzMb2bJgRRVOTP3BeOSYS124KcvYlO
9NYtdY0HfcXdncB5KEL1cGPIiYD+YDNd5kxc61rMZQ/c/Mnu/iRGVGbz4kxAiPEagnETvTyz9dvj
2pVSVi+eLGVw2HLDme6hGRHuzOVOmxhNP1ZHrixuMBtqlMZatFcZAoV3lVb0+ckHfjmdW723Y55f
RqUSbo8L3IWmcMCTvNB1jqpi6dcoDF+/bxBPgKEGvEn+SfMTh7pK9eea1bHXk63OnsPV0Qylbpm1
CGGjmUYP+eZobm9DPm8Z8pbxVzOmdJbRbb5sE8zshdc7+0zGEchZWUED+KuWLULm43xhDV7NPwXI
vRmOsiYR+b4aCl0SL18RLy2TnjxsyU9sguxsH4KpYUq1SUULGmGQVKITg5LiOMv+Q8k0mp9sQa2/
FpQKWyrxiZaZqK9P4rvOaslOOzO/zZZ9KdUjbnnxoYNeep2EYxW73PQ2bO+cAQxsGUEwTr+dyV6E
blXwzVgridE+X/a27A9c/v2iUD1Mobnx2/D+kmpyzluce6MgO5wxqraWmpuiSv5/XQneXQtc+cWc
a+A0Z81Xtd30yVTsMtMPTLTV3jv9jDPSeU33FCnKKDrYQQxM+KQXgllIP6GyKA/a0qOe0Fc8qcky
Nh6XJRXwKfv2rPVyfifK4JYZIODpsvBBgDzyM/wsqBzUT/MNpI263Pw5BtlNpd5838Gdxc9ZaBNS
pPivPzHjttfNWMPyyBAPvsJW2c63JputRUYp13xs7hCLaBnv57x1J4tzgEqTIZprsrUivLFKRzhT
heC/acrTCQtUdsrQq+zCN/uyGAjmREU4+jEdVbk0FdK84m0bGZcdJIXYGKgZ0zEgPhJC7Cy6o4P/
fBBTmG0g+zHjXVSFWmgOq33YcB1h1fn8nPwAOSp/6Pcp1xcBmOqXlIQVhora0tpV4NOYfLsZe7Nl
DgJzxIUCY63XaWwuHnS3vjiHEX64xl0dvlkCD+TtNIpXmqL2GkiZIlqBDT4E05U3kOWjeDwOI4vP
F3xGzcXaXZHYaGQaG11J6Ctm3nZpf3yd0sbDtlJy8E7EMw6elioJV+8C7eeaSgnIH9V6ri7NoGv7
MZ4ujgyU3miZY5T4K5iZYohDTeaOA1mbec5Cv0Y5oMxmTufNBhsKMufDtyKEl8pAlnVKzitjCmZs
TEo+/Dm8XOcVjU/DjVY17FQW/L9NH5P3vKrH5orKCZ2J1FtYPxN9WlmYhQLwLdcUnn7KiU5HsVDL
Bf2z2RNHmIHvAxETf2GKKdbupqpjINjTr+fTFcT/c8GcFNNooFIucpd++5W1i3EhCchclmn5eO98
hVHohYsmR5t9hURtAvMTBt30k5CRza2XSUzG236ZbUPq43KEaIrqJ9ZzP9LDEJGFyqCpAGpkgFdP
LxFnLi+GUsESng4VsVw7nw72skN11myoKgaYK3Jbw8ndIXA3GlTTkI/yPj5FejI6F3yot0eMPkA7
14J1x46dXAR+9LvbGL/YxtpC2V4Y6WAPUewCtyuN/8rGb6z4A/Z532qqk/uij5jAgAMp3rdaHDLz
zB3RC7rUfjiKWSCydkSxvrWZxwbqyMyAV8i5WEcJb9ODLjllqlAjaY/sFwcjHibp5+bUFaf7Z6Uw
DbghF4Ncj3SSjGwK4Z3NocxorBEO9DnE7mc80JfuDI2+PqT6Ld5iP+Dj4I5CgiCTKMo38SAofsa/
4zaAJfS3OPpeqt84QntZhlSrZi8YQROSt5BBmAyIIbiKo1p8FT0oMDhv0pHKkB4IV2pR/AA7ZFeH
YAx2RGns1+K48XQEzsUXcjp2cIzGH13YDE0nZv1iZpU5oIvu1Kkxu6vLCWU+OSOeBB4BIM6+St4H
RKYK+xkub4J2/speBC6isbv8cB+O+STT8RS7tPTqHsQZOmUYfc1ZGxdxVoEmJ3bSgkvZQLQuXeKV
idA4hAVduE++hxcplC21tyaQUqJzkp7o8LCAf8P2Qpio0mkSPLeYI8Wo+FcC4wFP4Bklbo3YUFNc
mtE1M1vaCB5KWFx+SnyQ/ZeAOFAhzTx3VTeOpAaoBJ6l7+iHzmj7mqc4hc3J+/Lec4pN5vaEmrvi
S9M1HG6NlYdTahxxJm+R+YwNPt6tVRSNo+aCD4foPUsOr+LvLhCKlSZ/Lt8y6NXH6fKQXq7ea0Gu
iyMl3T7pceeienGf2PlU1WulAmeRGPRT1O95Td1jE9IsEqezafMSOUFgtBRqDbaCAVwAbW9ldLB4
IMhlZLOR3EP6EvMmpZ1MbxmhfxkzLpyLmaoZSXaUBBMvKuOcVJec3BnwsaKgP02nol7giXCqX8WG
N4+7U2MMeomUwsX8K02VC+y0UzbP8hvE3D3Je3/wqPPyWODC/j9y9dCYWimdDTea8YkEFDD8I2n7
R7LFhCJbXSooiiXgZ3+rUi0MwNmap02271l1cd2emUXOT4Y9XY4fXPM+RKYL0IXx9tBi4VYaV/7i
IIRe3hY8DqXGDXdappZEUwyN9qwT4p79Ff4uzZ9YSOXiMNJEaU3Nrf4V66E/VVSEpuM8S2PqEMpb
kvcQxorRvBqPi4vZEvHslqyvf7HD98VwLilfRwJzRj0AtMkZLnCTEZdUSLGg+0SQkynNGSw3Se12
zmM5UyZDlQ0Bjn5dee/S3mvQ6m/z3Nv/vdDY0bk0qOcpopxzyuuBGAWBUncgvQj7T8b2GAnbttfe
u8QpW+dWrpNTretFq2h6WRZ+63RTV7epd4h3m0ypb6YMvP22f9Q+F0ey7ZTJNGC3q3WrOIl+ZRav
/ElzEcPXSQSuUEeZl9VCks0c0mvO0KepzAXL0Yga+XN2bVwNPTLZ56H0VTv3fJ/8Yf0bVNXRKvzV
9FOSag8MAeRyYZjcOGZvVBKBs+i0bUT9N+3S5ssijEr02wgpmCFzrcJSbWx78YA18CoXK+dAhBTW
Te9p954+7aac1j9yh3Lbj2VFO91AnANyXUrAp1lXS8qyJdgyV/Jo50r57L59Q0033O9mrovEnH22
XIvdYH+hkFTCfyzuy8W+rKQsQxTVKhEXGidVa5tp/CL3IVdteiEljpiS7sFQlJq6nUIOm4+wE/rw
KAEtQRPO2xyO6Hpf3NUFa9+3dqDoPv+m+TpL80xcGGJlS5aEFvK7xmPhG0DvIvEodZBkj2QfKaY6
2HkdQOumbimsw61r2qp+HqNDvz3WIokred4uqEKn7hhZXj/L8bNL0+VWFNnJVaQDGcKlj1vEvJ5Y
zkohQFIZsP+2dYmyTNhHQpE6XsmRTcZP04gGZrV6poUulbs2toDOUbcM6E5Za68/t0jA3KyoMsMc
Q6t5X6BUWUERXM8ypKbSHbTLlvEPKHu/X5My7j56H+qG8YkEbrWBA6tv2ihVAl8Z100XNZ/QemZU
btql3ct68SSa4o0KwWqMkQCxHdDwWB+V9p5qGA61SeYQRfOrUB6PNZj7qnC9l5GXWsBVpRha0wBx
OMYm2K2J4fI1bm6YX5pBz33zQQvm3X9rWwXKnbKnL8ZhX7mudIGcLuWmNt+CcRHcSWkLikm8z3z+
tmZW0gnYRqRnB1K1XMRmD/xR8GbKJZ/28pV7ineG5CpYK8FJeK690u6OCE+feQeU4ItxXDgil+OK
t5hDY9hV207mdZjAAJLKaWrbSWbYmm6ogWREreJIYg6YlyFWYhU/5LVzZnAmbLYxjD2unCdaiT0+
7/OuDjZLxeyHpEG2KdU4Ij8Zv4iwdUMhm8EHkmtQRZ4d8gYWtqRuBB0MCizr0hn4FEAwEcVgwWK0
MDNIoa8FzjewUhCVLdZjPsOSTEudistzBXPZt9nbOu80x8m9pw7rP23v5lU8bysPcj710fwPBlh6
AHw3qcikrBk8Ld/9Gp1getSgx9tZ3+UWUvwYeyH5KcC+k1z3WER16NUL/qE8qPFt7vP+00S/eBzZ
Ks/XKcCSjFb2XG9N9QRQ6UBEExkBT86zAVMkZscrl45po1tjGuPfycXMCHpN5ATurxLjs3uquxMw
sEC1QT5HBeMWgFLB2aLYA6+gYCbshw+plmsGjkgsuVqFUVO8+Bq47DUAhQzvoA/OYHLkN4MrUhnU
sO4+oskdnHIUOOwIr3COeMDxP02q/2tp28jRFShJlsiorZhyC7NG7RV9bs6HsdQxU8J8truKpExH
bCv1R1pACLyx1BESjM3ZMVWFxYZRq0ks6LkDeTdhm3qa70Jf6k172dYeLvSXcMyYGDEe5MSi+XLt
eDGnAtu48GSCKIdjv74ffBineVtK8Oh9tKKi6IZap/3ECrg9WkHSp26DIY9/wfHT2B73QZ8edXg0
FsQ/a18T7QQVY4dg9A+R30Sz3unzL9n8NiMtUOhuilI7kkEzOjy7DMniID4Yd2y3vKuNFL/K8w4i
keM+oaGDBss23jBTEsBX/wkWjfutzJBMCC9zyxb5+G2A0BG16LR1bpWka1DhDrx/Dfztvku4KK1R
IGaWgtkPPZZH1SEw3wuFiodtPzWzOVPc1wiCJm9/Fji40sPt7TUJoBJI/QMxr0Wm+oHWyjweD1Z2
9UNj5yXHFha5XPQJvrcCgIuCrAihxmLP/PRGGBF29rBQ6aMRBQlIFBGT9OtiqoxgVwt7KscVsGc7
bnrSsyBYMAi4gVzI9+JMqMa/Hnv4TLuufDsy/XMRuEwaPmDlGxHDDq4SRsD06r7P+HnfxuhFuj8W
M8a5LC6TVTMAj8/fjspfU/bnCNvvzqpUStnfcFZ2ivtjtcwCklGZGbDHwU8SD4dHSMPlbDqRrZ2U
7aO+hcjIGos7AHcNsdc4IvWypNI82m5ojbEXLr0e+bYJ4FjuLmZ1D1dWXm08ZRryQv33e3swyY1v
7LA540YmrPZTDpkThc9iQudEnykRiDyiPHZ/aBTIL/F2LY4PawClpp1PgJm3JYSna1vSVq2uaKRJ
z+RzBOv/TRMsX7lpJ3+c3nbmuAFc9Cl2+ydxhupYmwmpSAEfUE1/zN+3qhjqck+tpD7T0bJt5oVK
F6FRDm3/EMrl8+4m1t/vJgpqw5QccR8vCC90Pm8fntpTPGUt0ymnsNKzmCYTSmhUUET+NSoc1lmo
uvKAFZLUEq7BAbh27gVzu3kbWaJ32WcJqBvbxJDW9Uk3+XjcziAiGv8F2s1I0Yk582w8zg63tnvT
WP2riVIBvIJObsQCLnD3pbXA7wSOwbSoAHfVpGIaTLR/nQ8AlVb0SjQXzlA2n7KHm8SfJWaX5tEx
LlG4w0AAHhRrYzBMjuelTGnnDN1LFhn+mjFuKo88D9SyZNHstDElv78wLjxP3zkyYUPES9fom5mv
OoiiNuwVnBYcFlNgdmxejoq9pl6c7M02EAqPnlrQVJ85bqEqwOONLoFfYOwX5oJQ/c7oqhHO0U35
rqz5eM2HvXeDrEZezwhtkmD8xwknfdHLata0d94peVvuQFb1oF93O9Aj1WB2EE8szkE8lATECJVf
d3yTYDGChcnZmYWOP9HbJQB/hKhtqAkQGqJXxixxjgn6UcPKEEKDkcHEeEdmj+BMeHPqUVtptD7F
so2J9NgUzYqdkX17N2fIBby+KFLZOBtPju25lVY4oWs26wkoYjImpFacUDc9/v/HO7z7j2Hr1Da6
I+XPQt/vwUT4HIo1rOSChfyQ6FRiBcSVy4esJAb5qh3zXip1GtNOAw2dAAO17ciHgoQ8Fb8smxrZ
dnMRt6K3flDMdGI/jRoGJm3GYSXaTp3HuMehCEExBVh+gWugZvTdSkIyBOiuVwnRbNGhoLqXVnKT
vzt34Lr4ix2ylTU8WasWCxU4unc5x3okjtdqw/arfZVJdH0PBZkHpp0jn0ODtkT+2m0Oc7kuZtwn
imE08oInhrgjtES8n18NLfUM5dHhGVWVTkU/H4i/28PhlPNZdbIZTbAOjpn33D2ghKrtAhg685B1
bAemt5sovT0R/3EaRDH/URIQSe0Zzd7XWi8DOfpXH+T0xZdAwrL8vmFFGwYVtD8PI1dxq2TvZoB9
6ExzYF6iMb1gcZIvHtOA/o7DA0v/FkoYHCk1aO8LcHiijyohwhjOP9yf1JydAYJQcGS9s3gaje2O
KXt18XpuSD56zkLMqSSculdIknOPqoUqpQMbmwKCDteOX3XMHWUALZt3qw/pCn5QoAM9aMag87pU
VeijmNswDxHFVRd3trfMpRfHLrAX8Blvoj0mbswO/o2I0cFWLwKIhmGWypoWDis6e+F3JNAKR2eg
nTJApG+U0SiSAJURXqmegUuY+Gm9vyhykdIxIFK89dSB5wNxDZPKu+9gypzG8rrmOMSNEshuIGs5
qC0Oz2tVx3e08GJu2RGq+zh3U+OLkX3r7XgHYp0btfvjo628eOoJTjtvXHHaG3PpFiRiBKwDSzXo
UWwWz2ThDj7EwuGNNaP6dwTyJPerd4XQLFitnU8dDMloxio2GOWKXsKP3MTwc68LH/DiTG5z8jk/
jinglvwcOuMtPhuBQEtQz45r/GLggxX0+fiP2dVLE54vJr2SrxSbzaKtyzYNvBbmuQ0mVolBEM0f
LDuSsUFsXdhQAjUye9pHtypBpAWSmvqUBzAFJYbvwvEEIHMacJg0egqL0hEqBqGX9voHG0X8aRGa
4azNHxonYXDJocQCKnHAjCI3BpRJwdxwUrt7npvoTfCbCQvFM5vHKAf5DpNvVueG3g7liaizqT46
KDoI1OGNwWecKZbKOxdxdSeSI6VPfnEBEq/u7k9OPeAYgQq04E/BcrXN1ONOJxSjXyJGyeg6A5Bj
ulRFa1qa8nJOxOo9xMHkooomzK/Z1EaCPzz0IBVAaSRzlDiJyYbP9m+Ycs1RwyVo7gSAWrb/bUn3
wIxBPux2O3CY++OuTeSP8UgHTtGmtea8gO5/izo8a3ZwxAjU97RGIYQe7n5+K18gdwB/wzUdL/dN
8dY53iKIYRs4IadeMP81u+piej1POrhH6Wk3XLVJjSfRtSuLFOcTopbOjcCAy87pdnZHdV4oVu3f
aUhIL2tT8HM1YkPyDuHhyp6Z9K1XOCVCBsMermAodcNQG7as0W0Z7I4+sjIYviax4v2Kv1x6CHMX
SP1ee043UaPMAHG7Xk6qORa+1bOhTgtQ6BqaxXaqKazJBYkKljlBUGiP8hB2SiC60nPyRXmIPgOg
lQ0syCCAoKqcHh5EU8C3UuvCs6DXz2Be6U38/yLbZQnwaEQwgrjWta8vaxtl6mvhaxo4uHEXEqfS
6xo2qDRl/U+6sdHCv6LTto3511+7srv73o7piBz94qnqpYPX0x6rCm3sKNnkto3UEfTzO5mH6Jad
UwpNlPaKwvLb8auHXXuMlreH7SP8pLXxd8TuvrhQZf30RUuRaSSxebJ8Wwk8tQBlC9HI0yXNJX6P
gFZjNZB4Ycz/HP0YNgWnkMTF7EknoZr7bZbKG8Ez2YQdiowkkQ2MGGkNzYdurAyxjPUpXjR0KlrY
9cI//Dc5swiKxMOf/U3ga5qnfDIFRK3Qh2i0+ucuIihUI6vdLEU4MpTR4ib8kR6aLg9LDl91yLyh
o/BFXgd9H+n1Lx37cUzZf7TjnmypcXlISb0hGOKnEfyVmGK5DvdMWIZExyzC3j8jyTkohG9qOlha
5Ue+eFqaNqvrZwG0Ek0guX6pfEBZeVQzS31A0qT0SyAD1vEp/+kOOnZJVmyN/xRJ3g6MhlGm4lKl
Fx1J6L3u4HXDyfzkKwACl9Vly0zr6uCeApgD+xS2nwdUT6oHaGGCLeBDNRrFpHtxB/v116oVDnvp
ZZowE1JDyP7EY0D4beaWRQHxPLhv7Tf9Abo46Wd5QF73gy0uqmGo+MEgKpSJcAOovmhEnn2pYkOu
p++znh8pWXlEKxzeNrE2Wu5vR9UNHUozF2BFeWiCAkRC5YT3zqZGF/wfPN0yGCyKMVnzZh+0VLWM
Ny7+mg6bkbBXyRhY4pROzWaKRO8PkuUl0vo8gutKLzBkMQswyzKbHBaePpBzpFuCh8lWeSe7XMDp
ew65gtnSMMansmyLPS4B4VcNU2+ISQlKDtfMkrhs4IOxsEf/tJF4QKT8zwrcfLWWEc+5XI7oYsxB
3kGkp85BwCyQW5rmbcJy+8cLPvDVjHGeWE2EYHyne5AozHMF0RXZXf6/HCrknAOQxVP6q30UDk4q
nBpzCGAhOPxgrWY5QgWTnmnIQ5CatAqdpJ3WG4SGCVtSKF6bngsOEIAhBlA4qyhRzpVEK8mSabrV
CTzGrMTWdW8K8dkEPPkmOT5+zOIPMeC3vM8Q9Gnne2sJ5yBAwxZOl7F9RxbuQy8e1SsUc4AEd+RT
gtq9w7Nixqc1dDVGO+zLAiQdflZ4HyZmF+IuNMPIzB8rwUXFqxlhDlgBmMERoaCVMPHRSOQTYuMA
sGCveuugMhxD9RJ2grxCsCgJrmwiXFJmYD4ecvh4fwv1N5w3PXev7kJfYVRmKOuhAFXFyx6t84NB
+atTBK126dr7I6Z++fZpYhGqe+Wd76I5/o0z6r+fe3C47w1WfG4CI0f8tbleadmev0IPxrc1mMxM
wy3MLl4EV3xehUIH+J2ww76T5rQtJ3VwK+GH/negKsle1yprFkraorF5vJkZourDPtZ99zZBBChZ
0htInZZFoP1QkP77aBhtUiLvpMt3F9o/YFqP4ViYSvtd4D7hVqP8IovN5TPLZotZ7kBflOp7JmCk
2m36O+Jq2QuNRMWSSQ0fbOKVSnCDeYnNfOr4fnEbdEIdFMnqjx6UK/RcLLQMLBRo3snaaHM21qgC
ehl6ENdEN3gp6DP5DdtCVRR/kgv+8/xn1w2rJtc7bXfsC4EfztJ8ahf2+xmW51g63bgT/yV5mdpV
5fv+gLrFuUKvKWF/pQSmDnGKWo9N6NMTzKqHq1LThSHF+N7voTh2UIjsvQspeia4VhQxlFn4Nxze
rnv/6LU4YkocFMSEUtD7b3kbVybZtk07xy+iSLrO9IynLAGqQF8CuGPQsJnHboqNb/UTUf4DGKPt
ge1e36KRDKDu/3H/+w3GlZOAEsiJxzIFBa7RWjRIH3PjlnJP9UpDW5Emu8LKZuIFmZYcGteGhZmi
0mXjyDI/lk6C66QslhXq1l9IarWoQaq4zzwBt/OPHtgDoXgbMKb/GilI9iCrTuucK1pGcumBQDFy
Q5aYJOegm4qFGkeSaf+c0Eib5HfSsm/zDiB07aX6V7PLJBFq1vGcRNgi2Cjr99idgRaIhbhsZtLj
jSvL9nh3EuLwKMAvP9d/YkWuD9IIKEV5T0EbxsKGE3FXw1A21Sco5C0Fs2fKV4DTcSGlxO7Mt3l6
Z/o6jPoeJmuv7Dv227Nn0VDgwcKDR2WW8L0ghpYO8DM1LzmdBo0p9piSO81l8qIiMkQ3MN870LwR
PAZbi3wpE90a1ezRMwgWOmRi+T7GR9SVwVofWZzm717O7zh/1wG//hQDMcgwT37cZ1Y5ZdqGXuLU
4yVBJf+M3ANrAkxzRCEdWx2XT/+nYJTG0On3FuS5eDYM65qH9MsIwTE7Vu/DlB+4hl1gLOu9a0BC
qS2hz8IvxhwMGLu/AfLaImjVONF5rb5PR/AJ6c+mT0fHLC4Logn66B0ee+21pbc2MwXnbUtR6UsZ
qycIAx8gnEGw1lBpPZxHAUtrEwrWB7hKqIr9yR4WKOApufwe4Pjpw6FnsC5Rzcp2XoqwqgkuFcKn
GIkOOe9ZpsU45SX9FmFyYPqk32SJuIrLT2/ABL71RlzhhD08X2mUFyvV1I+e0UXiPsDpZLzAtFBe
TwjMgbvjqo0aFG9RrfKUR4n4+ahNp7vIS1q9FnsLFLXXmrapBmT6RfHDiwrXOKwmJkmoGWI4CSrT
TQ7WEbyw++gOZBb45PtmJ+gGAn2UNOzzeZUyaIPKP/2tq3G5dTcAOKw+OXA/0wvIlwFCNWjCZzT8
HrskCab2/7FHtl8EomTiKZ67HbRQJJpvYDxI47bsP1uDHao3bK1C2+oZp7gJbKCvVpPz3qOur1xQ
fyeFnaJOlV4pxfW8UcDZEN7V5GV5UECLLzYby1GF/VwWeq3kkuIjmOXerWfsbeem8PXAj4QnZVwn
ko0Wt2/P2ogPC/F/2CF+m6cmdsz8FTcpwquJbh/ePJ/HL0/uvayKSQo2W9mTrxP3OKzpa7cqJ6fc
Nj5ykV0CJA0sVCkRnUC6IDeQRg4j8dfOv8tdAGqJ7jWiJTbHsjt3aKJycB5AxbWlSMs8J9O30cVn
JkiuRjwHk4xQRVoy2fl95nEdBBzljRTon5GAwECCcKNiJxdxlXgMMGIbGqhds9OQs9i3H1JUfM6l
hIsxOj7ZWHQvOoyFXVWPlZ4llsoP3Wc5doJFbRlM3ujD0meAV7Mtv4zM6QAl2zbJdWrz4/TeEFl8
RdAXUt6DbNf+YJ/6a9sy//vbuqY430sBRm9gekuU8K48SPBsr+Lvfa4l2a71Y5BsEI0Q4X+engve
fOO/0GzHRM0w7wS+Q8QoTrgPCY08kDJPYf7xJEEOfDxdcZeKJwNXwy04aZZ0iAup0AV+BSQBQPaj
F8I0xIjv4+LW3G5YH5serJqTjKyxiDgYO2ofShZWpqrftrZMlZT3I1wVdOJYcGngOnD8lx5YJ1Ig
+6WUyRCNk4TFzntUCIBNMMtfeDM1YudmYpB9mcx7DWp1ojY3CtQ6koc+z9Y0oIkBJW1eMAvPC9J0
EmUM31EVrQ3oAOKXt2CpOdMROWqnflqEZxHvLq5fmM1ZGhKsDGtNQsBrVXiajYNUqKIr7a2VoZjo
B4esyQN6wI1/xkhYnUitM1Cofk11KltDjj+HxbT3lXu00Oxc4e+hoChoM5C+obQjuaZvbGNfJ15b
g+Nb3kCuiiQs0Sed18nTmClPx/FZj6i7ncuQVlQYrGJSKzAEnZVyFDE0Yhphc76Kw4XmQrGLESct
jSlRbuPUQyUH+8JreWyx1qfSoPPsYEhUaQou9aaT1BhuYA328J+rFHm2Dm38dzb/xXWuH1OcCKWV
HWifAlvkVrjVnlei5301lm3c9f8mn0ZiVfIWoq4XjW/8AbZcfzRCGcaoCZemZrlW7uEKkKKHojK1
dVXJ9+M4TUXIiNcammVKaCFjWl9fkYxCGE7IpqQRhbu25wMdO9b2Fq74NzyoSDYOKw5bkOAr8te6
nHCd11b0lDmQmYuKMk3A2/YS8HiXoJkNDMu+7uPZArlOVqKp9eCXW071btGZj4y15I2E+vKPic4O
NPUU71aT1LIbCFSkoDnOfQQJSVjNi12XVNhChw0kHev5rc9bntFCkebhMI4qjhViRId1ER9UjNna
PhCcXswD8Mmx63uJPLr/6Gf4b65K5pdvbrF+o5FOO+CExiP2xaq+AydHeR4MBoNWoT5xblijvKjb
RaOqeeCatwTabpQBXnPwaIDOW7X9URrAdu6lAfX1YErEt+i8lB/9mhZD+zYkTChDlHjemV4G41RC
5XGmYSPRNZA1HafhXq9a9e/OSanqrKsbOc26THzDJLVlSWF6f4YDYPEUwZfLYYQ/0Se1kyKrbRcT
c7EebLcS1A76cQwGYChthoQp74Tr3uvIQDfl114SK+fcx6HBlSC5fYWPIGtaY5q1VI5fWuU47ygH
FaovSNLLxQMUSGC5JmFrl3BZL4RvYbIa3VSAZMbqfY4MVBb7MaF1SbD45RlDuZCfUysQgizyd5Yc
3726VIFk+ANJo+QDcIBJIjeZLXmu+Q2gavP2lkcZrcEY0fEgKFVvKBy6TCsEf5nPkYDBFdcHNcGw
PBxWQqPhM3F+szbD7hArGP+ilhtw4jAdEo66dxDB+PfjZ1nmtg5NdpGKiyWsZm5tcih82v4r3hUK
shLBO2nAhE0wTLqVTTz94qSEDrh28XwInDUnG4owE//TF7x45mL/yUsIfLfk+5n4WTmZneOw9qFR
3NnOj4pRoaems4toUi4iR3GJqcT8w6aFHPRMF//rP8vYgPrk0GyZpf7isifMxJwtvmyq6+0TJO5S
503nsC1/o2WUimFnbvalYnX+f5DMUQ+tmIl7w7ZUhkMCHqDU3mbPYU7g5BNnfW65tMBEi4Q93P9i
AEgYbXdfdR66BSYL7ylH549RTph3yq1LZEwJo8bryfcN8O5dFEMBs/ZMflJdskCAKicyuaDM1MdI
ryLE0Hp9llJosluiyJ66U4sOJG6pOFx9yewUMbIuWoU7BhcF4gCqjVJkEAs+UUPm6z/BuakecIK3
XRP0K1SFRqcbjqS5Y5jEP/11WH0VYPt81lQigm9dv8odck60RRYBrZ065Y0yDp1IToOr9lZ9a/Fq
6K3O+OgX7XI3wRKP5pDukkft/gF1BsYtvvXj2rVceSB3FSjNCpHmYpbGHWgJjZGIXrS1XzX+6/tA
MlVfXOdJOyw0v7UN32TAswJ7GKaT+hOwoCq2zeUpwKFocteud4KrqSN/B0lbQ47VUgtBHFX5gHHm
e/rmi02Me46CEfWneJsmqb5ZhGAyq/KncyaGtKaY+VlH7s7M4jYdpKfFMM15uz2850369CrKdnsQ
IWJ7xZYSC6nBWFHrhF7geUyqs9c02AtvYnFh5pjbmgKRkHE/EQmqROnC6v6lWVe4E9aWyJyBNKVI
pmMuBSLJ921RknlBVKwv7J0YAJZvr+lEdZkZXcw/sc7y79FKqizVR8xPYoNHO3+zfUaEYvEgcVPg
XKlvnmUIvd3LA8aRHso4jqWYqnT2TGCd/cxLtJqe0EsX/yJ+Y2NvhWjnuK23oiNKEfVyeazmgfKk
0NK68Pne5vsEz6M5INzSCucAx5jdZx/zHSxH0jwLE61UBAErJcX4171Fy6kgAIxIlYQjJdScsYdB
MNa2S5J1trMZUdVtJ+0xgJFiSZAlrL803dGY2DhEveUSR2r15yb5T9o/6KsqwuHoeIsvVIu7t3yw
H9l2MwQ4pFW8VJOxUFfge4HaCNRGBiuqPeHCOAtzj64g3cGHUmnjNZ6hjky4AGu272RD5JxF2P43
SlyFcEvPefmGGOPCNhKWNZtjcTJbW80VvWWO27CG28qvmYC6hphlX2CDtxEWolmg3WZWjhDs8ba3
0K/IX2aYb1puN+JdpMgjkg3KkN/Yos2yjibsPKwX3GFPheIhXcxaQJQwzgp+No+YT70g4XyJqi44
Zwc1H2u5R6NzIN6RApf/C+11fAWK9WRduosVmE1eLwekIiRuC255lg186o5NQF+GXAbCeLhCmy2G
UmQGOXF0Dqim1xZAUdlIM04OnQC/nujmeZuY/mBdwdcU2MWKR3GJlQXOnUtYC7w1S085the2s4SV
J8WHVpwiAjnf+8VRxYYknrZGFivhdJQy1I0Ua1GfuP7It9l/0DsIAOfMXrhlQmzj8y0dPR3EquWa
peYRml4bXGJw8bBMxDNOHsi9qrNCpV3f4L0O+gQjRHZ2qtvJt/7PIozoHjzA0yDWC9ZwZY37QMZ5
T6AoETgDdlcAowG3O4J7O6QrecyETvO+NncrXZSXCqq199hqMKgWIzYwSPD/wjNg4jytFDaAGtta
9ie+IUviCCoxDZYytiBNzJtEQM1y6k85r+NjDdWJ3g1n6Ai+ORja4zctBG/BDCEOkXbOlRrys0SG
KzZ/5wTvdQcU2wV7peUMWoSbulMzmkyKMFodVDCIslNQVT4TLfYR4h5Ts73M5TA+kag0IXNrWS7h
IQr63jDgYwxKQKYGY0c1613dw+vuFi3+6TB2xh2H3Jzv0RLOTKdiG1XsrhjaT6PxcHN0rfJgWLBi
cX/YDJxsfih1Vo0F+FBvuopOPQft9IS1lUCC/LvgB/t5SpI8no9v2aaNs/c07WvJiqya1Hp6v+i2
xV+gclLIdCI46pEeF1OaiGfrKvupkqe9bAai4CNPWGGBdN7Eg+M2nylLYMTN8FkSM3YtD7RymBky
dxYNVzgXuN51LqBOUluT1TuMLZCbmkXutrIoEcF/X/xWYJQ4kaKVswRWWTSUGC0wFUXk7+7VPWj6
+8rwWlTIesHlodbYR/U9ruxaWM+TpacqVFnVPMsjA1V7tTXJxqV78TgCPTATZgUX9XxkO4AD/zQj
Tt1nfckTVJ8s8tbJQYo9I5QFmqAYgY942KrKhROIfH/IwngqZ5KKmOBeHBW7SS7WFtczPUSAUx7m
FDwL/+GHnWtvUKujvmxCQBkgIY+ifHBLBaKap4gtxBaQ4eKWM20RpMCgyAYA4ZnBVqVUuydcRX9J
/m7PeG/Ep7ooBW4H0NuhW0MLdNIvnAmK1mpi3+rRxpQzxfF0wKM786LnBd8JpqE3KKGgMFip/fgH
0qiTl7m/dk/si1k/o/oNkqmq0N+t8wNM4DsXJ87bQPBTv5Svg5QBFRzSOlLYPuKEx4UoerVwpBsv
Njd3raUb6RuV325zAHLeH0g5yTuqe5jle7WsxKIf0y3ejrpfYU1fFlDI1ZDwnHAWNpZEPfJAshWE
BIMkR+YHMtznfpiTXUDcqzsl1L9Cbd1StGAEP/+9tlSX0LLvscoJNudsJw9Dwlwud0lB/j7GrtMZ
S9SX8e8ZANCs6iBUv6GTI7JQYIOX9zJsGd9lfo4U0qkmhsOKbBt1ADN5yzgXsFDHH/DSQYBM2fUu
df6/Snc70lcJlupa1fLL4nYX0DlTy4fo0z6SOojujkjsamhpIDJeF+LFE6+wrnqNWl3ZbNtPN9ZT
qYqA8rmBT48K5EBPQ3rhGFGPddM7Ct3i06tEiXBLal/+jU8xzurRbBJs28DKiCk9YZXq+PvE1uEe
tuMNeBzujdLU5BfkIUm/K8Ab+cSO7r8TY3jMTfPuDpwnFmpoWPZ+Ujl99qD+CjXP724XSS0kUuf6
BZ2NNq0DLmzFVL652XtHC8G7hoCSmOh1unH0ztGE5qLSqyf7Qrj/pOEAL60yLth45tCslCFbPa1o
VyRiOAg1QCD5zlFxrcWxisZV0lmem03yNUHenrBDXF42DewQxlosdEcVk2AVFsrL/Qg/qP4gd7FH
7z8oDCsIl+SDU/nsJVqArkC/ypwSBYNVcJ/rw+Uk3AndaZMSir+iNzJBl92hWgUjpA3i9cK4tJAW
RAsadXFQDzNTNd9gRAaVnSC4CQKXbQt3CqpPNfaqddD3A7X7TaeCjFW0bmsuhhSmDezK3rxF/ksb
kxs2wzJs6H/O4ebQqKLXcbVcg3fUoe0+Li2UqJxVARtACsK3mpa21LhHIB+1QlmNao1AYE+fUsA5
3YuCeqUHUoJ2MCaXT20eoBzgO16MtZE/Os8KxGYroJomN/wxMpuPacPHxO7s3M9PYxmapcLvQwHW
7kOoMdeLChZecSZ5UoQKJB1EknJH2hEXUwKLXbIXnXNnvJVxiiTs5ya8Ey2gx1cDmlE2MBdguDe+
xqCXKakHA47zzhSIsbsGlBwI1GfbTdkueJhhObLaY5+UxZ7aabdS+0eFMr4wJ3gZX6VFHDmdGhwg
gPwIy3sKGgk6/fA5dupP8SsvDXnraQjc1D3jiwDPb51p4b18ugMd74SXdj6nJMwGJcqA/uJz+SsI
nfpRzwzFqM9qnaomW5ArAAzTOhMJjs2uQRo2p+DT2I6Dr/fIl04erOmjp0hZXYikBC1xCEVSVyT5
88+Z/ILt0uy8MFcaSA/PLDGoKMmi1E5gcMFAsMIfT0+sL8JjIih9ClruMPJ2Y5tM6qhK3BP05zGo
KnqZUhw+qeHMQFxbpy5i6BY3Lrory5kCHW3dcmmNKMC40zjdXyY0dUiZzrAS6LRnSrGnYqbqvzha
NMqNqI4qAvPv9PAKHpJcmZdAeCBmnXtAo5KJPoMHAMT65dtV7JS+tVhR8drnd3VHpcDhl6h8SWZ6
MOn6oaDbA7is47OtRbpeTa54v5QrHGprijZ21nQCQQnwI551omkRLXlQjq4g5n29QzKQgyE0XSeT
TbSq7vwbYZcMSqmpPTDCyPc5vWMRpVBLZ02N3PaDIcWJnYK/SeVlzBpaN6kngDF6eg1SveJdvpPq
z7GEtzE5ePcoYT6B9YKFbD1/cREp2pFGINMTsErkTfMTcPicTcEB2IrvB6vqr5PR+OZDxoO9o1+6
OM/nbqETV5aLDj8XJUy9p8yzV9Uj1g2a/zYAi2GPGphsBIqfXxrs0cEj+4iFyI3Qp/ggeYI/UxST
D/cAdEM/l+W/PBzZNDb8Tf/eX59vbAMdkn8IAnmk6y4V0UYcquMj51gTccrogNUDjWR0YBBV1iSk
4F9mo87TUY1CP/b+vzdhLx/UNlSVZTNo5HmN+9lT45NrS5UGuDFGf5Ahn4CJwBiX71nLc6lCziyC
smQzt0oztG9ZcpB/9PVO+M/FXFO6IXMbizbwwrRkWSkF8qikgcxqZuDKiyqS+5IqwlUkLm+0jJLQ
QaU1yiGo/SvhBvuOC8NhD/OTdm9p+fjJWRJ1FVne204vvJjDJ9nPjaYu9Sr/Icbiacb/CD+lNXme
MkDIp8j4lXRNDKUfQePWGwC57qPPm3pCmw+G3QxFb6s+uNZmZl026J6n4ejy0sJlDdaswH4YTL58
mAKOscA74E7wj6ReyH2N57RP2yskiqoJMdRg3xrQo58+MTS1QDKPCWWo4ek35ZpN6t1I+3JUii79
mT02JGIK4ZgqfNdvIsWZV9Wm+U0itQ7tehDVAE1ZD6yfQlPlR5KgQKOw1M0HVVQQqCkoy2nbzMzu
VKnMheWbEkuepbSykgVlm45N9N3LP6bbWepJ0E5fVu3s+FsuzsZzsFafTEF2GH2h+i4X0uOW09Qq
7S1cuPJ2z8a8BSLIPl5FroOk3AR1BxypyK9fcXoD0toaPtWAgkW3n+tfjIt1s9di3IyCSXtB7fX5
lJzQKkhkUv400pfjBhQYNajKMPQMm9eKtRLVSAux022GoKdqh+JM+3nkwJvuZL50/5Qopchpuh1k
gf2aiyTv1DACxdmv0EV42qLmFmLyl6zhWj21wTUfR/9s+ZjCmOWH4TjLeH/9AVjdzhMizAZir+4p
0cMxF477YIlP8iSDJaBjpYk5ByvtZYqNwMLtZ6zh7Ay59B8ljcDc71CY6IQCgROFydbLJ2ounMBG
izmZYzpSKte5v5mRSFvRSuyYaab+e1G0B/4cr06qEI1o5zuRq+/aiYkdhj9iNiLbMeFdb7c7ZJ5q
EODoA9AP+azqqusrurw+88AaBjXLIZOHpgpd6uHuIthWDBVEDDlNep+v3tEhr1V5RjHmMK594Uez
8Ig38iQHg5qA8zAQ7Q0YCR31gTA07vVY6PzWl+95Bw3tvnBsHML/0ZY+ggsVPXsCpfJwWYxD3+8l
ui2B5XSZFKU9EwqklsBQqpbWKb1p7tHuY1vobpTV3JMF2xMrqVm6yajnOAEJGAlf7qomBur5ujGy
HvuSxHTRfhaqgxEE89sQv613aok5QH/I+C7wbpy7boJu/V45jaDEE1sPhiPyhGv49BjVQH19ezDV
5pG67m4KfwOeFz/FQyh1u+ZkPFPwhlDcgu1+EeaJ+o9k2KTEFk0XUDcHOaRBct6Bt1rofpFLjRPa
0YqSKkFM5CAYKi9UX7kf92yU4m+VnE3O68PqtCqxoiqrQRem53VwbSBXkSLW/TK5hTD0Jz6wk8Dj
9YKD6dNgUNWd9HHPv28lCb/Bo8Xzu9u2h3/9IxNhO15G0DsO4U3tZMaL51mwsaEVquromy82dWQK
RQ/FRLfNygXCg5yTbeAieg/ojUthnEcS7IJ3ZqQx+Sywl5QPa05Pef5fhM5nBOPpGjxL8RABqZyf
eUWEitAmfXZ89MDahYnTIOSXNgCbOg9joffFAc3HlC3RONGDKeWqfHA4e9sy1Vqd8/OkGajQ34IV
CvkBkTsk8AC3HWnHmVi6PGSLft6/LapbWptiOuhT4kWYVyrQ0sxjuWjqpsAab5fHqpJVHVRxVEVB
C+SgH49QL/tGJ8aSpMV9IQVfGGycFIsNGqI7UonzvJsi9K82hhjj4Km9ML3xmTTNZfbBQo3BnsPb
+gWe+dUdY68QiausRPxPdTL3bUf/lFD9D6bU/b/pl0VLTzEzTlqUM3pQTjBdIHMGcvEyoU0fH6tq
G/4C/p5aMlic5W+BuoYdxenbmUcMGq2ruL04owgQ6jp3mps4Gl+1/LNPUZGGLm3aZh0v09JRbJrS
+A+TcHRbguT2kV1u6UqEX/NjAIX8XjqYOUjra7Jkk/VaD18TXiGPufDhm3FVwHFuzGrW5OyBKjiA
PBzesrwbUYBVygQfWACl1bJ8LLOqbuLaW+O7B4bhIyX8FszpiG6D300eiYIPVYrFpLG13rKwvQdM
dbnfzaUjJ0cn5EBNXyaeiWoORqeAspLod7Z47gOcBF1IlWrEOEHvz/onzELLU9BbvzcinutVWHZO
DHZrJH9jt3RWlg8HZjyR5Jmy22PzY/HebaK8/2sLoTYPvSiVOJL4V2lebmmg4Mzb3tezBkhN3QOj
dpZjGZrWroDGKLy/grsFX20o80kDsYMxVLGb+yotpUmEqB5Zw19HOJvAaMtyHytHkaBwLm2BlT3Q
46IxnPKZFSm2CEvfelG5f1Fn5WHO/g+c74XQmwAgpq0MJk2qpenJfLbB26z6RN6FTW3UqxF9Rm3D
RLKtvKxxeo9WmSBZBV4h+TI7oHiWGWcHR/EY98DZpBqs8rNu/Az9O5t1jdPjIxpQu4+q/Tk1bI7n
xc+78w/gi6W6bHHsjkfvNaAtt8MDRrHEFToNAVOUKJSpns8eeck+a6TtR7KO0wwlaJQpBXs5u2Ol
7VDpBPnS5Hqou2fqiGd8RjBmRnU0F/ona5oOTtF4mnQSg2mfo673N/4jh74mLzfyBddkaYJsIkHP
ouZ0n0obFN7mc//JwwBw5F8BlJucPr3reduPY9J+iTzmiGXn/7vARdOEW5QLY67q5ol+o9WWxvJR
iT2iB6zIOT9Uh5vxZ/ftNaF9iv1Plz+UoT69oaDYttFEhKXdx4hJJYC676xZNn6TcESZlxvyMvFG
Np3+lCtUc61uwA4XJr/yJJkgVUCwAaOYrSD+ISmeGCJJauq5F7tG9RYohAK2jlVEi+O/TPgYUxzT
zRw2ADBVNJRY1QqnqBy0QidHHjpPwHpIjMO5Wf84tnSl6G6UcU/1vEgN6Jo8wt+Af4VvMO756TmO
Llv9QWQrBKnhCB08LRc3hNApEPXPsERUWtUTCcyQ51b3/SNu9K8+LMG6q7s6WrymK9EzC9xoYLuP
B9Yx0kCfPzKVE2ZHCXlG1HpiXPA0bSIgwGhcMF2HbF1FljPGp5D/GhXAVE8QMH5MuAmYGasTwB+b
/Wf3A0znPFJojROAR2rd15RFor6MrwSc9s2ncFgB4U3oZsL99JBaLXeZjr3kn3TA9II6h/M5Tzb2
UXeasRrtE7jdGr1+yX9c9FjlHWT44mEIFPMkDUdgEFaKPQsgWRn3hMXLkhoD1w5PH+/coW1vsOTF
E9pkGzDC6FZwLszhtbaorqBqUhdDPE24JEjjK/ifVslI2RxKvMsKKbZxkDftCunF+BjiAIIItpLm
RyV0TIecQWcGQUyhskfPDvx8z5B6clNV5pxbu8eofBg0WNOC4KXTwaPHpv1Ef+sH0mk0Z+b9g89r
aAcQ/GsjTqUBhrt9m666w9GLuznQmuxYqvlzjxlVVLdc/tQm/F9TjCMXy1kiSBGDk9Gozrk5m46N
fpLW7n8/ocnVR+Df+dzAR/nCpdm1hqDHG997ruj1w7F/vAlmx64ul6qPWGr4HVu+HKdMHTtMzsrb
8lwWddfpCkURbLMZvJNJa+cJNdSzQpG43ff4aAqeWTDDzUVlJ4kxO4YknmkWHb1ppaDLmIJ+3eHh
aVvy0J3EWmpDS1dWeBTrdm+zFioWmpH3nlosoLN1E0hTz7L/XQQG98AMWBkFHMBs2qS5JiVomsrq
/rQheRWM9qPGuVahsIPs2OLzNQg7xfD8GruZI++CcCjpGiyHEdaUMBiohLGdrab+deSNsPCwsEV3
m05uCCmYcIdMxBS6LvVvyaOP8gp87wgMYm+6bxyyeLEp8i4EG+sEGUD+pJ3o2ZuTucM3iGiy0uMO
O0b2CdbVGYVWoq9zplMTbaNIOC++Yaq1ury4IDXYPUlsmtFnaSFkfWBuZ2wFMgqkiLPB/XBzkztm
op7ZCEPTgFijC0nm3Qx7yhpBGqyB5RASwq5FuDpbTr6WxUn/Jn+2jDEuJm6BRU9xPEyVlHGH7Qos
5WR8b00S4iP8MpjFHWd5JDi3oXOeAUM1fv2Mwz15m5E6C80VCZCeyBGjgr2t7XWsmLiPAEokuT5X
GBVH1Q/TVCNR+mhcYUmKIM6YbZ7VJjEnLMxdzmiX1XE53I5PDbZVUn0mq4Qi+UZ9BdT494oyx0AU
kWaAokPmL6d2FE4NjBtQXlmi3pJxcpO0e+GeIwGqN4xrAGI/wsc6nLdxVs2diBiGEfit90EtwpAL
ixyymcNCQ7q/6ebpaJ7sVAdxFj9ryN5VkpZsR8Ch4/aNW6DUukjgQc1n+OdQ7O+pc34dyuTQroZg
z1twRd78RKyKWF5BLYYI0wrxgsMirhBGE38lu9jlV+9xbPu45sSerlfBUtDZYJU2o5C9rn+ICkn+
gVPSDSoKxjljcSgJTo9sIqGe9Jq3OCCaJm3LdyWWRBp5iuLhtYvBJoB0IG/bT9wopRMSq+57xV22
KoblsCnaAMjy6zYxmdonJ22rROhnqjBZLFWXDzElbhZ7h4/cv75Om70Q8iYFLFJWuUy7wRKST6iM
KWKxVdijXPwMZh/ZMj2+pJg0GMB8MsCdLBW2f9pY/SY9i26GDAXq/rz/srUbMY++YKf9W7PavkOi
nOPGgm/q9MqxKOgK4N/tfbmIG3NYABYEOG9TP9BPXxfaxN3G6M6a//KKjppD/Vn5XZJB6IFiW3mu
/tKz12Lr++KWGGh50YHUBqs81viFkYSKAr2ao4yAvh/HgX0LxMhjv/sTmu+urH1+0ZS7PnVHX/nG
zs5VsQXutxrzU7HKndbapWtI4uOPqYMx2gY0afwjwosE/8baXkWFCReNb397XZGVZpGMzphyRrqN
5BIMUl3MQ18agipKMU/njdZQvyFFW99rsem8lU/fYRG8Gpn2yMbKw59hEQ6VKjy8lhDvj+2GCgaB
kTAFFdlT9jPtUXJKiVpOgg9JgB+yWwiRhLBxAPdAD7KtGQm130aMISCgAn5cbK2SSPmPf7GbA2RF
8+sD0wE64CQOmgETW/eNigwVquijiu0twtMKjdxq6UTLfOpQdo5dAX/kL3cK4MWZqZwBIUUukFpe
xWumDRznASUTlwFAmbKbEGj54gIC35yaJDCWbr83fvJnCJQdXXl+0lK3bHu6jdVRtF4pGCoRyphF
Bi+tW/6iKCSzXu9M0cadKzjFBrVfmuVQUSzJrfAuIgEfGgdnXAqjKqzMgxhZxQJs/0YdwlqVsL69
f+QgayBMd77lJhLKbFjntep8pXAn81n+XxQFvxllKkOFdcviZksAWkVqFBlG1kx0YpSSIWArsZAA
uGdPouzPNtbQeryOAdDPmy2VuMUqw75kLNDupret6qsFGWMKio1S8AiG7QqvkmvUh+PyY5SAyf+r
m3/rPRVywi3BMDTIFG6UgQOomogKkyl22tT1YKDgtIp21FzR1vY1pKDhOIhJZJQADvx3D1/AhdV2
37Hu2k0JiIrJioRkKiYOUyC299mrh7tLku9KGvTnhu/vLX4Y2r9N/s5GXPit029miaMK/w2vS26A
Hub1i0KgWGCUXZgfjotYaT+1/TsUUMHQfHhIN7929SjRDF+/EiC9ABECXN4xsarxyQB9yzlEFwJV
2w1xUP3Ykh+yx3ExSqA50l76cOIEQLn+xl7u+SgfHz2R2VkS1crgUk5/TS6/ikZPcKCUs4tJ+7Le
dGVyh4twubhDZetSKPSOHRh+MS0w0QHvtzbqcTH9t8MZ4eLBOrvg6fpXzajpAKJMT4HZNNA7h+MX
BcXt0yF4kVt12T+u0INK68TKWxmo+VOqvuHyTHnFJuq/AmORO8T8dLq9L+eeZPodTyxmD4gXurSf
DLtgqmEPj2o9AdnN1yw1M8xWsOvkiwEmECfuhaEwce17a7sdpISP8KgRgKsKwPOHtMq9GsiV9LYx
SToDmHwzJvIzCpJW+djoNa2z+JWl89w52inn7K/s6Mssql+PVfB4HkzVEHinmqmRMllzO10TnUqs
cUNIR0x4uOFrG5tck0r7WDz+BYmkw1fKjK1Q0POAdFn4OutyLa0/Br4qAnLeEFYYVuJK430eP8Q2
up83V7o0H8NgyRa84FvQ0CDce8ZtHR7RlyEEdZqmpBVQn1kbDB8vvMkCwowVjW5ukKa5OCibSUjE
aO7vXT283zNykt6FqpYkB1TGEWynVhlX7ePIylVnSHJnb174ZfNd00XTuLbqTV6t4lPNaqae3odW
P1xcVfFI2qWlLQ+z4K70fT23UJiLDjhuPLmztPR9TOtVh+nxv9NaQfmyxe7Y/me+0Amnyp88WBRk
fMBPYuYQ1McJsBsY94V22LA7kVVf+xj6iONwrEp8k/Vo7Q67Au+EI4VQbB+cg7YxICRoWv8Q+jEF
vetEWRwyHJSOFa0jTgTzo524eqtJlWTa6fyYPcdeSjhPV8VLfU3y9s2R/SFAmkIWTv4BCtimLfVr
I2ejfuN+R2JD/Ipo0YB55KYkMxtJSXHIBHwoBuZI4xVdHsHlEDfn8/d3sdmCCprFFaIgDcXjncEz
aqQZoMlukRaPwkwuNlstbbP8F+XGIPbD1i4eX3U0h9ItdULRPj2VGSIuobNorJ90S9MFJ+SxIFXu
fuERkLfpmMvY45JCWFvOoYi7nf1s7jmhklgyUTSYrsK7iHBQ5Ef57qt8Gn1ma5PPFdItjFHA7HlE
6iKLEgz4C7I/LVHZE9eNXYsUU09MIGJqnkYNMUEKnfKQvlcKWDiZi53RKet6nFNWHyRX9jOQ/D6T
g/7xX9drj4ZhZ0BQB5vImyYMQm4GdVATW3ht3gqZflPW5L34SoMi8WUaDJr9+4dhZkSwCnS4UKCY
+RFVTxgqoSnji8ILGw9XJGdygS8Ruap1IKskqU5vy228SCkEIO2jbFxyZTStTxz8AXdZDvVVbXx5
VThxqSYJtCGj4XIMzAfjAG3z/Jo+v3iVIFw6Ohseu2piEdhvUHuTW0uNLYN3GdggMDBZ6+dmKIi5
oG1iAre5+m8zMo54adUU2SDfuRhxEgyaQu3tnqhcsAk4lY5MYfRtUeYnAoz47rEflnq5ivRxjq90
O+QOyk0iMFMbb41UeAO9zyPlFuiQSfxyog9q3emeUWHSckMn4Uyfyky3o5a/eP4AVeZqSBUlOCFO
ZI2E8Ua3v2q2slqtfd8IvOkHdwvysdUUr5WgSS+oe1Vf7vEgWRdat0gm6ftuYuLtiRN7K0fhvpW8
P7FTBX4JdH7lqPkgaxgq8NRJoskMNJ3WsSJQuthYcMRrx+Rvk/fv09IUrZ3WcDb0V3QX78JtvXh8
N/EI8hWmESBJXWMCoN4W25vD2p9C7D49fBbAox4qcQnFhIP1ut/VlxeNU3ZzVtTDW1An0kwrl2qB
ZxTfBZUUog/3k26wCFne3YZg8cn4U1hxUqQl9Iec8OnSgBvKxXshaZpE4hzcfLPtU9QdyFiasMQb
dNo3OD+8pfmy8B6YAybhHEWrAAvM+LTPgvGSVpVp44/x0FaNLDnAielnA65IjcZ49NsP/M6+e+oU
gXHd+G69FRqNq3dyBzBG+NAvFBOCp+DkIUV2+2zhgUzvXlhYTRUgCWtnALyWpDQxeFKpMUYlb1Zj
zAhATkmkEmEdpapFxaDvEXYCznI0/Vda8sTVUoxciHwUrksgUUzMoKLrIbZLjRtHJFW4w2FZfgoI
vyTbGD7eL/UIJQsLTzsOVvsFvUQhUorlCB9jzN4wGVlG75jtkv5qnKi1K/lcsfe3LSBRICdVQNuw
SftU8uuq+l5yTFjsosSoZXKOZLCDyUX+Mf0JbBc3oDfyPe19j1pe30PXWs127kVcoelwrmeo/n3Y
er+I/ejya7mpF5cgnTw9eGoGw+AHB+xxDbo9THW0mIs9f3JtdwBol0CLLeKdsbkz6h+IVEZgUQQV
OZbxhSwO3rjtZVhL83KEqzzD2r3edlf2P3ygviVGpDthfixOxBtOMHdvCtOb5z1HbugIi73acEVk
t8Bp5p0h03HOndCMT2+hoxBAJCFm29aAOPYjVoM8vMyR/KUt/KTEaNVT4oHELfud6Xxffi5e2bvx
+JQhQq0aWnpPq0Z5F324c9PT9M4tLH1gfUFGFeefedZtJfl3Qjdq9uIXFHi6hs6P/C8vUtL4OsW3
I6mGDjqp3A7CwJEc/QflkurV2nzPNnoijevv+ynSgeXD5ccGg58sI88bySpkIyq99J6L2M9hQOBx
64lvZJeBqnUluOxKjrI95JaqiSe6Ey3sxCre00VPzkY96e2+ZIQ3t9+fIQaizYnOL+27RDcOS64v
bHb4W6V22o7e6A4KmDp05dPiB1reDWzqq3P0agprqzqR3yWWs75fIgMWI64jF3JGM9L0xrE9df6q
bb2jyOftK7oyAaLZosGCWE5AQ72aY7yE+OJ0GqDI4XIeKvUaCEPtxM+imOu6fxxOmR+jsW3F/7yX
uyjELj8Qe3P9viBnYSk4wsMvi12BgX/03UzgbN1tJF+dV6G1wZe3OqnggkFELa44D81mKVMrELYR
u61eXznaOxTHUsg+7vjpaaoEsdSlTaHqC7T4kUy2qJzRjrhtYHsADqzprC6Qsz2v4Z9Du24KwRkj
7iUK34PxH3UUsJhtCM2gAK+pneZ0y+aDjfVkkBPMRG5/mj82J4KC+sXvLCRDQsTVbAD8VGdM4Cl1
2uM136ePucBu1ZIwH/FkfzdxqsXhgRtwwVKJUgUORZFKrxRSVI31J7reEFgsUjB07fllxi9VV6KU
tBFIbNE5qk/0ARS4sHUWlPY5dc7vJIXW+KH+1Bb1OKSg6i9UWymnCK8nwHyo732XelyJwBln/EGf
nvbxZPXoVFE10PPF+aDWe1J1n77CnUk8zwLq3u5v8LT+5X4TI/M4fvVXOst2AZZJZaUzO6fJc2lA
0V2IacBo5azgWynV0S1E/Ijd8OrHi7x+Z8j3IZH++0nmWfsGxra94UhCcdy7gxzHnP7h5iXiMl09
VNxU3PMycG6eztI7kTemXSofikFOa5T+BFUTE9SGJMdi4O8hb2u6YrXOqs/Oq/7JHv5qnPnkROoe
BG9tU3rtaUi5yZCkY4jwJRp3+BG5jHJaeISuw+IOWq/REh1MDXoaXqy0yJ/9tEbe0iA2BcwHoJL0
wvTMS+EvLoDe1diAsRSyjfqNz6Ahs4roVDHHinKREHTbKGNTNKm1UVta6e0R6CM=
`pragma protect end_protected


endmodule
