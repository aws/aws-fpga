// Amazon FPGA Hardware Development Kit
//
// Copyright 2016 Amazon.com, Inc. or its affiliates. All Rights Reserved.
//
// Licensed under the Amazon Software License (the "License"). You may not use
// this file except in compliance with the License. A copy of the License is
// located at
//
//    http://aws.amazon.com/asl/
//
// or in the "license" file accompanying this file. This file is distributed on
// an "AS IS" BASIS, WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, express or
// implied. See the License for the specific language governing permissions and
// limitations under the License.
// Restricted NDA Material
// =============================================================================
`ifdef ECC_DIRECT_EN
 `ifndef ECC_ADDR_HI
  `define ECC_ADDR_HI 5000
 `endif
 `ifndef ECC_ADDR_LO
  `define ECC_ADDR_LO 4000
 `endif
`endif

`ifdef RND_ECC_EN
 `ifndef RND_ECC_WEIGHT
   `define RND_ECC_WEIGHT 50
 `endif
`endif

module sh_ddr #( parameter DDR_A_PRESENT = 1,
                 parameter DDR_B_PRESENT = 1,
                 parameter DDR_D_PRESENT = 1,

                 //NOTE TO CL DEVELOPERS:
                 // The below two parameters should not be changed.
                 // Changing these parameters will cause place errors for DDR_A and DDR_D pins.
                 // When set to 1, they will ensure that DDR_A/D IO buffers are correctly instanced
                 parameter DDR_A_IO = 1,
                 parameter DDR_D_IO = 1

)
   (

   //---------------------------
   // Main clock/reset
   //---------------------------
   input clk,
   input rst_n,

   input stat_clk,                           //Stats interface clock
   input stat_rst_n,

   //--------------------------
   // DDR Physical Interface
   //--------------------------

// ------------------- DDR4 x72 RDIMM 2100 Interface A ----------------------------------
    input                CLK_300M_DIMM0_DP,
    input                CLK_300M_DIMM0_DN,
    output logic         M_A_ACT_N,
    output logic[16:0]   M_A_MA,
    output logic[1:0]    M_A_BA,
    output logic[1:0]    M_A_BG,
    output logic[0:0]    M_A_CKE,
    output logic[0:0]    M_A_ODT,
    output logic[0:0]    M_A_CS_N,
    output logic[0:0]    M_A_CLK_DN,
    output logic[0:0]    M_A_CLK_DP,
    output logic         M_A_PAR,
    inout  [63:0]        M_A_DQ,
    inout  [7:0]         M_A_ECC,
    inout  [17:0]        M_A_DQS_DP,
    inout  [17:0]        M_A_DQS_DN,
    output logic cl_RST_DIMM_A_N,

// ------------------- DDR4 x72 RDIMM 2100 Interface B ----------------------------------
    input                CLK_300M_DIMM1_DP,
    input                CLK_300M_DIMM1_DN,
    output logic         M_B_ACT_N,
    output logic[16:0]   M_B_MA,
    output logic[1:0]    M_B_BA,
    output logic[1:0]    M_B_BG,
    output logic[0:0]    M_B_CKE,
    output logic[0:0]    M_B_ODT,
    output logic[0:0]    M_B_CS_N,
    output logic[0:0]    M_B_CLK_DN,
    output logic[0:0]    M_B_CLK_DP,
    output logic         M_B_PAR,
    inout  [63:0]        M_B_DQ,
    inout  [7:0]         M_B_ECC,
    inout  [17:0]        M_B_DQS_DP,
    inout  [17:0]        M_B_DQS_DN,
    output logic cl_RST_DIMM_B_N,

// ------------------- DDR4 x72 RDIMM 2100 Interface D ----------------------------------
    input                CLK_300M_DIMM3_DP,
    input                CLK_300M_DIMM3_DN,
    output logic         M_D_ACT_N,
    output logic[16:0]   M_D_MA,
    output logic[1:0]    M_D_BA,
    output logic[1:0]    M_D_BG,
    output logic[0:0]    M_D_CKE,
    output logic[0:0]    M_D_ODT,
    output logic[0:0]    M_D_CS_N,
    output logic[0:0]    M_D_CLK_DN,
    output logic[0:0]    M_D_CLK_DP,
    output logic         M_D_PAR,
    inout  [63:0]        M_D_DQ,
    inout  [7:0]         M_D_ECC,
    inout  [17:0]        M_D_DQS_DP,
    inout  [17:0]        M_D_DQS_DN,
    output logic cl_RST_DIMM_D_N,


   //------------------------------------------------------
   // DDR-4 Interface from CL (AXI-4)
   //------------------------------------------------------
   input[15:0] cl_sh_ddr_awid[2:0],
   input[63:0] cl_sh_ddr_awaddr[2:0],
   input[7:0] cl_sh_ddr_awlen[2:0],
   input[2:0] cl_sh_ddr_awsize[2:0],
   input[1:0] cl_sh_ddr_awburst[2:0],        //Note only INCR/WRAP supported.  If un-supported mode on this signal, will default to INCR
   input      cl_sh_ddr_awuser[2:0],
   input cl_sh_ddr_awvalid[2:0],
   output logic[2:0] sh_cl_ddr_awready,

   input[15:0] cl_sh_ddr_wid[2:0],
   input[511:0] cl_sh_ddr_wdata[2:0],
   input[63:0] cl_sh_ddr_wstrb[2:0],
   input[2:0] cl_sh_ddr_wlast,
   input[2:0] cl_sh_ddr_wvalid,
   output logic[2:0] sh_cl_ddr_wready,

   output logic[15:0] sh_cl_ddr_bid[2:0],
   output logic[1:0] sh_cl_ddr_bresp[2:0],
   output logic[2:0] sh_cl_ddr_bvalid,
   input[2:0] cl_sh_ddr_bready,

   input[15:0] cl_sh_ddr_arid[2:0],
   input[63:0] cl_sh_ddr_araddr[2:0],
   input[7:0] cl_sh_ddr_arlen[2:0],
   input[2:0] cl_sh_ddr_arsize[2:0],
   input      cl_sh_ddr_aruser[2:0],
   input[1:0] cl_sh_ddr_arburst[2:0],     //Note only INCR/WRAP supported.  If un-supported mode on this signal, will default to INCR
   input[2:0] cl_sh_ddr_arvalid,
   output logic[2:0] sh_cl_ddr_arready,

   output logic[15:0] sh_cl_ddr_rid[2:0],
   output logic[511:0] sh_cl_ddr_rdata[2:0],
   output logic[1:0] sh_cl_ddr_rresp[2:0],
   output logic[2:0] sh_cl_ddr_rlast,
   output logic[2:0] sh_cl_ddr_rvalid,
   input[2:0] cl_sh_ddr_rready,

   output logic[2:0] sh_cl_ddr_is_ready,

   input[7:0] sh_ddr_stat_addr0,
   input sh_ddr_stat_wr0,
   input sh_ddr_stat_rd0,
   input[31:0] sh_ddr_stat_wdata0,

   output logic ddr_sh_stat_ack0,
   output logic[31:0] ddr_sh_stat_rdata0,
   output logic[7:0] ddr_sh_stat_int0,

   input[7:0] sh_ddr_stat_addr1,
   input sh_ddr_stat_wr1,
   input sh_ddr_stat_rd1,
   input[31:0] sh_ddr_stat_wdata1,

   output logic ddr_sh_stat_ack1,
   output logic[31:0] ddr_sh_stat_rdata1,
   output logic[7:0] ddr_sh_stat_int1,

   input[7:0] sh_ddr_stat_addr2,
   input sh_ddr_stat_wr2,
   input sh_ddr_stat_rd2,
   input[31:0] sh_ddr_stat_wdata2,

   output logic ddr_sh_stat_ack2,
   output logic[31:0] ddr_sh_stat_rdata2,
   output logic[7:0] ddr_sh_stat_int2



   );

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2020.2"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
At9w/SOoW0wuP5cEcwSq6G4xj4HMbAwgyKNze1t5V0VY4s4genoXxkgJ8TaQMWr+lcv9JtNLlVIa
LTh6YXmRgmoTc87CvzFF7wjGUSCODbl174pmnPzQPzWvyuBU7WrN90FcYhK0qoC/9oDL+OUDyK8V
rhnwBAGEWpRqMjDO8zK8ut6tBMVfgv46YwbyRwzap45sXJu9AQo12eEcu+SkFaY8Ahddu9JowRDS
o25D9QMRpPWjx1BkzngFWVsb8JkQRANcgsJ+3CfxcBnYbb6SwW0LQO+VuPXoXwc0cuIXHbf5ctG1
eHtnxbF+CJm00JklnXS2ZkLsENXcJWFsFeumtg==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
kXT+m7VjDTiHDo/nDW48gAceiJFtxTEHbqzl3RxLsBi8qUPrc7napwDhOlfJ3a38agzyji8/ZyMG
f3kTlv9Z082UwlEXJROjqCx60MWy8xpliq3kfdZewhy8z3Fepfp7P8q7xF8UCjggPqkOmIGJ33nH
j24fw4vjRO334uhLEd0=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
BQTcIbLhs+naDTxW9Ptgw/MaKcaA64IfnZ8TsIVMQwVK9UqbW0Feg/8bffIXN8vkAVnIt5UQM0+x
cm9DXs4i9e5HBc3oFAmhFLaxRqp5aNA38mE8JxhdVY0197T8s3gbX/LVLM6mWCBb2dmlkGLLKmWD
HxolODHrzzZPQpn5FbA=

`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
enNtVfQaaLmakxVx0/jqN5fZq0zv61q/7gXujnd7Yevo0zRZn72rplCNWwxNPXi/7bA4ll4ueZBK
9CsqT99nEA==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 75616)
`pragma protect data_block
dohsirBoxb+CcKqeUG6EIQE1QwLOKZ51Q3n0IObQY6SI4efPXpJyIZnomRRf62jJqoesIDnFjOqF
h7IG/GUDk99r0wNRsrqG94CeWYm+WSd58MTfyiHIEO/dHBYkWL5uWie1KUrE6om5eUxIgFglZNGS
nnnkzsdv6JWreStqqF7YVDR0WGRLfao+d1ZsJeAeuCxOLlg48xlTHu2kZ8hqmF9CnByuP3RN/XwF
SLmzPAVmJxY6hJPHhJNuB4aZXVBteAZgZfmvASQ25QFg5ZS6amo753zlZGPVMAL8u5xEvR7xaPpe
S0/OUl7H9RCfHTiw4ZxlLVNZaJQsMNYDgk6K4emhskwHJ2lu8Omlo/0RqesQ0ez84T0vSmebfryM
nkx+foQznt9b8UaZczY0dktWbYnvN8GlQph60CA+KKYxxoX9IZjNHUxw5VZX279tqp2bIs6FM224
kutv4bUJnrFkx64Rut1+9itNW9gS5wy25pRt8nrLeU79cqWltmhHTcyp9B0CQ7+WNn3+oc+4zAcA
TJdHM2pL3wf37h+6U779BB9UUCEEWMHr1YtP5xxYVA3dR54dcUTZy3IeX3rIR3XlOcbZX/CNOORh
LRRbJs91lTnG3wi6zxbfUu1npPrqAe9RfaQEVecz6+RH/4dTYNfwHqK3/tI4Uq93bnKRbShncI7J
Wi1etkkwHV9HeCgQrh5MPDhL2+7ODgsyBbk3WPj4ZJl5J+ZgNWtO6hVXpyL2ERUrV8igcCMHQhdG
HmDnO3w6ZsmNbz+4iB1pczaNZ2zkQsna1H9M5Gi406D5s3zLN7tDLrR9VTKvl+WhXJg5jftHkp2J
iAPqbddblMAkX58RY7WjPZQZCMf9/3OhUnDTp+0smircGSNjWsDlHkwDnRhqPvXvfujxcEwCH7qx
M+okqR/douC0H/9VRPoZ8mef7Ilw2jSVb6e11M5eV6zB3AU5MjD7oTCbtYPuczekgo+s8SKCYtBK
w0m1hsSnsoaCZHWcn7EUvVT/w90Bgh4qP2EvMYJHbu0bBaL/CsAkSL57+cVlgDlIBxt9pI0htWiu
mYGlSzqn43xTdrU/IL1bHJMCGd759w4tfex3H9E1tIsApa/mvBlWJDXqpRD6TdMJCTySXQrdnb2e
4d6glGUUNDZe8SwVEADqWGSyBm0BOcUxRTdv7DbZy+YVg96gTtQcwB22iw9HeuGX9vmfC4LOR6Ar
hoO3Rm7bMWiOFxfCCd4OQqQP8GJJMx9ulrrN2PltJUcEKSJDr5EkKpchZqWhiQtAnDeRzLeJBuUr
IlK77ylIKIJGdOBG77pueo52+1HhWe5Kv4hjVoHBMKs/8Jgi8f0kv0/OvrHGkpgzThYONk3dgMnR
k4If77A9c3FkE0NEgnkEWtLCI8/LuGi9EN23UYQgT6qf9CWf5G1EZCxFEF2n7H8AwZvA6vtNmNtZ
Tm7WryV8C4kyI8dKO94GmzFFCuNFvtdSG6ABwsKW/vsGabsLjdL1/KbgbQigw61jnUKd605DvtRo
msCKQjMiBXbT9vBQrk4zwGtdmh+FdH/G9MXRXwpuT9vdpJF2Jua/wBgkSRUKnA+xSFxO9o56ue1W
tRr/F8n5XPzh3poLMjX4digW35oLHgqMimQ1LVCu2rEan3VuxdpcX/VC0HIatW/x7YPTQZLlMGKL
MBd+k07UmAEpTngSeDqc94ymUJ83EGnA30TZQ3ZZtOo8PPULCLJAVvhWB09H4sxAEU0d0YQ1TYRm
k+lC6bYn4bzdgVKDU+BDigarqnkcJwNyBSmLBia/tW81gI8GhAbPS43KCTBVGNSm98ViCiZWaGUl
p//xN4Qkas9NxXgvHj4FopWM3WZBMgER+Yf8L2J5UNO425K9AaAccUmCSXigxF4a5eOlTRgge7ix
1dIFWpc5gHnqMX7rypi9ojOuGHKGcJ4Fv8S4/G/iGSPnwMVSURm1WdkBVUnr0bwXSZbDlQa82QKT
5cYvhWt2kLjrdhfnyoEy0H+9Pg+OGoJUX1ZeL5N7d5wsxLTSrjxT62jvIVqCZuOGooeDMKc8b6Ri
OJD2X943vJz5KI92mEMVC3VG6cU2U1hOx+2z3oc54nIHxKodf9i9G9pBRGQKg1CKn6OYQU1I8jBg
+CuP+3a1crpdHb168tUcBpKC+3TkS4g8ME+zma5NhQxYMaWkt2BPQrxukBpM9QO8GQdukRLgxBU1
kiZGWlpgN0WkoTZAJHbOtgf4pO0PVGX9BI/bkmr0ZmsPwenTW3Vb1izbYyhiiwIj+VGozvN7zrZt
jc20kO6cVzvoNqKM1UdnN+NgEvZdGyD5zVQ8CGPbyrgw4RRJerKkFiVhQp9Kfi30YdaBKGYIdNvI
x5w7yo/QPOwEXi4fk9XHu15vvDQRRb7d903kff3rgSSoELYarM3RyC0hX+IWrmsWHnYXPTHwkQ6q
5mjB0KoQuC/JWhQ2yTthG/TYWtR7FOH6B5xN6kXvZZuBi7msp04B0Gvn8LmxHykJEGsXJj1qHr71
1dcmGHzexvZEvObqvtivmXADr9qL0N9CFqBJ6SAy4xw4ai1voeL8WTwmD57R3Md8c3V8wAFlQLNw
N2zz+4IBwZrqvDGebeGBpfE9KIYOBy8a2Mexr/EO/ds+G9EpOw0yxERksoBryoolRcHlausKYoF4
gsbc4xQY/MLV9W5tE8ZeEaMMtw6oXyL3GZkiEVdzg/g1fH/Q6cGUfyri43HXlxSA8WBRfq1nYMPi
ws+nNhH9chy8XDwMtUaYb6ZFAot7PGuYmkSSMvIoPzlTw/ZV1O8YB26/pEoyKwJxKSoa4hXd6ZE5
3o87x1HsllUE27LhC0KmwbEu5mW2WYRm/uLsNI2p6yBci1wzpgwZvsCkxOE0/VshWCuXVvdLUiML
02yeptJbL5lCkMCFTmT6I7LS+yphU+0hbCQKDyjZY/2F0KEQnpVfo6fdqCHrc/yHP8OclP4BOh1+
YmOmFrbFdq01eNZN442kQfzBkObdeUffUral/g/asfdRTH7rsYJSI10WCp8cQAzvX3MSC9tQI13F
6jy336dpemHwjnlF/W7Y0OKmB4a7AiSTtztgt81sSViWnzqcOe4kDsUZNNM6Vm8sO6rpTHiwbC4V
/3eIEjPGsHUJoR0ESfgLA98VFOlxZmJmiGNvuPUj87gEiVaAcDKlu7mpdXZn7SeIZN9qrW16awru
uQWCAxjEKohs2nYq6L9fSNJcpS516L49bSxsF5qMPzJvKCCC9GCQJ6/WRK/raxUFn8amDU9xD+5F
x2Yomvokz7rGksZpOOECwrrxt8CguwnpJguSLEcvSoGeAeaaz6SKgRvBgzNQ+4JF6O3AL+NZ08rT
CDxSjCrmLaM20q1Usvr8F0HE0JM98lIz4mAxSZBsx9iANho2a/32p3glXlQjZrDQTr44vlBT+KE0
dGVRs/+m+562aB7JfqymsCXrut6Zvz5wAEQrh1YuWpcisUszA9SBCtbOFYi5nNd07PEblyfm+2YA
Ot9eHwyRGh9VgJs6GutU4Rcks4CyZyo+nJd1hz75USGs8P8HqbAbs2R6q/Hrfvuc9Kk/vWtaGMH0
zaMI+pBy9OaD3b3MWgC7LP/GDKiOdP54oE3r1iElTUKWKf32BeP3N1jMY0dTCS/727KYkmndSNw8
IcoQTh+ouQy1pyYG5hEDNn7YcR09rpicZxlrV55+Xia4Qjkr/1EjjZJtxuoOxYEmXQteAqHrZPWr
QY8FOJ75woVmHmNnCD9lujQs1CnqhahzvujYhKn3I5zGJ630WiqRDM4go+kVbVt4I4YSZbBn75B0
OpPQ8ZHJ7NFLXBKoGgZy1z/1Im4XAm/Z4ypoF5LJ5F/ckhUhywcw1W/F2ATDUcJ0FmUOPNCw8Sy0
+GRZcTlFC4R2HTUjX+srIXTaMD/QuauOG9EhqYtEZy9KjnVZZVRucgU/71mlu1kM0GGwPkF32JHA
lrMWlliLBf6gqv/tJEG6xmjcHcS2oTYGBVz6q9zlrp4OByIXNdwMSENy1pQi9lcqDcITJncwV1fT
rHJaNcu6oGC7QoeL9f2ygc1Bv9tk/75v/OqjZuYRNlJ5UIsjVv8JjBCZ0yA1Hq5HZ3IigA065wY3
MTHgahwYiEYnNlDtVb32bKvkfce6PCbexRpTPCElB1vh9E2Kehf8bG/ZvBK7kOwYXhgC+fBr7egK
1usC4Eh65YkbUOVYTOJzSB4lXZiM3+fNUwAuVXGiiZDhjMDpi453eylEEdneaE4tcA86jj7q3Y9j
QzK2iSPoNWTgwJrBphlUD/Iv9kUO0pcA9ckbzQeRK3OxTkTFx2ZIAi4Uy3kUBaM0MmIXjv8xQUIt
1ofq8V+yLO702LVbq6ERMkizCIYIYPlsJI3izZDVaynBgqj7p9hUp43bTH7a5mGDRu13PG3HkH4E
c/fyDnskNq42WTve1YU0tOm/j/sxopYXa6xidAhnCdYms3DpMfE0LVjfGLasvYxq23Cb+/Piuki6
E8Ycs4c39jZGykaCzuFGRW8GwnM4XGA/YqCtNhBnOJYM+mAQKymIGr5hCd5dDic5ahQIHIUnAhZ6
kPbheHBTS/DRlThJ1XuUmc6fPZrjoMWstvKuomEHjMeZ9Lyn3kx76xU5hk+Q/0fMJMJKC2RnwFy7
zWuDtpZoascXM479Y8upVi8sQCIHnATMqbZcxrrilHK8T3BOGuvI/JFovVzLHdOjF7i0rJ3sz1Zz
55arvV7wBRwrpY+Cd11H5hQT3spXN8n0cvi856fQu1sWGR24tkYbpy6y5N5AMZRyC9SvHglH/LbX
x4Y86V8pQc6/lsRg1NcynGYH4Q/nYIebl7p69P0ZszaiCSNIT4EBGx0EAqzplFNDM8JxUaU+CATv
/2D8Quz7JashmP9o0Vuun4ViBse72KPG/t5r2PvCRlLTGQ1OhIODYQ/MZYvFMcADv5AHPkdVwvkk
ePi5WnRTek2nBL6xcnC3jZL+8E07OgHxY/WRNbebWmuHy22Oj9hSIiZY4GauWaKy7rPWX78C0ePq
WNCDd3K52UdGdJ3wQT3CUiWrYzpE6jQRLFbrYlCYJ+s0UAkOccYK/9dCkESan3tgM5FXf/TRsTSa
FcbzRWdqqDOt7mLLV1QRPri7B5ErOvoWOcznAW8IqRTcnJmtYP0qjVdqdZHJb09MDMxfYnCAZQ1k
9QiwVZ40rTFVKHUILDPMKpxYkE1bGMKtCymwmD8ANO5HJhyworYx/Ci81YG1b5P7UQKNGJwQiSVW
yuY6S3hDF8mKDc9mXjxrwA+TwaWwDH4t8r7zedGi0oT4BqOAc6BfGcoSazUpqyhv7tjiAWFgxrhz
Pa6IIjyc9JvRWXuI1sxEnz6we6az64yZpZu8z06Nde87AvohHQ8S2Nrm4uOjzjdB6q9SuDCKtCvp
Y0KAK1yadxbVgtgqbr3bdzVdTnyiBh7gAGJ8VkG31BbW01ZNamHIiOcmnDvCDSU5KG34aY53NgMV
haQe2WoZVHK93w0gkJrqDX/Q0EB/Gqp06BY5Q/TPw3MPik+SidS4AVgEmFsMM4K0D8yBONM/Huvm
+ohWh8x3CDFI6e7uA0NxKSNUNYbbMzUShcDvI6if1UBd4kZf0DUHvKMHb1znm4Gzm8gPWFL/IcGT
mjTwsaPfn9QoMBQtOnlT0Xkc0LybFu+MRr7js8VBmhR35JcHva5GsWhWeo42zOTJOqYpseT7rMn7
HwpksgMaOfZScQMrA/5h7Ia1LojQm4gxBCe3eQIHBOWX66kpHzBgiRK9pfDN4H63zdaiO45d+ALm
mLOOgUxSPJrMalJVj5YPGYTIYlzYsX7/r8saszw2DKAwQOY2hkd69kl4PlW0mGu7yZ0dchIhqSk5
1ytETHH9TE+8QOkyxV+pLWalXZ1AThrZklgXSjQheShkZICYFmm28kFm/Oh5du5Qo0aSFOhDJx3d
c9EtCWKykbMmXX4hvORk1hjwVob7D0zFD0rtFD6ITuoIXlgRnaTbtT9D/L9LkyZRnwJIaf0vZ4Wo
4Ezo1U3IW1LlH9R+gNrLDbmaiy9pP0moqboxa/p83qbVoZe6ZMIBcifOULTeri1H3BBZD1ekixiy
ZG3oVAcvHFg7JTZ6RpxAOlRXXUcUh+3UcZ1XRcCiHo0WMUGwIgspIFwHVNDJXF9+GH8COjhVpIkv
CTeUN2VgihnP8jte7YI0EW+M4vgWHi6o6qNN22E9snoArzFN/4jDtvzZk6kCqzQRt+bz+SJBRK1M
pMM6z37PJpQW0YWhimWL7gkF9IMO3/kEHcNrG6WRIKsHczTZ9hvy7sbLkpkqSyM8ji2vdmnTLsNb
R6rwD9FLcw10b+ZHLAf2R907ncgnzTdgApq4kmoS4z4wHJjnBKX1D7gbyr4jmGqCYslXczWbD6UY
vMrMfiS9G6SgO5/XXGCEQCwVr7Qns8C3+P+vmVIseHwswc+6Uvbgo05LT7Bkj66T9OvBoAeT5zZJ
AvZb/XgpucUXJ/Rf0rFnf4o84qlN6A7LroDAuCV6cl3/Vhr7MbOTh513EHC91URwevWGNLLDJQb/
IHRWjmrWPpu98GsOlQQiDwI8FsXSarmzWwnM1tF0LsRQzByrswZqgIGX0JliKNoHY/x1Bul5xuZx
1reDrdgbYS9M7FfMs5vrm7p/lsv/j3FkxYbBswqHJWxBSQURghSm/z5dasihF8f1fY8+5rmuuhqh
5dMlx/urApXTAgM19XQP/jwWQTIJKKNYeB8IrW/mrIHp80/iOZNXTvKZDoI2feaKzi3IE41lsObh
qbS3PXj7IJGLtTitXuUpkV65iIOzRRQaxEDP17kzEFmTmKJ1poPD4OxkzGre9VaZBa5WJZ6mXkf7
GTRGBpuGxyvhLQBCFs0OUVAojySGHxAxcnACzygPhlKr7JHHYB5g+Jo4YMr225RkeIUivm7Tj/WY
YuzI+iKR3KDa3tha62lru9xySkQbV1j3dM+QZG47heXhO7eDU4vC18vnotR5g9sjdNSmsBScUEY1
i1M8TGjiXIbEBrmwwFwyl/ni4Fpies81y6zVcktP2pdr1o2PCCvT7z/Ami9elvtaqN8Zj6TYVDEM
i3PyHWLDhM1BeBTHgrtD0YOzXqcc769ETqvFCj0LN1l2fV65uNCqf81junUR060bb5v0pZQH3E/t
+IKtBC1cKKyIeHqWtc17czXIg4+9OiA2yL3eV/NZ2xcnZxKhgRwJ9ixR6RMz/adHBuZNup6VZYHv
75T6ohXxLdygb604TZ6f2BTFNNiOhbVLEcMeXG/wuGAV1/IXA6hD+z+egrhFycHpO7BZnoPlZxtW
OgiYEMw2f3fZEwqGXMSt5dmkhc6uiYqKxABXI/LyZRRJMnQex96WrxperAFjKinQpCPMJ1Gpmiy9
hJwozX44xm6hBmjMqJTeRpEyIT9aBjN5VWYsH7GRG+NklAvrAnE/t+RfAeP6ZgFy7UsLboLj876z
HIV1raRCgOOyAakq39kp2ihetiA4W7M+BceUkCZIDLOov8Qp7vsVYNXMIx6RpGavwT+35V2MZePj
OmX3VYMjnV65VXExWXEOTnPB1Nbca0P77MYi0kphCvt5fni15/5MWtCVEBMZCWkvlTrB00U+9yrt
suGZbhKtHrQDbirwa7cqfoCbCTl5DbL/qEMsbcvZa8QYgSiE1tzVaPv7Vm05yDPr4c3lYgc31pnV
xAZpvv6v7yRGi8xF4d18HgZ/S+0TQK3k2dXRVf4E03GqiyFKNg/HLzypw7498s6wjqXw84FORT6n
poXKYU5DOv4u8h7zCVmoyBur0uRH+2OWXEOUQLwHEX1C9BEfNBxfDdzooSciCfM0bu7Tw5EJ1eI9
F/m3V639THI3TYZEZvP9nZBZWriVSXlIu7WDRp3Ughrri9mJ6NVDAPRlBuxrlXW8gwQLrFMBWtPQ
WIQsfIgXVFnlM77IcyupPLUG0oXYGSPjAWj1HjqQL06lei9LNqx37un0rVLQkG7bz8yYepwMKvLN
80tIUh6KAw/h01C1WFpBMk4og3e1qCdzUrmAS1eUeiAo0pAHJJYwY200eErW+Hhd8rkehsVdH9YI
ZTxIIo1sD4dm6JvHwWcXFXTZQarb+6h7sRa4lSKIDoXbIXjqrxGhDVqI1FzjxDFVxZGTyhamRyPi
ZFntj6QbCF0HDOzybhXZ7FSGSDK9+mvvOqVP21BC2IglpvrdnrwWWiQQ9025P9UWGjXnR7Zayosq
XHIns5wWtiJxZkF/DqgUWtIG6hThxhX1CLbrGMyvWaYIDgloEJyaI7aq4xPfkk1MxnUgG0qtx3gx
x+paDC5jxd/J1McLTvyThkmqGV9AI4U68PyiMbUBjW6HmtJu/wTP/LTDx1vmZXIQDkE/kblq86d8
uoxhyMClIbRgcBXEZl6Pno4TL4z5R9ccrsP9QK2fHz6FmhOR59T0oHTGmsYuC/dkwahZ6y/D/6Qz
xWO+EwSjqRdgWZpcRu+AlK1aypodIqOx3oPL1duEK3iAV14PCMhpv2HkRNLv6D7u15d+8Le1dvJw
CzrfkO+xHL1aaL4MB3grBpWk773+EIv8KfuuE4bQPbPmISsD/pI3h9YtdW01DBRjO5UeUIdT+Yjy
oI54oAPrHMrPotjxI2+IFMJOIV7zYxWD5Zl8rYQSw4vRa0Tc+lDgIdraDbJX1APtqZCowEJx8Fxy
lbRbTCsAMqh0G2BfEx1s0KsGStdxrQreHldeaYrPiF8hx3j62oHmA+xIYD8fCzkcQfIMAt/ygedl
pMyZD7yYCNa8j2N6M1tvMmazQGuZ+wGRrOOVBifPiQKivGdXlMo3awxLxuaELGhIUktJYhDTfY7I
NDcwo+42XwTtcIX+eARxe7R4Z9CGv0NlKbOb+SNBtPhPxp6IyeACQrsGwKOvL9LOkRopuraMVYgC
gEfK5L9zAQT6OFNvkZRh31X2sIaCCjK4PNvZLbZWToSs16pQQ+ClRkjPgwPoIfy50+5DeNDpzVoL
NRQSmzOwrb9pat/XS3atLT//2G4EAe2m6cao1Oe6IZWpu5PiRUUB+yDIlvcpLYSf+KQCr6mgI4v6
phzgJinkNRRIh+TRj3YHzar+RFF6f3GzZf+boa1YnY0MX2Ld9WtQ3HbpGgJ63A+bZANj+9VUK93x
czp5ZfrK29TQr6N1HGsZFPxWJaiLIh7vhLmb2FyTwVRiIVyx9rnGtKTchz3ikw0atq8F+mxOyFTo
ODzq3q96/m77OwE3NSWdMw+FB6BvbTsPuBQOEM/IsNelsZNfThg0pwd07YgFFh93wLnrP0glRbKB
NWvtNb9pC0KsDXY16U4mPcKhILapRrqF2vhbWGvPc4+Hi+uXw1CJVDsMx8WUItmlt5HUOqTWfvst
NrB4ZZgs3rgvqHUGUeAT/1iGDi85BrXNXwtexLVlbgnWGe13Pc0WkyOd/9JLiEwur1gN6+94Uo8Q
wpsfeGkWO4HRoMhf0jxM6Xvwe5i0HSXdiJDpuvlhdAaDvd0Dg2EGBJnyW7DYvWSIfoEtse7k30Ph
ioPN/v4JbmYMpD0JAqne/VbBq7rO7BhRjCFUbxjO0xbr3HReqrHTBU/iuFF+LfTHQTxr8C9mq3Mt
hMiskjuGrDyGzdYQ8Z5NPB9bTGjgf+H62AyO9/YuIczcHn63SqULoB73OLf4wE7FDuocQJ/rptB+
Sdxeuu72eHFUx3VIew8wynNkWp61wpTfJgInhP9f//uNguA19wOoE3R3NCKWlDhLUvYEsMOAAzTb
lWSBqVjwIXRO7HgekENkIrk3Hme27E6LVX3qi9EClVQ9VSPoTYA6NX6Tw9ppWX2an5+xIdx0eoOT
W1rpDTSeuwXSbDweAejs8EH4nB0IEE56ymG6TEr2qgBBBkt9o1m+4orgjtSGesN/uOcRaoeu3ETP
GzTyN/922dRKNcEbt3660Lamx+g15oia7rpNdWWu8x/i25y1Gketzs8zptzlVlxjZxK8xyvLvgQf
4Fd510DSRoCZBDaieKtmu4YYNBpJ4SncNalAzefrx2ADlI/TFDY9pbgbTGnuhfkBb42ft1ThPWUZ
+yNwk1kLU2qoW0aSLBrgZlH4L+QQqmNWfYbuHurdGE8jCAObppapdqgy0KWrBEaaAJhNb4xOM5JS
aNmqRifowLlLUYfNI0c0qirrk5AD5/50YITVFUNYTywj4CskRormFuQTS69/QzoM1ombkl+DRHvQ
EierPIHNgBGHUJrbOKoZOlmo702ieJty1Yv4vzz5Zm8jke7tYRTfQepbcUsmAkL+YSovy50e+wj4
h0z4g1gXebU2OjTSYYO6DfTl4Vsm5j06Nt5reu6OeYCBiIN4a/gw45p1UROSTX81yG/byJZcKJ0X
yFIO+Vtrdau0Gec6icsBXRTzQ8Wq+MP+xb4zFhlMdv6w/LMoQ2TFNjL1vnop21SvNHBfkuwVPq/9
w1tIaKzZ5sO8lCTuESfwusiiWyxLn2dtHuGOUeZAHr6DICuBJ88jMuSakNlGB9ypaB6kT759Ykbg
g+LjXd6/2yYibVrCbhv7b9X4OL9ak7vGNLJgcxrB3HbugMi1YfeRhsbSxykZW2seaipr9F6a5a+0
PaPtSnVqoDZNy/1X2R+S0S7IujicW/d+llI5aYM5i+fO8xoFFZHh++kqWJlBzkB09TMG8MCuYUYA
BS7+NJbLDMlyaFbgYAKFkI3yWrErlObl1lKzQWV2Q1jRe4s6DagtFb2fVn78O04gZNSCp6OGPMCu
PMyJUcNN8fOrEyv/t4cvBlQrdU953Qmswt0IRZwoN1pbOHr6ODW3AAHEhzeNyaEF18o4uGr4lgvm
Y77hnCcBZ6rUrgJq/jErG3d+mJq1Qtg6C79HjZLMNHLG+r0FdMiapkg3RWDONRuOGDPgjjY4trz1
BQyLGkAfel/wPems+jvmG88G2HM8AIg1fbWrs4NS109rv0IGDSFxqsfqcNvW+6eQMi0hPaUzdvhV
phyH5LCCEx4KxrXqrYZWzG6FxpAgEIhHMeBLARbPQRQwBx+S2GgMgFaj5HIpNKUomOETGvVybblh
3E9S1h9BeJ0ehvWGdpNl0iLXymW8n1H7BIk9UGS/YKKH4c1RksN0D2DAJQLJfXdGjMC4brlIe1l9
0BQIslzO43+bMIAlW5P5WPlo9xVl9o/ASb14ijNYwf4zTsHWEkpcUXMZn8UKTON88uxMoedpsC1s
GlK/EkZuvl8kXLXoqCt3xp718yJLyTecKyUsP3yFrQJJtmGVHYIOxdQF7+/keC45AiE8rkLpNYfR
faiQeRRG/o0wltvURyOc7sDi/uaidVQDHyW7Uq8crT5Fnv/gONOlEqq1vI77/T79LCjTPi0P0MUk
guPKhqtc1hGhPBL/ZvReo3e/RokaQZiTAkXCcduPdcecpkS1Rff/DTrBPDaXTzZxMlXqBj36AfYv
nEkBn+dNAAQXxa4/fRH22QGyxRDVwYR5feb7dDQJvgASsXl1wZ/wOkIp7Gr97cvXB18FqtXj5Ijb
IIQgjPGRfeqBJi6/6YoH07ivmN9joG4f8CBchPEhUcIGw0Mezd0Qr2mNad4L+QJT2t36vYuRmznK
J02NK2w/i9+miBb0PNRUykeG+IlE2nMzsGnO3xBKoZ9ppU+y+UXF2Bw4XKB21P9zL9zjyMHalskz
nTJsU/+/MlbMMFZ+X4F7uws3s6htlz1jEYT6YKHi/3rW3wGrY9ooltZrlkR8pGuo6PcL3P9pRI6O
ibGaMqY/tsvd7lw8MqQbyhp6dxrys+KIhSC3VFTNtLum/0ocHuYzCE6n8Y8fQMCiU3XHYufEZThz
E9ykezxKlAZQ3DnLjUB2c97rWDqSFykO5Vc1nhFCmnjiOXIIsF4OGh4B8o1p44JP4fMtw4ipln8V
OfYJLlcaESPb4RmSzKperLSZyo9AyEmlx4cWDatnBnOEZCDctg1zKIs/oQEPFdxdOHgI4Kkruy8I
jtNI9psYR3vI7TNFWA/n/L6BZQzPvI0AZVkOv1VrXSHN+7io28YX8sr04a77WnGV+l5s4F4gSImi
TvP7XQD1VJyKEfIzoaz3ZGbKjuqFglrvykIv1fSxb4SohvjYTl7F77i+qMuwfQyB9GpoOUTgZTxc
1EswaFGTGq/g2NUl31k1qt461EWdeDD1oj9ywEWxunvnBnEoFDA5L3Rm1tnD0UsgdQU+5oGQOJLQ
UB0klp4UurQHF7YHhNLbh/otVIDaOlotykwlDsQ2OCZZU5GjVyidiaciAOw1xCohPqCDvXSq01cJ
gs7aykg3e2KcMxmVEgY668vDx2UGnz5yk8dzew5yycxF3UcfG8d7ZH4ap6FQHM62Ns7NFlo9SBP3
5TnaoKt7flvA4NK0RJk2x7nzgQDzdXC9fnAcjV2kwUG/wkBltr6AfU8LVgQvlkCjpKB5UHRfy1Wu
OwMBpG6FUYcUgaOtMH6GquBYBHpoRMmvaIkwuJbnSfLRevfr2G2FjcSjUvCkGi/p+mufRH6Va2z0
S7k6EKxjLFTSe5xIEzqO5wJRwhLEk7z6NxV/3hRsnUxNugzCQ+dSCV8XZ7Wx1ZK/MxkmWInrxx94
VluaSTgVF2M+6W4hw0VvuyO2AtnCMQ+LW9kgPCKU/kbE9bWQAUt+GY4eT1VvPPZYO9lA8GdQfQ7b
CyTQo3ymvXnJnpNRHJNG01hlvUvNluy14TQle57fJYelEjaYfAKzDB0+Uwx/9vN2Bh5VKYSYbWgD
VBJawVwh0f7op0+F0HdmK0zEOvpu/rGlYuYop9NcZrKYvs1rqlJ7plahU3MGRH/lMHtg/8C4JZv1
cqJZjxwC5CyRhrvxjwCGK0QPqQHJhspGdP70Xy/irZLI0LgrAergSY61Fq2kLis8QDbP0zNRiLu9
EYZMQABGsSqkpn/d3iOO3HH6TLLu/OqgVasd9tGvaqZFJrcsV8pes5GiLY0QrfIuhJO4BOHGssxN
GS9rlP+kQxPjwmOzkqLfSRhopCXWMYgveyltPG4g6DM0eB9MHxKO9SEBz8/VHyKtGYMYEVYw7V+w
Dza1BP3Sq31jSB8NhPMSlS8O6g6kxr/bJ+qsIV82JGVaMdHPjq/ata10ZaXfBcD8C5Ue2dKumMmC
pLO0UHxpQU4+kRdwul53+dt/KdDZg0Qz3ii9VWsUZedWccU0w4qBTfEbOtdUd7n1t87hpYTbuhjx
cAz7UK9lYeeJFXTf8RMqzydJeQL7Kvb6gOauNrjf8aCfy06MuKwf+2TmEuzEKqP6SPTaCfZ4Aeuw
wxYZms1LqsJNq36Q0eU+5jrqXY34TTX49jz61ipLUA3+Hfj0mdtsqehgO7JhEEHzU3AV5RYaftW+
rfVEwl28WB9ElsKBc34mEFGWSzZAWwQAEuFIgJ+GRPNjaUHBhGfNtG0t8ldhjk5EalXtA2twrGgQ
3C1o4zWlp5btrXx4ey+2WRqmp+Z9GXj3FuCR8oUGDuGlnOprFB7qglksqWFSs4PkPeRJzmpr9mNp
NMie81ODLLi8i58X3XUxH11E8pI8jfB0eMoXdZeRoK4huz46Iy1fcC0oXJ0j21KsdeVyLCwlqYd2
RM3SrWivkyZxlNiM9FBWrR2kH/oMmTufspCPF+2u1bDBTZGoQFpUUlPm1OVWXMai6irV++e+3NDM
eygApZZ/63SpDjDLDWTXhWPMfQttl+L5garj1sYLhFoqKa0F0Bqsi1FTOL2kyYJiByQdLoDLrNgW
IUVOLag6hjSPSOYkINreiXQwxj089AZOlP6kwYW+DNAkWOTt1Ry7fmFgmqV2OENwNOuXTu5Iq/bK
U/3fU1Xwox9S5As7gh97oaTI7lWp8lrC3JQn5ojfkI6u8lb6jYkZHlU7llVHsUj+SgF8TXJ83TQF
6nmXJlNS08DZMtdnDhp+uSyDXGn8SqbzXrQGJCBkiSy3TJaSmxraFVdL4Z7gYipzHQqTcbQTouT2
fqLtEDxvoNl05cYLF85D7JUTmCfzbDay0duoj4m4acuvYWIpuBu2H8DMmBHLAuTxwpmsVx1A1ybW
CN/PGFke/zzHrl//TrT2xcFL+scZFn/dxZS0l/pWQFk+hdamIAid754LVpboAHQjRoN9OeWfLJkK
vMO7i+Xubk/8ub0VnDpy/Bpk5yBDwGSJEXgcx2ASjFjzLewMr0YiaLj3Qj25owkqDKNIzxFupqVN
wdzw1ZlEHpmxPfuNqbkXoLba2eUoeqDXWNpZNTDKpHmWs9PpuhSo2TLkEryNTbYfx4zfBqU07iQJ
H4N960CzOKoIzDnoHvCmx6ZhdwsTpMlSfsEhfiZPY5iOcpz0WJ+elpHxDdEhzpPSgwNoWGjuTOPr
Lsop/+NdYMoKpnPoCCAmo26c+unhhiqC5eDeDte0O/vWtbgSrLfoP0NZUse/9b4xvlXJNfkmWzOq
D284pZlB4X85el2LsOjsGd6ygQIk+PQJZY1D7AVsdgD1E5Hz9Hvj6aJszD1W3lHra7vTb/3lmJDf
CUXnVmzLy/JV6dxUeFL2EYBsjf/QWYY0/AXsEDrU4acgm+2riKyORB2Lh43agNoPiqbZ4pkBXc3d
H098vza56hzgxiGZTuxANtB8zKw+FQ7lfS2m733nV972Nqenx4w5sRaOt8/OIl4qgoEixdW522vf
wRtowbr4OAkG4PxGeotyUqjeyNCK90BUiZmoNunjlOOzK2eO8Gzvc03wksIXbsUMT/cT4pc1EPOY
Ecj2d3LkJG7Mt/5zpuxulRDB9oPRcJaokvHXuTvx50L+PpBmqyUbo8CGFZuaoOD5+zaBqmYyf/0Q
ZFmTDn9qqsJVDhO7WPZAdxnIE/ns2zpbSXc0E030NTMEm7X01RBI9llgW0qZdsr5+LV+0lG4PV34
Yw+t6e3emkXYqZRzUWctsTb8jr054uTk9D1V0rC0r2ofNKUQFbx9DyHmOyFrZsq3IcuLn+DW4wpg
vio/7mJgGjxeVv3i/MHDk+aVDsPCXCd8gvUrqJGID+fckl2Z6ycH4Jgpdyq36zuZM/g0Gi2Z2ev3
wDbu3jOvOlmYZIcFEa7rVNzPDWfq5yDsAUwEyH73f7ChkdnaHMD3Bu73s4uCOPoZoqNkas8rQRsG
Zncb88uhiDp14tvZ50KeuHdbZBUWWaUgzuxrjO3qFRhn6jp7IrjE6FRX8k9Y7G0UhnQ7RaVYh5He
r63PI3MtTRDh7gpHyTgU85qEZ8zO6q9wSuMVhCyUsiq1kTdwsGCmgMtMm9Ups6RWLOdLMq/9RMxf
LnCcfo3MT5ra8LF4VqswQ8u70qBS194eL4bU+8KzpULVXvMgURBWzthuNiD53WJBoXvhr/F0HQPM
F7S3Ba6LFRdSOPJMPlR1IkMRddBBhOlsfk0rCGc6stGAnVXPzK2hj0pPjYZ3V5TNZz7iLDephf20
Txd0++Trj36uZr7GWxF0hQ2Q4+aIV+1/QuYp7MSAp1YwIhDQljfGMpiBwgZoU91nmxK9xGJNQUAY
tImN60t024Rf4OO/THE99lLTaEir7YfJ9awtJgJtIbt/dN3qW8WdQ+mbiMRqiFwOOztfgoKlkUjY
NuMlDIMIJOM1sE16EyHqjEJG/xMy+gtdlDBj0uyWLdc8SonARggR4p3e/jjcdeb1O5+VJ+5ieJfs
RdwttVLtkU0nT7Zs7oO4dTs39iEMqvqkb+xrhs9vyGlCQkZy7Mvgym5mX8mXk3ixkts9dpETNlle
SPgYK0J9gvNqPCpbDq77LL5Gb4sF2bfXCmKC6MeDfHIXC+r9QUPu/NbD7TT3aqnEhI7jG2Qyla5C
DOKr23fS7yhJTZGOdV8DLfrHDrRevqgSFTwZndavHI3Sjg0czoDEJotubIXEccSsyhMQkWllt87U
98cYfFKHNCa2HAMTI8PEs0qF4YPlzJCyH17QYpCWY/kMuaNqBWSFiRIEkI/6deQWm5QKJs0sRJOL
Qd+pIhfu4i+0upoV2DaYctoHUUGfOHUl4ZyMIw3YOX/QI+E7/b+QSvJUsu9KSzj2u/35ZQZq1ivQ
b1FNT2p4Y9vAnc//H9xNrPNMhskx9oJwUMHlBYIPiNedFnajE0/H5a944ClSV9qDBdX3yM6z+QWW
LStJ+qUe5QSY3ktAy/BpDVp4EGv9eKkrx/RyjNGYk43ULVQeXKzEahywNmWnwkjkeBBzrtgHYOYc
A88ZjpZzLyOCVrcYzsJTn9iD0I11hahmokGc0sbiBXGYqD5TLHOTBo7klHFD+u07lKXvfJ2HikuP
Ss7jKvoaQ9enrIoao9Dk4MNLuXlopEvnsBsgNTNwqq7RZGtoCYgrkpAo9WbvnDKMwGRQTNmZ7Kj7
ciRQluTBYOZS047UuJqaWuG60/w6PrHKrjwxhvZo+VCGGrWetBDn2UscO7ihX0TThEbN1epvA2h8
5Zw5LOw9qh1Okffu6tn0clc68DxQK/QyXSsLDLDSLHO5Mb07Zes78MhF6ImRLUcscyr4BO7N/f3H
nEZDCIUk+sc0BlDogmWvtwfItOoQhmLVb8FEdIiFyeu81bTJvjSPYVuwtbC7VI1HydVgKD6hQqKR
o3wTvMfbojjpVQDJs08xcRROtayLBRJ9Ij/9TfzAK0pHZYYYehrg2px5PqOeJuMkAswaljAa0PjW
6JRQruN6ThgZQJ6YOjOPcDQCARcVwXBW6r40TeOQHzDxj61VxeXQZvR4rVqRRLZgo5pVTF5zkKVm
t6O2AAjlv1905497OHSMi829aa3N5KLH53z2E63oO35pjUwx6P7cut7ZMqEHzhhk2iBOdYfbQ/a8
Ol32xucN/Qa3Y1hdclVrFZwLbhYvNPhZ9uSPTbN4FmaT//wsGfoHSy/iCVZJPbh52bwSa1VawiBY
2M8teHAM7ACqTTfvqvBv/j+fj5DV5diBUZJIpGnDPiLlC6s/Tov2nr5MV1KY+Wf4dPrmYILXIIyJ
wOyBiW+o/BWi5GWyxZRR3KGXXMP4uiR/9bYUWNWv7r5Ygaf02VSkLzBiawcRJBLO5WL+uv/f/HzQ
ak7DMmPfBsRvRI+DncCwj8CsLLonNefDMu6IuHXcH3IhWhNR3g7bYlOoslYRqp76CMFpHVV6soub
yd09tiPaCtBj4IBO1+NpOoCS2+E1xbn2E8b7apDy14bduVxqLwF824akT8+1b4BjgDjZUmxQUx2+
0GusWlkH6HFEp0xbjtZ+d6e0pPk24LCI+nZberEc5c6A9OtNIbHuAFZxVvVDhJCRox0RWJ/2/PN7
sAlkt0MvmTKdZn5bwI3ayWvVEfVTqiS4z3FbyYyVw5+4pglQynr/63rwNCfzL+GhFPGIU2ALepRf
x8T6fBc5/ovwSySeRy3i0UgcwG1Op8fBMOhiRUinHRA0/HZcP2VOGtknvfulMfCfxHVytZXmTXxL
4HrZ4J1+bmFXE1va81I2XY1Vy3VzGhAFsb5AIgyfc6F6JzhLRGPPaiD9kYrM1IYE8b5IqjUzrvr+
vpZkP3v+CJQyzaRnyVODZ5tcElIvseQgK5dC1wqWJl3Oz4rLmr4RphBY1Q5PBynt9s4LQskPwUKv
rQY1InpEmKO8F4Btd4G6vG4c/rXrBqVm+74jvsH7vc2QtEUYcMM0TVzK5o3RbIsMYgLckgrfjype
iywK8FjfqlYRMxR1wIiNE0JPZ6oDmMRzvLWHlkZQTwWayGlVptXAUxhMdKy6zc/BoAsuj7uDHyeC
LSA7vofYmISTwfZMqJ1bhdgOhoaEyp6vptM5562wMhtXec4HcU4WVkhjxCezfb3VKH/FA6M8cn/w
iS/1WzWNJ6UZdyyyPf016r6drS+SKAVRPE+nUPMuA+1XFGEOLL88LMGN82za17wbyg/lSm3WiPt2
M9EW7WR18TuDVjv7hiyZUYuQ4lq5b4mRdLiB7okUuEuj5t0VJAUhAVKRMz/EKCzfPTSyiLuDZHhk
a2vAOo+FPhOLI4eNYspKBGCrHZxiwG552VPOAgtmSEa3jT9kfWadnWgAkGvag1Vc7DK46R0kbBXk
Aul3lBsxCFv62pw15a62ww8GOvLsyKvFe3taCNPVmUtfF2UCz1+JuTd0JISK6ujUlLDaf2WwGTt3
0fFe7WTKo0uAkyjDpFCdeINwBs9fKVeqw75u3ewAuF+U0KAHGfy2eZGtEsEc1opk2ebapBU8A8DS
Vu4eX98N4xaRg0pkocx2V+mZRG7gq1LQRgX54mwZzPyKABBDSF5N8pqlpCMmCD+mu4x2ZYCnE67c
sLMjHaxDz1of+VvEabn5/LWSBdil2dfrJ0ygiYMhoE5HscDUpv8JeIUufNEuasekUEsrB7gjp7j9
LT349MuE+F34Mz+sJ8LMCIgVuKAXh2RLnAVBGAwO5eRNc6Rcnu06Mq3BtCGIDTCYIeYh7p4ro+lq
vXkRgS7ojaxl+Fcj60IzNZbnvueK9LEN3/Tz8toMcoIck/yjyUdOa13eCLWnThU9XWkUcN9EnTYm
c7BNMpg70TsNvzSOrKDgoQMKLzeIydwm+/LRhak/N+JFPZyT6q6Lflv3Aoxr8z5/46DYp0tbWPD1
DBA3egLgapE6qo/deS8MY1BOAzcuiRJlAoqyTI2JUd2mcVu4WOIaZU1BQ6sSe6gm0xJjPL+HLM8x
btRHF+7dpQTugzrEa5RRIKBYfvbI/3kTP2M+u/CAm+ipFLuSjGIAOfuLk4Gy/JopkDUvgzqTyFGD
wXfPNDIxgH9Vl5f29+ttj+/0kCdonYunSfL7EeDLbCE7VuZOIpBy3nbZOZdQEud3gA1Z2A45yRL0
GTpeLWLxjKzOvH3VnS9/yI828dRHc/qyYs6MqwMjuIGJdV6c81hVwHT6FSSmlEOSwS2lPckoJGXk
/VMHelNRvC8sOrJX5RkuBCedAwFz3FGNR6xeC3ipc2J01pIEOJ6xE4yZs9AmkO9KWOGj0HKTEYNi
ODkH6qkqlTg0DX0/MnOXdJKp1xGmeEMjtHTKFEmLdyTCWMFtOi1puZlo7dxvksYzJMIDIaRMb1Fd
w6eebkYvKsyjHYBohhqzKC5rX0m7hV2qEl/IIVk6XOdvG3RhIRjDyova19eNx/nh39HenefBtm15
dDwZmWE3Mln3SMuNxvPU/cyfZON7kfou5UZil8pCDAFc//msOxQAYOZXsaZFQoMyjMwPFBkDIIS6
irNqNMIFCYfpSAEv6pkfNMao9LBYWP7b1SZnkJeu4Vrk95hfMfAuxtjqlVgo1griy1JjnxoaMMzX
lM6J26gff4uFC+uEHP4Y/hmK0fPJ4BjnmT3yPK/+dteQbqQoUNRkC9NLcXrVIWStgmbnGdvATQDm
oInOGp9XXDtqYbQLKCPcYa5GLROSiXywoGaEQMyf+wiBuGQid2ERvfFvJubu2XbofTH1jbIEM8Gx
QaqakZa+caTt62tJYys5HrMrk+BIuFdC0EXP+hHCzOK3Ai4R/SSIFX8wIqUTJIf6p5Au+NltujZI
phOL9IVVhi+1qjNpr/0TKI8tLRINS4xe4FSJgXAkMEAacEDAIEBiGgvG0gw+cQYD9T0kNr8FA67M
z4NWy/sJ12bdm4WgUUr9LH+aT5EgwKDBeoUsBSUhh5kcqpREaLXh9Mk4XXXirPhY+RYj4SUOQU4B
fGmSJRYOMC2eKhBDYR6k3FSL1QsA3pak431CLiwWcJwvegn7DPQPU5Ky7mAyns5xpwr9FvkJiFQE
8nSXQTIvtB2kN153QpI96yZYqx3HILdXyYlWlAdmAyxDSLYbu9briBpvFQF/jjOwYdN6fQhaa2TA
yHV6mHpe4Z9T1U8DaTWrMMlZVMEtohTZn+cWxei7dzpI2W0221HUW/VrZsvDP7hCOgZQ58krEmjc
3Q+6D8cuUaNfz6xj0nGIkHsTt9JZP7VmKDqlyNGlVUY0rt+TxuTfyJWbBwpb+wKTLdElL4B01yUm
seZkt3VuciSeytR7+150rfFwb8BeKVJEz3pwaSRXtwUL9E0SyDm7eeK7auTv4xwB4pHDX9V/Knn+
8uX/xgmBfE/EOZYvq9TtER4QOutI6NwVYISIbbVBwSYmaaNCb6lwxvLHXQ2Xh9FtSb84z9Jl82Wm
LKo2SMSAmdOJi+sjdApIO670eZaMaqQLYQk/4+jaLTAfM1yqGJmzvENSmVYSd7WJDABcE3O6/d7x
45P9VGAlIm0S4bLXIybKVDoVTaLynNNHiO5hdWm4ECTcDEpTFzF3JijXg4MTKEPpNpGnFQfY2ngB
AdRUwU+m6nnyQZfrlk8RcN+pSxC7u8Mh7FHukguG3j6ZYOFEHDNkRrOScE3L0qMjz0WqaZKAbtz8
oPAOxkwhbe6dRKUVcYoZyFP8/kgaheec5Xo2HZ3gnQDvRx4VmgG4v43m1hVUNeJP55AFRJ/LrzIv
plk3zQNqp/iZ8YrQc8oXsuZlx5V2JXi5QybBN/IILH905XaNTWQXgveSj2+03l9aH/rJ9vCwCa5+
gO8WNYks0bgFmY1be102EWOMXnqDo/jUAx2U6hckq2DMaYT8a0hEXhX0A/vke5xBjbWQz0wDmlvM
CkWL9P6Ep4ldV7PnAvKY/2gZQidhcF2wzRJIRk2l+5tB+KLITQ988NTJGnBrmBthSh9hDkhZo8ba
/MAeTpVCvjvuAf0lGyfHWuz1kbU1S4ZpAkx9IG3OZzb3SMLgFbbqj+Ely0SEu6SuO6cUrIO1UOEW
mREEMxIkz0LSr+vXGoPYIVc2CNUu43XBT1VnZRK77UznLBsalSSXPUI7YvmYLrLe/rXdZQYnAdS7
Ufo50aKCj76vVWXbyFAfECs6HzRu3RIgOgkp8XQd9fuoFU02eENP3qy3dvMJ7+9r6pi9hk5lMqMk
i41VSAl/HTmdXOgOWgSEo73YPbjMUDxLgb63+M56yHZKfPSDxr4a7flXaPjs/u/nB6mhTJkKj745
pi+zCHUO6+DYECmNftyP9Nh0kDeo1xYwi6zTE+Ax1g7xuamH8kRYUYBxwX8jH6rIxDMFwX+h5odQ
cjFqVsrAdq1rO8/Eca9W9V2XgTapwQ3QUtebJUlFIYlLaUsuKBI7+jHDSvXofFYSZCiMUJSjePvr
lN1w3ICymlWZfigKqI1mZTh70ALzGUTvyyrLuEUdubMfEMLApiN3rYq7pJmNy1+oyx+ZBB4SqYmC
NAUeeX4Si3wyEKBfZaKK0YG43Ew/NZj4SVWScsF5JgN++qvLXrQrK+sM5ofLquKXl0ogrweUYxpn
TbnFzu8qXrI45cKqx64gY7pZHUbkRtbs4W4YWjtNPj/8zK4bwH2HxBOZcSC0CnKNdIq2XYG0y4vc
NO5cSYHZ/Prj5EHP9Es3/C9hA7itB/490AqjRDtv0jpow3SdhevcmmgMOnQOLTmO1wybcmTo/oWN
YQ1xbwWguBrB5YF8YeKHDuPKOicF4itDx7AVPPeebI7IG+3pUMP0ehoL0V6RiofZZqqUlwgnHszH
1RE5Stsx+UyT8pQc26RjsxOSFMnOLlnrVHRYdz+2ZoK0TkN5Dp2aEL3MEMzFrjZONoJvHSJYTrT7
IsDpgj7Dlz1YNDsMvJvymG+CdyycOCCfYJysel59FapZuZi6IcPhryk9u9Dc+wA5CzteBLukUOfs
W+2/twXWHNfq3Tx1smGtNEhHDiKOJdR2c1Q5pWXZ0661GlMEb2aiA0qrpJA7wpsQcz7ciAkyRGuN
Sj1SexiZBTfy+gdMEVLZPl7mKa+NkPNkFAjK74/AaFMvVTf9VJFC+zu8ReKC4HLDOCjmI6GbIqqc
TmZcaoKpVtAN2qhwd6QFbU8FeY8dfV6hcb980jzTKt5dZedbZCbbH5KwI7phv5ecEIPpP3uPULl7
+ij40T+qRhKlI2Mk4y8nz+dJ66N5IPGILzPNX2NJjToi6lLWL8BhSuCguxCdOsz/ZZ3cXk/aqZy5
BrzxIA6HwBOTTS66D7h/H8YQuuOCJQyNG58WXP20KtZHrEA7iGSJ4pRlp0/+DPCvXxR4C8X/+hop
qsmeBOd/JURb0EMDfD22DSxcbD5pI47jTD0Oy/PJtQV84GpcaSZnyP8fbWjvIiqC+Nhz4egnQvby
i71iChN3s2jqNWzFJpIfrDxH1SSCUGzOa/zM78K+e1DXbiegZRrwDyqaOhyqimlpy1WqQmn6SwbT
47uqzjku8jgYqaN8HigC5Gb5KrFesuNaDB10LUBvBiMpphbw+zkEw4gAVgo5a187EG12oD1uf3CG
H020xoQfS33Yo8LYxN5rlKE/KGMelo9b588EkT70qekSKyLf0JF4UkDDVWxyQSYKsbvKSUjobjCz
OpxDEnx+6NJUVjKTpq80eJ6+ALAMd4Lt6DgwutRR/H3BqMiQG9huPp+B9gRQsd5FFILTK0QN3LgN
s/eyZPCXJGfYQEAfd7VMA/LsOJCuQrnCfa7fvIvBG7wbfmWT+uFnj3wVbGOYq0Dk3SAEc5YAG+m5
pxQS+JERMeyHiyW+BTvHSLqT/qLuael2on7s91QevZuQpaLj/QwDTVsFuElXwBfHo70GVGk8Q+3M
j5kUb/R6vVLF7pDe9Ne5Ri6KR38URcdfOfxA7NHzxERH6AFZatS8Uextjlp8mN09UYGif3mdOGb2
8D1MMMIod07Pvznd1HfmoaD28WF0B6GCq6/5BNapXYH/N9+BHOTPRRQvpKXzJUb5+ta+jp5D7O+C
QeO/7Nh+xk0Kl3orSpocPKFHO6+ORKsxNtoQO8xuT25DhvRGyLpVvJeKUDS+0TPK73uhyw+uOjc+
bMp51GwZDkqv/5WqknPACQdrVlwLoYqnWTdlOnuqlmdPWVZ4vdmTF6v9ALlLQd27VI/ASIHUk1Qy
t1C8g5Gb4kfJtSpFg9j/QoUdatrxBbO/qYpzkBNFSwvLApLwPqzlzmGDJG+YIV992+opdHDcfe3E
8Xlvz6IlgRaPKsvbWRDS72jKSc2/2z2+EZB9UbbsIq3PFxZQ9aPqrCfZYxJpn2aY+dlHYZL0rO4C
S78D+Iyf2wwLU0pqzuy3+ORoCdIQe1j/ah4zwkuIViC49LUHc752KooqIrUDYqjXKcCkbE1xzCwN
YmO1dvEy5Whvc02n27bWrbqdJXrepa4FguRmUMCKesp1/UPIpGfBtGyDpIcbwdwvdZx5+FEkAush
qSm0V3Bm1r5g1oPuukyWxilTWMWatAgqsfr/KHU5o6giArpRMHT5gHHy5edPMiVwmSGkkaeK8u4Y
NKc6RftPvKn0wddHAIyspS95J+XqFIqqg8ZB8nwRnsd6rCJuNnC8yB5A4B51jIVdKgXU+zzovOKc
OTgNe3qgWPva07ojqSnUudJTScGBcwH6BlxsIlMUpxs3QWROywwprbzRQn/ylWIsIwRvGcruyq8z
FXJ4nMCSSbQvpr18pgNKMNfKPLsr4gLUJcFxBkIMa8nfu3XevO6fpDr9sVzROgfjLxrU8hhxBLnd
FcLXRuoPrjxg9QyIqu8urXPW5Tiawh3BT8lnin4xUWwPAh6I9jHA1HYdXeM6y96Y1wuctSYOvC2A
h93U0oUEO3+q3RMuzcVLwgRn4z9sjrD8AI9TGAkd2KOPar0BLyzseFvo8OAIv8QVMztY9M9tS80n
vENf0y0tyLtznhd3hS/xaU4jvpTQu9QOO0QeLqLv58OW5VEGd/kjl+qhOOdzQG5RMPCxFqBzWyT9
gxqCc5QBRf79WeRes+acM8JsFHH/oNenW4NWhX49bGcPzK8ymUQ89CapuqQ+prDJwhd59PNORFys
pBCMp86pP+3Tm4q+hnIcWXtxdE528LEXGcd4sGyaKpllInSWy7H/9D5/aypfBe9NwtzIEqCnX/MN
UdDo91MSpQzVVF6YVvFX1ih9eSrVzgjC2JJMmSZu66pFUR0ZtXb58gQBHMFF4tuFB2KS2DpSZAKV
3LiOX5xZc4O4gmjYKi0F5fck9TfWn05vpLgDjdTOaZze406ltfd/aYLTooZIU0g9U7g0InqweE87
cj9/oWSGigBAN0gcRRRl7dJyc4CTLsivWCoL+koSNxw1+D9mOCrZGNha2tzHin2v/AIk28+aE8ni
v2t4r8v7gTqBHTCjxXOkfCvcA+EByBWW0O4K6N6l6FiDjCaweuDiPeT9KHknzqw3whEfLkjT1QbZ
HhTBZ82tCotm5LNI2AdILlFloT2aIiSDOHaT1niKaafYy8mdGi7E9xCNTM9D3ZBbKjUuYkvM83fb
j991b1YYPsjSypiARDnl+rHprVqEzZBUck5kT1SJ/MopLuG4w0Q0YUZ5ZVt5Wg99lxmNga7s5iW5
7h3cxVK3wWpsltctX7PkESE4OViyae1XdMv/FIkpbauplfWtZHPdD0r8YhLybfdwuPEHJWnuMiLt
FyDszaJAnPBnQHJFqpFN63olPxCb4Ul6HUui0VriI7fyAj/TLDZqFnYfMXXeSuY/rtNfiiuvMhEH
aus+Xk9ejSgK2kO02usRY9ZhdfuWtn2mG6HGRin3vRzGXHQKmQY8jrdyZQHHiGdk64aNFrr6G5Vy
uZfX4qt/a93i5/7q2HvWGSxioxkE9s+tsxfY9nGFSAT4C1SQkuaoijdfcZ4BMMJOY0qB0E7RaWTp
gzjK/AU+iEq2LulVcp/fbAqvi1sy4h7JgH8LZvjsQr/vMJ3LXcCv6fKOe6ZGTf4mpPEcUShsKDjG
132bE5vPLyz8RKlmFnXxnNVB0nbmN9EP08vmOWYtfFkmBgZbE5Dc2kyeEDl7anH4n/EtqjKhU2Bj
tbbqN/HJ1MRcLxbX48nFYR3IYWwmHsB+TZpd+SrTQ/9IRxWIPX0wnkakTWC/b6c62sh5N7onjKOu
w0J52otnoZUg1Q+OXATWUdldwlpkyHE83Zj2VUdDJv/qwc7RIoczml+vCNqiSKeCAN7kq4oqYRW6
1JxLtqnyBrTkMw158xWhtHdUQpBRjNyh07RhZZDM9B5e4XQCV4k5GNDVhuOLJk9aW4sW8CpafDqE
m5yvZh64wPbBF299KUncYBRMZDZaLZJTxFD6wbXQtkyH6ChaUc+7/B0QXv0gYbsD7UvYqZLQtZe0
80dVjhZti+ThmVFzGbiFs2cca+AnwyaMafS3xUZTN2R790dxog1ROfoCnrKYJFWDVuV9EYU5eKGc
QFJ/64jc7JsOs8FUpCQwEfs9HyFwjGEMGVA6diEPC3NJg2qGk+ffJEG9we51YECfxb9TYOQODz+2
Ooyf2Pdk3BYUY8bg0vZAOKOLDM8f9jWv/qgE2Myb4yEAeu8Cs9d5aPwrAMwdFwS8imbQFCLB2F6j
pFxi5kqs8f3+wOLmJ1RGUTOnqCmJV5tDnMXHKZmaI9pYQoEb5Pf6npx6evr7HYVyl3U8WurprWgh
jeFrzz95sB3urE+uoEmuqXO4N8Fizx1o89De12uI6IPRY9xeaztt98OkUDc2PksfCZ9rs6QAWlj1
n+2V1tEBW2o1XXmWVGTNiF+d0HyNQStrF7t96EiM3Fosgu+HJDYNilKbIqk1GMFfouMxNFZ7GzAS
7CmJ0XhVWnRkn4aWKlP/NV9+4wesaSDH3VPL97x3NKiczivbtV0fzSFcmaHetaW4drHDKzvfCyUg
h3kHoYskukWy6o0U++SxahGaqA6c91fXV+tfV4U/UFhJxO6Fa0uUK+qUYq3ZLRWT9FQb3F5Kj0UQ
jzmRqCl5MQtk+t0z4oLT9BrN2HsZLDZJkFqFogHxV6XzyuuEbyb8+3r5OEMwItDmvcahNh8MQvpQ
Iykmdg+CQ14b66J4VIvjck84hL7vm20hfjcbR1mwwlVbPmyr+SMIMbIYqxfp8z+uPl4PJIxXtNcA
2Xbwxtf5UbaD8j3PdpBeNsf4rjP2rdm5KukdLhq+004c//HR00LT7bnJenrJEl4JcNFWLhV38psF
MgXsAih53K0WjJIXgeFSSC1klkCzTe75TiqfC7KztlP1T73au6dw88LMO9fr4ZtBAZAW/IlhjRU/
Ogr8mezhbc6SmtHNvbCfh4yPXrNZ9f8aDOIZEDbXJF0tdI1sHR6ET5UaWvzMH8quGP9FYBhCCc4a
xxVtI14xvkZzX+WFuqhMCFirLWRZOAv891SI/0wlvHdoocfpgqNIZNlvaOXtBcupKuGhL0YVhflQ
3j2c6ETf5GuYs6Zg6yzoPl7yrTc0pVvv/ewaRq7fwqOxag3xvkHnKR3JONXBxrdWM+UuYc1Nr75y
4Jb2MZhUlheuula378OVCBm8XBbwYBCc911wwLsxqzoT3Piz/7ZQhsuutEbVPcceJV0tI1DJrXy7
P4MVcKcWTLImr6Gty/9wI6cbqWqQYvtmdD3sdjTh815cNJzzHpeX7+HnVdAMmS+9Luhtu9kn+WzX
36g2E4ZlAnj337ZIjTzLO4/Xa9qLkYZ3JqwdLNWYQoK6k+UWxJOyM3YqCLqIo6lh03T14uozkoMn
LM4GBquxaroazHbphtfmOD1gYqwGnPNZwrEa/XcFzywE3l86uSnV9Xg6vV6KD1FOJKOEqCgeabTm
RkhUwX4W5edYxIk6NKRCrEG4d7TEnSKRFthiNWQMtyP96Ldf134Fk6oaLF6yZiLXSsWaVLWFQiMx
Ah20HXC5ZluaMV1JLq1FoCyrIEpBJx0dThA9EVRgTX/jieTWy6aN1Kt6cRm2iCt+Qu9cdEUP3nhh
J1lo2lXsl06euvMZCq6csBRwX9ERwZNHPVVm5RgjE6isNyU9ZW9xT56+ZWdL072Hj//jZmcoPR7R
E5ZwrktTyA3jHv+Kp5ZXKbwCEypflHHVAUAbvAV4HBnI/cg3TFX7M5YVQR/Qpt/qt31FrScamGXn
TixR9DQHpcbDC2Jx9jK6ANrA+chXat9HXOAXarP4gz0FYW/5NUbniZl9giGchnFnl5DKECH/JaaD
RFd6v29ADi+DhVmvMDMODjQtyHdOX0nT0bz8B1y4lk9olb8fy96k2BpXW2qlxDxTbL0Za/imXFSZ
D9C9C5qLmntqm8flPdrvkn9GtlAtO9F1iY5m6YPcXBgPtXAu040mLaaiDOPVxmzv7Y3geeEBJdCL
hEwq77Cg45JrK7eW/B2e/zYrGGwaLHU+c6799DElObrcLJn52/VYmyzn4zhLe9qCx3R/MaVPM17l
Fm9iRBlRt7/lTW8BJHIISbxJ1Azvaro8aGFq/pTQd+L/a3m/6Q5gq66CbzS6yZ2qpMHBpRpESQ6v
od2HMpsXWdTUyxSTC5us6hJwI668D2x+iiYfQBeVfg++mCqdCEBnThH/bOHBi4wK+uXt9fBKA6R/
9AozXPtTG8YGZ16keIO8/oP8Kr4NKImA6TsERojkUD+XEeosFxPGT8D4ixvGRnbunloA3ewum8FB
91xMSPd9sPgCJ1Km0BDn29Tl+4fE4MVBbClR/WdkPxtLLTYj5kO+dcNkVAA4tcCbUB/h3WegU4YR
uEneKuJUPEDDLawLh884u6CNXthCeC4fwDSzA4jlY1rvneFSUcocb09UKy26MjbjXLETFETV1alp
yPos7SkbdFIrQ0XJcV5f+9fDXNDcHV96wk0DRj6zR94q62nD7DMbkyEfnKktbTQzmZ3+CvUClPIL
IPAgLyZmavIqBQ/SKnb8cc8crAvhcHws5UF4pGh+l6t+om1XsSCL5d+wnczCnwvTn8z+mD3cw3fo
FUcb/Se7YqiWuMNFfAdyKKqBJVLWBXWNG1XiuBN2vw/jcvMfUvVepCRq9BDD3Q1SMEIXpzmWir0L
tYR5dmmh+vNWLUSB8/69Qcx6gFVvUe3rMaQjwSk18hZi4hjdRcn8NYw6T+Mw1C4cUyDBLRPtcuMP
WTWm/55lYdROFWTle7um5VIUTpHWV/qRR3u2qYzBtfUdMgniw9D1Mh4lemggkXvoSJawe20yzFsU
Eo7MvMbb8i4MEOj8dGBER3Pi85lrIV5wA0+8R9C+qoCVyQiLCgOqbSsuaWLzMTFzSR5dxrDAV1AM
lGRyGnI4VvdNwXHjzqbYmdZ/Y73NcxVyiuhgzrmBCswJFWGIjPq2mIrqUfGBx2SCRbfwynOWd7q8
Fg4ejQQHKiYeS+uBbRbAeKLH+2YIuLKcJWj9dTuq6Ichq5nUW0dz1c11edWa/HtLbQXrPjhx732L
WkHjbu4E2cfiswxiLTF4cAA7ACAulDyp8M+24OY9SwzyDv19mGUTbx4i+R0VJYr5Nnx3GW7JJn9g
ygVJB1euJ5qCwpJMh1HsmT4JwdUQ6SA/ZDg52udG8+X0yZqPHXgU1yy9pgmipqX81A5Pu/U393MW
Qnw9g2wA4jpwjxwZWY9KVM3CkYLgST61PEnuS7fnFSG9Qf2nG7tyQ+5KCFUvapirqcj3UDUDmNr/
YmMRhcclUYToOnAJhYDZjM3+VpRzU4RwlhwpNKjU28JM+E7mhWn6BAMLmhY/Xmp8lsaQTHRmqk/j
b0AeS2m61Yn9ulN3yf0XinNCsSc1xcWvMNvYEkIzIFhwsUn/1yMIhKwynZF/UtMHmjSGHGZkc5KE
gB2vTaz6jd0Aa0ZkhoEQW0n2iOkU3mTHChS7xzCADVebh12wlEznBLFsWZfbZSeJteLUbThbgkQT
vIjDPYSozqmXAo0Nj6tzzz3LEcypRSJIkI4EbMNDFSuTO+fRUH4b1SMQFSO/TKVpnJHwNJhHR0Vz
sFp3omqcuDixAwOqtARNIPGYmjvhfyzNe9qHgCUViSOcw8RAmID2JUPKZMoDSeMhMAJEs8jYIVWo
1hWTO5w36wFhWRu8jfCCs9tij0PuPlWBplK0ZwfjM3nNYTW537Ogz9Hm6Et7ax5i+yr6pzZ/STFv
rsNyXXZrIqhxSpA07G9Q+EqLzv+CbO0tiMjU8C0x15tAx7b1OhqHBXGoXrlp+bxgV3/2uHQABnb4
iqJjcgU1t5iSMkiAo+ElbE89T952zC9cDL2htR8jigGkB1cpaMdQaeiqjXI/XNtrmxccE1zqMmR9
evMu2q7UP5DPhitkNWZNqVyhy+B3ctzkOWFej64hXnxbqYdzvE8n9pBlb8WAjKgooJVLOmJt/q6L
w7X8o/Q9RupvbUt90sVV8PDm9BmEbBlO6LAffVD/JZmKE1CdfO5en1gztetsFHBTm9fS1Ohv5cm5
XVKw/c2hWKfMW6FvWJxKBx8Nsf3zF23xOgTXjvh1lwdy93Wrk7Dj9sNP2c9xiL2102oeV/1lgb4i
u4eyqAMbjVBtBTCf53BGNDJc/Rw77MN4kF+xse55s5PAES/MdT+AnvTCPcR4BwHIK6B21QHc3MFN
xwMrphJ+ooRibsjA1zlUfHrFQGjQt6fSXcqaXnAxLZMXgAO8ObEZmoXDJf99RQ0hKbFZZQIWaWPN
AUWap0HfY1wn1nvNDIPHqYlP4hETMXMfLXVee/sqzkyqMzdYgKLr0ujFSBmJqHDytMcO4j6eQk4Y
+7JqnI7Twxe5ptKSzv/h8Y6ig4J0JUjBdO1zhO8hPi/4B94/LdIpLpkpMxT01tEHZAFjA0ZXqyXr
cmMEi8yj9OIJxmHaoXgAr9wSnFU0nKIpuSUr9LjooLMJw45135U3TDGuCMbzbf3F1wjAUw+w2e+0
eIfCEvZlptKgjLMJkBYKIq5HHXbv61dQ+OqvscN51vYtFppyIWKjx5UwEaJgG694zizBb/lGNCaZ
7kiUXPVjxu/KLBe5CKEFhAvH6b2geqgUsV9vsFMJuVdLCWVMNXU1GWuUguJR8B9XjXIQzhlI+sZD
FTrb5g3uojX8yNlfwcH3iC45rn/i4B/399d3lrmyFP2KeXdrsURebDtokrpvAdTJ8SvAlFk4sDIb
QaOg+co2/7BGMZhiXRa6fFVpWvOGQ2JJtJ6Y7bRAYXNyy1gqvdZEKKcxuN9Gw70dtT0dkFwebHEO
dhW+rON3YlOpqSoT2NrjQiWw3TFA6EdqjqxBsNJ2GjxBbQk/IUvItbO71KXwigGqwmORa31XbffW
hc/m08HTsaHMHCR3OC3jmj6uGQUTdl2sKolo2jay5+/vpxZlkTnNo/zZfghBHXhTYRzFk6gKEHVS
tMqQlWFHWOESTDWKG8kYCI8zQdj4RV/+p3ubngK1Ht9lMDZwgaenIROf+3l/hu0zRHxOIY3dTBX5
qk4tQKV9X7Nwq9jpgoiMZQvP9lxzLjx/gyJbgzg7Av+xwnGuF4wODDheUSaFEBlzyvXwDEFChM8B
cR49Qxat1+wDgyzChPWSqGmkAL9HSbrHJxOWIMlJRnQcurBkVIYp0Em1xhmZWIKcWRLHgUuZeQxL
mqZjeAZBdT1y93pZzNv0ucFU4VYSzpeIledKxRSSeLAoeTStKuLAisc6jZQc92vz/oAB9MXaofIw
tnY1OqOTCKDQqX5uEnEDprApzB8d6PM5KuP/AWNN8KqwR5qDC1KwVHUEJcm8PZZKh14/Q0YnFE92
Rx1zfzLeH95CTULNQjoXdcSsYk5FeuBiADv214fEhedU9BrbbXmnjPbrCVLGVBDeXjqj8b78z/eY
SDEgDYTyTP2viYzw1K71a4sh0QX9gPDGBa06Xzgh6U8k9+qr/Cc5EfWfzBW+c63sP/WLMk6atMYD
GOOqF7Eoue5maVOKS+kp/SosqF6pb1MNXF/052cdA7oa9ek/Uxosf4hKNSQhaPytF/+bdn86vHds
VxXVG+rPezUHyiT19KzgfBsT7n1GImCnlj31orHWcXk6S4QjfkiwqrQbBMJMSJ2uacwPWaN9VrWG
xZDo1vRqM7V4l4R9xOdryfQZW66NwB5sB7GSB8rffjKpLrKY/k7JSBUxUaoTXbM1VqlQ0v0kmoMW
KpOC0VYeZNTfSNZ6b5aJXqdZtsYRnIg/7thIG6gIQ2NW51WgYhsHrOStNpZBub113+/cTt+eEXYK
4LEumytUaj2grLC6Cy5dWdIHpguRdevWRNSkOH9/M3scDMs8dRYpjcq3rgc7XFF1kJbMlBz5lFyw
Cc2wH1KBsDFlRpbq1yLvoddU6Ut4xuQlxfA077Md2f2qH390qttAHEaBRydPcdAQYq4i2grXk+44
K6OWKTRvCwukE0RxG3roWpyDDfYUQC/rlvdwSQdh/NZa+a4L6YMmgHsUSqOnvaFgtP7TQONXOvKo
2wsMbTdgSYjWdQ/d5zkFHu54j4XNoHr7nAMtjUPGBq9PWJd4OEGZyAqt4k9hx67nPb/1uXIaJpT4
Wt4E6knMnOcjJCxueV3/lGlJzHbr+dKHt40RAl9M+B8hgG/Uq4WpFIzKIwCLty5bo2hJZG4cbUxD
0sasBrFEwW63gLeicQIPaby5v1J9Nx3E2WW9QoRK2sNIQuht1UtdpZhJJ0XpBIBJ4/L8q49hM6mv
dYkpOJNxdoOSqNLTHqTc+h/Zszon8i02jS/o/gYGNyEZ1qQwFXriEugPg8XXgUZ0gyr9TTCT2Puo
CAPk/Gx1JYZn8JHISFbgMsTBPMuWSeRaYmaaKFtmvJm+Eyy0HAH+AzU+5NFHb3/gogJh9ARQCM4l
lRd+Uo7X8B4GmK7YxKbkQ4IDAtMQ+7FpD8cqhTItoQYxMbPLd+gvF1KVd3se8mfYW+vG9O5iu7Vf
Hx1lLXHyxBAnSubNhYrDLSriE96ETrtkMa1GeyfWeuj+r0vKwe+crqaaZGQMKKQxV6cvJYtjinP0
tN9XvKI+ijMgmMpuzXvi+++YqrGG8I3MiPuGeUo8CAtRbu2Kb4N2/Kw/NvUEx+WgerTm+AbwmdHK
ZvPGsPEYDyAU72jBaNxCP2JD9hjbKB68Omczcnc3mh/OZ51+uc+gdjsz79pELEl6c8vMaaDdrLqi
gZ92ZX12SaB0nMzFwcok81eAdpXx4rS+YrPFpRCswPHOPBncJLfEP2D5PP890rFzWTK9rGjCFXlr
m27zgDjcOPftCKSIpgVA77aPhKxT1w9jylQSOvF8Cb1F7cDYipRg+rIAXUabjANZ0zInlBUp7YAE
+mEC1JzgRKVTbSv5/XPng2dPsdoyVe/TQ6Tax/yRLINRJgkfJzwqn2UuERyqkD6H2lVhDKKNw+Ir
oEOJblHEAHru/NA3LCOOOMS+057NA5L6dL/MQ+glpqpvjSiuh7BEzJIQG/ayVzly5zuabQRkYcp5
ma5QU0NHzEHKn2w2bqo2yhz3cdUaTwx3COqe06FBlHA0rEAxsYnD5XcW3Dw+7/X1vVF+chP6aCCA
1mkeZuI7HY9Ff90s7qF78OaTnhuyiapywJ4eaoFYZjKtWv3KXSnCNpYjM3L7/2iDfOhPjq2/pjZY
L0NbTaKtqR669XRkyR8l3GODXp0ugBr8W50Bsp+NhN+8krwpCgN11CaMQMFcadDZoTV6uL9rBFrZ
JbNaKuAg6se3ge3qVPKRyRPx5Vct9+NcGQUtzIu26ABothhc1KJBwAEmzigu9zK9OTW4KX+QbUI1
K5pEQcfd33Sv6Ralwv56Tfvls07V2tC1R+85dvnv053GM44jahM98gZQcCHR9F5CYUqTA5hk2NLD
EMlEU/KJ665tjn2I2phwatb47/HHUoBhtHn3Lryg0jyv0nXrzGrAYcBWEttfZtjTvYa/E3GsHH3J
5L1Aw/FrjespdTulBInqiu1c0l283cC8e1QGKAvLk9nsVsAReGa4WVqlVkDhwM0mfGy8t5KA+lhT
l/NWU1ArqtnF0MGo9G2lRDgpk3ldM3SdRMDVO2lgDb0nmKCMk+nJeTFYvcQk0J5eG/YGpQLuDVaX
s5ErTSjlifZkW6qeYTvW8KE4esoNeveegZLQM8g0WIp7r1Yy6hrzHH3wG2cLdcZZqAqdti4Cey5/
PepRfXj6zA6HC2gkGlKxUdIIznl5jOP52AYu4HnEB5TLXUnd94nVf4e3vri2XM0++tMCB7kTP3y8
p6gmnFcSR5qaZLA8fi3tizPTnZIZyopjIEXm+q+FHFmSeMkbA4PQqbx8u+IQl+rjjx9NcoiCZ0s3
x9O2tSazecxJB2oDY7GoIwIFGhd/I+O/NyeA10BRlSWNeqN0zRgKyaJEWCSh4lp0AVtDij3c3IX6
c2ON2w485OgVZF3A7k3bOwowRO80hKx6P3fXmancdkVo/nODhn7v0t0dSW/7bMIwITw29wXbtCvt
1zAuV/Gm5p6Ba7c1/lPOVpgGLoRWlWWtjcTTDdXEh94wmJnIW0KVkOXyq2Um1Pr5Fh3P98qHELbN
y4W28lkzdtLcqdb6P7lhQ2XaEEbbOYypFkAbs1+q4b5B1QBoUjWMP2LfjtD9pBS16mXbp3je7TMw
YHof0SdvdmpIu7aCRFkMe11DGJpPzmngHKWa0eLFvVrlcMkjpFMJYxoJLnh+0Zwm/wRvuY4//rj+
EL0ln57HL5+eBDyemjQzPGYoPybf4zuVXCYLgiL09uTsjf8fosZjhxx/c2OxLyD7JG3ZrV31PKl6
csnw+aV78k4AjvXSfSYnazMD8A2JkDwAAXHLsMR8DUc0hZeotGioqPwVw3Np6IQxHpa3nBmag/rc
0Q7sNw2rJzKgH/U+niynFKaNctghEvHhwL+m/2V4Mjun6Jd3svIyVLMDZKDT9mk5x4A/Pknn5AEc
zAtyVPkQ7Ijx35B8JWsswD6J5v8z+hwqlZqlWzCm7Cp3IXPMswd4rg2WqeUXGT07VnedsmW6YD+3
Gg29KQDSyCYa/y7Iryui9Nlc5PcnOSuYEA+PUj351zgIB61e57bE0Ihic1Ql2mY3em16zFq4ELTL
bMH2QvtMONadJOOYhqq0VVHYlk4bvLGPMWq3EGQ3100eZMdB38tzOR7BVhpvmWJ9jwidFOIqLZq7
j02fifd7VhCUuZaKRU/c+kbUNXdWKjpjgbZhjHk+BCc6C9XygIoKWC4LydD94zT6Xa2O1JDr2vGN
z4y8KgJH29jpPRWHa1XJu2seTTOt73cE8Efi7r/b7XAKJ5XB+B9yTHZG7p2yqf+AAqJEJzOpR9pR
sNyB+81B6thLr1uuHDQLC3XLqdxh+hBniFnNUAANaIHM4ier6JPa2y8eBh7ye+Bha5oGVY4Y3RfC
sQ6nPa8UFMubSN2CUe5xi1wOdGA4YWfg/UwYLZwDrm+wDoq0PhFAmFRF+qpy0cM4pg2OqvCp0rJC
Z0y6wCPcJK1ogkoGqSmIlQJh/Zm2d7Aylv1SF6zBVUt5GftkeDXZSzGLqsJIJ1xwC4UtRsctgLnx
lEDjSvi1LE+MWklKGWcv/TMDf5gqn/HV6o+IyYo2oYSoSZPezSNYSc7ZAUEqwpcSsT1uk4BDDz1O
q5GFnwuA40l0at1EJt1cZhEl01t2P4bAgiSq2vKXsmtQ4KUZhqhfYNwBTdmXKnsuD5uCWm+WzWZt
pJt4WLHISVDVtc8Z72hcXXDdBxm/Njk39wsfVJ67jsCyWMg1IIG4q1AlgZggyk41fOJDMpU6zFuD
NnqISWqN33DaowfjGB4YYSHNomBlFDJ958mkrJd1NOra+Df8C1djfcpFXiv73oN09YEyERquleLJ
MG31vDWPJiSg4VHwHaGoCorf2I1v5l+epr199/hRUDXRIlT4Lypi0GNhB/fDPJUnBB+xm8u0FPFY
f8917MQtO6WKwKQm4Oa/gYoWRaxDVFqwvgIonbHuh3SSoCIxr2w2nikno8BC9ivfxTGljxXLlKQ7
oZVPvSVBwCX+3wtYnlHqbbDoXJfoMvmc9GMBcwKP8kbIw1pFt9OCMhLW1thU5V0NIcKgiq0V/JwQ
G9bt/Gf0M0kz+fAknzaGplYgMoYJvXyz/1Bz8forR98xNGL/GVmLiZf4ZFddtrkArpzeWgbriV9b
7VG+WeFhwIrFX+RQbLv6XWknT77+SdNeyTa7j6rbNHT4h2PuuJZkI7KJCgoloEp2UcTULTrmvoRr
RLIiFgnvQSUEXPuv21X00HLXuxAhZsk2rynLFeSCVkRBlw4hyhXlzcvC9egkizvE6RyuNVu5EvwP
2fk5z00VG81/fKwfRzg/sdDyotd4XHJlQga9yFNfftn8cqfedT4Qn+bw6LBLnhJIZ4F0wfxUuZRY
YoyppMLjtK9isqwdNR+kvvNttGH74EQ+UHp7ugkMh1lK4F7vESOiOodA9ufCDq9DvWCR44eE+4FX
oNdNBDs85cTdsWg/HRN5qH8qMRdGYmOzqlQ3s9fOhaRHweXNNBxi2OPXxQ/2sK2K8wvJt8iw0Vhx
URAru9CHIJLoRQJYuRzMyIWcKLxzxVd8O9KmBFpUidAzq+gMq/qIayLodJ+hIaUv/2dO/6YoK0zP
WsVGE35p9XGkqWL5t8/oD04AoxGey7iWCzjAQGmSXyhkyPeNw/YLbiosf8TnchzHl5bCKpsc53+V
oV8eKzbV1Tks6AEZUho9U1/o0xHsalSE/jUq+vAPNctHxOJLoQtN0GHRwP2NalyjmCBbjfYoNzQ7
pN/IEBhVVMZcUQbIRYIwiYdxtkVRrLCiiHj+Z4cLA4a1G7f7x0ZXQ1xWV9fn5xsUtj4q35iGZL3z
q5xuyMhnHmvcn8l6ONIq6plIKn+j81QTPDXRysvSUSkk5F5GcaYnTbYaG692yWEcYEIz1x/uyOSR
lLE7T4PqW0zeKmczXwgW8//A9s101Z2ZkchrCIyPOJ+xKmMr2owezwGy/fQZXBGh8pSDQa8mZZS9
50Z6Je5z7PUiA0aaiQ0rrRxyG9wIOMFH52OQ3g25Jh5c5xmn0uBGwV4nUAVGOzke5a5KbZnbe65L
i2yc/Qjaor1m3PowLuluR5nAQexVy0bP/lG10+droxF62qJ0auuiizaGSqH0WTFOmu8NpCs9qXhV
VQ70BohNXYR3bfVHH8gFDvfmwT0uEV4bsa7kUeDa+8GeMBrG9QSW/BFUwbk06ev4mgKLmfrR3bos
MYgdWgEoXNv+H+cnVANqq1HJp+19N18+4+ptDu8p54eVTtuDw2RMHwNRFj1JH0VXxqG2SeiASUG3
AYddrlJcA86EsgtqLnCjGsqCPvbeQtx0eKckd1f0LBift2ZtJ/4fe7k62bG0Xz9L5LiXRiUPCNdv
Z/3VFVFRT57t8b1k76vSA0Ml7CiTdgeJnyyTkTyomncP+/i5eTxNA/2Nl6p5ZeqmaIVBBEH/hnrA
q8taHWfiDQ1hI1cVdTQ2OlJm+kxNV7tphlY4pCUdjlA+VVYKErIrYsOYSHoM+DtpJQfJNKDvTfbq
ZXH5b+17BxlpCWBnkRLN9qolAb/B5xiTSqWLbgHjO7rFqRDBm4gRFiWhTa0JJ29NvLu0C9we9Avh
7K4Cgy1iF97SBmrVP3oY7ZRd+fBjMSNTl6dCsQMaBUn3Gho6s4e3RArri1yl2uCNRstRfGIBAnbZ
zPWu0aP+TtFzK6af6EFK1GqS3k6ky4dt4nnVmf9aGI0S7hQ/IpFV7/P7xwdlHFVeIc9wrJurx0Ic
fHJQ4ptaP86DqUATm/r+1+qBz/qEtNnVPSRodzJADBn5pVkyAwJiR2k50C/c/iQM3M38pXTRqZoG
g4+ZobM6JSmaCPC7VyFqDUeOb9p10VUK9/D3BbYofgG/ZqITXNK6z0J56WtH4jlTsGNEX/phnzTy
TNtDpAcrrEf+0UUw+L6t5lAu9oZuJh75POZUFO6ew38SnX/gKdOEWJpdyDNka7Eivp32SixFPgZo
XyIesHNwnUT8qlswJ41cC799SBZx0FUwE9r48DFtq1/2XU/EkDEHYAOHvzv7KwLqfz/fqttqm5E6
8Juk6hvAVhuvjSGvZz4S6pcT0AilWsnHdaOGDMt+LPWZOEEoISM/40RKaHBUHdPpDQ8JQfcq/+kD
s99jthQ5JCgKRY3u5HQBobHVw4dYn7BOtAMcg7ncd7FnoQV+1ANl7OkMjm9sypCaYtdnnuF82FH6
Cdk4fTnarJyw7H9hQvu4j9u3N2hWqupn9nhQVtZEP1uxc1+dTVlBVeZdk86mLT2mCCvGRE01Xg4S
3RH3CacXNPbiFHlF9ZWeCbXfKhehn9NFCoURpCvrpNgNHwceIrnB60Vl/nDeIfgktMgwFgDwi7Os
KznGsozp2xtJ3E3L/2WpQfPULyp+TP/BRfq6IHttqfF48BkgTR5yXdVp2k5faf88YlKlOltA7VCm
P5QfUuWZHyjiqZ59DzEpJ16pJTb0G2uOIglTS0TxhYy1mh2xsmdVOl0SEzxdYdDxRvdZjuTenFv3
GlPJ1ljzb1Vd34V+zZKbZobbWfVXX+5p+m1Q7TJ31C4o2YjN2qE5DAJGeX9h8ja067jnfWvSXLSe
QJTlUd6AcV6Py32rDgMME5uO4+CtgQIEAtqJZ3vzXUOUOb0voR8RBVAw3kfPwX6rXwRbQKFVH2Q4
VYcLs4WBTuVlGEJH+/hZaj6DlwvH/0RP4FgLJJfCz3B/xSwgJueJkVvQI50kHkdibKSpy+ktD521
/gqZg2Q05TkaUYwhwTYj4inE35NEU85Ep0E+E4rBRwfPKJZbn2dPnatBcysSetX/oNqQ/9K/DP2w
9l8nRbsutH325Zc4RRONwD3DEhKaje5EbABIdJnpt/pyy82c/rIDGO/k4Ypw1ANRvRGkgOrQNqzX
242DsINn22WlxNkPmzoCx70hGG00MglHCoE11CWuoonuOWrjcPQ0iQ76CjSpOziU9phbrccNMSfk
/NrFegf06fKicx+BQz9flfua2TfVH9OOYNsKFlexnGb7HzNvZYhLfDokYYbcnllHYGimKIvMiBeL
tlkXwVViI/LgsVzVXeCViUU8ZzJAoIUQeNuaO8rnIV3g5l0OCC5po9WugZ0CzR9ccofNn/HT+3LX
po8xmHVsx0kwzK4RrE9iUmJQyN0DvBcOOvMQ9/nEnqVVlPN44PYQEuDHQgfgjrs5Dx4l7ACSXS7k
aDeoreybbhlyJ9VddF78oLAZ0H9lLin060435VbJKksJqCSd5QFEsj3DZr6nFfjHy5u6DycSdo36
YXEN10qKSPDC1Zp5VajojTbvX8XjaSmGpVVLmKt+j3ydxeAlxeODelARutxMFOsjvMhqAvXdYxbB
JU/HNN5TjDORzSkFwNjwTQJK/xKMZrcFY7Yv2A4nSxKFu9pEnvkFIib7xiWoSV4D9d1LJldqfUaL
dIuTF6NSHO/xXqIx6eg9xAbX1srYN1jU3aVsM90FSPva+sZ+mK6cEeY7vE8lcES6w06j4Wdovd1q
IIIV/j8lRBYxfP0plSLgMjk7CqEE5uDVue81srKpMzqPZmIQZ9kuTULPtU2mZwOdtt/Dgl0fwnXb
/SXvqKum99rWLuuWoDnX9TA3E5M2m/z69KrEe80wt4TJ0QTybJlHBLI+TSY55Lgt9r91GMm+PV1h
moFXhiKKHDJgNhodhjd8b5C+yIsCaWRVThlG3nNF1K75KQ8XrZfBQ8j+1C4QpTEtQmcuqX+9mCN5
6imysm3AeIgkjxofLlGWg9JK/K63iErXVneZ3lIQmWkT1XO8ndJ2KftUD2iASQuKptvTnXikTmWP
EtCj3rfhWxkORu3BxYjYn8F2CL/+TYON7sKmqgLdxQNMPWimZZIKYEb+bHDfhINBpvH6WGQsFLqj
b+bYopIOnKzY0Nm84bikkgIf0yD8AT4iN+aPRnPY1iaixUVI39hyKR9suAuMQSWAFy4Nr1UYAwqK
4Xs6fFTHtXCp2w9x+KQKLrFq8ImB+8PeMPHB6SKipb/eh0fO9YbqgbjA+Eb8o2I2BCMOkwK1n+bQ
R6kfP3vPrArb7G8oi223qfB8lKE9ym1DjkPB9WgYj4Dg84PwNeVvTTDfcoXoN2D8jUdSTcAMDXgm
Ix0pTM0gZzRs3Te21qul7gteZHxy4/Wi+lmhlO3ukqlbElbtFPv8Jsf6qx81Xzp/DZCKLprgmJ6M
6sW9JBcUCVG8Z+OJHT4gOqXWS2q1u9EXT+WBh/HZpcNogLakaMJ3zHx8qJfDP1Hgy0yiS8Hs0MQc
At6/SSH+bWT/bYYRfb9Ntn7UQlgaoklkyFQt86P9K3Vtmh77h83Vjy3YMl2fm4zC5K95HqTCSXGs
ySdIYyzqfz8uFiIZDcVBFnbSvxMbX4EHh7cS2NngqIrQ7cSo+LxQOawlPJy1ddAtoQHe8QUiYMII
3x9rKV00EjHE110MJmSjQdVulBqEfoIpQPu/2oG2BACicTo9L/8I0ZsNAJCwLPPWf2VPowpSnV3c
cQmivMAa67jPPKhGyTfmi7pdtKEtzMHE0wG9ygvX+HDcQQWW3cUYYSQx7ZbAwdF/xKInteOIr5Le
29TkxIJ4QCa7GSrP5l/+GOdrtPLHYwQ61xxvF8Bf2XpdO4K+e0hNXxHPXGjpPsEtgU480hVERCRq
dbZ2/nDdrotenZzPK9dYX29OowbUW176rwQ0lipnLq2JtV1DF9MuIBICDt0HzQzD7GtX+UGDfT97
qhmkg6JmMl8/VPn8CPNF4t5IB45dD9khxKz5TNvGLfu/9yfEn7Stw1R2XLEsQ7D0NQQJe3eyed5+
KO0+m2LC4x6dunOXog6B8mmW6gYkqbizgBfXCeT5P1dFiLCyz3Pxoo3oJpbFIaTaPOMNIbzUTq0U
p55OU/XfSxjyg5m0hTQJriCesiKt3khrOynFqPGTWEl4rlkTRyXY6+GYkp/3QCdk/bAAKyb/kb2m
yw6QJTtXDFqW+JNO+cvXOqwv9dHufYSYsjglE5ec3RUnTa607A6Jzs9rzgs35Imv6F7ateEutAKB
eZolzA/jY+fAVcD2gOBhDXzzV88nsk1QyzC+tAf9iWQJQFuCGf5XXzWgA0hKvSgluwXo++jqe2LL
Fx9cv35lzfllkkkQK5LTyMih5/A0EG7v/PJdd30LYuRKImRFwnFZutPIwwSMPQN+xtYibfRXhH9k
UKPrxbPxqGrEQ7/sWv2gKr40LW9HeBkJMCvFvdz29UhBdHUufIMPiWR5rqV8yJI5xN2Dzn4Waxyx
50x3o7chDYLV/PQ8KMzvH511leFYiHskmy0PMfy+gowS47WzPV2JT28D4bm4UMZ8gySpkaJAk4Zz
jat9FRJay5qcq/VmNebdHuVQXIQt3whiMLe2HOiQ1GHeRY46gmDniIh0oPeFs24Cqm6R1PujPwVg
fsRoDgzmDs8IlWpgxL0yogH6d70CwpC4BLLu8NkbS1Ed8hlCz+CVPlWVJgKiXm/jpZEuefOGiydD
2q76SF79Nz3LB5oNZHNquXERnuH3m6KztBXC6QlKMiV2ZAyw/WHZMaFOaHbr5HZ2ZXlHM7WeT7XF
sg5kfJzjNEdhJeIa3kV6skCI4iiAfDvpYqHmqXQS9QADwC1aQhjtg3y+9/6LgDMni7fYY/d6pVSp
Pkxy7SZWWDp7JrZodLFvmzFCr233S4wrivqXcmJPTxDAy7J6y0fG07hLZAJ9avXmqjlxJWMuaK9t
nnLkpK9TD67qXMHBlXO0O9eHfevpq2gEY01+v1XoPua/UFch9B0cV/YTFK3dc2X6s2/67Wk2fJNi
rNHaXpAw4rhjVllVDA3gKVVzYhPcncJWI64DXzSQstVx2dr3x4XQiFAiI0uccjFWJ5OAzC/6Jx8t
mg+rfw319dinEqrSuGcEMCZFODx6tVH2NkNfrY4y4Eyi6yvqDx5Y/BXwrVG/wvrS0bI3TX7BVoVB
e2aG/GHQVgDL/cXhdKujX1sLHKVRebVI5ARbRWAARYDB3JkE8PSzzdLQhVG/PHaOTaRd83MCKciD
1e4tONchqU6Fy7X79KDyLYjhOd7zJ4VVm52aPTJvMgWh5CLRp0jqlrnOGuQJ4Q0AMqzrlaEMli5R
n/rjM9l789GqdPUeaXiWSOcs4Qpi7UnXUZZ1YD8MZZ4p1hdMU1bM/iKMjwJt8oIYCwwhIjImtLgF
g7cM1ob0EIqO99K1DRn+dwQt/juMf4LY+dj9hoENp9HOLIm8PhriR90pQaPQJx4XCex6Dge7vLL6
8RD5lxEK92Ecdre04SUJ86VWKVetv5PHE5lRmrxyt6LoMEDpIviDfJWDy+WX2eg2qVhFFLuvMOMy
IjSRmVN4q+7E8omP56vYlEzy2qm9Cdd8eeKRGl0PORT6jElMNh+l1DIIwGaEixNYtVygCrqXxFc8
rVfgiGGEO/tA8XqDPVF3n/Rr9cJQn2XnVgSUIe7XW+ax2wIHCzG7yl56SgG/jOMh0oWITDugJIha
xngv2rvWGbOMQ93gpp+406XfZaFevpC2UaFZ4/7Y4s90JbsRveyETb//XKeuLtqBz79Gd+vTkRGC
POkyrAEl7o/0WxRMNNpW7YxQ1v1i6cu7qznhc89u8/3ujGXQufR1wyyNhUPdX3JnyG77hncroJ/k
UVZNy+VwScJrWLmkkWgt4Z5+0j+AnmB1tuLE1Wm+ntFRhGRBGGpGvfONCxfS9GjS4I4dDGcWwEVt
i++t4DLRMMoRRi+MiUF6lTlL9THhb7p8N1L3wDDLToDff3EXLFxnhTeilzFckFHG6pSFo212E9Ck
Lhm0Ttoz8K/dZChTMTccjXsQwaRsPYvWrPhTCt8Mpe5MjiDBncm+34MitnApb67I97UKuvsnuOWT
lLqbeFeQjuUY7yI/Z9VMxoQCslT+5C0zaddxGx1hOsFv4D205g/VxMVyI34xee8zdWiYcULi6F7/
ZQj0VGirvro6BBp7ARF4869L/N2vZS5BuCr6KLn0T983L37d2uUXr7tdhrpTXqVpEU5+lhBLE/b3
dYjvd9o7f49hf8yzTevHgR3SBE5vCMukHnzFWR0VD4+AYMmc7EWGX1Zn9bUyntaK5qB07bRDckE+
Wf6L9ZQs2GJTqVsZDlHXpKNYjfGy5fPbwp1LT8vNO0NAK51R9twYcJdF6uo7eQmYywb1CVZY7Aq1
Kyc2RB6JWofGzoCd52LfjXzr+dn6Qa6WcwtW1fZhKdIHFKzjcmemWAHdaM6SegpsbPl9ypzF1nOR
jacUhx55po7ix0ptNM7aZoGC0128kmNEbM4Cr2CF0NdCXEGbcsSUzCF8XwYqMxmPxqZPXxXPFyZZ
fc3P791GHq/ok0Fn8XoMBOXlQTZ6x7zQ3xjzY0m4GpioK0fBoovcZRR+o/vytIhVy/UVC2IySnD8
dcKqO5jbKANw8TN1rCNhEFrj5VWom97u2RyqgXwc1NIVv63W195Ty0wcEuqWYl1ubdk189pkAEJ0
IG/Is8nySeObQLbHakcejZg4SCFynlb/Pj2f9iZuQttEuK5ypBwVJYK4TcdVb4D8GQXHtMKrdHpb
AGypQZlIzg561M8ghF8HrIIJ9vGvlVx7l33LlYoo3BZa3paJl4dOoIQAq+J3kN13b7m95W2wpAPY
cB7eDzuxURrrIcFF7PMG4J4J8qeDYKeZs7GGXtI0Q/5eAQ1G1xeoCrrfmajOwPrielf1Q73Ski2a
qqCIs8wfD3CIGVlRWdftnf0HxSR7mKAJdtLD/tJA83sulPlmm/0a1KbYBz8t5kjmy+G3UpyMiSh8
EGInVo6g1uXrbcEhOGp6uj4hZZiCQm6YHIO0upi//wrau+YIj+7a5IHprvjoWjyyDjLS7pfVa9Ml
1O3MPqfu3yrHNvoEqy7WY7IE1iKFxjARuI00LkvZaNaUNpVgUAln1NQTSPZ2q0BOkoKJtAKAgYEj
JwQ0Ya2McMOP75vxanjkGYWtS6CGRBETMCcpqi0qhU0voiQz7rSNxe6nMmTTB1Tx4kN3wo5xrZy+
FcIYEh7ovoIzTjhJQEoJz8N+1ie5USAiFtEyiFLqMeo3q0TAyJgiqotbdrQJz65k4TNJ0hOLqO3z
tyIorvsshBdr9RmVmwsDEsv5QJiFC39moDUamPRefMFB6n8FKPXTN3LRa3J46mMog+Kbo8FpiYxE
E2OaEeVz15E9JjA8OyBtfkTacBp6n7feVIyZMrs9V157OdiJX3biUoc1D72OhfQEvtvWO82SIGr6
NjLJeSMozuxqU+5uYbAnEhnWRZUshMOCy5bJf9emL3DNNDXNTA7oFo862oX+jUSp0Uo1zjmPNdC4
YNTsGNpyBZg/fekXAHzdB+vUrYpoxk2OsxJmz4mCWVcCyuqM4s/8Gvn19zJJKeXkyKqDs/UYIBQW
zpbgtz2T9lIBo5Fxb+ZCUkBP91YDqXFAZVvtpDrajIPB0PUnXQfH2Zy9awyLT1nmGty7vfYGJVLs
IDiPSNV1aS5AGOBn2KcozOd9OcZpog7NevRAqWtUQBEOCNmrk4m7PVJaZc93SsVioqtwnHnQEzK6
WvAbBbl0/Kk9Jp5hCLidYyvqaO0nVVzhgTQh+40LaP1syardW7jNasGIpDK6GcXTj3j680RWJRC5
k2OW+9CZF+VwMsSKrH+gXlaEPnWYengi0Cyo0xl6ExFA9Eg8EsB+bcPkiWJPG7f/uFjl3ia56wir
20DvmA/iUQ9eqGl3kWhay+bYtUsdji7O2z3gt2dIASMJEVd4WGukf4HmZ5qnjveQBTdlph2hOPMO
A5TpJ5oKQJjzeJjaMCTZ+DmyfUkZaPRT4q5ZlT7CvsoBXZ0zD795H455WTp9tbaqgqKJP/t0RKpP
vQTDfmAo3nYuPwoZvgayKYmSQPOayXQjPvLNrr3vB1vHCfV8RnKOM2HZ9ciIxrp76jZ+UsEmQmgs
p37bS0xqVPtn95wBbMypjJ/jzCeancfbAeBuwcKNOTH8R9HU+9JGFIWzw8tdeGfO3iQFxa8R8eV3
6PaMQHCr2AVmdf786GFx8ES41RQf9qNLG1S9VYV3h956nVurqjN7IGJFx6F4zw2e3t3eAAhepGw8
RSZh5dcW+2/1hCOFtOEkvJ1rIpGpAyLetazywSX5EOuS9J2aYdTVJ+xmZxt57RyNAPaeuc/ZBtWL
wymSSKPX18u8HC3+C6dkFGvipjALIrhMBZ+tA6IM9Z/gPdU9hLaUi8BmLMUc1DQCli9JKo+/KQUs
0WwcmcKVycuIGKUxMCiO6i7tuP6VxYdLKr/qePo5d7VTETiPXW+01JEAEKNQSgwANa1xQQ6qfBXO
kSkALJekByyEYImjuYcO+u+zvGGDLr9j/SovkZeWg6HAx7FTtC+aP2bOQtvDW3GRBOpQ8IUvGnXG
MmiIA8xhEgrLUH7G1z0IR2Szf+fnQljDdbsTc06uNpLCH4wAMap0GOuMGyRN6jgi0y0l5EAVXeUx
bOPEQGiTR7s4r2a1xxk+qE9U8+5xWSoj//JUO798ugyUlKhfkCqJtPNsFz1g9G3W8bP3zex/FO75
5OBMa/T9p8iwS+Y5pRDwtDc+ElxUNCaQSrV3/P2C7G2YYHolf/vBHOrk1ZrB1s9CYCC8S7tM38iM
rZeOjoJNXOhAkET0sF8FM2KlyoQvbr6HVxA5q/ntlTsy5MFjjZtGFwgbjOFD/IcykmfhB3AbM/F/
YBdpW7Gau0oih2IfLNXaTSqboD3/0X+QgD+JppUjOMy4aP5JhmpzJS0gftzJn5XHYSObNGaytyny
DF3VXiIGiY/2/c0oOExNEGSy3ZVHwlioMXzHRN6Bz8E8z+CX4vPAk5aAtsq9lCOBZxxiWqYPfhU/
pGvbZRzTRwE6D1Hih1fQwVrICgBw/dpD/BS3C3fl1pmkd6Yvn8E38xR/TPsQ0VZjV2yTndSpslmd
LGkXFwNVxyGpMJ9YEy2ngc6G898ZhrOKR6GkcD9l2pgduzJlQD+MIJwa1Aca3ZBGS6o0/UVQrhvf
BZfboXh5Y84wjOu1hEDKAOBE2/MW7IU0nUotA11hNpJJ2Ym/xz9VnasYhJePyRTjdVmlZuB6ua/N
EFGPSKcSWAMkFPeMMgRlImp+hgbXPRWicVUJWGwT93xI3kxP83X0Vk7p6x27CAwFkxxtN6C8zrht
r25lUuwcbjZZBhriKiJ4iqmQSs3szmEnC6Oz2O/a7VXvXiN+a1QQ9BbITrQMosueUfkN2DUDpnJI
KrYS7Tnhr3ajyQDsvhcfJsL0G1b6+77x+dUf3ET3b4/UVU/AAQQwMpAhaFET8DVLPXcZMWg5VLPf
quDBnn4WKmQsU7MKv3slrX+tz7ztCnIDscPEOcu383wFJY67eBm6UtxU7zGzqH8jU+xExoy4U00P
ADSBO0DhBQh3ey76C2dxh0ZH8H3OUCVPBJMwT4cILJ4WOyW9SoHSQ9u6ulrPxDss3iFeIKw7ei4U
QpTnb1pCrs6iuR2kaZVTcwxsH2R3RNxj5hQZCaKGXfdk/aGcOF7L+i2IHGhU3qPRzGamvvgQC4Lg
paqeNcms6FeyRR6Po0p/bEjKWMJZRQLBH7U7jUW+pPrJ2QsFO9RCMHsLvZ0ifAop83HoxkYJSDTZ
C0OfHcp+wxmMcisiyQYf+RdEcK5/A2SNu7OBZjv82cC0blTeaVM77pEk56cjFDa2eXZtFCmwLdjC
WgDAuUD77WIbi6TiRknGZqT6ILFfrPaQIjRcmjvBI3U2wljAZRzmHbKuD1tQ4HE6KP4e5yovfVuI
jtEwpg20c+tLZA9eluckrZtILbL+wNNsw5o1gAjUR7MP8cgjNSqHgtNF8vqVd8zSu3Mbr+SCqvDZ
kv7mSP1RGfbs97aDIY6U9VqvY9URohRaAtYZkgyUNP7edtYtbr5w0f+7JC0CmW30IUwPYO7Djp40
9uLA9nrAmUtm7RgUx9DmE4e84+uz28dHdKdA6FvDQj0VkguNdpGMMn+peXeUbtT1akFyHedAfxUx
tIhKrOBsZQESKaAHAk1/vp1/37DhDw31bwiwF9PG29Pi3g7v6l6dx+rTYFTG8LrjsoXg+7Ivoa8N
ujFzSzv7W0gI+Br/PZi9+RtpMCdFyHLQYn+g9EfPdWT2iR+vVPOEMk7bWupoZL5dGpscZ6AZhuQK
ABqKYYoNZXDvERBy4e/akhOfXDR2c+H79crhMpifc7YSdlXudqAcxKa7zagw9OifefSjRKhqCMnm
QK2trQxzBbeDE6Zq8fQ7Pa6mvhpn4wyZrYh2fVF2n/oyR8jrJviI/oag1o+9ZlMG8DuEo1OLk30S
+c9Q5119D6AvOjkCNBe6/+13Le8DrX7v20dWACEP5LCDrzm2kDckxTp1+m8dqzLHTL4/IsBI6JKt
fXP/m4UqUsZ/zrLQIr3Yv1OSoCwZfkRUL/9Hp+MT7BGz1lUPdd0fU6MjoxWoc4o/N1ZcWh6+dvOE
Hh3IyfJK8x3AJFF0iE72o6eyRL42DayqUwmCvvheGgYCYbdp4uXSTY6w9YQ34wG6wdG5iqP3B+t5
DdltxJrN1gIgLFSPH/3/8VV0m94U1FFMufky6H7vyzlmWdCADa7zs+Uet0EyKs4lDHtUZc3q23Mn
+JG5qTEIAwPXJBpiQNeaRzpnxRzFO3LDT3vhm22bsbcqjoUVepHt5j3NWgBFR8BUtM+KzTX69mjv
voOzLrhF/hsYn+WbqfyA5p+K/0LhMCwoi+zfCgLxGva9hnQ/RcrOxYd29emYvF8XMfM9F3vlIemN
7Vprf8z6NvI+87s0FRvAhSQvr8LZca/TzFNBDG+ASWiTHdmk1tWATjTF4fpzbavNdnRehh/i49Tt
JxLV0WL4NRMys6wmmXpiE4rPmg3v5ClJg1kXeOLoe1eIMxIs+x+c85BedAQID2NbuxOD5IrqPMEx
axGCdJcmAiHyaw8Eyo9FlMDjFD6zahfsQiztegQE913Pxd+mvBmiEqGb9Uf1djyN/INTzJAi9jGy
t6TJuTUdHkdx2a1hA4ulrPQe5QiIKHp0pSKV4kNqvjjK0Wkm3MvzbwIdj4dafvz5qoUsNjVamCFy
BmPCyLUsrSNiwKVJ6iUttNQ9bMib8VhRSVLZYDZto0LPsBGB2u7QFhc12NlT9r1y2yw+YNO6h4I/
25WBI3AlacC2JVKpiM+Xas5NEfv4pchLUISy3uuSiA+qWWxnRSK2kDnAWDI7dWIeSlpS9JBD+j51
VDUwDkZU8iq9uI7tNnqnOEdaD/ssrhIARuJcTvAjkb5RNwibmnkq7MEYlAvP34IjjUEko9XG2x/S
AUrX7UC3VhPV2X+0bHvvaVUHu4CRyEpZFJJxwlLptNJOXs7NvanSI1f9Ft8p13/l+82sPEgXgWzW
lw4tSI5kBhyVgl2kMPjLjaYXYwMzNQ80LzR8GgzE3A1U0FSms17lZ/kcDAGTW1EMk8m44Lq/4swV
52HV7+jPLi5lBRkxre2jsJL7UWXGXfs353G3ObCVx2qGiylAhSf/R77WaepHc5p8Ls4tQLvI3lPz
N6tAfVHx+0JmbjQPo2NWlFIBWYl+xUYM1xhsaOJEeJNF7Zuw7u/Ob4GfY9tJPLmMmnPWjdeCfSn6
MjVQ1Rm0JHdsFcH7ilD9Bgzka1tUo9J1QUEc3N7Bbh+zKrtugmAWcpBf1HnnsUDHx2aXdL0QtNxW
sBKFrFl0ixhNH4weqgox3OKieM9Gqd+3+oMPIn+qzJy1TcKVT1Tm+LK6n22MpDUbFNXE94/+A/Nr
Bs217cE9ZfIJ5qiLep5VMb1HwTWg+3SepfA9Z23H1D1fZRBTl6mAGrf/bihIaHYgmK8ACg6vmWqW
Ui+2jhvWl8kG3D0owE0Jj3W2FCNFZ6N98rdoE7ISZZ5KnhzitJ/fccArLLCpd0E6MAnD7RvRK5Ey
NpsYBrah4a7PsnfNBVgFCWf4YIyhDh1nZLeXfRXzjuvptbUf0cmqg7wy8e6z/4IKY30nyT0FdCBO
JP3DqHAxm8BgZy4+A7b3UpP4ZxpkcuMe6sLqJpp5EeYwqUORuZWLuyr53ZIv5GxOG72Kr02Ofq2l
J3oKAmMOnX+EfVMZ0E1cpSmTzlvGeGlzHl5Mj5fPNpgpzvqV2J7chlb2SdPAe/rIPcKespmxUkII
RtuxqXfOPov6FqhodwQjmFfRdJ3t8IAObT58vXqfQVTDoM3xWP0Z76XRtupeAc1VoMAi1O0ZLsZd
0rv4Wp2YPmpZJm6TYSRmQZ0IxYK2utN2YA6yS5+I/7pyp1TMXY182hJxAgBzaOR9tszEwZ2DDrUF
nblFdi1ByF9QKiJ7jFbfDcwkVYJB+VDYTYrJ111BmL7bqFf63v66R1dcdDSoQf9Y7VfqSvKkcIyp
H60ZQtXPo/a/Grnnsi/83430ql8p0fG4a0ksTOS54VsNiZCOEJDKMJhKWw0sN91Z9+s6d+D9DXHn
9iFzJWgCAzCqnxJVE/0KL6k+cn4xsovHo8gsGTNRs0oox5cRo8EEZeXbTmNjaLANXnWxJknnG26L
7ZJJk7iwzhW1xiGr9vhqhD6AKn/UMbdBoT2pBwKN79H4NYGg1+eMdX0VUjGdGLtk0rhIi2tBEezK
/kG5/M/KOTHXy8D3Dtcld2ff4fI15CvuIsMTXYzOW79ohLuku1NCnabmxIcU2Gwx2mq2JF7Zs+ov
a76YKHD7yrMn+hAjV9cJAmqMeN8Gft9DlLZgi/cGdld7a03MbK1KxQPcuaHX3+mWFCWqbHFG26iT
c+XeI92SCRL0UyGT7TtqH3blSkNpxnOT+jtK/c9q/G25Fi7ZRx1IoJefjWLyfwPaOCrWg7Njlx7a
+38F1V3SA6hKHmqTz59RNiYVPuGwV3tWGCp64R9vSHFHCnd5ICMkrlxY4N8hxlLYWH39tB2CDyIG
kVZGNDymqIj+THo+8xPMwvmCgswXFpepz+Oo+8go7t/bHvjj5zAC/XMRRfx6JVzHWYovBQHd8AyO
LHc22nmOpruIQqZzDy2OWIQ8y80kQGnZi2xynz0DmpoNNRqRL+s3TqnesmlQpGXyoppaeDNWtAMB
4y9qH69k+s0kYatE91j6KSUSdBZBUIHh5sQyKd2HVk+ljWwTaCmge1nyW7VHjlAM2HxbguJPRcFv
oNyE0QFGBn7PlIACjOLl2kL5MMRD8fnwVK7rFP3upEUpVs5pcJzGchEqYsXZj+U38o8dtyEbwA+Q
DkPlBhtTbMn7rp3+lB8BE6RNSliutPMqWXv0rMIYacYAWSUR02FmWXXYxUovNmD40sB7PYmTPOIn
wNb70yp7IS6qzCpJgWzIEG4gtdFLDKVORtgLjqMfJJH0KjtAlCw5AAajmKYVrTyB1xORQ/0AbvX7
F5bIMgXuaN5NIqhGFUixT+AlnWyFxSzkzR7pd2Bm/wADAssnURgUTjiIksI9yoRx0mwXWanwbsJV
LO3xlit0mALeBjJWHe4nSFQ/v3IB9//LUmZjeJ6bB186DECMn62xf/BYtGuFMefEfQDweGRV6pFW
yan/dQfEsEcPPE8gvF6K6PKm2CMd/NhGZSGXbYbR6w0jyw5gxAho2r0hiqBwyXW37LfFf3/ahA4F
vSLemLr71+k/qJET6WRT+3lh5/yOfKHiJ1ILufDkGy49UFOf8qaFbJJK977PNK2x12V2Oe4utfP8
z4Dw3QGgtdNolNREoinuvE4pa005Ec8R5fZsHHCxcJhRaGEaRZx3ENEyWUmxauEERuiIBk4/Anz7
psMg6jK16AmgTfmnHTjQ9gNsLQ7V2PtGtHvft6TK5Nj+FDhj3mmmYiXX/GTEfa/7sweFX5hPVM+K
OmsyUPWMLS5rp2dBL2GA6DDdOtzNZi6Au+dfUj8qLzybTC7+UBpuEWGkm5PDzqIBIjhq52pFnwbY
NJSXXWYvvwWzYrVdaRRTqtOL8dAr0lP6hCFlUZncNvHmAkxojMuGID06tYJD/kcqkmvpHVxkCNCX
I61r+4973H+Cel8HeaP+4yUiDgpSUH78yJItezBPTk3DEWCpSQOJc3bDzMJT3vy2rJLBrp09m/mN
xQKC8X9+QSmjsq4IKSxGImMMNVy2UhnMuUbW/FDQLwkNJo05YUw8msMFOdMWBN8jjGRL6z2bc30g
rVPr15TL1Ct59VvLcw1QXgNxpK0Ll3eJQgzoR2pQvIlfehaWETImSZyv5ipRYRavLWPOAeyJE8+F
c6F2Kk6pJVZECPy7XgSsYUhpFQSLFTy1qMyWoChPzdYR5Rbn6TEBrFdWBKWfSOojOvZGTJIdu6To
aYOwjIzIIqKthH2Db5rggV9gntpX3e6D8szMLQLJ1+nQSS4vwdtZ0puEU+xDjeF6Cm+RWFCvCUoK
kXYhOfx/e7RyuXNDN0k6mCH0pC3s7qKjLHU4t8zuQCWKqY/tfSvvs2SQ9Dar2VsBGApS4nGm4eQx
hUloj7LJ24JpLAH3qcxiFpH66bE6RwQNb05cIFiOSVBhL6kAkjrhY9tF3q2rnRApilFPQ8GLnSTA
OHGS3UqfVvovFFerUsrtafvN9/dhmjBGt1J5jLwqIfmB3ZIiPNvafPVkvH9UTaIQvZtXgvlPCAN7
Rd1VQ/8+bV7znqwdWQYIgLBGJeCJCrbQL6N4CQlnn1Sz+ck/SxOSJSiM9NOFG374S9hsVpKTkHJ4
d6mfWdN6bM5rbWafn0F2hsIRJLxzGa1J8v2higCayuiKixyRy8CFQuMH2Pg74TnyoZ9qzoh7FgcY
/9B7t2lK3NDy+Sv0jhMKg2JLRp5D2Irfy1tBeO53bFlAXCeE4s8IoW4Lp8RnDSolwzrNacmhPnEZ
BxIEK0MMGn0Fczxgyp3Fea4QS7UOLENO0hK1AUSHByHJOZ8eE9fReSwIT6ZEzujFbYbNLzbooBy4
vMZOAAsWeqI38FYRe/5P3nDZ1AK2UZvYVz2gclO/+p50J0h/OLCWo2LW8NmCUt9bF9Ooz9jwkYUj
iYKXPUq9UYbp5P8BtwQaRozbvpFjg9mjBk2c7wUvR33vovqPKAD3wIcstV18vlLNtN3LVmHY69dP
0Gd59Vm7FDvSSeTtNipGNpzxA8O6DKbrikFCx404kUX6ltddsdSLQxG/UZhfTzxD86PjrzPw3tf3
fz/Ry8oVRD9V8FjxLHNIw9fg+oJ2mCshGBmajbtktUyKl/m66qQzz5+8tOF9I1U6o8ECdqosQNCH
PtQuSil3A7VSn2E3cguq+hxDgoycfFbx5sZ23S0mJCk3I3UTJXc9NcpH+N+Bepkb9R6kq/oTrqEJ
4NT0FlNlMHsKJQJCkShbG0vN78Q5z7uvKYX3TpkgGlFd+NtFVLs7qvZtNDu4p4eSeVO6uxx9IsWT
pU7v/OSawGPgcSDAGpwFb1uOQEs16DLBLwpaBe18EaDpI/TaHBBZDXlp1kDPbZJJUi1njqaAYv7f
O5P9aJJFC7L7Q1urrpJZu711qosWSKfgShDueYY/8dGklu4SpP+J7pGPk2R0xhrKTbKDr+6aa+Js
sWZJUGL3k/l2EC5ZWHou2GRMXjUo4O1MgehTjbPs+o07tcFAWTgZHq5KUm6l7lsqAP8DHkAdvQJc
Co8ykL0r2TsbEk4bNOucWYDKomONUlhMzL4Ca4KWyquOn3mRTM6Zw4uGbBT7LkC0NOks1Ga7FpCw
edoBglEdMlwaxKIgIvLvpLNaO0+GuAEu5FXnUAZSUah8CP2W3PEYVc/takNwwq9h/Bc/umFCYvUD
Eh4+47v4OxNSJl0jS+ik4ueYqqDIsJsy0Wzs85zepkrjZSy6gaiLjRc+FbUFRl/UWgmmlBc7RoTi
i6c5sLHEEFsBAojMmhK+HKq723GAktsNYdvlKA640OHlhyxcAg0rLnmS6Noj5MqV06ROTga3uCo7
uRUNd5ywVEvPU6Z4fdRKNQlfBuYrtkefQ4eMcCo3zuw6MzwssdSVpGip1Bo9dKOXOwrsiqFC2G/v
EFMWUfHOOke16pj/DGhYAkyhovy+q5F6Hmn43F71Hd5JWL8mc/oRZkpxfHfnL8nLsRy8c4by2P++
vXaxf0vyuXlLtb9/otZ48AiPRoU+ahnp1RJXsRlcoI/czgBLjxJeAJMVkoZbL//Q5gFEjCJ7UaCa
ayfHU5rth32MJ+iGqs+9ZhXN/fzEuHPP28gqWoZBLjX4lNu19nyz5rwBwZ2DghPmuE5NWU0QgWCm
q9qpP593r4A2Hmcav0hzI850IyGaTRzh0s2uaGWpbob1gTKnFPkETWdPSA2M7Xnh/yn4x7oSC56Y
dupgEs+YahJQ2Cdmdgc9pFcm4YUvWMAix3wAz+ZaIMfWj8v1S88AZ1z50XWMX1EDs0/O1mnQpXqO
nzvbjr2BZ0sT0OxrdkrnXBzaQIMYdH7FntVPGhPZEJjfvF2LH3ttiS+W0H20jFnv80eI/f4kuqZ5
K32eUI1Ty4/DPCEkY6FVORGSsY4mU4ZGHdV7QnYzf4sTwpdnh73oAKxKTnFcujjWc9hkg8hiteAZ
9C7Ia3hBVcj5QYrD1Ugqn9jSJYp+0fA7xvX3HRFeZaUR96aI/mBCaHQEKWIjYHiG7H7HN9N6AG3t
LgmOxGAQ7WzE+T3gwyFHBcaIJjh+76tM7EexXL2LY5wG2oZtqbOaSF7xr2fpqVvbJwJXoYcZbPnW
82EW3mm4FfEa9rRyX0BQJp3ffc1yvq0gUWiOypWw6l/hy4cyLOCC1D3xlMiV3/4l5Qmm0WycJpFw
Z5OftmQitTXb0RxQv8AKi0cK42irclZd93+DYBzO+O3jeO/rwHWkie+FfXKqQtPoOCwrDXSBkFoP
cOtgest4jzsFN/IAcHkhoy18AcLDkKo+8xGjUYz4tx3F/9vsPUGRiTrlq2UALl9+WHnLlMxIuICx
boklmtjFfvhjFMEYIrtLyliAYImIlshwdB4EVoYE2IPPs7QhIO8PLCP4sHmukiwTaelpDJY9dTfM
Ny9gFrTX5jH7oNTjmtAVY42tNLAxFb2bBAFd8ToetnBQES9qYD8N9EPy7NlLH7ic+srtdX/pitNU
VRbXJNFyX2laf5CQbEIcydEYKgVVBCgZWYV/zkj2jGJpqzQgCevmMi6yiDrjqZhmRMRVdggHzRlh
rHOkDGDDDSjgoWaOTSBhon72LGuv3NcJwc0xNGd1+xIp8nIChw+PwOah8G3scKJQLcv1ZBljrCAg
166iOfHPKcyxrlAvfJXRu9Vy8RqZaGPiHuuT8v7pMckP9NW2+v6t2ng6X+F7VoczfPCVLNRlN74U
Rho++dfZPsBTmB/RFG2dYIWKgzPbaeuypw2jRoKyOD3ULngAK2bAdzFhym6S5v+OC3TR62mP5Am7
7bOidVBZWSl7OLy1ank7QC1XeRFFIMF4lw8cdo7CpG2mu3nLq6yTyMOmrJNR/xzb0gvNYU6gRIsJ
kbmVz7z3eIUm7/TS/Gf+k0OUH72NeDJaB/aFRqmNzQ3HN2QntacBqtKPPH/Bni5Rzg+WSq8eD2he
CY5tU1xDgh+/D51hlRw9RWQT2VUcmPjX/rIRFcDznHGHeTS5LkvvJB+WHngW/JP9wCb9yFZI8/k2
T51vOPigm3W8wZr6i+dNklB2nhadawWDj5ZetlT5KYqvUZGUZQqORyOGrtcEz/Cf8d17MDbILA93
1rKXFQIxekl5OE8nJbZsnjpnEq0KRV38HTIAN9lKknUa75rEAbro/zbOfd1QImiRNtY+bMAt2YLi
07+RfFx72kLH+tjly7puKoWYKXAiirjOgfINCerClvYkMvewWTZXZs1p/TNJXdChbFBMwX1gP6AV
zjdAP14Lfebv6U6eqV4uP19adEx5y+UWRvqsE6b0tKDqURAys65JmCNyDkQ3dkIDs47YEudPWceH
1gX/BSMrHCqqun1qz8dQBtC3GETpDfFUFA3PRJ5Ej3Svn5hOIe8rDH9kieQOt6In+TGithpqTMNS
SoL1wTmHbc8qomf0fUyFZ1kUtSjqbkO2fPKMWWMV37GdG2P+VpfoYZnbNjgRzn7DQTd/+2NiwfhX
0PmDTBTTc14zuA6KTYYpKhEXXmadoCuhv51FNX1BGqDMMESv3YSubw211XjDBAAmJp8LbteM8hUb
AdTEh8DwCdsmsPxihk6dLHbEOUmukeTZr11hk/LIZ/Ry2Msg03t1sGKHXZCluzt1CklMCvLr31gA
+2gwhcc6IkmZNODkZwCvIi9RWbGQXCHNGO0YER3D8TenM91iiK8cCHPnoILPOWG3zX1kLQ5jRFzY
vK5bAPCKMxkZ0r4vkIxttiAanxddn1c8vBG82YePygpvZam5dJiaqmr3LzVCCUb6fXdySgiqrVop
BRPf3HtYZ0a+Ue5QC0m2x49RENKUN5Q7RoQuykgpXwgBXWUq0oUKjURoqGgcY5brKLff9h3TUxpt
iL/JeCz52W6BjfxUm3M6BmIFiWBxWOj6r9Bm8ygbHZ4uBwXF2V0pJAdo9FQ4DeCG1sr1Gh476etV
1HC92cltg2nTq4FZqJKzRV82A5nWb8H/ooDENq3daCu0wQDvGxEGksMvw7K2J48FQ7HE5g398rsN
PpRJOWy5beW1TTM9tnEFKVPa7Ri8dUEKi8sfOoUIjaQyWZuc2c7hjUF/Y0vEkOPTKGasCdL+5/t5
ZRsVC+GssyVw+Ax6pA0TTWMsdc2+YR0Ww0J8u7H16/aUjIQsMjhg/y3jPOCAFr6bMVb5LGtr+vJh
I/MVdBNyy6o2aKogc9VGTiPduembUozm1STvwQTr2ifG5DllROnqSeqJAQWNTx7E1DcUXrVBcGZp
2TjK2oMjSb554aPz7ZRzVACZ5hNNtTn15hdYykuMXiLmChNunWu/1dqW93fFI1XSqgIOjYbjkz1D
79Z8QXq/JGv6pEWmjcF07FESFC70oBd0vivCRKf8cgsaNAouEdhsohHCtHOOfQkWZTp175MVoPFY
WwBaPuqgSblQbiO7UCO+sy5KqFtpdvLMe8uzG45cIhSKTxpnsWQt2HI5XYG7LVnSsrUKxaK/bk4s
UsxHUVHC3yN3IziP5L8wqwzT4ETQF2L+VFWbm7zcSDTcc6UlxGPfLffEk+hzV71cEuOA+dgUa3l9
MaDgGhNu21gTf7DYTmUvxsn8ITfjZyDqJm+Lfmou8egaiPDv2fNRe7rqDvnMI9hJeI3759ULBoKg
xUB3q0i5lPAQ7JF9LGkFl2jYrVgL+vaRvBPasTLDNasBGAbdpBGB3BXVrKEeMi3KPzvmKc/Q9jwE
tt9fwQnytwrNkgyS0nTdjRdLWILCCCx7b357lBRRnaiq5IzBIC/SZf5lbOowDIRVLDcXhzZinRTH
W9JHF8wb7gUP4opAsVmE+p5T8j7N2K2R1L3aIKGFsexa95SJMY18Utry14EgONsluciy2u9yUZ00
7RRmhWI8MF/nfDYBMHYzYgTcaW/uM438ClNsbYEgdUBirz2lKVrEnajgE48XWKMOnYvOPVOVGsun
DVpheHZIv8rT5nx5W2fuh+pxG1BRuXBSP2WJAMy07dNTukMCDATV9NQ0WUdzKrRwICuyIedPsup6
/Yx4ipqDgJYN4U23CMKo7TY06/ZPRMXtvWCWTrs+7t2if7CV2lC/5W0PQQMu64bcXNTTV0RC3qS5
ecEc49hZzWDbiA73NTl3xuT06tZlHEaknEGLO8Pc4SC0d6hAIPmkzJQrvAwdgKfwMQB2aBdo/yjA
IbnWv6wubrxP28fE2MLw9QhLjJ0PbqAInBYjbMvmNiYk+9LyKrqrIcnfEbIzS5ZQix7Qcn2t6c0q
y658lP2dfQz8bh9RY9CI3G08qJLu4DIQG061pg0x/oSJAsGuYwy6SiYn+ToT7bu2lv2zUKGzvhVC
TwlmpwsWMPDlwrjJzkX89pTjKm+kTlofMasglJucTHLIY12qMCtqO6XU8ypr/lMXz6agQkQdZ3Z8
9JxtowJuodK2TAqcJd7uqfGHRAgxO4duu8y0PIcKojFhQBM0Gvaaj+3CtJzaERRgIgfWE/bmP5O0
+CulkwO5doKKFi+84MRPgsG3RlUS4lb/nddW6VyzM2DYojPnk0hMezXcm1x2VtK1AT6kz0Tr9TfP
vrcIgwZ10rT9Kyj+dwA1NZ0W7kDyWy908mEUzFY8HrbYqlrmhMPiG03PVW3dK9/zZZP0JyvuMM+E
ADA2+w3uvra5E0p74z7k07bjjbziIy/6b9dIw0tlkiDenCM/bab+qlLLMRLUsaV7xfPkFR+Q+p1u
IaXdCLmUy/GkMNYbTsF7CgufWqgArWnCtFInroOhj7NgOYcyGepleeYUSfpdp0xJ86ALQsumSdft
QCj7aR3UixumPzPtiZT8yOWkGsqs/Zt/xe6dBa5IQe6c6gtoESnKL3M/OSrlLKnX3HgKReBEaAf3
BFksrhT0F2A3vz4Rf2m9t+21GPYn5XbQJbRaZhf7QftPUzidtuPoubf113klqCZBJoQlragK9Gsj
/FWMsaHBr5b5aj5sfOpmutEhjFExJAuuqls7nWPk5CPL66QEMarcQoqqaH7QOUh3Et40c8+qqsll
QZUq6NjJt+zWgUzO8GGxj0fKIuDeF9HaKXCgcrVGnNpFApxWfc4avWL5Sop2FGq6sJhu8QHhvN4J
J1e3SUIBxuupJRGMU+r/vm8BTA+AoTlxN7EtbBOKbIKqkFdtFE4UXJ8gNKbNhTadYznSA/KzD0xg
PpgIme266pFK3mKLhI/BvKDDBspTufsz6qErowmlI2XYQO0q2hXzkpi156yhV3fwS7WZiYhq3vci
MKBx4JZImNHbMXtziAwxumpz8Myk1Os0g5s/FnitjB+xgZXppyKG3J3WEmtRR43nZomO86q+9yl2
h/ApLHG31LmtdQ2fQ0SYnJGvpVsTUn39K5jo05Ebb7wWtL2dHcF8tEsuV2C146VsH4Uinn31ExOW
+loO7vMMz/kRO1Cw4Q0Z5LZ+gmFitS0bt0x3PYoOB9Q1o7NP5VnmxGbUmkA+UWLFTMkrxZZCmTk9
jAhL/L/oCVWh2JUNs82K7yXvHk7nq/f/IPipPCJU1NImMGjiEmT23SYjut/r2miN6bMFhaO0/GMQ
T8LH/Pm2mA6IhhVH3pXPitcws80B/akB/frWFcVu7oZytL1vool1XexmdB9Lin1HgwQU4xZjuYy1
RIo37ZT4baFGIggAQDckcKoSF56/25ZUxFifKpRc23BVUhtSKT7SHBv/qdPI6x2o9bXyzyP7Y0sf
f0K19YXDcbvGpazzcQ3VFyQbZTWwauEKmxPvDEYfsvJAbQGxzkhgI/dQTxlY3206u0yLHe5sSdll
3iAJW0vFZyEivYu6knX3V6Wiyb9vqI8EvDMbpsx9yxrTual5noDUrGu/Y3pmXHor63Z7f2dfbfdu
ctyVBaoPMBuX/aZKGdbYByCQF9F7kXO4DdUW+q055eQQ+qPLyIuFG2sG/YE5GEY2BT6NBE0JHae8
JLNczqVRK3hJSNSwLJvx2pSrNxYAiaAv4MnEjLUpveG80aFWL4HLVEHxfyURz7pqXdBIltmzQF5s
o6cjCTwRLdFOXWufGG/zzHtrYvEk69hp28SF35+vxDslnTZvmdU5DiMxXVM6HsoCc8eCIrfbDP5M
zcKYycQzqzXpMXOojkP4X50ZnkDsCk53ygooHo8NQt93pfwjJWZZUPy8vyM7X0cSJ0ZOz/TQ+G12
Yw8qOYinncR9rMxVwIXhOvgKW6oup+ZgcExhNj1BUHMuJoY/gQdyTvAdJgcI8LmM35IZUc+a3r07
xwWOCd1v6my99beT1BFfAzqI7q+tSZ3726IMqSnBtji9lLiKwtPnqgqVFhrRePJoiV5v0xLfU6Pd
yu0DRhjy5i94fk/CTldJvkOYGWt6tcbsVBYEw1Ej2boJaZwU+FTq6eOp4tmuZufjJAO0mPDuF+Dz
qbliEEIq0G8f5zbjlvaCPQdLYRGy9BW5rFLoCB1RkDDeo5lx1f6HHDXmz5ghEczqt2SJsHuBhwzi
ni5+4fOGRBV7WrOSY4WNAiaov8+Hyq7S1GXtBkxhJxSLeGO9uGD5HC177FpPuuTvYfEb0uoA9MA9
xDeEvnrIQFX2nHIhh6ppZpcC/m3koHhvQlNziNdnxEhAzLQAHaa4dudmU+IUv9M1yXuEkeNXDS7a
/jxsaLzN5vHc3/loM7mzR6MgBug2Z4s4ZlBkaJItt8pdavgAlu/vhWVOB2DbuoYXazxmx0qoeUzo
rv6SnrwkVXUc0yH/N1yKv5yU/BGE27GrXVTAM3PSXH6H1e3OYlFkIkJxS/HM1N+LpmgP/zmBtjPs
PvAWoc3m7llSXknf9gMJKjG+l+51NDQH4KFDpwQoXokz82dwkQTZ0hIZYHQaLIR/8FMgxHOxq4ao
y5Y7S1GHz9SeAw30J8l8nWZ+ZE7qpAYKndYklDTsfC8v2BOMsIJoHnktkTc3c34hF2YXXJG01lGs
e+oytVzrEHPBwoKoNXG0Egv7A0h/FeySmD2Xw0pd6zFGS24eg/b1opTFflhmDSh3e+Es6ZcVbXqc
tcK4LVcdb2VsrcMukGqafDwcAcI+clYFBZ2VxvaqO3XkctYE9wLPB6CnAYf4Z16vv8Hgt8SBD/7X
iwhjS7gRXzyeV1sH75Tw5jYH8gI6ZVEP2FynpK1ps/J0cV5Uce5Ui4Mo3KiAkjhph8m3HcmhHfxd
osRZ98CslI3x+rKa29VS/4Xn7e8Mj3glp8P5Fp3Z8tj85pj9ENpg1AXJozZH4NoAgT0iMRWTgWRi
uL7Ncf+bfV5cEIw2ohKwbW1rjMWG5pZpHDZOIFWTZu94YPOu31SZBIeTi3ttUG+VHEhqBKjBWBSH
WM7mK0gDX3Ncca53uy9oYE1dssLLYHpc6FT9MX853sqaNya83C3NbpSpWR+nnqG0ZyOf31z2YcG2
hAPfb0GYaOa8IIrE2MQ3HLF4qw6pTq82rvxhqeJcVzN7pq0lwLRoyT9KOFB7qtUB/F0OWWiN+Paa
lkZYkLo1sgRRsM6841gx+vRkh+f6KLlXD9NYlVipt9winRGfVC8iV/isKpHWPMPU2VvbSQFTVmPP
hHUd6UcDksQEJEim8/nBsOOlJaV+waLM/4NVmIPEeu3v1UWklITwbJvRkGZ1T1fyCrqj+UVaiZPJ
djq5CFINsc25bDIUEwlVHGHoBIIWfwfiF7O8qBVk+nXaegSUsftEwTg/FueDU8hA8ZnDn2ocomPJ
39WZUHL2uGQfLkM7mWkSt55Pcicue84vArEM6axSeBxOp034aWPscg7hXSaGAP6zxTiOe3h5X0DT
xAidHPtARX7iFPB5QpiGQCC5taNw5wXN3R4DM+7Ird5wOKc0hRboHWHnd0trUEH7RYt7cPn+J0Kz
KzMuyu8AG3cqaSSZVpCbDw5vN1Zigx/8XLS2DE+t5H+cIm1O/a2xbdr7b6DddbvTI9rD6ydXFbgU
xVqT1FcIymWMFS085xcx2vpYyjYvWoki3BHFVsBdK2v6lp/VebIvTizcD9mprtxNNIP6t7zVyPcy
k0YZGZuwj9DrFV24Csdh+vcyaX7aUAZZgi1GIdGePTD3DNgVTa/wJqdMXH8QIOuR1mWRW7kmKUXI
MTUkiN+rTiYKrDxYl9MPmynVmUofGT+otDGP7fsG3ZPl4iuD5mUQqMYFtbS1ZlXeghgLdw9ahSsW
hvbH0OLwC8vzUR6uHP8V8oqZa06Q/8HBeBG/Yt5dACDqbsIwwW4ES0ZKkUY0CnE85U0v4CQKgXnc
ZLXhyCA02l8VARaNcuc0GTujxp5CyeSGrwEQtFHyNL0x+UMRnQ8kRcyCgSc/yLPFRt+1X2rOJrJ4
frDfTBPx+fDm5mvsGr9UOW7GM+SfYEmZd1bcl33ynfefiIPupzGfPQJQZ2lmdoHkB9MefFkO4ag0
VXWE1KIfhfJHKCQ4abasWgM3avru1er5ITr3N0VBkQSZm0JfVLcSeHmFA3Lpe+xea/1tKCQM3f71
dsxXUiMYb2lqocO9BtyVM6E7fwCFtssayW6oshaaVLWXeJ5hFeC81YoasrGvRGJE+kfJRS7ECkgL
gej5JD8/y5tgufXPMjf4mqWwSz17COllC+h+jq7wKyXR4zR/6mpec37WI5iWc+udokDuYomKHYxc
GlcR8P5YmAZXoCNHGBwpj+tn4twzAFfQd16HYB8KUKFGgrTvomolMjDQr0++sA+gcPCfSUxPuv9x
qd5hcAaI81zbgfGF+xOAtg08gdJqkKa7ZGmUbdaoIJmvVfDFstlBLs+ZjgMfj/mJT4K1SgnYw0YI
M6rsQcwSYabGZgotuuaz3CDz1E9dVSdyUOBHl26GakQ2d2CsIpkb5nkvLycyckkmNFm/3MkSoQuU
d95Se/y5l9OMRAY+5k+eFabKYtuRD8QfKBs+CYQUyuzTxI6p08tOPKhF0HfkCNLueSpCdKaimmI7
I6C46aTgHOTaebN45aHW4r1GiKWg/tQO09FlI0MwqLryuzfeVez5h+ehMarID3aGmD36YHRdhYjH
Hy9aBJ1IgSmQ5TADQ9SmVYqJbKH83jVmlagTbg0DPBGHPCdc8gWp+IPuol+JBLfbpVqBn+aTsgcz
zKl+vQ/KwZceJayzhoY6J8x8PU/ZqugaHKXGJpsuNmQZxwy3BKGwf1bHHF08UKVtQ0nNjSjQrhLB
f4KKhFgjCD/ntC7LTMdr4hNXGhPp1CLmtzMwFtK11lyeXqjyuamlm6kpnTFrfNUqOBaMHRS8BpoT
tHg+yvp1Lt77S1ctH/YhMONSjQhLLd4Jjn0rIYAuBJHISlNUd94ucWYct0PL+YNmJLFSikz5RXu5
4wHLq4zdCDDL2IUv8wyHr8X4hl7RdNR3JM7qLqn5Ik1av2+TxsgwzVVbranWPv/lvQYf8J+VDpzq
rtCWJlqPZVqRzaL7LhfGtCvl5T6RdzB/Lf1dMouyqV01vPd7ZP7LeTQ8ltsj7Q0dWI+GgGyp/7d2
eHDg2LmAkIshlBYpnPyd7V7leaFHYWxAo1KUktmtq1176/qHoWKTUBztosqYoUobP+aw6rO6zTDA
/xy+i+Cdj6bFmQVEjvpow32MV4joaaCvaNGO5QXHH9Zivo6TYYlY4fAnKGIk8Orhb78irjNtf8te
uovm3NMhZfDUfUVHDeSBlomJgnyg25/QUJpZYghsxp/hqSBAHfdVK3k3Sirs0SoNakkZ7uWL7NQc
aTVymOUMwHsnqec+fZuyTh/2iG6a3au10ISBJWetsyOPy+gBMzomk1V2IAWbzSrKect/lTsTODgB
TnJDrVUu+4JaPfLeLjsIfcc8psQ3P15xI+22FEtdjYqrJ2C6w0nN9j6TCe1nR7/K9d/+HuX1RZuH
HzNzOW+TMfqVeDH2VvhToDUz2T+uVDKBZyQvYpYjbnJ+T3VdCWtLeShDpkgCyhC6zrNhMeVmC5MX
Z/8KE+SNE0EdBTAD1owH4Ym4+y746jOFLG3rUD6Woi4E86z5Nj6VICqSWAqkbNv+gQm7oF95ufJ8
3MjnvCCcnm03So9ZRwMwQqE1uVPgejNaEAev36JWSWB7VjBqHGOuRXNx/SEQbob3gc1HPThRrXHx
XL8ml6bNmjHI1K2CKPnFR5g0p66yDodM7yuvV/zgdlum5f9rfgpYAWUleEHpSaywD+cIWH1WkQHK
GF20MD+I3Nc/lfhLNYL6R/l0f/50Chja2+ghwTku/o9lcf6Go67Wfs8Tb7ZrAulNT4S2YWHClZx6
cuhAQ3zAT8L3K34Q+POevWdPAjCDmjY/7tqzLVPDUk9psFIdFj4WEE52njcA8uWMbHhxpKJ2NNRs
xkqaIRxpmRiW8JqLxRiN3Osj0iIAii28Kj0IO+vvD0Y9Np7VgwNyeBSPM7V65ueVq19p7RRRYtEE
eZrpbDdlu30fN3hBiNwCAzETttaBg0TE4J9s5CsNu5slwYk79YL2ODXPqqI3mcZdkcN3cWAMrzXQ
aVJXWNrsoatkiLxh5TAv6EY5/zomeJwjv9J9kAkSPZnZlZ1WcvvRKw1FqkCqpOfbOY9cTI83jFUI
9JkZ4vkfgcrGKAE2MlrbINtN0y9ERnzUq6T6YSdyaOEUDYqdRi+aBUmeKbQ30Ny5icVDoviU4lJm
/V+xbR79x+tKs5mIlI29bTRQqN4izGjnAppL8vjJC8oquZkr+TLgiwY7ZrsL+ZofVoscfdBD4XjO
H3/Kx4s1CYhDIQWehMfS3fEOFzM+Ll5SUjONh8ck0dlywX5IioPzyD97BpAuALzcSZieVd5GOgcq
G8T3eopZvUyI35H84NoHR75YlQQKlI+uhqQht71kma7HcLHvru/+xAEuyfcWxJFER859KbUvQRPP
OdPZeI433shgPm96F9BeHC0/lUboLKaB0SooZ/8cnwsVzmbkz/yL8ot8wZqAfEjyb11b6m3xj3Iw
ZsQQrFPbiQrjvYPTly0dUSsxeDrNt+RYnN6j2O9rfuLnr4/TGYXa9yV4Tb+a6pzC7ZC4P++xxf0y
9wYat57OowD/OKPDUjEO3CPhYrtZyA09428E6QjsNj448vKmSXQ05tIGuSzTC1RkQ65CoWdV5BXH
h3aqTjhkBZu7d1bxeJQxsJufpC/bL+lV23ufzy5UMZTG1CL8Hrh+d37rdCiFR8rtjRAIcn7LrdEJ
Y9S4akb8XCvV/Uo8iyFFsUMlKGZeL6yGY0sjYhk64JsqCwWGNHzBU/NppVU421xvKgkil47TaD7S
+D+yad+da1tcYEyhizpa+czRzj7adAIxcOiwh22in/HsHbCnkkNHXu5eyfBP53zG1TIKQSkmWgjp
O5zHPngzkFQsGGK8Tqw423AagAhw712gl4+ipOcqdp7CEzquPy2Cl18vNjbfgQpscBC+7644gLzd
r4GAaUu3txFxWJLLI6h3mSF1XbAkCxpvfx70kkgCpuh/id3CSYxmkLQG45nDeludn3FGYl4twW6u
inauqMAl2cadPxTex5mYk1EjaV+lVE7h8+DIBl2rYBBuv5m+2GDtfepw3TMf1X+gOprMp0ofFH3M
mqiTbgRcRY2Ss3aq3j3MEr7blJkdy7u716csfQbDL2UhmU6FsUKL/TqYM/l8bY3eAr5NFVi1A7c5
89IswxtUBMw3OOcHT8HdR+Ky9O9JlS4pOlWKFJROYHVzbqa8uGwMNkU4i5llhq1cgkPxh9Nx1TSr
pzlul79/6YbiLhGSmL5xfSYbaQhA8FjCAJGUPosSu3JpQnE69dCy+Tj7xp2+jdElkuLfReZfQC4l
RlrwMEvaF2tYkrulX/PIuTxRLDm59FwpzpWN80i3y2nR5SeF2mJbmXiHH5D58Sx3Q1xcNNKw1Itq
D5Xzk8VmKTuY+nmzAnVtf7vOABM/Ruxm4VstfewRPLjk02+vV/sVtUfJdcJaeByGN5pcLfcm155E
KtpmRXWTUw4MWWzUEJZV21umikBKSl5VAWX99VJ/8iykFT+m9+sakcrkfqg07k0D0nx6mn9+wac4
/JOM88pMgxDuZX9zG0h+j0SkmeExL6dR+gysXUNX1zWZ+0/QqaJ0NqFPggjKJkJ2Ntck4xQN+v8h
0Kqcq6dqdOmDTtPfl2eVCRFehDSbq2fapZkH8B0RbScaQ99yBZm5UNLrIDbqf1774FR3cZ+5Vbzv
ZdkYDM9pIPXCGehd/yqs6ZKEeI3UnN/C9FaV61VFtRav11jnnL3U8sifu7IqDN8brveqXiCo6dCe
tvrfaw/0DRxzVha3jbynZXST+1JRmO6PsTwhGUdPFdi+It4E2f8q9iSyxmAfosdqwI7gQQcLJLoS
FXBERUp4cu6QC9tlOYKFEgmeS90GiLkhjvn1L5gJ1Qwx4EQu1UkkFdB4AtJZm5dXCcT/FGwB6Gjv
vyO3lVhHP5126NUrlpI46ZEPZpExNmNCI6+2vOtuMK3emd5WkGBCTnFtLxKHa/xXRLr1hYv3KlMK
OxYjlbSarHd0XxZgLoi9j+CbAAopj8G9Z6va55qgXilm9Lzf+6f0jKBaQHncMZRy1+dY6DVclE9v
EfIHFXz7mo7djstXNDRQuq9LMg/aX2AO9o8WKvFve1Q/AsB1xHJpmJlCsyN24aywDp3gDxqNqllN
JhQoKNc29J+AkHRbZkixW2mbIXwVexL8FDnGScGex4V7ypJq214bHNkl0tvmGdV9TY+X/xwTlVzi
FA9zYe5d+QERSmme/J+BQujoIwz7ykDhHS+cHhwQ1bNmjDypAi1N50oJuLxj/Dz8Wtwbe77P9YlL
EzR9dEHU/nrwqhxPYtd3eNiNMEg4VJIrwgCjjXCW0Balh74tmeg+6yaQBJuI6uGSnEECJzI2irTg
y3IJBey5azENDNP+b12aXQuzwTNJoPCV+lyf29E6xj3aEJTw0W7QusI4vrfucTKaoO9/TrEG9QAw
g+WsZRDtiKsRErXmtrtvd1baptbT3DLnan2JmhcxLXwg82GjwEBHKty1pHAthzg5lvJhScOHVVfR
MWFlzex3yB2YsQLWvnGwLuuEWL7crn+xnAJhZxOcOS4vGxIe9227NAxPUQWKuevpV5KMSYef6+1p
uz/tZaX88n5x99H0JT/uiXds3R0NnS+XA2+F5FQXJlogxFHqjY0G3GppObwg+61+hiALSO2+wlUK
Fn9hgkc+bnTLM7wqbryNt1Mzu8R7DyYYtvvzhnF6oHFUesUED34bcQGFKqcfsuXGzW1IuVyLODVp
snYW78n2MDWK43g6if8wLhuj7aPe4g8DyMU/NDeRncnnRbs0BxXJHOLImjOzo6wEvPxBTM2RXeU9
YMLD/h+SQ1CfLl5mK01MehaUyA2HISMsGLI4SM5HyqHp/zjX5yWcqwoZYYmFgFv9w/5Vgz6T1+Bt
Ob/rZ5NHXgFsrlslY+hvm4CvSMLvKEeVSkCAqRQfgvwLrImJy4tQWmGaXnx1hxoXtLJwVXwv79DT
ivRL7BrT54OQouteI//7m773dqw9DOP0zJMuK5MiMpZmllrGCNSYS7rtAIpM07Uo9gpOflp1t5mF
9UPKEv1rgpmCYz+sBU8wMN1wn9fMQAVuVoYBvsFEj7ietSrrVdgM0swI4SzYVthyyUbnfsUA7wRO
Gk5LSKVAYK8QBmF1XhJPIufBdRv3HHbRgIvVGCaCLioUm59UtMKXCSWcqG5TloTzBniyPLyKJidl
5zKFbgfccYf9yCOakxC5PoCT3gKChoeHNMNas4OUkK+qR1jI6fxFJdYnRVO2ZCFXPryQ0jruKffc
jJRGRcS1Zx/E6by2nM1DKMC+x/ggYC4AhrEJyZyJHT6tgA/n/YVDvfAWfNvUP1AC8o8a+bPfsv5A
vmeuSWhzXz3El+4LzuZrIqzlh91Oumjt+Y/qIElwsW2I1oFDc6eHP32SacxW+vg96aCAbCipLUzL
AcZUu11itorZ0RWNFW1CHMFR+OAnbGRCTJuCaT2jlJuXWg/lroGhtxZ6xsqFNRru+CgB6HrMkOsL
myWM73ILFuJDyXC542hjVPhe/s7DAyW07QimGQXwmfiHbfV+B0vUmFMzBWmqwd6/m2OTgu0zRIFD
xm9RUVeua4XaGsThlrmMb6Nx7Q52q7MRpIc2LZFbz9tnnewjAdg6ICxP+v8aoUwXefEfWJex9uKd
evJtVTFmTWHjKMjXY28HIxaiCYxqxJ2IOn1Wjpbo+BAzrgdSkmPzv8svjXb2wxg6aNyk0Dn3YbX/
x42l7CkcSU+YYoIAGvSHiFgmAtmVzKum293j7GTIUvZDEUg3wskYrZmbzIUGHcTDjfgyWot1/UWg
8fyYYQUNo6UJ5GwbaqcO914/RIosu7dOGfgTrQO6d6krdLQDWt/tnV822K9vR8Wyk5ElRksk2pCz
a3cG5YyQ0R5CLtuz0rIWvfjGYsvc5ZIpaB2qXy8v8b/AfXcckvG3RaQhqLO11sO77Aal4LUhx8me
3usqjVFBWKkQ4FYajTPzi8BLUolFZXf6RPPHy5nxJySx0GvcBKRngbjNf+kieG77dw92VK35DYqV
UQ0YzwYW9A72EDje/dOa0EGYBpaQ/NIc9/DSfcNRyQ6783CJNAQR2KPvBAVVDGWd+Jjyf/UC0GMQ
kp1Kig68rpDWVP/caNeZmo6YTZ5XOIaHui6MjQebJayPSkAOEbCjAifUfJ77KWwpHW47xULe7WtG
HNdIQskZ1VnX+vEDo8P2a1VDk8Dpg99AIOFeOxM/8IyOLUk0dHx1lm+vV7pIA1qassQ8AcJ88jJv
+zAbQ3rKdtgwOuuKQwxybEO6s3sLZYLsP2TP3zzJRhjo/dVpuxVyyW5hifj1cwtuV2hu3XwX0Qzh
RHk8iC/i2oGQ0VUjsR7WeaVdIUb4cr2tIGOWp9Dt5jYVrc3PFmMba1uCu1caXfr5ZJW1M56d8lgS
YYE+FJBIpjVVfd2zTfQtDGMpRQwzYHY+r2DKj97HY71m++gi4wcb50sW254pXKo6ASLJde2yxLxW
RQwOMEtil7d3pEH1A6BgQgT9vKZLASMEFMjxnN14kd2ZjTUefZ1NL95zBWEI6aFSW2csGqMpDoUP
9VZON/PCKrRFod4Fr9tUPjy9wHDWQHQpX2psOx/J/KfTxBiDTOYlfnw0Ml7OTUUUraKS5gvJ6ZRE
Jb9DBg3Z4azSfbCyVHTzXFhzoKik41V04HNXewHzhCYfQLdCXZObLWHkr93AW5WkAj9tKSZfXQiv
bOVfs0lYAleBpww+So0M7tDB+ZJzQqPMPvwfKW75TpXUtfgwXP5DiiCc9CVnjvuPqb8LJbYVUHiX
OwTsY83o9DKgh4tHgN8mz7+kbrumUnGJyNbP7i2RgQbir8URcakkffLXNI79xbdwiXmZcxKHkJc6
Ig7Yn95lEZFyDc9j70blLUn4NaTEQcsZYBNIbUB+zvT0anttVtZg4WSQtJ8oy+r+nS9geLBwak1O
DlNB5iMzcSAACWYiH5KgzrtF7x86RjIosuJWJ5J45unprpoch3HhnT6hi2GSoJuQcsn27ASQ+Y0D
oXpxh3ylsiXLyRIv6CC7WrFDZQLef2mnhp9cPn9Vix5U040zapK6gUDgz59ALPg38sr2sW7vJA0E
NFTUQEXMbWOgZJqC8tcSHhgiG5c1nJ9uwvwiI1kZnXaxVtCrOhD2VOHjeuJI0g0nEXUSCllfGrhQ
rDKsAhSe3lX0yOHu/VOYSKK9Gose12zumJ3s15vJraKKK7UE0vGPA9sx3hsTeE0CeDu1jfdbE96B
EUARe/s2I1YbBY+/QUf0WWoEDUrQ2iUiMTIwcS3zEHeMFMmy8Kez/p6ZpSm4sk/5e3vDQJr8okJO
1x4jGUttLeKPvzBsaNdEIkbQQIB8I62dJ3/La7D6qmBFDeIgP5U8ldmZTzeqA1actjjo999DfAu6
/eKGIsa22UG012vebEguxTplW4j7/RSizgf8tQ0zmzzcROqLfDNknCez2miHVOUBKtgOe2+4NrFi
naL2DlILcT2mchPVzW79+VpEmft+TM6BVT2N8QiBWbTD5mA1rEuizExbPd9nh1Xe1MxJ57RNN/ru
V8vMOn3UhAdIbSSj+qQH2SMlbup3bpF+3ATYIG+c8qbSOY1ClB1zr0Yhvx/3UAYlokirdiMwDc9W
mrtM7i7aGET90W6Tl2rmm/7GCffGypVKWWXbh5m22WTMHQzbTdaqOBz4687Vsgs98Hq55uiuW0pb
9P1EKqi93/yR4qaAQls3rN3CjcTV2MNdCMReIyIzN6VKF+rOYI5UUQAErndFlLqJkf2sHXrw+tMI
q97qgasHtS6QJmO3yDo5jfPb3ybznk0g9tlQEMcx+lfimK6yM+/UjFpD49mp7pwQiuRayvm4J5zx
+pUsTkS7PXMbMvwOP/FuPKxXbcwzyq+NSBXbCeDeBCMa4/Z2I/ovt83buWfhr2AopS56q8NNmJhB
AnxB4JL6py8b+uXVTa2Juji4P0SQQ2Z6gmiog9E6F2smkv58klg5k4MRXjmxhzacl2yRckiOd32P
NI+0FvRVdgE2DNDRkhN0ZR0E+m4Wk1a2aMIsybtqkt1khOBsrQNzhSBPVOV6GBruUdficC4A+KlN
ZEDMln4Way9s15+CDCwAPX1QLgORt5PMosh2cSJEOzYkD9yBaW8izPIwoA3/uKn7HkvRjRGa9CBQ
g3z20wCQIBZM7qChSRhgOXHJ3sAW5M5/BjlrP//nRZO2Nx3uHwn5Fx8tj5WgL1KkRXOmLR7L1BEM
bN1xwv8fgM1OVSvE/Dm0zlQl8yZ/4AF8pRADeQhltPCrXKGNX+hiAyW3RAqGi7RQdFxOmr19gdbH
quocCpp7Fx4ak5i2AgW1CO0RrSqCCvLyW/Qc6KgIQPWcXdWwaNBr2Vulasyvzq7F+onkWfFy7Qdr
i5JrOirmt12lM3HejV77qpAFJT2PmXyTGCECW89rnaVeK+TFzNbs2YDVDwLJYXOcJpx2vHGfBa9+
kH8a1zHNXug7DhoRQPRGcjj0YoA0/hkNz8FsYxPmSUrkCqKwal/hCXmkZyQcPJErBb76tmj0fYx4
MpxOkGdWARrMUtuuM3PEzREieoZ+Ob4ZgjLXl+QL4RlzTA1YrJf14pSDnGU+yZ6kXdeilUZSaOJd
7pC4au4r5r8b774SwIXX6x1OyJkTZ+LwEZepkdxdTCH3hk10Els+Gl/aT8R2CsHlrcAiCtxSJfd+
kWIOYvu4Oxj94xF8yJ00Ekv9bbe7FAPkyRg6URARciWqmYowGw3+3FDb93TjQcesQGKsjo1bcO/8
oCeNI3xg//VHTdxJKM+p3Nz4gYRURhCLvPNmrDtLfUbOI5LqoC2Am4cLCS0ukJntSBEZ2ITjSnNy
/vOyRfsUqVYOqk5i02kHZycJoIgaBAXmDx4e1g3MCmlY724AbgjgVxnkWNp2qO/ayE3C7opWGfYQ
u30DqPBEr0Pnm+hgagUoe5J77MZHasmsHUqgxqqVSDCidZTrdv2b0E4+fl/qhqt+FFSlpjHihD7K
ni+PzCNZRkbuY0tcf87/bJUed99Ts9rQyEppZEC3TvLSrEMKQatrLuAfwvnZnrfKoG4cSoZ+PcPD
vgeuEk0+t3OTtA55XEu9N1nQ3IjGNNUuVZQw20RC5cVUoEDQ3W8gavWQ2RzCD/Az+jgpr2iYKYsZ
bw09NsaQ3UYKHKCdEexo4JiHN5Cmc7CJEL40FFekM1h6JgiNnV+2F367qX76AFFrT4NxPXIh10A7
qiQ8V4OK8D0x8LcUhhWs77uq348JAThaZPWYNxLR/p9BaKS16+qtZwwdjAQr/ygr3h5GMBAmXHSE
hG59M0wTkl7942jncmvi1HomItuqI9RVf5tuTplZZ265B0llFo8NmIvKJKJly6tXUfyaUvFZT5DQ
4jihWeZZorly+DnLv/bjz6ct1PLXpbhHy2Bw/mii8N+tNJza/NyjfrLXN8xaTCa2wQqagIWiwbnB
NhFRCrl6NidOONvPk6tqpvLmHxxbAXs7qJsQeIdeHgf/F9ysbx54dC/lVTdSsYQdr7mSwuYiPByW
sYTQCinNv6liLqKo4Ul/weD2xzZvqptIZ66gFq6V3Vhkzvi8elgwxJFH9G1LlToed1+HinG9GPXw
gQmGFzY/C6UTFTN0Xg9vcViFXbxHoy0NYWG6AdpceBE4vYJyeu88Df4OAqgxiu8KL4zvumUZ62R4
2CxHqu2UxWsaY+tgfGKNKHdxcyAPSOPznJmMs4fDY1ra3D1gR6qUe+f+IifIGE7bd08z/wYMKSsY
2lqdop8zxxdC04Sjo42kS+G5DC4WWXHoCD/ig2rpNxXdJnlbLP8f0Orfrtz3nwH1v3K0jIdHI7Rw
Re8L00+UqwK8soOdsCqBrMo4tN17Btdb/OqZvQefLQMSRmhMuw6IwRPdNjFmIngwsjOXOWq2QDTp
PVeYLGyg1ea+veUd8fMfPzLoJegHbiJOTLKqJfyTG3BCUASwdbtwMDYNYpm14nRBF9Zi08z8x4QB
4IT6N2l14aCjvXB3yjRIMcmzMWHtSz94nBeeaGH2F2L+jkrV4fmVoSciuDcumrlc/yztY3EcgqkT
iX14o+hKHsuDr3gZzrss/5LYNBzVi3U1s61w4NDJZ1BtdCkHgOhBr9Wo1kn3xzOrnZCAEZu8mtXn
61AqqeVaXSMBauIN1Bn/tdKTMdJlYG3m+L8R9OlrCbEItcngIVws/ABWKPpcWqBPYfomb9LEr35m
4g/fOEUBC+T+Lf6SYPkP851zXZC3sy+zKrt5QK2Vhdz8marKArRT6zsnIPWc3adLWykPqsNRahhH
J1VT5i3CDy1mvf5wOvdomoVj5ytKXIXIefiGp5ekSSdA3AJ9L/4Jf8nxlzS49z4uRJicwlX7r71n
ad+K72zNdfT8AlVNdorEhG2wGdJpHvEUoSm03QddmEuwEAXbkc74nZwpPvCZAm9raxkLV7nd35Gp
13JxIgQF8pELUZUIFzxpMtRpSrq1/Wrebpmn+WKKcQu5pNNEHEXwS1BSXvwZxIOpEy0uaaSazShD
xS1Q11BNMfmMcENSdoS7W/Nji8i2jh1fwu6QiSHLR79X13AiD+1oZqnv0i9jGVY+fAKXP2L0C+ed
uLlFzhex/BKZK3Hr2yKCqPPyhWsxsXD/39L80MupMIVCkkXJUDRUVjd5jbg7MbPmdiQYxGaUduNy
V7buN+5761mHrCnY5N8uIxHBfkJL1exXZi57qy9q2re9cRfWkT3WoTZ8XgZDtBa5jBWp2ikG7cJ1
HMepEvIb/V0d/X2xRQmbn0/t/5GiNF1kEaRHpWsKjaoJ5aZN9wsZQF/m1sPk+ZEkWJpgWWbjRRPp
o2wl751CMcsnjBGkn/jRogwBGCoeFGxbOd24Zquzs7oBczlZ9lU5JPRXbQ2c0200pHTqklFnOOUs
QhtlHisiN67UFqChSpck59zo1GMOoaie9YBHMczw/jJexNp4JB6fr2I/1kQyMU+DES/tKDHoC8x6
LF6FkFh0cVc1p0xjpN6ErOrrx9z3EpA5epErvBKHceKvp2hmtAqZsqzN0BF+LCsWY+744/FmE7Cz
gr3M0XovhTbkFjmuPiBIkutYTtb+ZRj/SKo7Gr15NYkc597sG6IuMTKrWzfMqYnf2Vt4VoqogV6G
VLsGH1VZfJfK6OigQmFQCp2b/bRyt7515DnNN7Pfu6nKLacKjF5Wdl9VN8FV7aq+iO39PHB0rL6M
wfjvVNDl2iVMVXqPFXsRcAoQH6ca4lguPoREGHucKXBi43w9Orm+yZKWjvJjzJvOz6gfZrLKkSOa
ar1nK91+W2tmEGV5WmAx1YSeFbMxYYIIsJuPjpO4p9PloAsRYyCUNYTjxuqMHMSbLp9/ci/H7/DC
Lnn99FGRMZODT7TGIPvAy33AlDbn9egX/xz8FkrxfeoyRIn1EOcJImFW6PS5Xf6+koWgbYrPMZYP
YsKw2gWcyu2c4tvsUmkyhYrVRVU04qQTdjvEAnQZhPyPNhOi0bl5U3pD5gQ+54R8vkWbNarn0nSP
9AzXzE3SBNPsOGV3pxTm0OJrgRu3RrHZQyXvjzn93N722kAWIkdOAUoBEqccYW8TYKHi1hvRolH+
HQUuOtEuKwiVWep/jF+N64zB/F6yp9PtluIc9XEE1G2FzfoyBKCk0pW2a6uWT2udML+VOEmV2+Ek
e3e/oDEoq09SrI7vEGbsbWSN+ZwJVyIyIhalTyWd/jny/AiTmctLHbYJJUMpmBkKPBFfXiKCZfm0
5Z3d9Mvt83KwhMordz0xn1RIWMr9UwGIzlPyMNH5+Hp+PIMuU8XqdbErfwuEyFiytJPddWjtOBVp
/UWbLVNtpLMM7bphDQ7m8tDD9jxC6nViw84xnRkt990SvRwwHQ67Xv+q9LkCawq/tvtg4wt7pftZ
SxxLwJYlklHh2L6rX0oK9E1gRuMGugn4B2+ujtJYKR7eeHz6WdwgX4shfQ3V0f9at28UY+SeYRZW
PePQ72CHvsy8NAOts2qd6JaydLaO1AF9lVGhsfnKff3j95QBk4viSz3NsRrXA042mVaxnwI0tdUV
7hfn1hIhDznJpe+NExReuXIgzaD3+udXfnE1XcB6sidlS0W0x0dqVJpyMqs2714L+oSFvlmtKm0q
yDJygVsWX5HV3hRvrR1WtM1ifryeXyh5lwxo/US3LbRhsHQkbx+4Bul/xUM6BQsIs1I0Y2sZsI2Z
8uHcb5nwn/lKi6REX+c5u5mFsuOSZyQPbR6xzBHEQ+kPwmoPpRAq9ipBZRHhmiIOpxvf/ijCUyX6
jyX+NB141KGMkmjRIpjZLFBKQEu4Pv3NV0hTavCdNyBptHprh/IytvsNi14oK72zeLtSl1m8OAnG
iQq4BK/+uqvyGaszJM/q1ZjT1+BQGodzNDx//76i17e0msrAZwbmFjMTwxqIXUFD6RyTw6OINTTw
kS1TGTDQ07uNW55SeKMwGd7T0eVJm981ols/pOUkuVK9PVnxIOJAjk20WYjHwXfssXto9pfx0S1S
QTHVPw9OzQJBYagQ1ajIRZx1thT9d/KfqSgGbedYHyhZLvlOPGiu9ZhqRVSYv97/0UeOFlFF742M
kUq+P77VtRkwZ+kRWZSJKuQctLk6r3/7ao7ij1UPqfLlCYFJFGxjWKisoCl9j17PBSQ2ZtNp1D5k
IeZ1L8HOWcZs2ZVfwBlFf0ERqWHy4hW+RJX68tVFLszMPLlVRYGZqbLelEY/L1i0qoRb3ZR9bbrD
4MJEY9Wr/0Lysi+3DmFPDDxJeglbOC3KKY9wma++pHUOfs7v/0vHSiYm00wg3mrV/pb8eLfVvt3+
IekcnKOcmzHjpY/ExinakngKqX/ZhvyxkePQKVySLGNEQQpBKM8B+JDpL5qzCZnJgg7S6RtWnlA9
DXtMNvbZAHFPBVXOCdCjxY1Qaj7cPlbRu60eqTkRj6M6hxb64zdCZcQDUHvvF3EGvSU8D2vqGOlD
6/uEeEDh0C8JImsxmsuJX3zP0JEc8XG9cbEoWtER7GeyibAZXkjJvs+FvCyeBba/b6d8+9izlo0R
Hop6OOTXpQ3C6OSYHtWp96lphSnUW9NAQJHViQ9HYPtsgXjgx+ztG99CaQSNZveo8lkJQhchwSPM
z/5XPRyxkyoW8hbfgpylv6ZJPABlv2qAQfQVALm7QBPr+b1V08hsh3ssfjpZUmE5Qbdpa045VEwJ
zMFA/+oSltykp1JrBESs5WYPaW0uZzeHm4xIEDLJmEbmByZ+t1ncmd3dJUTcY5LVsAywTmlrJG6h
fgdmZRH+eo3kj/2Kg67huJyOlITxvgbjpC8tW20aa1SGAT1n8h0Coq8DI4EMtNit9eVmuK9baaIt
73nFHT3cNJTPVJotbpVlT9zZlZx9ARoMWlha1DX8rfJWbGqC7onCPdhANUCCET1wXaURwEmQpOG6
wxJv8EKKk7x1yv0yniT3FcSvDFXa5ADi6UcSfUj0x+JT/TWYcB8b1+mrfDW05sozl4Ca3wGDo8qj
uPx2qA0Cdux8VBHJYHtkwAM9CjvkHyuxA8VTurFMriIRf4iszCaDGdlW9uCFh1LGzC8uWmyWOIyr
oX7HPC9Sf4yBrUHaz1ydi9rP32Baf51uqavn4K6VQ/Qq5BRnsLQ9hFNY1aNE7IaxiwwENJSkN4xO
0A+B/lQmjajibiScmp/xxTyCZpSf72Qoc+LBliT+7yMjDLbP//P2dkTMS7TBOd3ZygE7g03XsZjE
ED9RyBNiQlrFezMkFmFVHZnn29/NXdLAZNFBUEzlmcgrVequCX9AFwOPhEg0omyDmp0HcAlZnJLx
OrCvd6Nr72f29RayhMFme9NadoVwTcQF9iLr8iFen5qryolSe08N+WL4u7Cwlt6q0AXLJDyHd0oB
z4ZMHsyYMgNuzeXmRP8aNIpOPhLBPmJy17dWwhn5Fc6MDxjT7KmW0uJ8qQoIb35j4qNMbdieOd3V
EGPZsV/TkY5eftxzsUUCM4lODXwhCL6wkCH6oFGv02uK1TJBV4s4kLE+GAr+J++JNO467GFEcb0e
73Nz1sg5hSXHEyO7hJ4nJD102E+Gro4qWMYILUJRbSxzb+b+OiMMFQx4dx/QKTCRQ6GtUmEtsqki
+1xmsKeTw3P5gVSdyX1evl2xv0ojoSp1IoWCTcP2xeXW+V+VZrw44kok137BzgvOOZMn0Jap8SvZ
updfD3Ji32uBqALXB+E6cpiDMBx0cDK/IL71Uvm2kJ0ffDZieNdLmlXuSbeKh1NTYVD9BktrGQCA
tU9Sk55pZIIFnBcpVnUbjvwFQOAeIp1tKAfDFyv+Cx5p32Cu0WISoliwh5gie78bLGw6cYwEby4k
G5YRZJfC1BXJQJEdVbbhUd7SwTDWM2G8dmn6P45g5xE3/3OUtGdbdFOopCdM3BTrcBggNJjgjP5e
zklqQ66/q/NyzgOtkw6gUlCOQBt6EB9RoyFDEk5Othtb+FaoJY/k6EF7tVUpBtILSq/r42qiEC4d
IYuKKGgcNrw6gLPyHRDr5Ty6FNDGrvGGbpTrJ214Mz00Os1E0d8ppthdbGQ0jJn8fs5GCH/PWOBV
Qj46SHvgxRH3/JiE4A7qIRe1tJAT8IAzBpZ2W63x6d+kCAIcqaL99OkAQI0oP0F76d8Bfp07DHvp
eKNLcsyriz1/uHv+S9PC0YvPK+JDak1BKUIyvkUvYaRo0Aj2jz2oEutBEs/Rc7d++zOq7q6VVIIN
ZdN2yizxQpt6CgSDtYWJJRyn7oeGPMgInzubc4JRW373teid86vZfxDM9PeW1B+1sPbEUEHZzn+H
5Spy+fJeO/QpprVMTXg3KBLMjLci6N1cvQeyEocI0zf4ZSs1H7uGz1ZXaaxQOaJcw/kXYUPsdH/y
bc7PF5p0XOZWRU7QHPHEeGHe/wI4XLs/SKTBxeUi6nNXK8LRhQR6aXPfW6Sxi9XQb9GXEggn09Vo
tGBknuZirr1+bKb7ycaxK7qrWal/0A8joETJKqtW7qLzVmDv7GeYEZZAdbtAd3Pp9aUjbIb+W5z9
s3MDrD9kKyoOQiE0ZXCZwjkr9IHS7o7PDVXB2OxmJkS8SQLSLOdCU38ihc30CX5U9CeTgR1zrzNg
Q+2WwSN3bRPBgV9BLUdaBDxWGcvlRD4UkAnZ26ZpNf+XBT8DHStaE87B8OPHuw1ukeCaA0QJpbcR
lVSs7fNcU9VKoFRDN5r+81n+7uzZWU83Os83tsTO8p2oetarU4+64Hh585vSJCpUnX+q+cPHK+ga
CUnTCFKCf5RoyoJ3M5AK+RLsglFdF26O4ErzNt0v4HZ5/QQrEnWiQk8Vbfn/685BwfNmTOn9C4LF
MUJfhFVFEGYldUT6dWTelDiMqpcHg76vlgG/8PQHWzAwbYb4v7niILNE75xCUD7X0NHrb1m3wlci
ohtwtPR6gLQtfl4B4LbXu3BSYrRHuBhsR6ZE+pqLbq2K2LyXN7JAcL6w+Ve8nxSaqX1nzE8z9zl8
c3TfB8W+EWDcoOMLHgqg1vQqYIGYrh9qIE6OkKEifV8FDfogl0DiUt+ky1TYynUK5nCjac/azzX5
ZYhCN8rvfjQv7zFJa1iNwKff/h3rHSH2cQQj9So6xbL4S4L4Qk/3e1K37YY0VRNRQY0MBO+h19Ib
yH96qgrB7Ibv4SyKYg+KSilxUZPbEfLZoZbjtHVfMHOv76GFMBS3f4fHhM29ssT+4k1TWxmp/sT9
MFttF1XT+N+uKgs4TdbF7Giw0MH1kU8PkMA3JzRXD0ycr9ikX3ueTqMaq7p5kJ9BfLCNJPXtV/zb
pbDMl0IsgfZ5K1hgeaES56os94MT0DFzYGWgZrcTyuOR79I6/z81UHzPZHtt0vODuHN+fNo4Frh/
Xz1krSV+VTECcuqwz1/Az7vtVSQiGvSaY9K5O3f66tlhVnzhpPRDlextTzxIiL/yYhp+sNyhyL58
8mtHXVX5ItGDSQqCbLb9iMWWTKvsqxfRQKBYN+8SyXMCtWKYngoyMZxDmw08nCBHFaiafDy3psDj
mtmC8ySolr0odn/q10lT57azE7XlHZm5pvNu/A03Qa0WeDpNDSG5mYC8XosyXZspPdvQ2bgzWCVL
hKTs+F7Hrg2Z2C+gM4fOqb8MrmdN0lfDKRqRA1yqHUPoj+6T4nQAiWpXg3jEoSwH2x12cNlB6XSn
11zMDmcQviQPcyy5P9nXJrTWhIrTjW/mfqshqs1shT/Q+qUFmUtcIxQBLK9livkbP1KdRCLo1g59
789DYr5mg+uYMTGah8DDxLz/sYi2NmhXTn0OKpd7JUvhkk0utPcf8bDwYmf6fy3sx1Q7UXh0kLkb
dE7c9JmdJHIlAOFeLjY84nLOWbp1SIvtUFKxZG5Z9NuuU32AjXGI9KlYbHDWNnaXOWbvFqzbOj7w
+KRDcCB/lIHRgJcon6doF63fgSjnMf0hEJsSygdHSfsFqMfOXkya6xGW5uEyl0tDXbyjAnXe9h3i
o9k8eLi7fGcolrPJGvqVjhXMs/A7DbNzOpCua6r0Etts2xt167elYZUoOxaazVZqLDgSZhVIFasx
KMae4wBc7R+6sAGT/yEwSTvFlBB5KoXyNjPLyAR8O7Qwv34g245iJcrRyXFyB/cSuGHOi3f72xUI
+h09rZXbyp0JCoKoT/GMavr0+Ho/JFR/I8ePpc024kIW+jBSpt5i+/1VPFcWVX3kjsYBtOlZ95uW
qLQ5R3clj1IW4aXVjXurUABzgbAmPzFbnvpMu94V7e77xI7XTZsof22ElRkVWVeWSMJhZlqjUtJ4
JhpTJpxc5SJfRzUdxdBtYPIR26yCPEEVCkIo9zaPVTDQqtxRJvaLufgseNFzGA6qyNmnk9rxYLKL
DwScbzzeJ5EnL345J4nQZsiOzLFnaEKZoemQSPSQRedEYRrsLUzYah6OHuAEJzELynDUpWykQgpt
520LOq8UrZklO4khnmBRRuLrjMd5UKHa+EAg+HQV0+ZgNzu0x9gh2lMyqgNqijF6T4wkfynKf8iW
wKCv3mejmZecwo1I4mJtQV7qGLnteKXAXssWKJpgwRnpQMCo1FElmV9+L0X2cFR7nx9FrzJ2tos0
+FUSRMP79x5RNS5/ixuYy0r0aEXtJV9Nl77kG4pjw6PdNjkEI5lDr4PvPOr08zDfqFkR2lkpA3o3
VKJfEZWeMmd/cjVv7VKoHjDm7P0AdbQO3x21v5ADCtqK8U5T3da/olXQbXN4XOtDyI3mNVcVcJCn
OIDNLl/DKWknEQiiNoIIRi+MmAWbuSZ7LUkF3lnDGe2IGWeb3lvEUSX6iuPnjNwqGi5+Cb7t4QxX
0KeIludUJON8h7envXD0FOzy+E5lnXhtd8ydH6TbwTXOH0YDJHPd4yRVHYMhwr/aVvgPqykn9P/F
WXMs3mmTFuI5a5lLfz8MP5eSYmWfGA/MMgphUxzT+mzgxv4IZIrSFdVBdy2wmEPMgDtRnnd7phWG
v6ZdibUKz6rQDSeVjXK6tjon0CjLY5ofdrGUINWJJfW9Pp+iDUm5kODyCwwxpWVZRES0YVb4X8uv
TI75FZoT6g+2cPYPeHNqTjYjhCpms9fCajOKvAs73Tuc0xu+A8VAURxx5KqWLEEWnbv4SEJAk7CR
vKd2F2PxbYwTNqSWeiethDS0GlvqJmNPjOns/VHNoVOKm6M8hqHhO4KVsr6Qp3+0MbZYNrqsnNbp
utR2+r8DdRzknAuNb4c9qUoqvn/I7IL+brfKwF/x6Cf53KuyZfmn5n59ewR3n3UN9WBuY0lOWRUX
1fFakqUYJ46CJ+ml+VBxMvUep/xoct5SUGuT5wgRf2shNnyGnoli/KgCJk2pnykjE9R9NIJm6qdG
TqJ2npOf9AACgjW7osXt/8129DwiYvqURxh+mlSkIsh5zUmvr2OgrKOwL7q6hjRmsVSDpi8OPI85
y3g7KmV6c31fK5T/T/HdJBIxUgL4PIo13xalvTjzE2rW/gne+9I8rOoSgWEPhb0PsIL+3eSuy/hS
YsxIHvMmOjGtvB1QK5RHabW2I106GbeshvenoVktFrFAlCRvC8Ikd3ykABbXhUX5Q5sQMHIsHq8v
VY9suNsp0yy8eAXsH+jCQHNAnwKnI7Ali6DIzAzXdiauBw7eVaEf6Glp3kw1vab/Apg97t1aPhY6
FiaEwyNlr4M+LrqT8vlmgO4Mp/DODGThZTlvQczDT2lZ/Hgw3xkAq6KJq49S6jt2BTNgdbPhx6eG
CM/9XjdLkbjaOYDZH0dzmpEz41ASr7HGZK417wvIBKwkI3KMEpHtFyyyYdjvziEvQCo3d1Yl/I0N
dwgoibN4123NxAabEiZZKg2bafCAroKgeR6xWHEz6Bn4VzcHg2Zsf7m8k0wYtCqjk8EQrJZExgD5
ceexc4TxkHItDnRjFm5myAEHNtdkJ9+KL22LQaf0G7Xxlz3SeSDim6KMI1txQHK+KLIfM7K00u2R
92m1TQbYMxV9JwwdbOmUrXlV63xH9UWgErGtgP1eZjZlzA4fDjlfaJlaFcOPUAHXyK7jVijWBpD2
VcvqWNWssWvrLc/fLOcocjdLIr1an403947xBmF6dxOkKco0W/MfaCWK0yIle+HxUaGluFcaVbNq
gqkeTJWxlNS2sNyIM7A/fPf3YLOmsHCCq4gtQ9D6ywuKuNBm4ed4gBjKFX+sJYpZVNRybeX8Gwbf
FuBXJfwDAN0nwyY6DVIZcLvN/+N8LKeXhvRf2XkWd1hkG8Rm1mEwil2CJP9X45cANeAUGvbC/SM+
ORVNvn6gFYvhYCUFxi+ro1H1Vs74P3AAoLMpGADXjWh1txA8sk0kjzyLgnISxm4xPp0BknjVegwH
4teUR6f7hPl2hcgZo+8BpCkOgYbUR8VqqrIirhJb5boojTir9kIggngI3v2bW+dghcjQRdX7vlHy
twF3zEMFajLIV3WvuXmmNQcDcIIqC22TPcz4KIjChs+UxXYSzyPHb/XyMWH3Xy+PgXehUrh3kOIH
ibDzeEssT0P2yi/SRWHa7IIMlY6BQsJH69V14LPZ758+L5nFQGNlaQvZB5lQO0RL8kHekaFyYjII
6JP8MMJwLK8Nq0rLDJDbQE3jWT+tMZuZjElFZX2/u4Jd1F/Txhx0upGfaPLVM7aVCY6xbNW2cWos
zYBVP9MVygTzRo6mLRkS+JaGP/HIfy96LvUXLhKsER9KvwhhezGB1LZJwDoarMHaCZP65Q7I4aDy
YTLKWaurTFk5i6A4r30UcqcOoVecAZq8TNClYIoIQD7eIjxrfUxHQFafWwVlH+FLxyS/kEWtaWNc
kLOn+qerQxVHjyiapyfcFtB8f9UxLamrog/Q9tHrzEuiPtny8LvxZFyKLw5Sq+Z6l9KHwVhppq4z
K5he02NCSb0U361uf++ewjIKL7AcB4Igzv0LirkTDLBJwshNRIhZqVxZT0/L1seG77sRKQS80H8b
D5G6SZvrZFCD7TXfjAbzm3D57mWhFEAi2q5YnDQ2Efhq/U1mRFW7Z2DUSB/c2K+mlrKw7FpVbFxN
wvuPA3TJd0XndLYvQ33D/2EYJNEd6CSUjFUFRWDlfIo3PjWlrheKCW1+BTFBvZwEmY9x8Nybxb2B
rSusA3tlS9MJfBbu8R82hlW36lk2OCDgKL8VlEj6bn8O+bGOwV8Bi8Kt9UlezqD08JzqZpvwVkCw
y/B6KGuGYpp2A/yUSJa6Hm1UeSIYAF4BLTVUIDX/4qbu244qCNTiG3PS1UjzhWVxrglcdE/xpSwR
NsXRj2Bw8Lo69gyF0NSeOGhamxA0TYK5l2+WRub8+mZvym2/fDEnrDikzV4VLI0T1TEqpOaZAmLG
atB6gNi8jkquYa2vpcXg2w/lOrL9a4rReIpot8zZjICb+Xj+ZwE5afj1G3AFT9j0v1KPMkO+kOV1
M7AAkNHliSpVXqvEAF6UGc9WBU0hEcKvFr6nwsAmppi2Y2IEfg3nWRDoR7Q99Myplxnz0+h8b86J
hdchk3NmyBeWAdz+o+na0cMQohCntoE53HDoypzMEp4Si5reHmZP+Kg7sh+8CQVKa5ksgZSSSqHJ
5PlJ7LKpuf2FGoIQdN49X6WSn0zVr4lEbfswC3vNT7tdyANEK6f4uCVx+YNLSV6DrNVF/TvxljDh
9AI5/cwe7i8OxSTPbkxpnfUNXMh1UK+CIiFJum2KZJcqxqhpBroDv6zk24tjkuej23GVVkXwT9e1
/A90XMinxiWopmAWestPICp7Gj9cGiA5LKtjDjfIRWKwq3ufmLTSwmYLkuHvNqC4G8lgGD3Gwp4X
eHvOoxJaEOfLyDEF/M69Ev5Tk4ZsO+vEPmQtM/M+gFlkOHr16wIgiePE5QUWrOTcXoFRp3Dofe3C
ampQ9/3UuI/YQm7bHmWBF7893R7nPc11eMVkElmrbR9jx88xGJ5GazDTV8nFg6SvRWIjUsC5z1so
OZa3GDjAxkd7Saw+bcWRlvfATYoVRQuPRpohNtvXslhLCAOpqAC2nkQwpSRuX0HlqvTwAQ5ezCMA
sp65K7gdWn+HDGv4uK+Fs4mHFBgh8lOzAP90y4jNf0/fAsVcBruSFHyeAW+C8g2NxwufK1TpPX7M
6VZDTKZWV7e1NvkCtFCaLSmCnjbd5kmTmmWPY8axmewewIMTaozchndCGUrtPQNNcAnkAlyIRJ8f
iAX29aFdAEpJpMHLA4l0QqvJboU+Ognr01uSIZsboiQKsY2om1siR5GaWR1r2yxbFC+PyIsTsIGa
HylPofV2rQcRBaizxSwTyW8LS72wU3iUfbkoTEbKXwaMODxsu1yQ98/QByPU0yIbGgfJ4L+sS5QR
c3yDNE6dU5sO3p3b4+Qyct4FTfHIcKqvPHh0fBhC5SR3Bw1jPxYU3Igl4Udg7biil3Gyp8lb+iEs
Jtc2EEvoYTPU4m9i/NXlU4fU+PAjiCv7BiHKBdHP0KIBJx2Yqv/dxtG0f5XZQFDVX2INbF2EEEzp
Qr+aqHDAPw9TYFa2yTUjFeQih8gVMhYEDEggRYtpF2zcuU9Ibgn2qOhryxRiCOrkVpiLnQkbnzlV
G4nM5/+aJHcRF2X4qYFMzj85meac1N+PgAWH5sHR3VEUSqdCwQ+GdvZAiIBeCZyvVNmzisrRi7Yu
oSPdCFB30jCXcOh/0JARGZibnifm6qFmRB0m+J8/E0292yvRZJHzImqAOl5JWXVPvLDk2k5ijEcB
j1cacU0UktvK9E4MKFAj49ZXUOa5dz1dacXAJP/wcA8Y/rxmULYCeXuSGdgZS2rcRGY7BwoQ2EqN
MXYP48oPgL+VjHddqaHq7kIcVPi1Tsy4WOy/LL1viYxMEUH5uqE9Q5wxdMk15u93vFMtlZ8C44/x
u6+X1kc3m/PQPsANL/+wBtTOnVfC8OOPMIBJcSAqYZp1KsZulOLZtA8JQUk9Uuf4goYxQ7iVfncx
7sW99xJ4iatsY5P+nCWuqJ3LLbON+bI2oVj1GI1Cp1JwkDaFIz8sPJ7DfRH9qrf+8EcV9y+sS3Nl
MtjSBYnaO9j51xt3Nd7DxLmLPzkSFCnShAZufXIxuM3hxozFPzQNhIuEuYMYAHFO8+tYQjGBZIwD
+gBWQFlIbas0GtiyDT8MbcU4sRvjZTYdeXzTgAe9iS4ebHNoA96yWW3ZfftNOhjoWicmxvNi6o8B
+uX+xcAT4fdrotRfQs0B1Kgq2qenn7rlTbQ36bIryfQxPd9xmyEJDYx+xd9JiBtMSSdtAHOGAroF
HcZstwM0UfHbFDCxGIDg6SRXKwBTML9fYzgkaG6oY7DWUuI32H3COhSZ2uDftSF8GsILGAgxM0sP
7oeYB+ra940xoKhDE2BCn9Bnf4wWkyLsoHmDprkr+mCRvfpGsE3S5fKJHwA9Btfc0df2oGYPBzga
eBuuAPvEcEU1Ev+YeloP6DgCFOtYk5j8M4IOiGqI91vCqJ/1gSuLyZS+hum18jiwsLMaMBQEjRvG
r5+uOiaopxZCaLH90lh0AnLoNtYZl8runXStt5O/QRZsrPRTx6lE+HNYSykcEujuJo76lNJALgso
OeD7b1+2SEeYZJ0KuR7cw6xPRy0gyVgjrFwS6sohflo/+8cI1CB87JstEEAXq0ZFfmSQzm1qQl8c
7kEJlbhGYZg+rt0pK5j7df4vA2QaHeKqO8s/h6IxoV+66AMQ01iA1za4IHkqiL0lofNRNAH/8iAM
x52BY7+NOGVMwg4i3Q9MFyRx0lfrGwaBnvrtCr5F5ycxvUDkQ0/X55dXXjml2zpJea3u1mnqJoeA
6pVD98f2alTrjLXCmHlR8QX+wvBZWsxaw4mcSXqUNsenCsJ21+bFkw+gyB3Vv8iLk/weweU1Oqo3
MKsrWj4/9XJGvdAjRqtU7pYS+j+Jm/Y/5hMpvnhgw2lXNvvjZwG35Y6aMK7KCkZcqPAeKwkZBpMH
EE2x7UeSmPwkYP+XAX5VYQgnDjeyQnZGlIyFtIgLdZ54RV7rTA6MPQO9VD3nUW1yYW7XaE+qQH6Q
LelceWMyiuM3KukDHLwxpkuBdum2ooKLzWbyvE63ADthuaAPWcBpFvF+rsQDknPVDJ/a9su/b3ak
BqNGka0gM+EGBR+MP9wZUEbeggWZ08d9aZwqiCdCveJaIa6ODCbdfTJZCrKXolXHswHvgfgmt/L3
J9gjAIr1T5OOXkqJkeyobqsEYgclxLFpm6DUySwADJO19xWWbuq/YltBCcyIKDw47n0Z8pnPMlfM
A2ewHNf5yua4/S9hm5bsbZEe1j3qlixVJqXdacX6OiCllkxf/jDl+nF/+5jq89SkLamAuCnZkMXm
NnxXBPP1OiA5pKYb7+G6y+9eTq2l5uVacazcF6hme0YaIkVUdDoIIW84M7NWLmu9/cs7OmoweRE2
nv8DZFPNON7sUbKN52D8t+t3qTSOXjaMFtjZgF+AgnWAIJ59g1fVnZZI5Dk46CdRwqT5vmJ/SeuL
7SOEoJEK04PSAopF0Ao74SniOPrs8lwH0UUC/nycCiMCHn6T3oII1p2hqX/ei0yTUeLIwvOlPOCU
A44XIcYqBhc/EQyGX27HOKH367pD0mxUCqmqINxtVZ4suFV3WeuAlM2a6Et2ikpnO/xILDlp8yMj
440D4XqezaNuC9XUFyxwfaIm+bv8csw/auk4EFS6EyenOq+qbpFvymR1AlfwV32R6jeqqc4VjfJ2
UrsVri5cSnv8NsgrSh2RMQIxw5qsr/Uq83KVqWo/5ZHhInDBatoDTyurBYYZJvqViXlUQORXK1CI
yfQEh9LWZ/8AaBy7a4SIxThL2Ji0vqA1IP52FSMhSvzobUBAQngvf9JWuBMNOn4F1x1Rb1lPChdT
XhY8VVmnTJZYoGQXFYobJqdjq0MUszKktkJeXJNrcgQ8nkrqXNXZNBlTxeOf8Elrbj2o0C4eXKEm
OWDKYkLx/lwb77V1Egtoa+/RmDXvvgILSxYgKMv7USbu79rZrj/La2Ous+AYAebu2VV3xMnUFSqr
BeSzjgDLAETZ7rB2UN5PphTo09uzaXS4XWPOBefkvbJAV4Ox8Am9Ntpt4tkLVUSLcvxfSTwDjazY
0opp2F41HF0AUDsXqW0SaRB+MNLxI40vGUOuJgCUf9qOV+6nMRoSZPD4PokqjCJtYaj74wiEyl2r
bfo9d0BhK/eshkGlBDFAmzj7tiJOn3PGUFutMN9YeOjftMl5PrZqTjoOId8XA/FS2Rs+f8D+sor9
qzWg/kzlB8j6o4BP14ZUGqRIcSqNU8rgT5ntldqwsU/b+CtWRY2whzZ3PA6c3yRcQLfYTFdp5gdk
eEwM6ilZ8pa6F0IJ3w6fkbhRymmZu4wTY8LW4Jl4994zwKh5MRBlrXx0awTk7eXHySyoUEODq5z5
FbYXxgIDa5eIXSP1V4X8LAhmK7IurKsj9pYn3Gw96rc7orpLeGXRsnTGrLqmioLuIe7a376n2Ajm
oKR+jYhlopYvfD1TmtPZsjVWmFoMnGjA0m7zfhFRPyRNTigWvpjw86aaCyCJxDaZcjLgnq7RqujZ
KwmCEhiDZ4gu36wbofCiodwVGuQRxCxAErotLS9CU+ueP9U7MiXEfvKKgS3c1PGELPkb9do4QWnp
y/okid4bhnOPdIJiebd79B/A/UGJMvCjNiKsRrHppj43oxD7y1vaSvCywSaDoxcSOM0J+WWhTkgo
Ib9hukZIjADlPaWEzBOQI5yaAbQuLle1zxvv5abqugGuvbkTv1f/bbbNImlPTANwQHkzY8LOgy6P
k288tLUgjWJKIqjYKhAPDDGmYA4EnQtTm1VRnWJbvBqz46qypYbUNKOpjldNpqjjSZ3Hvow0OpWK
/kwJmw5TfvLGuOpx4R853MBYwF8cg8VIwjJ11OzNUNmRRTLqa1NraCFrLz/cIdGmF0F7LBWyy20R
IXtlJemYyc+NlVBOCM5PaTveM4OefstEN3ZGas6BbQcbFyGfbltD0UmRCmEV2d1QlsMuvY0J1R7R
4k5ixPdMaJuRnm0ooA9GfXXS8Ukf3gtyFPbSs1TCVrRIZ+Sq/KtG5LK/nJrlMKk9wJZil38kSgBM
mPdIYc+riicssy99xk/NXybZIU1KO9AWIvFhx/h0z0RURkD3pSmewWOQlEi7WMpNKBM2c1VvozDc
bZUZjFFkIKPK5mkw6CBi7ZFly3rjE1gBrR57SfulNfNhzjtkLmLYRVQmrUQ13iPYpOT5ERo0atFq
QruRrFgXL4BqiE55gBo739be/orap731VCS7fISHZLT9RdXWPVSX9SLPZkmIyBNIsbZYanXsvWhq
mmVwHJpGspjEaomUGwCfMIQ6p6D3Bz/DmhoSit0Rum/cFBhkwOMDr8Ww5udzSt4h0B4uEc51RE70
CmiqpCQblocfipELjLGDyhiZb0Af+OoTFX84/stXdm/54WZXBivjWwBZYPFaQgsVIHCirnrQrv2L
2W8ZLglKUwx8nwuk+X+39WTNbNcv68XpTsyYiDB3k+S0pdNRYHBkgYCaZP24Nb56NETTTNuQJtKL
HHYQzRGZEwFuW5v82+Y3W5MCnnYPvqEMBkHNRpU0MAeXetSszpgWWn8OBVaD1xIXSDspkQ44LrT0
cEYBld2VHLrwwsberi7d2T4Fg1xeuj5RV7n7OTBsXZtJg8y6ULXpuNBUKYrfB0SIP5HJSDWa/jU1
5kVU6dDj1fca7C9+pKv2ejDvmQG9ZbOSzl15/A8aLssCmzyhG4c8szW5R5OmjKV5NxFrtdJyCugs
DwiLZwJb9hC8LnTMkLI/zyQLObgBkt4A4OfhbV3Nr3pA4Ivi5eHivVV6g+Lr1/qFZ8nQLpUJ92Vk
uk46WqonR1ic9d3eSo7OdbStYV9bAKfyUWOtLpi1XHp9ISYv6YbVXPe3wQaugB/EexcGmQh9CHQ5
xa3Fo8e8cv4zhtxbQNdOp4Z5o+uHTXiU3Vx1XZYX5uz8TMq1Lc5dgPBz8VMfir+/nyBE6JJf2fHx
XSeqoUNzjdAdbvMa5/jnQRF9mB0s5TaNMkwVzNU46ybFvCqDodAgoxrj3mC9kFIaDOCX412kr1SH
XzPaf4YeAGmOatnlQI6mF3WRb97yJbfsQTizuybHUcrj6PbO33sNbw6NHm0bk+WLS+XN3+HWjhs+
kcRKk5csrjs5hT9CT+HKSKgRkKwp0MgbtEByEUk2emLO7A4LWmJDokAjVT3p7XdDYHS2iIbL3exv
C770n2p5oWZ8SuBxJWVuFMRTAFmUcdgl5Lj20slHKvwvQ5tfKjzhAxf78n3obhj36yCx+l0ruBbb
Eqd1HbMqQV7+t0LwePEpg3UoFSeWZ9CZ2GDTLJNIBB+A8Hhfc9/9FBIfKTWVNqaneppjUbXcy0AV
+MBvRTaqTVeqn7zETR35fHTNY+9L3aLCVsNqr7mjaa89LOu3eoKu4jT/JHT6xKvLIQPymKTf2WrX
qBge0TznDaPDRg4awAme8f5LAIuO5d6oUSykNOsmlPUwgszjOIus1ElQQV43NWPaDsz8UB3XzymK
CSUcjMB9oCJqFQq5ZdW2f22KAVlNpgJi1p64Gho+kQSMdrXU0Ds8J27IZrsFKLBQ8+8li9qCKZzh
+/RYnlEUnJ++i+PwOgSC+cPhD2neD0td0rWPvk4TdZuoutlfRCoVqc+mdB+UmNYYy8XBnU6TgEIm
FTNgRNDWtL2hsSuPMPFnhUTWUFV//tSfcfvuRp41FgXNID+48BbkbVyHaWfrNicP03iF4AviNLSJ
Sll294pt7ZH+p2vdGPJ/oB4f/9yl4U0ijd9jfU3BbJHySTNcF92XdxhHpR4poZEtfuHWoG9f+7Ko
VUWo25znZHCs/SHyjuk8nd3lgtHuNtzhysvgzFOggE0L/soMdzRDfNBkZS1TOUhD51U3m15/+fij
YL8zIXBsvpGjyN/oZp418Lz1lcAynm2lpXlyKSyJ3OPMfA3L2Zi3lRTfw2cbKBZhlVzlKj9FkACq
dtW5BBbVUDtvWtyeLhwxfgIOjFCkH6DVLjQrueEmiHUVGhYnWZZb8egcU6ypQ/0/2O/WnAao4Ceh
b/U+VhYM8orHPzJ1MhGh/zk8ml9T3pfhFKgegkXLSI6n5UWRkMbNDjmDZmlG06ONrMsQJ5bsjGI2
JUZisWKwFS/n3OjBaGvH3oFXJDORx7aRqHV1/XfwV/JDXH9CmHzsZcKceSZyP0SlpQJ8h/MflCps
A9F/8eLE/uagI66Ayk111OTfR03Nezkru43h0PALK3Fp1/miO4GzZVWGKfs5SP2jVl60xnCWAEC6
h7ceviFJ2k8kJKgLEXEuJbFkopXJTG57CYPMa6iQWMEx5wG5K66Q64/Kh3eIVleC++wb1DowJGTn
Rc1/WQcS5UWGjE/BS6/6LiaJpkpudI1Bu5KY80i2TFbD28qQznRDWashjh1o3vu8X/74GVrMD5Z3
UlbJ/bJfPg/xOUK5HyCq4yl7mwbVWWBvHVAAOq9stoo7u8XWOyHJfZyq/58DE5LE7X5SNDMj1p30
GM1twh143DPmVuTC4y/UDJoSwXhP8mdC4ZVQFTIzScRBK/2LyJ0DxzzwQj2dy451JmckYwnUm8+L
/laezjnfnJz7beYglfGRAzRCUpIzU7B0QXG+/JPxUssjdoI5K1ggL0CEH80thL+dOExIWuLQJtX+
YL0e0oIvyg4XJe84ls+ZKzaDKAg79/AhIUrM7tIDEMlA7g88klreJM408okISwIb8a9LysExQ/Lr
My3gKGkTeWTktKetNXB0WJTpkgFdUVghWmGP3jSmfCDAwThkDgKyrMscxhC1pNIhEg8n71yYpsq7
hpJl7lAS11CqvoxwMrrWjY7nneWIKe6uQHWiYj67CDHrDPSJp/WgSUSMOfcz27NAmjlKvlrqMEOV
VytsCOJJB321F3WjfdcW0DCL3ipgIxorn4xrrdljgzoBJH7lXl+6jG5uExgHqxA24tZsWngbmncO
q0QYUfJ0rdxgesTbr5nKt6wYTrn9Q1BtdWnerw0mZvZ5F0Fw2rlsQCckYWC325GhdBUpefUPU/Tv
MFSEYpj7tM/mjfqLw6S5W6c3kJZXgyXjJgfPB1BI1J/jwf5DgxpRn9H/m+7574FPxjAo6jmvIjvD
4ZFiLWpc5mXdZ/uOjzegjWbASJRnNQyM0Wvrg/wldO1AmaYs7HcbCcLEpLLqLjqrudusOmua9TN8
ZMsXJQfmLGlYRXtP47WN2IhXAWkG2w+ksoR/92s4Sll8RxGb/StqAI9AltxAtFf6Ct1KscFKB7Ww
shOSLUdSOSskvP9LQvVdyrjDsK8B08J8SKE1cVF6FVuDK5N6OtUeZ3bruvatyiuLfIYpwtoHgu1T
97SxA3Bu+q9wxg7S6kMgr9rGVwSoKQTxRh6lq6xxWUgbwkdr9GivKq+d0aI9YkPFMv4tcER+HWrJ
GQJeEvqL06o3Dw7LV6wJPv0BM3b7g6D64Jp+PdeCNLsU/gzvZhPkAGFdq5O3ZBE+uRtZBDpPw7Xz
KeUAkXMEg38CNVRIzSRCh3MrB1jZ+oOb9iscJeIVs8qW8VsvFlPvGU3zqHl+ozmFtCz7Pm5d/zEo
WIl6Dg+uhMMlyIikZrnkZYQOJ6kTHx4ZEOfaVuEq2bz1EUbUptKGSLBEjmRBN1JJA+tzEls6Lztz
cVnsYNQh46zWbNBwvZPZQIj6ZO+rR0ZO6kW1ewho5bCSxEdvWhFdKTnMW+veAf3bNQefIHKP8/n6
d52LvoBlJfv4sbGPWskanfI9I6F/B6iZGw4Ff9DUMzFWBH01YIVcsMkGMEHMWVOe6abzbn3bCviJ
qEK1gSuQKyXgFzD78TtYzrJofbs28fM9wTnnGq+0tMSny3WH69efuCSKfGK83j4Tm+5+fjsE4VRn
tvPZR1ySCQtFL4MePiyD+0O48nXxO6b9HhuscZlH+e/+E8SE1nUQ7kryGQz08gZB2DPGOvT16iGN
FzaZgxvVHiFM8B3lmZCTmv/7eE2/NIG3mt6wZbdIwkVRSI9W+kbRrqroLShV6505S3wzrQWq+B/0
+Gtttx/3WYQq6kQFqXFMCIubakylHdwsdOnS3AKC0ckkeSf9bhTIR2IevNEd3g4o0Zg0cEOLsOOO
zWMECqbO4hpyMv/JJc+UNalFiLj8Rltg1WTIYo3UF92iKZrxpqKQzpqPbpp2fs5ObbzKlaoM3aHs
GApXGD2XhFdsYEgxlKR3zhgqvscd8y7aB0UoAFJlzeI5pevurKcscd++Y+e4GU8+m/mRbiv3YND+
Nl/rmEtO8SLirQ/7W4igU+C8h8uJecPyf1isglx1m36o5zmutNVLXmeZMQDKe53Dtd2/4DTXaeWk
zXbiqrnIMTHRCguinuMrLFrOMdPlBvr7ecfTWoKI6nytbqVN8Ahk9AUXPPYj7aYxnVM7luCe2vAl
p0NnbQqOBztLn8E/J8JELZ/bxFmwr+h6XMQNCHAyLflzwJPyfhaPGbajEh9GyeMxo88ORs+m87SZ
STq68hBSAN8CBctOPaAG4LEQzdHWTJq48HeGhNt44E7WcTyTyMaT+JKeSAAxBUDvYVQhYuoKaPBP
wBe2QVmwD5UVxoaUKFWFaM4x9ygLncyZtgctm7uMhpwHC5UHTimuzPXNxAvKLqt8Iok+XP99iqZ5
gt+5qNqmlnsMOrmCTdTmR7pdiGpQCBzu17BwVPjvC5gFQX9P5ubihnkK4b9ILnBsoKQeHN4Ny+uH
dh9NGMQg+XecI3K7YP3NxNP4A5b1uTgxhdMAB2oz9Bgdt5/l0QdR/YWdJ++uJNrwlcb8cG/AZ/3U
gDXcr4pT2FiMNbTuxNp1D41avO7qECq/z2BlX9xyWzwpNH/2ybNd8o7sgdVToADNjoNd5LRuuvow
RjSrl1gjvVaqw/wnCfGFdUi870AytA8r+Zro+Wwo+xcK2yKpC33Dxm1XWi0Jftj3ye+Byeh1unHX
hP02TJOgT6YEW6zbLjyQj5v6fV/RkXEOqDFSJ2/Oosm4m2hfiKoFk5ZxhPulSb3C3klgo8xUrM0c
J/u5UDPzKfRcktoge7qY9WS8mDY5/fli1ZhUWtiJZws4TaQVSVqQDMMy0vgyGJFX7vSQYJpcTUB7
V1s11OXn/H2odqnoKesr8N/S48WLE6oCAMQ1JmDnDYyKeOgF6L8F1DR28m89yzJhQgroorHqLgSC
ZO5IVxYUhsIERbWv+Pdlum36A6fU14POGUKahuESyiJTb5WBIHQzu2kqeBTN7tFvJz/3S9R89hEy
h/vX6Kbs4sPvDCqSeS3FmDg0GZ/2i18PkNmKpUc5ghyU70UJVvZHA7g5bnO83cfLTVx327jcEyWf
D2OP5qR2lNoqJ37BQrhTAWY3vKIK5BqkYrbEkFQWx9nBk1PzFmx+5s5m6zATN9C/iGMcLz09gXRU
CtU8BshIaDJQBQvWKZ2BQih+Zu9Uwvt8zoKYpCMgiOsoczKnZcRVhDCb9/kDDdp5i+13Al5jEmKc
GkQ7qJTB89mYy1czjwC8k+UY+uO0wGLxm7hEghKOm/+TPig0pVpjYr60fbK3+ZDyfA8oJtQQWGrK
Uz0Lpe/KdAHZ26NOMXG5CZX1Y38Ql8T8z115YYN/dToTW+5u7tqEWMO2cHXtE+etaZ+lg03w/cMv
bMEeI4sDtX2ua9g6Ww8vIlcTBdlOGGWXssbtlz9eH6AiKBN+w9xyYbV3OqRK/G7EFkX3lMaHGqmT
9wHm4USpuFztwpGS5UZLLX7l8fLm7Zrhk5YSI4Z4lOYXcrFAqD76/LxAcQpYU8DYn285ropU/DvS
mjtB0ZFWUWJxCpja0OnwxDE0qOg3mhcN6thNkqk2tAYiofN7Uw+PdnWGK92leFfIcxL/VnACBDhX
KeFZ94BHwvnQXw/4za8rtO4aPRkJKLw2kGT5rPOA/8ETsYib6UwjU4BIx9qhBcYBXq+pL8arWe8N
uMV23L+kvZS9HUTT/iXUdvkTDUuNoj7aUXJW11FP8St/3awVjxhQR3Ud0iRTWsoiCAoiV3AqbWkh
uEPLBiDqZQgPxz3Z66Klk0IFf8RnL4IpWxsaOzzBFSGDiNcnE3BOuNiXTc7GDJ4vx5Z4zD0nIvb3
HSp2N38hzvJj3cz2OntWwU8aCXkIZ2pfl5t9XiVQJLfpetZudY1y+qHcCloXtcarHltFiwQ1eplc
RKG4kX//VwTrTih2HP6lT1KInsKYD91pNiUIJ2ZcEw16iPWQu0e4GRJxPq4LtPvN/HkEumZmC54F
k2XeAmablFnHKzMsN7161vsHp87LnIsiTGNYCclatYVBjlDqFEm5THlt6sD1x1EgThfObptfzIBx
wq8M29s9fDbRvSFj8oN7UR+pSAhu8vzAo/XnTq5+ziGAg+Fm1z3oiuoYvCMB9amf2zYqgNgInL6I
7+b5bP6NY4avAjn/ALIaDU//Y/4BeI7nHMrm7/LOpTFgskDWp1yL6aK77qyxDxCK96QPYdP+kfCN
zQVIMln2VyrSGMPv3Ot1FgEMIzk0cKi8lt6O6RM3Ui0Bj3aMRpbrQcuzp7qEkIc0ghkM95/KXC4I
fsRgRcjsiHBzvc9+d5DbdK44p7Ss4BO7CA40hAxtwqlK5oidSVUSbLwRwgmWCJlJwiPP7cVJ+Z+s
nTrQ6NB2abQiaxKbKpFSHCenzktSJiKttsadnfsK00BkxcGOKUL/pJIS+eyQwUzZfvOEer+QX++D
jfeWUMiwQJ4yDxkOKJGWWRAJj1BuJtYDLWyarZAhwLoXuLcKa7Z4LmMpTcKdM+A6ppMtQ+tJo60g
cPsIH9HYCgnr36lHMdrSukc1G563Us21TFmSmPULCbaf+u+H+xeI5eV70eAnvuv/gyW0GuupejsB
Q/tm8hw05L6I8Jk89LsRwPgo2a9i8P1uDUDXsvTHt3dBuMd9t+G6pVewRoXGR/Bk5vG7nOREKof9
GCczJzflH39TLREaLHapeZ9nbZyUk+C0dxzeQMvl/UOEVIfbLWzL3SX0kQhzDBdbf8RmSPczJ5Lv
DIN8m+kBlxqcMmAH5a9RbVR5zWMyBsiZP8tHpF+8AmZvWR7oudCIa84VG4Q/hJjzuxWyzOQuPhRL
GobLBiYVT3vaHmtRc+KDxKm8Ojbx2BgCHpiU3SaGjkPlnuYmApEoeh2Uv5Ek/gmG++Ci+1wqz8Cc
RzZFwBgenGv49m6ZCdfek/jkh2aineX3w9lHaAy79PXQR514iZYp56tS0P4Tu6p5wPKwLthOWw7h
lPOxc6mCozofXEEqITRXasqTEDqdCo32X42qdSNRLvYLAqLJh9irJZqj1N3MVfWyx+YRBW074tT/
Bbhz+R4xYxEO5alJ842tBexai3uAeQQ2akpblA8gkbaWm7kk4T50B4zRxZlFbfsEwWurOivBdfmk
xj3rGnGT7WN60QpnrFfJLPzjQUZgEkv7iX9rFWsuRZUyDHVA7auQc/qzV2q6ydvEoeKwlAyQZgAc
kR7dohA3gijyRXR9JSPUMTIrstfuJJqFCIl/4vPhknenD1k5o0a5a6kyzlVinKxas1zlecXtJiFw
oM1Eozeek9upXKnVOfp6ae9GTR4rXkfA0EOc5ZMuUNfmAEBHXxyuG+pY64uSS3n23wKLCWSoNYXR
UMr3cFLyog9LU8pocEcjibY6ImRN4LyEzfiTjreLE970GbQ6qhqJXv99cc8JG526zVFk4fyUwtDl
eo060TaqdC+2wcFn0QRX1CITUTF0IlDoPZxwpNZy1aJfOkuND+ENm0bDl3azup/8Nd052khgRyrH
wvZakuqHXKqMFnStSpZ1fZMujONpAKsD+pkON6Q8B/8i7r0/4MMCvw1Att3xHEH4kBKfETe1eVAq
BHtAmAVOonoTdG8Lwi6VoWZQXVoMIu5XkU/RB6VeZin8jtCVSjFAqdYPgrkCuhHLkizgcamG3LjM
85UAGFdoQQSnH0Udm5dQVjNebfJQovZZoNIOtI5mB/M/ywcqkw36+OIyNuxIFtik15aoSw47IL6F
IJHSYhYL+nRo4gVhgD/J0uc4nKEsq/c650rP5ZDvxi2EPeI1iP4PpcInHZNjCIfGorlAvwhKlxjI
NPw+kjZRhVLFrZPYybbs0/rSa5hjeU6IanIhT8UEnn5UbeEUSfMEh0PgtAlNy6ldtBkCv28qruH5
Mn3P09KpHdnm4B0Q5Rf65digDsx53mF0uA3dK0a2OvsNMql0TRLgujc+rsPtXu7HjrQtnwKbrwLJ
lYucGtZnDOEU0G396JfDMEKWXpoSbA82eoW9plWEogQdUlmDtdOueTMAElRRJV0NaL/Dns+/ur3p
jMSYLa4dA9+T8BoOWSyTfViRCaziF2TSCMrway1WIy6aHGCyjsp9QufFlZmuWg6ZHZJBIu6b2ePY
rFpclC1o7KOGN0mVMKIaKVZNKqjE79qiY946ejBDbfYendLQJBCaqVp5uv0gZwr2J3bnBal4WqUb
EBUAQsZhKYXwNoU+2q0s7ylQ9AmLOodeL9tYymxZYRpLLTWHjwHJXYpbNHhBvITd3v40m/kXAk82
wiDtV0UsIYKlZhtzO9oooIjTyxIJpXjaUIFKI7oXNKXx90auYurFxqHmegFTXbTLP40/nUTW2U4W
Yqp2qzZP+bV13BllBwJ8lSm3oquoLjCxir27c+/oDd+2ixXJVFlZbI9WKhHohx/3YwQGNr6aFQAa
Bue1uJ79G63TJbd4VIxKRYu6rJA9xbdQ+BQMCb3gVY+3uNJbm/HWuVxHIjSdC70TMt9w9TRQIJit
cbGRjrbDW7htTbTjNi0rgVUL4vDC7nKUhU63U1X5evNDafydjNEU/XguNhOO01hJsTgUvv9gN7tx
KQWqpxN8NswfUndK6bCHl3c0vQ2wEE70naaHhd+CtZ9rmk2N6p9w8nbqZeoGZ6RyMS2SqHU9v0Gp
qlIcyV4dFeIYq+mwERIEoPTivZY4oEVa1Q2d7Bcutx/KASSMb4lL6Hm60Y1rRbQpbTJwL8LOlnIV
04wmn3iK2nRwUkj9PiWy2Uol3blsXgNH8ZEAIHW0E40sDEdNYKRyPILT7kTXODUp2YZN8j4lzoiw
7qRCCMBNzLgPHT/zAkCT9pJU+87dd8ipcmw/pBfRJ9LWgXwNoYQdlcoNdl3M5+QX8ci/Nl0/x2kw
Ddzc2EeqdQl6mmJ7WKpi+5/iOb5TR2llFZcshdMjpUnai+HFw8NK0TTQZQJcGPyDe+G7hDIhE1OC
XKq2U0L5IgXBSGsFr9inl4uvs3EXMWvV9FqePmm2kVPVLEyQV+lsecbOOQbz2Ztndcy8/eZ5egqe
EP4aUEPgjuTrDNfCyFn4+Zn3lW8KtLAaBHudRhqyMAWDVhGNP9wYhqxBLYPVBv+pJLZAV6d8PBBj
ME+xqjXou0+A7jJY2KW4zb9k/Qjl/btwVJfQRRh2Qn47zDHGCHA2B3pRnqkepDtXTvMb/vhUwDjO
7lowMBiU/nos1a9c68FfbGqOHs+tDfnXSSw3D5+pIcOkHs3Tia3i4+Rj96CqI1pu2wDmBncNFmIK
cotN4BXme8X5//+RUgFxv1eYMVC5DCRqxjyLMnZneocSorM2IzIcEzQeARpIekjeCf9X1cBua8Y0
V7rrfZvqe/U7f4PUdADZOzDKs+q8XzYoiQZ357VkpH9/OKMunZK9uxxx6iGYJizZY+hDLJ5K48I8
wfLlnJ8SEmJ/iSHL+eTZgyrrliIu4mpdkg5ze/IZnD6Q30xKTSxdHpEyqEvSj4zDS02wHE5vvTJx
9qMQnKQYeDIlSzJUwMI9VemAa/SeeojXTyxZAJUsrgELoLKZ4zgq42bdPOsdjWhGB3JGeYSuOXNk
YX9rBPeCLUlhSSHL4OJn/ctfz3t9eLjIVo/OYLJ+1qwH4kxycUPPaQJ7CwjVQ/gAxF52VDtaKrEb
FQZ6qYbjoip0pgE+exqhBZrVU4hCCOSdYUb79LH3TfdHnfyelJDfrTa33B8XsHglc7CLVx1+hkkg
01AWrIUisZaAUyAUvJY0KHhyRTA7Htp9KEDDJtxKegHHVEuierkZBWi/ZVFGsbkEUyg/IVY0yfkm
kirQtXiR8FQdw9zj11zFsDTqP1NhqlhNEMKJABdwPFPJ7/9fV4l/Luw/pWRWVzQL0otOpVRM4tWJ
DICaTig7U/WaZHDqoG4U1XU0WOBcjDWoKQLLntPjeKrT1S1KCFLlimNtCzHrgzP+LdFXbIGiMJoq
KE94PmkX2OH0AALQt5t3ukDrntTHVPiuW1Gjra8paTyVORCCEiXcJ7YPUnXDjxma15hDbCPb5V0a
5ApG3NLL/0ArqeYc7I+rso50z7SQ3GJpRbOoLDboloHwK0aHI+7M2B7KoU/vr2klxQoNAeDV8upJ
SUH+mpPqdcUgDGpv3i8efQlq3U20aEE1RvPjljX68RZDtCKxFpSPkDBVUjW7Y66VilbT5/UKnSv1
vVqfeS5l7PcgitrxTTJ/lOEP9itJ9oddhqfNGvQwzxGg/0VqgIEEF20UIJG005UYkWtC+lom6zEv
d5+2LYm+gOsvdUH6ApiTA+j7L4e1DGtc8qi+9iQEJl1ZIpRe6oy0KpMVNTuRZ0qKtdEURmi+P8dr
agtNYjGxi6Q/E9ZyGUoLq2VW50deK51x57MN1HsaAjBufmD7aDMKbLZRQ1w7uXXePipvOKdaXZRy
DtrQc+w5ZbdBvGhYrh7dHvDfbEjnYwIDOCW9N6Zf0DVeRyh8fRMwFOs963ROIvgFrhuORo6pIfXp
8dBP5rQgurnqgh8DejvTmxYOcDfK3NbNVt+8rc+iapXdkb64OND53ktWHSpcVPP9N/6HJ3C7CgyK
pSYyC32XVj4b7/O0T312ZLLS+y6k9kAw0zk16kgKaTmA3uPhehE0/eLXiOfbMMpgHvi3BzdwF8vy
r1z6eQCI0Nnn7NcFfHy8k3w8Hi3WtS80V5Mh30zlruvrjJTx8xhFZI6MAkNdX036q9/udySwMio+
WzyKWfWd102sLF8NUWNZ3eKCzuxE6QEl9ivHhb7FMNjsI/RPt+Ux0kiRnCHJpGBDFRz6TG97bnny
6zRBS40EQYJK92Pc+ltfc7pxqHKQgJPSZkiRuEX/VIh2ClFduSmTEc0+b1zdSazRnhSWIq+9uOlF
GsRX1BpIdfnJlPZ5JoKZxVgvi5W7e/RMP5Jr1dhFFZJ7rOe/A1bqzeEYcIt4w2UfI2wx00iTCTeK
EvJvoLuyF9oHRRfx5pMUMG+62Pz25pFdMJZBNW/fm8JQudcvkPpSGsRZmPzIJYyLPzkDYooOKwNU
Ch0fv5NOpKS3YxIfy5fAJ7pMDzAeAFaJlqOakl0kY4U7s6iVDWE+lkgpW/q7tYlhUPBEBQCRXHd9
iDWcyeqycaxP7cosLNKSByAQtvQ62nd7qHy0Ia0UQBVgTfweAGS6EJE2qqViSyeTPFM7I0Gm+ViF
SCS6ZY/LYokuwzKX/LvPHLnvQAJHIgml2OJuDe1Nf26z3/hR5Yv21fqWUxcD8SgooKnKlERinR5Z
5X3SyhNImqC+JcCMqlKlR3gWYTcRKfz0Ul6aEUDTkwqXsxZy1M1I/N6Dsti1zTC+MOXgl9W3+E3g
qpEe2CZ078TzjVih/Nth9lZusQMmz4m2Ssj8FcrsiOd34pBTisywrkNbVW+FVth5/KX4qURe6Y2w
oce2cPFX9taB4bgF+mBn4uqczXWEG/gG8odQhD0xJK8wf4FTNMzZqC0yAq6WM6sGKXwpMWeKS95f
qHpDk3VPYt+Mdm4aJXraiXttnzJiCGg7+jnUcQ3/gZdd93JUCB6Ok+DlgFv8E4Nk/qfp4Xi2Esgf
LriMiXOkTE5DtF3TxVKgqg418xBUsXpnG3LYVc5z0FAsTAH8IVf0376rvoYd5S7ORVB/qw/omx8f
qs7Xis1FUdtyjN6QsFsPBYQSU0xgPD096+l+CpGV7Rcg34SyG26W7knSnVvMPvkrqJMhlPdIzBTH
ggnqn+9q9pm3S4GlPyBwtqG3mkVuqOknO8uOBksZxgQ+cPucsaWgKc0aiT7AgKCI00qm4Wu9V+BA
0Ibmz7YEWBae61v+ThePgv83kCnHXtY0eo0iihimf1UoTPd4pBZk62DbHC53AyvFPgUuta8iGiot
zLJ/NUDufbVkwcWI9Df09LJhnwx5ytOiCelDQ7+J+BO839fokR0f1M5aJy8xGp5kiJP/jHf35vU1
VObtDpIZrTxkmOUD8alQOlm93CNOa4HPpSSfbbItf5+C5h+GdtczYeRPXvw+OCkHrYMsu6eCPA7q
CcgNr01WWvBZ23kWI/Gb6sA5NcJnZnTQJgUlq6tDl050EjuOWbUGbUNAiSyppc9JSJEirvmvyj4n
amis4+qIMm+fRIvWQxg89TDGesT0Nzs0EcjuCGqt23crbpvvJjpe0MbJm/2tb0WIuNs/8uPkoVVD
uH/xwbzr90Idythj+cMtxKQpeBHWuzz+XS82W5qJ34gimJGbNj82YB2oOpEaobQAk/LhUXeqMPWg
IYjDU7pagHzcpk31ru+x05otOejYbA4BKbc6CCKo9lahwvcB+s6g+cUR+lwN2y2ns4PiyGAAmqQg
2WYjcTfOau6g6le5n4EBIcBoZ5j9aDg94+Ik0MvTHue33+a9dALVQe1BYs+PiPFLaRNgw4fmU1KC
+c1IjxaxE6mEkuckZHsLUM/e5+37RRtDI1w7HM316Qq1LuB5v5zwo/FNPcPIP6Ob+wKrzYUBCaZE
EShWop2ZDLsfZ5vjivP+Uce9l/2UXsTOJbh/forXOb1peVx5K05bhD1mxkCRyjngEa3gX2SDasY3
fjRXoUjia2HIvBuBK/ZhliwcDHPf8VztvA3BcBWCjqpDUq0NVvABddjrdFwekw83SlFLivLRRdrl
JGUSSRbMR7xXs1A+iZ3dFoNhNgLWsFFhijz6eZZDAPe6B+CO6KOZlmaHA7OdvKQwTZIo1J3StOIa
h1eevcxDIPbWNKtgTpMyE4ODZykX7Q1L6yo9o9FctaFWopgv1rvOeXl6HWxTcKiDKOMhSmiILH+v
Nlt+G2hd8VV70giwzLDcsP1K4QhGEhZO2uYGbHEAaHt+oVgaL+w1rT/WCYnaTdS5odSpCAOhyR2z
A96Pk0WLa/vY4MNIeotPCbzQvufjmLgcdjnQrfwgC/+tHQeGNszvcbznOyeD6WT52Vd0Lzd+3eEq
+tvBZIQLtSzWdl6EE4iZ2OqxFRE+4YSst8ZpjXDXAqkSoxqOhDUxyvpoM65K5LGqOUIep/K/ELfD
rbcJxOuCg4Cgz62G2N3iJTCJVsNMi6hHHiSeYpSafq1WMPyUvVZbs/uHLY5JMQJaveLdJl+T+Q2v
0i7zrHVevAghjxwddz1Pf9HHZ5Mkk08sxYCeRMn6bGXpQevQL5LSGRReJ/dfNXdX1zxYsL8f0inc
zEASEZJmt0ln+IcuyG/9YPLkUCXezBOmW5rtUyhh6kW0N4hO6zVpBHOLC2grNc68L+69Pgx648IT
SJQCGsTk1vrzLR2rnub9dW/E+NfLx85TE2IrWd6dYm+UbSBN2xFVg+Jupdft6qbxmPQjhI17z8y0
BQ+Ru9wtWUGFz5ZL77/JngpXH38kxTxv+I2lOHhJq4Y+AbOoRiLPymRi3P/WQhi6CdTabTTy9Tw8
tMNA5icepME+w4BtBJbeRgJXoy6FE+wFfV/r+73313oh8Oe2SSaid30N129S9bmanIezpXm8ZDrz
5jOD40lrAKJHycqrB0TSxs8bXMv5Fn9+m+6itIHuXhsAiI81W9la5TlBestEIuErj9npj0gZrPDl
gFAe4hSINrQ+NpRUdIayIlACqRhhZM8BsIXylhNeybzd20NdPF7IB6Q8xLltEk2OIOKMBRwc2A8q
RAZ6QL9TwR7vhqq8mHyw5T8rmoDlfNTLzZi89BBJ3lISDjybvHdClFKkJRfYL8fhKjFEYeVdyf52
zU2GTEj0n3EHoXw51/hTqOcyaHBy4qNNj2nQDUdR8T7E52IX6NnelqHI658ZXLt58klIG62khMk2
O0sTqR8WWEv/Wp/Xnp36TmiSv++nohhbfWE3OjPsbgXmW90a6FtF/23sXSdrwm8FR0/3u2qbpqCS
VPXD92hdpSMROWjQ+n9UyH6dxwGj2YmP4bmNmX+slYgVL+e5ZMJMq++Job2pJaowABjebJGHjCS3
owQLNiYxLKk0MvYActG15XqkVGI1Z0nMEsV+CzzlGJzBgGeyl+5ZM7a7UhscOakPJwomOhQiUVPA
mcNpz7Js2dxmEl45yQdHAfwvTts6gnfWcwWfnmz74/8213hxABYKQTBfVVLWOq9Z3WlZkRB9sY9M
W09pWhnEqHcjlC3fanx65/6U3Jd2jJgnHbf3ENXY/JykoKK2VRWPx0YlZgGErhrW3AMtshGM3aDx
MHLvoNv+Xksc1dDhQT3JVgIB+gvx5yNXWck2V5iyPf7rzLyc8v4fqD6JITm2y+kTO6pZCs01Qys0
xuBxmSyHz/pt0mYwNtqiCu2KtCGt0jZHKNkITTYZEfrdaatp6cnvy4iS+LfxfQZab9T4fodRmmTy
jARUy08jL5sOO1lw7TXcmhuYLgoYCHVIw1SBix55MvZnNf3n+edar47LfAzh3CzvwF3jy/vTohnk
wcibaac9mj++g4YbLBL/twtGsL33vOWT2zV5NwAmquHd5hkjLeCcvfU04YucWsKI6oWtP11faJ53
LSDU6hoWY0nZMo4hGG6YjHLj4ziietPOI+XBA1n5S95Ljk6Ti66h6akqTroobSmUxfVb2IqzzS4a
eH5Be0sARlxNXavPO7vMqEM/1RScrB5BRrJJ+xuQax4yBAnSONLyKNBsWyKmmIm+KkoI980uB06i
EpEBEePMHKJnqLHemIcN398cdhaXJGuF+judTFvkSOCdt6ZpNWJJXCaVX+JV9j+J1+PII7Ky3YAr
DVbpaUh08deLmaYtmwBoviP7WNXn+WY4TJzfnOZ5peZ9GxhkjizyEMwO2B7SWeT9bxiS6yVY4INo
0Q9vt7jynPo/FUdlA/ZpgKB80mZEg7KuYhHWtHbrgQH+rYkxM+ax6KTWOIfUtaGiTh3kIq4eo9g4
UKMcSsvZ2K5a+Ka1V2WozKjZolMH+KX2LIfuVSE9kVKGK7bm7q4zlupAcmBjflKbht9tfoBbWl9L
0sxythT8IRIEppcTYehojsWUZNDbia76qyqCNlbg4MdPZzV18VUJjTxXvDghf4g/e2vSAE03BPiP
OoCfoh82/SHUGjJD8TmqVWtowQ2OCBKklUb1lUvOwAsFDDSkospHkX+/INhMd5PMXjLqjl4NlOvU
v7nLnL3gPT7TXOVBnMlJOlJ9g1Qulf9D6iK6fRNANqX66eiJf2/C9pGRjIl2voMHac9BHNgn2aZ0
NOYkz9OVGQTl4Ul8EHt9nO6EP2Cz8eYSeNd+2RtpP0XbJg+xlZDCnKXAmY+R9aycIaZbUAtocf69
Ybpe1qYw9r69u5KP8hDpn2HG9+d6XpnZGiROCD62CEZUwiqs4E+SZZyiZbU1UUjnBFQUrxtacLSK
YtIv66NskB6cIO11FZlS9UdBZdJkTb5cf4r+bmC/8WKlZ6ENB+XU5HJi7gwiDX9NtN87sUS4XiwX
yA/RRP0TcdFqPxWO7GbvERFxy9YUUGvnHF6IdRQERjkLJdmxDzvXYxTOXliDFW7rMqL+QlDunNbj
7qnCjhczbM95yA/YvxQqAuCX8mOy76gBB5TMpaI6d/QtlJ6MNU8zcmA3mwU2+3HMh6gS8DP6pXiW
MT4P+2CrNLc/6uJqHCG9ic+B72y2oXNk51GrXmOnWdL2yjtzwJ5HoEgKRQUtHIFZfr2UBDM0KGcD
DvY0IaI3uPriYPx7Ho0QfxxB2iGDFYmQsWQWP8rRkAipcyjYq3UJDpqrcroerlhFXMGIWm/nIZAD
eIm4x+hAYv2fPKNSxl36DKEPTHtafPViayYfjGM3LB5eCD14g/4VOVtheRAlHmNce5wodXNzJWPH
nkXs+Z0gIpbNL6z9oDpcST/sghMjoz7x6gDSy0ChCibp2Yx8Im5OONkkmsCZ90zagskmDqu47LRR
7p099SZAH5Ef85xkayhlKBuCvJrFW/PAqy9FgEQx13AeC9jG76t4jO0bTXdlA6CC7SK5/9mT9eGH
uPqWVanu7vjF/l4rZJakRc0pPwkq4mPvVOpafuwCK1z+mBOz7Z69LW2g1oN178gDuTjXmFdRX+FH
tcogWVmnoxiAtAe8aHTtxgrIW4ddgWXrANjnKuLm+jk8RBwSalXSA5jMAwf0g3p36DunUSpIl7ZJ
zGKMvejsx7cnuSp7rb837Z+nbjB9e5Ojf6/UPDckFq+WCLlSoDSOyW1XXN5aw+mjDY1GfwVYyJFL
RD7LXnOyEu3GtVhopo0p6SqVC5YVpkQgUcx8PAwqKm3blNzgNpgcCdekp+5OjleqCyzFqHQVt4Ao
DgB7zdKDLk6hp73YpA4uj0/9zmcBDvbcWvMl8aq8IqHRFSjIeaMvvuS1H0txPpkXqN+/ZyV1d5l8
6QHwL0i0DpKu3rqeijAWHHkxwTZt5Lks2n87ShdTfzpgIwpeYhY3mfNL/h9elZn5fGUQq0ThDQpV
O4QJKrGtUAk/wgB8BwdJFN+OHe3U34rayt+izGPSxWrpKPmKBiilTnh/0CUM+4PzRkqQ5zxtdNMh
fJfgTq1cqfAs3qb76loQqPXdholyPQhx1GPSge1LInpUQ0RrKVrepUE1DrJYcONwDSQ5VHLrA9EE
fPwiXGSNpUrG3zdeVqenxbsLfryhmN4bwKn7GXxXpUtckBQz987GuIHxKztNRF3D7TAGJENi31o7
0Sl34iR3sehB/f8u2u1Z3ICPYvAVrJVh8pgwd2aQJTIKaSvsEjLMKPb6y+qhmCNtI/q1aFCLM79P
YfwH4ILLqERJoOncq7XpAPHroJNTldSQzAY/DABpqHZ0q8zrpf6JNAKTLtNuYhRaczM++5dqOIds
czNciJ7AVk+mphiltNCr0NmbTsI3mn7QZxsQhOMP9ITKR/NPmGGJokqUDxhqMkZW+todGKes8ToP
VJVSKzmF1hEbeKS2M0K5YBB9U84YtYdRXq/yupYcW6MFVPMKrkSU/bwPZSdrAFXVrdatskDHrNUR
XR0OcrHv6XEm2UxIgyWtNzrZAz44kKucCdg4QQrRtFPMQw==
`pragma protect end_protected

endmodule
