`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
FTsurPhIDeyqjiDAXCfUe2lEdosuDSUJMXNYHZUkZ6pw9NuRqQmnxOSGNmvVo7gtQZzwKM/67vwO
j2QIgkcY3BUTpOpvXdR5cf7Q2gzCHqWRvBbZS6BQa0YGD13KLJTE34PTP7uZusftFRdV4o8DgGrd
6zmYYhUhqVyIcneuoltJHl49ScStUC0EYFXhRlaFs4KGWWM3oYgs8CY9C2Bb5my88OEjJXEdjo8K
9L2ptKOyVMEqJ/e27XRCUMygle02mfaDBlLI3mLL25+y0L+pOHBJB5csH6JejDxFScbiYeHqXfMy
8NPBXOs2U/eDc4j6QithYT2foqKbcLuaWfSDmg==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
GCOjDgqgg23feHTe68z/YUiGfmso3DqWeWSjWQ375NeLXMz+eGXFPcTeQCMdT7oj8/CXeJey/00u
Oyao6WTRXY63cmAVBd3t/4yGyzOrFJ5fE0eIGQ5m1X08zsBfwsRXtgOTVa4aWHYyfDbuoxSmxfR2
tkO8/3pgEAwYDGKawEg=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
XWMDye5x3spUhgDuto034wp4xPfCX8aJ++KWviXb+tAnoM9ZmIK/uahPhtCq6diFmbPV0546MOnk
9uZxVTmSTFgt0ds62TxBUltA/2RtD3SnhDWCV+Br+CuQFJuW4OGszmBeBWIhnfsM/QEidEIrxTGD
HkCh1E9QCNly35NuZPE=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2624)
`pragma protect data_block
z/u0NfnUPZ7mL+DlIx2PTTMlRCfSgpgsj+41fJAPZ4FcDPmSE0EjE//dBaO8Dq/f5XzDrgUns23a
dDYJla4IafnSoop7dil/l4A84zAG1v9KkMdogEt8oKv2iugQTT+RZZn9EzYEAuAE1HRiEm072OTb
hTVxOxRYznXNoBoDkmIk4z6ucZopSt4DYF6PC5iX1yejK1nDMJ9wO6cUubyBujzy+cy4ynj7MV1n
jcmYWePagV31wsp6in2zkRsj/4m4CBCxc900MuDiMgyTysXfbhSHx2MwQxbVdJSq7rCmbdIfATGR
ZMAqa/7i7QVQLqfOIDqbxXs6iEO6TbbAit9QX1YdEh3/TKHcoF4XZMxw3FwxdXZPI+J4+7VH+wYa
otiSGyCnWcNqPxM4vdChg/FXbUlKt6DJnhJ7qEEvpaUALu+tsC+27xdnV4xTncW089q69YYgluYu
3b9zMxIN53YX87xEm27lid0NrXdfYNiB6+47TbuUemUsEsTm6yN2Es9b224YqOPM8utRpuCLs+wQ
3zfNan735HQMUF/Hlic6IW9h0OCPR4j/ADj7suYCRFLaBo+QXPB4upr6udjsP69Hpdr/BCRMwRkM
iieTqRE03jcJl0MA6Ll67wApp8bYH3mvIJCsuqVEC2YLYl8WzC/abqWPYKclRd/lcwhj8PSQm5Ru
TXS+1DZpGLqbL5fXCujrK4ucdhHSXYrp04TkVw0LXegdqR7ZmwZbstIZfewOnUS0iwWSYR0mRJaJ
8lm0zhsqUxyEgbw0+ytmqLDOm0X3+8fiEroH5SWOYUQtvbZmXaF+Zkv++k2fupta+jcaIkdVdIHR
pG/UyIeOCHMzs0dXU8V57azthsK6Xny0pOfD+4X5SwP252vRw4aQAmb/PPgejyLm9Q/MONG2xr8z
agsNJvHZmS2j8qbveDRLHu2zuoYSmRc/augZUp5bD3MNtI7oN9Tc8gkuhyw5PLSJQudbVPAk6ttK
mc+Vycx6MFuEtkB8Ty6SeW91nIc3N9q/t+afd2WZeTaiH4YQedvd3vbRVcoucjDonkytLt/dFeOM
4IGs3voD+K7Uba9HZAisYOyR/K0fYJYpXMb/Qt+Za6OvuuG/oLdTn25jSin3f9aWJ/2emP46WCC7
EfjoeiBR5szkThtGzAyClxCOKbajwUIh6VI5EHQOEcFnH2nWYun/rZlNzUSkkunu/i4BVOe4HOun
eNuszPUhVPbWP1UIIs+NS+CtEGn0HaFfPnK/1xc/q1TWKX/WbapwqK5Rr0T2B/6qX93j8s0yHVld
G0HDX7Swof0GnfSmxwwoH49g9QsqHqBMyjWdM03Z4dyoiivRW6oE4mRhrVBX77geSoBQVG2L5YwJ
ZIghedKaSiXrpaprdvgZZ5P5xEEOWihnBDAM3DYBMGGkCZBVS6mquwMPCjZqMfTcuc6LpXPasDzW
oxLM5UqJFW0lNlcd+ad0CGNUxLpZgL43yjJqkYr5RdIz7Dyj/Zk7DrHim0A+r+R0OMWjcSUiLG33
QXNSH+lOWMzkLop+V9aXyzdsu6+pZR3lia4vvXV9EuwY+cyPVTNQx5LT/xuT2w3RITb9gK5pMYDw
XZd2lUonc1FD3QpP8fQCxXJSkysVFYdxSoE4L5e4H4oEZPLq2B8AGZKelJs8gLWBgmeVXW4/VH2q
MXgdxLop3CR/EvtE9tzJl9SvtjZ8sYTXuuNgJGIFmiVjmmXnvrt+rR/8kqfF46li0tsLb+7SkNTg
OZafTsQCdhzDVBb0EYLsYLVBRYlVG4YSVZRJc8sgml6IndXSoOrX5G8AadQXkQ9cpyWANyzBhfm1
YvyZV+CXZmCkfdRG4j/MoQod9mOZvL5p1QqmtkJ87b9uqpoWNMiJwIII/0kB86IdOd/hOetTbL7u
7IRjdcjVMNcr9W40GaLerW4q1PksX91U51eM7bcfxPueeWAjeRNhJbJIjE7WS1xsFDXtfLqCLAEj
FFrk661oqqaJXFLFNl6TyOWXPW+OqJF3fy5Z+nr4HoL9x2ZJhc6N+6N2/B6zTSLue5SmzG47K7ya
zrLQJTXfexA1MgYAoTBAyI7GrwOS5VS/EwX70bwz4Ubl60MxlU6gQwCv34aeK3BjDuUeCveJ4GuP
BNkkE35zcnct2G7yfsRcUYsAbxdik+kFdWg4yHDm1q10VFwyx8ZtlqcIWN/GB15DdVPE6LGn27j6
sEXOkSUr+es8Fm5vh57wsvZsd1dyr2D1ivaZYS1vwGmzDD4rk3LbpsYGXt7X99+V8fVWffR83h3U
FxHyDRTcKpR+BaXHJChBf17EcUmRCW0UDWUMWq6MAF2V+HvPi4pH49HrWXf7Lq3T/5tomgpR9uAx
dIkgl3t/h9jM4B8HC2aatdDNh8DB5x/jm0I84C50WEzYSPXCkX4OlDJ8OMoysKRUyXB1tClCn0l5
OxG2cXT6T0BFYHEt6YYAUMdSFPLorSJ7V529YcEQkMquZP+p64czt7K2PtvckJyTWkrOFIZC5Ndz
TYlHZV7q0pBfESmYFlU5V5hpLJF+0fXanLISuei8APWae4vwuGSAZhm78t5uCeSlU9j7AWlwFplE
RFuVTHx9NrHXfbh04ILSYTWFtNMqZ29PkALVwWjsIdJ2NRZcnV3R8VW6gZPllDFuvyrvu3TuA8r8
xkP3ng0fsYQ/2KebEABDvJgevvBbJK5ot+Txdy7Nz/gAbPyC3hLIUn5SCwW7GeiUNUFdNapg41+r
E+XC+bN40ci27eNN9qIKTSRuK8d8DvQe/ec9dq6ZH+DRa2Rxe6RZwwHfB3rir5z0Kj/35Ts/En5Y
ijr3SZB06kOjI9j5lwClfXIeHQ0R5d92L9Qdm/zp4fMu9CuG+Og9j3EnHYYhtHX5p4mORZEJHLDI
jKTPma0aXDEfl3HsKc+LA22kT6MHyajwDieikH1dlHkqj9GaiH6gsmhCQEBkUQUaJUU/DnBlmVIh
Sz+pazKuNorSMNQsZ4AD7g8obvYbB+mnzpcRQAdOcnobAgM0u1FNneicCgXiGeSq7n91rTZbTEEf
0db6lECRwUeHlFAyIduDQnRhv4rVB2+Sio63KfvKOfAu8V9eT8g4dRbrteM/emjuZYeGUXujM7rO
6ZzL9CQXsjbkjhj2GMIp/UExUBX0d3yjjqx7Yix4zeIYhPd3ywocBASQXy4a5NxpiAaQApBpj+QP
xInqufXG+TvPqXiUidCAXjehR35mQdywlbeuI3UCoHD4qNoM0UXOjkg9w/Ivg/7H1YeTOUd/UosP
dzCQ6AKRC48SC2Xk+R/Qh6hKSmkPL0txcPr5aLtXsQrhyrquWMvU7HvUUublLWeIEH75kMMP1U1K
X8cm/KH9379O0XGn+WT1thR19X+VahuMINrcfqqOMoFo5Kf9c5RevmT60MKcPVeF8qQR1DzN+Xnf
r1nvriif1o12c63GjVlcLLHLlYC9390YuIrJ7NQg0aMokI4RrB5U25lPkWcJWKt6TJx9SXY8BkwH
RMY=
`pragma protect end_protected
