`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
WOJaFdseDCMpvxev8M2U9fxlaWiAYMebhg7z6DZhg1XPTsrHkj4zJVEvhi3LY/ASzmHCbkJncUyi
UxRVBi28u7NgWAL4aUvAfcW2wVNTWiq/NWJhDcKxdJX21eybD0Jmpe7f/ie5cqtH16rrXcXZJdEG
iBXH9kpfDXfyE6jKvpoiBnoVaiR2LaPMXcX/kgttzSMENhfVqIIeg0uJ7w8ot+e04DHQuSJ+jm/t
XAJSxGwRHI7tJYLNv6lElor4gukyaewvko0f4ia3SHq1Pr5AnCKAZkyV3WCzdfdemnB0NXEyMLor
4M0s06wW9mERQxHtJocXgWhw4bNKKn0pHupySA==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
1nJPDteDqvBR76PNkErQxs82K9T40mMO8jGSWY2CLUoBqiwzpcJLUX/9/yp7KUy4lsqUZ0j1iHHz
Fo5iPv751GE4qizHl0noaGdf89bHhcIs9KxnZKPgvxfSo2FpFXMvx1DsIQ3Ab0KIPxChSBcNKIFV
+6Fp2HtI7wXmuNbKriI=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
FdDxpEdUYKvQidgiOVrqQAf6qAYcvcjT8JoeXJNE5whKNbUOfI+xGNJYsZlvrcu/FZZukrd4q9Sl
Miln2zbWraf5lIskOm9ue3UmIkDY7vLmVqckWXfoEKiLHfnj+Wp7zUR2KkWGrNYCRdB1kHsZ8EkZ
YsdXyA5Amw2vTWrNC5w=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3920)
`pragma protect data_block
zPp3cmtETpeCGhGV34FWOv7EyN/Jjaz+Az4w+ZDOnflzq8Ma2Nad2paIPxf1rTNGn9RH6OEt9kQP
/UaLco6eoSZ1xxGDY6Ki/UVW2gRif3uN44DxtonNmhzWL2Iac7HnB9xAvbMkA5kct/1bPhxsX4x3
PwG4SV36xNfhpvP+63CLOmcXbxbshZgSMclVnfQ7H3HE/5V6Zf3s/QXtgj+/p9UBS2ChKpyoCTk/
7IhiKtLOt5tHD+lLt1/HoHfM6QPbcjxaduB3Y31y46Owj5siRtvtakJ+RR30FnfZl84yaHxOyXeZ
N9qin/tJ29WmSeXSCKurgVRuLSlaZv5HvO+55b1p35QJec4mKZEN/a+Qpzdi4EGQwpISi8bghjZe
jcDhBvT9FQZPQQCCOKn+bCZASpzdUm03c4GrBXz0853LwJ2h5UISI9gxXLosC56gHXq+h1Pw+y6S
pnlWCqIvDJoJ7u2lmtqdPveUfBrnsI7irCt/F+lkNSQSI8Bs1zWm5J8DNwN+diNfuS+MmMv1ENeZ
fS4GKiQjdQhcPISZE4WcHmk5JtIb6dBnK6oeMBsR/aYXJCZI+z+UqBfWS+u0BsVy5Gu5x/UEDCLl
E+wcVVHE7tDIHSmbOHnBNwQgntVCYMUqReT9aXx+iCbRkGq1gE3gLdkZwG2zim0lX3z+MkRaXEaj
PAeFj7hJX/sj/Zi+mWRH+Rj2bPcvpQ85GttNXsrAwWnN8f6GVZr0bHvGtH/pH1ICYgMv4TFmXel1
rtpFqqpViVC9/DitfZIlbfnLCFE7T1kybU8pbNFpKrWVvAGI7uArRlpbeh5GV0xWj+IqEd1GqSXa
WnTa8auMW/YXqGDCZJcASoBnpVehTzzn1jKCRJ5FDCL11rOSpIo/w9c3hagkqYq+pQH6pJePIb5V
tyxVru1vfVFqZziOBEsHTSlTq//useNy7Xr1DwF+k8e5KWHR53WS1J2zVvl0ZoKEcA6J5WHHwJuH
GFDTqaBpkuT1s0dm13HGx9zbFXchDFpiAuJbSh0wEa77xTyFH5fAchdGp9wHpbgAf1YPfuIKHUPj
vgBubs8GagNXOGvlWDTOWetmFcrB4TbHCnFT5jMunfQZSNwBoxAiCVSN6/7GImLVJwR1mw7HQnwT
nP5V55yL7OUTinTg/34gUM15kUm+HKCL4+IFLvNe5MdrMoI+RaNK4m9jwy1gdJ7iqBIJRP89NF5k
a62fpsW7VtkWgdLbpKURmKt7xl+/CFRlxCKpli6mlMO+u+M6YKO/Ue3u2WxrXlvqjXIdFzqw34+k
uPpObV4ZVJQJNCnSG1MXWDwNaO1F3miSwgNOJVyIfH/vgAGh84zRxqdnd4brLEMVI+aC54Nvx1hI
lpggmrslffP/SPNhtdoCCEVayH57KX1WFNHVxzr3PG+NbIa8csEAzSmSxCeI5s2VdoNnbg03OjXo
nON/ALtBjk7rcAgkQ9z48yGtREaijjqA7fJJ+W8lhdgmmWQSz8Ge7K1lwIabCCZkeMDFSxrR3La2
1b80no+ZNrwyU0ze5Omx+xDoWEhF2P88uzjcYpC1mX3t8ZSOHMu6/TdRzqpMAhq+VQRewS0+vcW8
4aFrG4cscBXmAXjZpP/tecboPEi9YrgD7BwtOKp1KzTtD5VJ5AmqiP+3u6SbUHNNkLW8j/z/lmtG
XlZCcRf2x4KHT/snlRIFIXIPcNRLAWFPDPHZFdYz2Ov2It4svWVSOlGnIZCQzp/qbvLdw8OSn+n8
UtcxiGgM11MDJbLytjMQ/CtaaTpCk2RiqMSGwaWAnA9WFEh8EVzs2mQB/mCES43Epy66FGb6RUhc
WMQSabLvAT0FelOTbqhpejs4DHbyDkj1HGxHpLuLobUF7D1PRvo+mQkWLRE5j7PPnszMT4UtiPvj
zLKM/mvgj7f5zWhY/ExAKPF/riWp7eO0Inm3EurJgqKXx7u/Cv4M4jxTFalHOcQwfO2hAPM3Uk0E
7blY2hwMdHeLOefJuREE+XTrbJGDHlre3PPfF7nMk7BAaOAlI0BrF9660pIgHSrlfzp8g3A3jA7b
fsOv3tMwNpr+ZWZktd59Kg1Si3n82xdphSvaZ1hGwsukKSyaif8LEOyXstTVmNnK9/a9iXCqPAi1
JL6uAMOU+5pJo3e64uPfnzURgq6qc6hYYX3IK/bKR0eBfDBZ4R+lhjyIx11oJgA3qHm4pZz+pQtV
T2GRdOwWvFmKqqAfqbay0XjMSdc8XTi3uvPty/p14v8OT2TLetPJHm5UPorArnFztsHWOr3DAeF8
QUO/sIA35GW/u6LCRoHEN2W+YB2CntPeGcqAuKVHxGarPjhdJyqxc3w6Fm4gZBCbOmAcLY1l0VcM
7N8ujsiiZYa2is+JQDG0J4GlcQZ6rpNhUou7iH/a7dj1Q23pPOBix5EstEnskfOtqH2UBhiqljM9
Fx/ISb5MG88qqeieg0FWGq9cEdRql0R4zyt5x55PQj1eftPyoEBhu2FI5PXCnCPGbvFg7pz32+lv
JzZWnLpT0xyGVx0D4d7hqlf7P2h5AB+JusgsdDniInH821+DWKu1L6IT4hfWquhSWVw9fIex7myo
Z0eK/zgMjSNHdhUEaw9sQGbJ0XsSgymvj5bix7UcyIr0MCRZ6cAwdBhPyyRpezKJ/Rpy1s6sZ3PN
aIGXdQuEARkNuciddgjgaVU3gV2bpLBU9S5KzYRVq2B7b3omcjXaeDA8cXORC19mXz8p3L8/eFGf
CwspgG7HV/dsp/Ds4Eu+sGgHA/R89VEmV/N0bTZKLzVVe5fVTsgXc6L/9vh7V9oWzQPBSiyFuLE2
Cee8mw+p1vyV1XaGeeTu77H6vsMzJneY1MFZoCW73e6fi8mjLSBiQ1xP5+Y5fpk9kWTNtbCxjpEs
YuqSB8ZAOmVNVFl3sgZVFwRjMKejkkqCLHmK++FNMTcUGmXOIaNYAfOrDtv9JYAB2xTLaA1IvwdV
aPIwLTRC6/PpKMb/3uFDgMfSV5VoO2lyvCgbf1ew6vWXKyYuUQHmMCrcJ5OD7204ttAcEs5NKVDe
QG9Y8pTqqDEU/zmA6xLW+Ksx8ubb4R/NjzfQFmCLLpkUeHw6u2yzIefpldIlCqU7UnZMOHBtEl3d
PnLeSsi3BxTeMo8sSh7QVZu2pNr6iIVHWx+J/o5NgDl8LNGZBt6tTuMcklhjxxvrq/GuU1mFVqpE
XZ439sJXMZSoXEgFoekCo9a/jpz42P1ItwX0ldyPEP1i67sZ1SnYoPmpKZbJZ2T54nVW0LkARE/+
iGwnAZZVsatyO3FiBDkHX3jW6oRFH8EW6gvYko+iVBUR2/mi290gmXumH5ZgptbPiRdJsR59lp53
ZgUMw7N5HCuhX+cVGPyQtTxPa4HwDrmtiMGlovnTvCJF2zZEGbIgU2jNQQq9ITYuyI7A1rwAwPdL
lre80lhNFT0SNcmXMttc3BhIb8Kz3tq8cn0A8f+z/fSXmtppZD3iSCImM7l8K/wfN6nkN0JHMX0N
qfNujBVDRfGGc7Z2ZRZ9xdTtPmkSKQmvRXXZ5Gz31joTi5WmNc3fOIbF4vhx8R5J/ZZvdsVW0NTV
2mX7XYUrFiMKYo/SBNm9K47f2JmgLItwkKvduRinsb44YqAyy9nDqwX2ZfdRbogcgOeAjlz1kbVC
xMk7p26Wb9f0HDHJw+9+MP9NUBKEYQrojZXc/6zchD9XbufEnoPyy2/yXlPJaCj/RA6N2jFFqxKh
U3i5p/TWbZFPxW8L0H1LSCsHYNIS+qjmVBwpb+9Z99H1QWWzZ8w1cyXpw1XGJYwSoWE6qOIN3c50
K41YpKEncHJ0EGbr7wRZTHmTt8M/tTIhx0X5JRsUgfI7NKtcVBmf3pSBLwT+2WEe3buQT7aT5JGm
pWBQ/4rMth3eKEvsptH6xHzggo+gkuxO8nOftxpxofieATdnZmXfOifmtsFhIK/e/EB9VicJKC96
Bh5Es3UjlJHfPtNaXKy8PjJQTFZ2feluX9PYZ5b13M26WxzTZ7jWfozT/+14VyzhEPtrGUH0gI1R
dBAKHdisk4C28NK6PhHzoUSZH2rq2wziWPHuZZ4XuS3Cn/tozn2MOXBs+/M29egcfLh7iiUujuPP
5oi0lq0jVbTSIuJobuaMyXHaoMD+/593OiDB9yUUvJGomsVrBwEDClCDwBEIGjVtWsMoWvY1PcRD
Cs8PCSWJY6ZPo2Rh2PdqPsc9wijqzSkXRcoN3RNvgMfkjA8KhXDcxHpsdxqhEMl9iR2amER/HXS4
DO1HyH0C5cbx3/wmJfj3+XKW2jtjw3i9B+nbveBWGIRyqA5UWXeyP3twDx2f3Jw8CPAghtEh9DQB
WLp6BWHn6ZchcuWZXgHGIzvl6/nLgxIHRxRTmJSDnmV3b1uxaQqofoReOLQSA845fMFDA4olyi0S
z4S/lYqunf5zfNvVyzx366vGMzlp26OfyyIWV72HNuV4nZ9T1QaDUnAdj43goh2c0EOesBFbwleZ
8+6x/wGVP7668wrnhflKj6eybn7SYrpHL3HtFv5tqJgxRPD3Z2oorthRTFXrRCiUDwly7/RNTx8u
Aq9XudhF6UjAFy3kxnI08U8kCZ+b7JNwttGeVtNyA9sAVw/NYF6kK2kv3UnHE8s21btExVf0p1sy
vHbJdQID88ASNi59ekY3cZ1Pqj8Dj/vbyZmHsCgQk44q2fXUBoMOstD1g/WiDfrjW6qTDCHe/gyj
gc18xGT7Xj4f7bSx9tPwEbSDi/Tk+fiz/gfJRl6GmgXELvxlH6n/brEnZHU4+kqpznWvUtMsot6S
HrpVOsQpHbET6OJqd+itIqJjnqUrMBu5H4Wjz+ZihQnMboUPYoCvug1HcSCbFuflIofc804bW6BW
rtCCrmk6+XPhC/XSNwyZfk6tOB2Pp4oDVGXHcnrEc2TgFLZD1V9+1tO4z60Us8/7+e6QQBEDbGpp
ohO1Tq9AFsgDeWGS/4whdkznY9IRZUvsYQXCf5Z36DTH03uSwMf3UyLc/cTvl0i2fpAF48NnyotH
u06QQzHpKILFI3wvevmAFTBi8fJ6FQ5depa9kBLjCDNeGqT0uTc1XCwbR5SzhuhnHrChlMMeXXDU
sa4ufLciTgAuRj7HxoBulCOmBIkDTT+O1VkJ4q0HbwUdJcYr2OQ867/75C7TR26ObddX2W8cFZvb
hD+aIh+MQMz760L+LwCIRYzcZMFIkDIcqEyKneXS0KlMczFC8nxYYGPBoS4=
`pragma protect end_protected
