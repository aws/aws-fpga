./../../../cl_dram_hbm_dma/verif/tests/test_dram_dma_align_addr_4k.sv