`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
L9fPX30k2WFmVT791Noz6VJUhd95FGmkibXVBYGjCxCgmc/fI7o2Ug87UXqjSizp4HyGMBN9JAL1
S8MWV8GrcBMBRPMT7HN8iekcvDv8ydVXA2Kw+aFfdXaseyOQh2VopOpip17913RGMNOD4CsKrpgU
2/CWN6RKUJV2XMWSi+tfDjtAd8/JmCrDAMGDeNA7HF6OqhnvfDRuuw3e5j5AqijkUYdANsrhNVvK
HipmJMMkoeNuk9MHIzew9X/45WS7eQCB5LUaCGsg1hkmDsY7xZuJD8LQQAmzzLVR4/UuCESRuxNC
mjNBH4ZkGXWFJfjjd0i6O9Zes3hnI+K25f5gsg==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
JNJjm8GhrmtoaJK6R6jFAdTtb87wGJyq8F6U4HiEbvvyGzMG4tTTurQa9XP3JeMvleIkiqIM31xK
aK8YcLHFq04BUCAmHn9RuG+otq1kDlvhHVdpx6oRJLNN6UiqX6hsRE1my/UinFoSGV8LLiWLRYc2
jq/bcLGaPyQMwupgA7w=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
LOISpfV5GG3Srr39aCEEJMeTgYrjXwfFLZLbfg+IJ5UKPkbUplMq25Xezz3B7HwsVY1B7zT0t+zU
19PLufhL8DwFtFFfetmW40i43WiqmY2yK1mEzOROj38svEUYk6EnJXPv93LB5VxJBUQVicgVZLMC
srn6htF4l5qlFdsimgo=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5760)
`pragma protect data_block
uWKtcnzpVv6f+bIk281T7X8yA4hGD0BRSIh5nwTwR3IAWepcaCbXenVNnamax/HEThwC/hkhPvDU
+Hzp8nev94RBGwhfApWrUprSvf1txsMZeE4OslmlZ+5RmGxYQ/fimGJ3wzvlZ8ewy5gLEpkTDc/B
ke1mrBynmyBaVgya6s7KXbeYn+4awsI4G3X8Gtfx+j6aOIH8K2c8U34/QaB4YcgmkvwZ/kMYTBSE
ykSLDOhRL7ofVOcglZCQTYR+pmFLbX3lJzV9CDpZAnRSxjhUlr9QAXqVVJubZqZkgLoSjX2eE9+2
92y96xypgqfqpbe9AFj8zv4pnNPOXGHbLt2le8BT2vOQmcd5zo8rVH6zOArgywFtgZGU8K9HCVuF
Evj3U32jgjlgyvOF7zxuzzpyTjtnoVBoe+oODvL49B7di3O0rO6xwAhBAaCDlOMrMl1Q97XYI+nM
cVWnMgosCwHAKu6Mo2RycINaaq7uorSnLiAW3Vn3IFQVY2hGX11Gnhc9FTi9BmRwpv4TlZqUXpHT
4NpYhuGpiWjRcSPq6p9meVjZOY5xPZsUfw1kdLR6aVjmlNIIv09rOzS+XAm7TIoiTTTTlOZICRqh
p4/eTqu/uIaMu8iaq4hn8kgLZUeum7mSO+u1NMpd62/BKWFPzGEVVv9N9sr/9bEZJVom+Qg7mMBr
ONkwlUNn/ZvQKGF1pkxPyPRgESBvoI3tHas3x4ryryK6jVZbStXtPQ9Qh2WvMUDDCfRSyUkxwb5/
3cxmSyPnNHMqOHYHgM+Wc8LIohJpkMx9CbqaQUoTyY3PeCqt54CqYl1rMFvzA1cophJ+vVXXHiMG
7fQv8Q9BXL894tGxRsJbBOqaKGO66t6qJotONM8zZl10v0Ob8zrUhSf4AH5oe52A318cdYuuuBfW
cib/7wwItmsPMFvIE8mL/moD1u2enn2vivrjeH2SqmmQdC7S+7lkwIo0LGhkFSoxQ6J8kYyXLVSL
WKfY/xjcaspA4EuAJINktz2CVfvLcfwWvqFTIyNR1Q4+OWeX3KZXv/ToznvBj+0/aWO6I4RNkf36
ILl+XdIZsPd4G6hfTi8xdvh1g426tbiPKVOZCzof5K2l1hxHPxEz9n0LcHm3fITSt9Zj77nLaacL
nVTXmP4WWSPcWAZe1rrjo0jsfiatG5BWwOTRV/fO9rfmued+2tEJ+SSTizcWawCtjPD8hXRjofvv
7xy9WE+BGr/1oFH2DGewvN72+d3sOxVrUvho9gMZjEcJ13hYdxy+a89lmot0qyN4Kw07L7fIwPme
i1JkhNrtOJIFoFMVZUsRG4UVJwhnkEpH7UVhQ8CWLYVSP09OfRSXWsQte8wZggh/xQMhF6DtFs6a
Dr/NZS3eYarzUoc+EHaANcnUFPsO+nm5rmGMm+vX9YnAprroOBJXj1IwrArAx08BlmpIQbYQwHTY
U7aY7VGcamCEb25R4FhqsrWgvZIz3k2Iq171hWag4A5B4o/rxxtSmzznFcFu4yKawSArTijgZ0PP
gNxq5vbPcgiHhKP6b3QfuH97OSU2EH1X+LwJUV7cHWcRQJH3msjHLgrM2/Mz/Y0XRTzIrvAQTPBZ
yRHBZzgxrfIFrSVbN1+NH5soQvavM2NjdGu4mv0jScVGTXn0UoohNPeL/8B/vJVp4uRUJcz+ZAxK
4XkSjQznEy2uz7NFMYw/PlKMmTa1o2NVsxk/3uPJcZ+yYFYEgR67kKyClo74i23lcXyve9W0QZHz
t2wxchDLtsheX8qHUnp5fkxrZmGDHtLl/uCT3UEP7XmJ+dyRBQ5/HFaVtQ23EpHPOPgOf/ghRKnH
pvVyWHl5XrjyrsTagxPKm314RuW9P660P8/FjMDU9LK1jm82xfVdAwmJs/E1qP6uuQzEBmAmETjy
mcVUOvUvhU4S9J5a5ykOgij3baRW0O/6cGL0i1sCKQ9OzR/QPItcUt92p56OEscz2A3kU0mAv0lC
Ksr9pn/97LnPwHnGeUE4vwrobBGMAQXaBcE39kpK2m+RtfX6cb+uo7gilM4n/WFF7v7sq1dy1VhO
CmuNV9zHthckqspgSeZl6NC4Jj4XZN2sS7ZHKsuahyWY2Gov9kUHCpS8nW7EtMJqt88Wph6ODn5i
sTig7JM/89Uxclgev2PbCWiuzAQegJ2+iNnenlTiSFkN7NLgGBUzII5lbM71FZ5aAUi8KgmP7EYr
D5PP5wu3VF1Xx/geYM5TiAuCYopeqKZk9BgpW//yE0Kjudt6GijAChdMYEolwCGkEDTbLQf9KJRf
R6X1LRMtLh7CJB59SujBpIrqIjP4mzdY5F8wFUDUswExf2E83EZWoK7dxWQ69NjJBx9RK5ZzehUT
kF8c28k+9/MngzDUeAOXnDgI3thsLp1RVVcqrRp9N2im6GjzQZe/6wQVlKPLAyDBlbxCvuyH53xc
Fq06pV/q2J80sFHDhJiCAlVSE+56b93hHgPv8zZ3Wq5BQlWkxief//M80RdOL4SCfqvraioMIv/l
e7PE8ZDQoVq895oqJBDPwEfkgM9olEJeG/MjN2siqyNKrEZceaQB1bB5TpjzpbbNXU348+pX9jM8
TYPMDbrQEIGQwPj2/5rJ61HePu8WMvFxYkNpa+FQtkH7BjQIcC38QwmfGqFjxVsH0PBSU6V+taK/
nw3WM9eBnylGF2c3bQI6CyXq2mTlP9WdfFgS26e7zf64fx5oa6co/XSrtucYh3FzrSNE8Fob7aeq
CVdAkI1JeIKy8gbzqnGPNKWsi49pdWWt0TJgNFgPx84/XYvMASS8q9yoN7RVe9hh/ZdWgS9D4gsV
htznbPfHLyZRj7ssGztP8Spte2YPtEtdSDW0GNpjcEo+uQCWh7gv999iadpc/E007EfR0H9iy9ci
NwHCju7SM+8zKKN0+yo1NLVXlnikohTPgu0+avm2uQsu7Od38SjgQJOBTFTskqdiy82JqbT2dieJ
U6qiVYjjd9HQDckk2aR+MuDbk/9ETCBPzOEmD+aqzgs8UvQjU9dT907S7XKcJAiNN1kfPsJ3Q7Xt
4Vifo+1HGOsvICmglrGZSx3SNdMU1sLH7GPSCmVhtkYrNxxHwkMOCKVpuGKqk9+K+Jk/z+iksOMl
hOpUwbzraOODTX0BDBuXNstkHxIl54CMCbUglGQ/ueWLYpTlV0kxjXfu2F71mWlnCKFgmkLIj7Sh
fXyelSL8YoJE5W1JxnoKmOlNtMiFIP983jBtdMcDbXvadwo45Z/TWEEuwxuaRkPWF7Vte72ZLJqY
NnDxB8pZmSlebd+8lNV1+gYNdUsjOSLAExlKLfWSQnans/0KzuM8xPo3PjYu9QK7dBCT+C87M/VY
IGbY1mT1lyjiWO9DPwtSs0l6G4cPZcVXrr3l2eII3xVQZ4I5OhabEfsoq21P+2siCPvoEUU5cdk3
mLiVTmtfqORkK5AXPb68nVqtNXY+2f8JmPtrd+8ksrWzzxNcQA/sfIq90xhIfCfGbACTD0f/Ztz2
ihOv+mVYhf8gqelhA53nJ4cAoWGBGgTxlTttvj6XpxyU8Vhpw5gD6OK9bTuX1mZYhVKutfMxQnf/
1BzSgdcB95GfdlJwSm9if9oeZRzsPa/RcZzE7NhpIODIg7HetOuCBRAHZ5H4itTy35jaKswhVQIT
zkyzEIZHoWexgj3ivt9vKPCGOHQJ3tYmA9MP/tV7EQAh+yEaSRWNl+NAQ1LuHlWTmHn4GQWM2OGs
gUPztDof9hNQN5hXR2uAf+cghAruUDO+R4DnS/64RvnYgU/T9AXbaYdNZvgUwgn3eRvSGZ+uFDbM
gG/Y7OgFY+Xm5HRBM4KlsNtWSscc6N+Y0DtIdYVBwHWPJVKNXrcKZsGbSqsiNBv/4tMmNmy48MiI
Raoy2i6CV8UE9k0B6WRmM0v95SyVjAolc7TjKYiZCBp30J/4g8v7jmdnV1Z3nYdHgMnjDIkENSOA
DoL86Lcsrlxqh0v47POKO816WV7WHMZWHEo2w9ogGJ0lG0h5Y1a5kD6SRBDr1ZLihQpD744PbmRA
JiI6ry/hqed8FflPDNb1T3YbOksKqLoc/Ct1Xx1Dg5ZsQlHB26vnOnnFsQCuYbPJVwoU4MSGxQ2q
Z31WDnQGrfHlXRwinnjhUsxuX0hvmAH+Kr18tZUowR2DsaZi8wIiuwfPFHi3+n123CJ4GvECFbJp
8BgzFkCJ2aPC9qey7guI1p4+V27M04qr6vlURW1X7ZrQAbwR5B4H7RqCQJ+Y2JI4Hr+6zsOsdouV
TYXg+mDhktW9UXPrQLBi/49P64K0wBbwmVoVP9Xqmn0FcX3RqWmrzL5iITXq05C2aLhZI9El6Be8
W89rZ6DA5Cw1LIBKWFEK+xolAKnBbriQhDpjzV8Rt9sZ7+pMaeK00rMB6j0RpJGR5ROzhhFsOK8l
dsMVK3X14n6Nw3wo2K6ejmCIj0kc65cS2S552DF8+M0NXLVPAoGpBRIS4MW9mLESCCrPoioE396V
ZtcDDwj4SQ3fpLc811fkfhUqTepkZsqe3JkTzgrKYAzvIjNZwbQ2TXLLD+pw/x1nrBjITXyIvI8a
YjCjTLwtAFlG/NQ+X3fdrcDFiudo9E1+uGeM3fB7M3fbf+JFcACmZYrdPE6mA2EBYf4DYN/CsaeA
lkfWEMXocsf8Wsg8edDhcqk8B8ff0m7ZRHglV6/oYc8xaWz7pmFFGofmXtFeglLSRZdLIxm5ZS37
89AeQpzkEsV0W8FT7MyxsFlpAQBc8ffUOsL662VToHnWcCU5ojPNBw13D1Qavlq/2QbjfJu5hFwm
bcq50VoJcstGytwx2zCIo4yjbknSVQGrz0TB+XXDG57dan8CJ0YH0+WURnGnFXIcd+WuIgfkGhGO
j9nR/Y6On8VRe9z1YllO1oOqPIjhwNSPKmeMsM7yslmebJ2FaSJKPmv2Iko2LJ2pGRTz6gSJatou
lNsTULZe1+30VoGU23ASPjt5hd4tHTZp05C24oEfdMik0UY0JhXctk9gNzesw2qRFzwxxYDOCTVI
n6iiLSIu5oAU8bsXm591Nsw04ffrJmaxG4Eldeb0c+SI1EG8P7JyB+OaUzQTpiHJYvwmM2oY8tzK
73Pp4Psh0HbXb/M+SFDZ4hND662iFmwDztE7nEYVSk1oO/kOyabVanJ738cLYBWX2a4yQGTXW2av
5fGaXDNPVcAnqRyRGTKzPFYlAiUp+HQVHi+fJUd3Uw3BV3nbBaHI0mBIA+pUWr2Uv9kQpZxHpeFp
x3frcWu9m1dwF6rSWRIO2D6PWpGQGa8y+sh4Hin0Ueu7bPuC1e/uyiaSaJhq4APIGFQ8hda8bmib
ZORxIYt4P59Qx8MkOFCCup/OpDuw8Io1C6SQO5YgVYrEirqUwMh0k9f1+Sz4H1BReHI9/xMGPgBq
bNHRiDCg7x9Z4l99WOKldsVjBZT+ejKFm8Eu8v5ziTGhm7I1HOXUfl4nL5Dq8P9sn2+n4EI8VIr6
jr5+z20Ly/EzxYERXiLpLBKMOXby3Y6u5HIuHlXhwu3OlutuoOkbYczZT6irXc/be2lWOGkDra7b
W0UU+eLUts8XVX5v0Dq4VpjVZyIW02ZF3Bl2obrnMCx1e+iD/rx9/kayePK749ADLrcRMWMTetWI
Vsu1WxvApziPEY1aIPAX0h3Ep2RHN8cH2HO84gqhrPPnrHBmEj1kLidk0Zq1XRfOdrYWlYc9sABs
fUYoT9YY5CSUnuT3bbzAzK5UYmU/6HPwyzNE5kH13ltjzb24OkVRIGsrBBmIGCbBfmoWxPBZPDCE
awLwobFDvvWocsb9sbN3NI2DmzzIl+1ZVrtlvZv2aTb/uvn3be0MPId/M9PKWBuJIZkk0wlk046m
wPSw4YCGW7Xg4gopS5cKIDHsGXwDx/496/nRC9fJLL6Detsuz0oW05JSvUppgQr9i4SaZ513vyKk
KKxO3+82kEkVNCIJ3Hncp9Q3oQlZG811bLeTOJ5WSgotEdA21Fb8Ts/Vw+r9+vfXe1cUxiRewE6D
QiBI11NwC1smj9qAufnV5oIi0yXijvr/t9p1WCJQW/2j0UZ2d7EOmRV6Uad8pWc6jMLhuufg8pJX
vlTLleKhH857KQkuyLmUBr7vNDb5WsFIRmKDlElEDMj0OAu20KPJJpEN9SnJdwHbHes1IdQ+Bx37
TfRn/MpQvTJq3neN7qZLQsvnln8b49h0dlsgqhv3Bm/Hg4QSCt3pTNiIfesv9jU1moFr6rxS8SLp
UWgBnDibUN+rwi1xxvygsLIi0BiBaL1w2bPA+oJOzpODlI6mYDhKX/YtuoiZWyHZNgFYCXvT9LI7
lNGfhJeCYZ7SGjxRFgYC2w2sjpl5Zk4gZzmdDw20Cv4XOco2hG3fM01hz107ko9lzIqjSPUEE5AH
4HN7f4HtlKK/fjjvwuuKfjT7IASwI7vlBTMLmErFhJwEN5wyDNHgSkYgsVrb6Jx3ztgU4F9c89m3
Ra6vWOS9aAy7hhQRybs+9/9Tz8/YVgZAiCYxbisUKyspSE2Y9Xg1u1eT/ZG/o+dE2NEjhrzBQoKj
4KnoY0fBOBuam3GjGabh9t4zZVHqna8CH5blr5IOH8WO5DtYXC4xY/6KjSEBhLa+BMfpzxGVJbBC
DyeM5KgUGO9z6ilca+hpMwDAZ2PUh2ir68Jwri9XHB2W3mqcAB+TI5fNFssD7CEUAue+DzigRwH6
/+wCfoku3j0qjrkHkYqNj3OzBlKcevy9kHs6UO3e/XX7NUogWz/fCXHzzXGXTxsZlR9hKQiyRQF/
45hoYXYwF6EYSFteXEnlYe3ty8gzqjjsm5ylieb2dZPNq+8kf1mkeWmEIUqmsPR7NV6pYijm0Lfx
y6V16oTAG8MNCk9B4M0Ze+w/VpFYd8IDWFUBWklt8OCrnrq6/SCDFNH4ZBdy5bXbxGJ2DmjrOQ+J
0hAQ+G6Y0wkZ9ZmvV4giLJ8TOMHsr3afm4B+3lAWauV8vegdWkZrBnL25mUmoorOmFQ92jaAz7RD
yiDVQFH2rOkRWAX77eG07Nq2SZQY/rtoOBSU82RTCy4/OmDRtuTAbyTGHl+cI8GUhEzmrSs/e3A0
xR1ClCZj5tzn16XKn7AQ8D1OY/wNJe0R5M8cAhGuUia6KHvRQAwwT8lTvwniMjzcaCr1riZGI4d1
fxtrxbc5OcfKApA3lLk+Uum3sP5iYYosxTFuqM7UqJ0g0YIQPXmuJZB1AYcV20bFg5Q6c7YiQy6S
eX14MtGDmSRyrj/F3RKyBBE/RgyFpMmU1BDh2wMYRNIzxeckNFy99+Uin13RkeHcE+93xJ2TUh1p
OQhZ2IKHZpEkj0hfF5BkIrc2iyJRWSVm5mZiT8q08MUhm6l6MDp/JSXEOmJGZjN+nfvRCTsa7lnT
lCTTYr5N/lugNlaGPc5bKY7Tih8yNA6+Np80gLGVxiuwERhk9g/zVtVfvNg72jmlNYWT/z2wiOE7
WmSI0Bg9yzFWJgbQuFLXrGf8liCNrElKT+wAepk5xq0GVw3yxrbwrRbu/QAuAScqMx+aAMHe7TQ2
d9VqLIpeWu+qQcS8mnVQZbtBQEWU8Qf6Je/JMP62U8qCMSFVdPW7JqivXZQrN4OMfMHUq7HeeB5a
EQfwn7Zt7Br2DsUcYNnRia7Vh30JFW0BKL72dlUZGU4kLlbxpVIfWSGQwMzQHgT2YxCwXWAaTR3M
uNFR
`pragma protect end_protected
