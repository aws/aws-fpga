`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
foJ95hTmk2gIL1mHadmZbQVpWm6gdInvLlC/ZhQ9cySWnuW6WN7UKGvm6b+r0yBogUwtleZ9Zffa
Vw9q6bgyhc5k6BP0o89bq+JjfezW/sgSlArg11LPEHnswW35VfMzHM/njX7oNHm3y3/p8GmFVg5l
IC6AewbNtn/VgRXYQr3DYx5AZCl7D0KLqc8e91qlj0gMTCIHquEFBwb9//WR5sEXhsiyp9jS5vju
W7hiX+kKvQmXaxmYHB0oJZwpQg2Wn7BuWJCh9jEUVMJOmW49wQzHA0+HYODYR2nSMtH7z0dguhGH
qF7eAAKXwSbG95jFDZUuIlAQQllqTVHiOarsQw==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
R4ykz9y6fn9oAhn6o1YbpeXa8M1w2U2JbCPKs15HHidwHTI67Icn1/gBzji6Th0UwEo8slWm44hp
NjoBd51BYLaB0yhM5oL0wogpjsiqeKXHIcoJgD5BTDMdHSIkFn7uy3nP0bZxxMCHjhsBTSe2TAMr
VZRGiil99WYiEPtCUN4=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
X2jLhwK/XwxYfbn8kGICJX2OIiWsAB2XLKkS6WaAvPJ/7uZ3kHZkBKnQ/UlwJ7GAAtkPSgT7TQkZ
cojVljIRIFNJALHqeDh7ZFXKpDQpMp73jti2eBXRgRV794eXTVn5Dp3Oy6789b+n35xhgpInqVgb
dBF+Bskk1a6kp7uGBAE=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5824)
`pragma protect data_block
M7mZIoe1zu0L0ysic8Eqvb7ma8QZQjcyzfX55LHchXK2Jw6QSB41c6bFybeA7DiR06Vy7TFj0cMW
JQQvAQvn21FAkmBHQVBY55LKhXX4JjLlw5Per4/EtXuy7iq/n/tcYqWA8jjSZzORjv3h8TOloUyL
slJ18kaVc5bZAbuB9OIfM7mhP/gPqwy7qbIhtNxIiD/wZbxd1ICSxhDQDrR6sAoF69jxMPdiYdl+
Wh7kL65O0NevV1K1FuFMXNv8hDGyCP4Tsgge9c6ZuBUdPPXjeHnPofoT06xOrDZVRTSt6NOBL0L9
qGe+vWwG14TVSqt+54nqU3w23TxMkMjDkB2g/bITE5Xie9IoaLM5z7DsiXd8YuTTPEWOhc7+w4SX
Ul7GM9h0S+C9idUrMM35HGfosEbb0O1Q7pNjtEmzRkW/Mr6nPZT9Ad2gQRDyenUrkRfA02psPcpf
89Ksfejnur+OUPNBNaz27+9f5Sc4252X3tZ9vdYqZy2feUhAj8/HIpd7r51EEOhb5JdIQSUM4qN1
Dscn0mEMQgjJEfzDQ16jbEzzoEicqdsqDJZV9JSRn2fkzL1yImTjUztlQOlI98afxE1SSm7CHtgn
YlH+q9X6WWIrEAT+K/MejIw6+RzoNdC3RI+2xISiWD6Kyw3C4IpmrSnm67O3ODhF79Phum0fqRmr
m3LvcgDHMNkAXV4GPlc/nLtNmf7r1/t0e+dEKd47R7EiV7ocuNX0EBmGyDjaoxdIeC2WrXtqhZXf
3g6e5yJvk1XtotgnJJfGauRbr3Myr3/8L06yGE7APeSXZlHtEOak5w4mmhk2jsXL9SC9mFMLfyY0
BUTL+U/56pbVt3XPpQuyp7VCeEeQiPSSQX2idOBrbAU1nnU7YyYL9Vitkd7OpzvB9MS5/xDzHEqq
02Qc+YJwTBOvvjNm90TgMa4bmNiFD/7r7K6Ys5eoLkjHpcMK7SlMbWtkrcd7fwuO3EM/GVv9HJz8
SWEvSY0wpoWSMKtWKE1A2bbi7E5V5yrHRtbVxuOOqJlP120nxVoQQXO7pQEla+9Dpu6Duex5LFDN
t63Ylgf0jfYR4x0KxImMnwAi0RNIGKCtVAVYczGsGXflLsB+6sNiuPKDq7JbvqA6/yAkSVadmhK5
s8cekk3nYNnO96QWPJQzoTlPgIpQZAxuC44ro9v2uNeqcKTKsqy8H8H/Hh4CvGlwXXW45EvAGCGQ
H8Y1tkqtUsxuFHYBY9r0N+XvcUGnRzGIdli6Mg8sSJCPHk+bgOZGtTRPi10KU7n94XFzVXc/7kd0
KdYtZ2maUiVX0kdwzUJEweUUD+0xCk+6JBqk9Mra/GJPOa4w+TDT2d9d1e54SzqSyc8gPdquSGcX
wNs+c0iD8GdNjijJvxdXRA47XdrFDOGbWIlvP690imIVnZU5MWR/IPftdXbyCyfG8EwpNumKcwX6
LyOwwDC2+yrMPLYQYtJ3ncLqBWj5PJpp9oRY8RsCATfx0jk0q8Cg0+hYQEmTqpiQYwUTP+WXugIH
ne1lDD9SSIX13OJGpV1dDUAdT6y3mjkxXbQNjEGtJ+POnLforCbmaK4jZsAmhJreUzf/EkqYoBoq
g7Hr/M30R0GtIPaQnjnsGMMOy36IfNE3UA9ZTuxA8edAPGiZYrLLpM9Utwu9IiKo5mundfBlPo4j
Iv+GQBeWNcdi5iLcd5sHXDWu53FQmGyC4fbVH7HrP8VAMe0sL9WdNhj7UsHVwcdVjqIe+9n+Rm7e
qY4eGbofDtqFnlRLQMntGoq8+XN3nwnRHoe84w5CRpkHo3JwHEw1k5O7z8WM5dD2rv5Yuh0Iny5r
2tD+RHHUKeqXB0+0m/DJuqCC2EiNcdFtrYLVNmzLOnBtfHyqAgTGJVzlHne8rOJ+MaMVu/WzUYTE
3rqClc/2PoOlEOFNEtlAP/EI5SDXdDdZzEnA6lJC+Q+FJg1dy872iERAwfCSWL96tX/73sqIlZmy
w3BmYou4Bj78iUialmVbkJ1cZtQR7BmRTuA48t2tSMKylaT9/HpgZLMfkDFduKxYZa0eiMVuu/W8
Xw1VVWGlUB+D2Cul6mrPvTp+MYQJP2BbH6rPX8KNAzkv4dv7qoXQ1Qp/I9O2GiKeGEQgB6CLSX2p
Fx4hSlr/sqwtS+SKyXZLeBDEVqC28SEKoGCzR5vwjKZhiYpbEbg/vy3mZ19/ekILAAg2QvlboRA0
QOtEE0givZTpt5Op3dfI+ThM3cuRzDJyKd05Nirzw0vwTP4O9r0bVborpBJJnI4PPjMhSbmJntVN
RHsbTFnOk8zIMD28WYbx0CPwE7KUjIuFhvs8eGzPq2Vd7JtsaiI/788BfNoMBmplQPJnPC7nFXP1
BS4/gcYrQqPvC209cAi4MLCrXxCQoLSXpLh6zEVlKJv3juogQz3/uIrYe39P60T/HlIYtDurxIGs
NEosngjRxlu5TpttR3cemlLA8WHC6EMYyq6ycvkoQ7YepcCM3SIqyvQVI/wIXQGAodks0b2vIsR8
MKdf2mile05ckJIlXGkxIBUYxRTnNVwD4m8QfZpgdvoHQcs32bKluQ0lzT9Q2ZIkO46ig1B8gnCi
v86rBBrTqWJ3M4c92UTXIhsPR5aC6gqW5EbqE527xb41fpP6n+ZsnfLzE8zzjGikUAKMsNlnc7Of
0CGiCQT2CQ6E4bzbK4ypTqbbWztSg7kd55gbdAeQYkG6Gko+WAC7iqFff/eOmlCsnsDak20kCN6D
bXr0uehl3Rl2i/3YxREC4KtumzAXzSdq4yURPhzPbC8aK05daEHxp7juGWHUPnBFzbQbXhekmtmI
W7VmnXFwWyvUgQ6/wlL6UvGLVyE14P+Jsj1q08D+cakLWBk6UiEYBK4g76POopAGQD05nn6d4X8w
xU6zc8uLxxyNLYFpZIroxy22Nyzy6ZqJ7aQSBoB80tPedcbPv+NgcZP5WAMwRm848RU03+CXEJ8W
JnXCKufBT6YHuyDviEctxT3rwSZaUm8r9wmqDmuG+b6fQVhjRp2r4n59ezzT6iShqdahQV6bGhgZ
SZtQbT1luAKiiJQdon/fRio7y/Nvg119OhDfQsgnhp6JaOy5Jog/aKW4plytcVYMQ8fH3ewD/UYP
Dhp1nWCp/AvLUvWG6AWqwc8rdU8gmrmcfaY1hUQrQAzmPdk9sXMhKWJy0P0Te4iNyKgC9naD8c4m
t+wN74thUhJO+h7w+gIU739pANi653xi3nvf3Twzk/hJqQP02Jgxfz6mPtoI/4eBQVLAr5GRyWM/
4QA8iwoA1F0BDnbVCEvGK/EXjYIkQp0WVuW6rhpPS5oOhj4r5sTHJH2bcpZ57YoPUU5sH7bxU/dw
Has+6gXRR8S48R4lHCaFaaERik1jI766hD5ELweG7j96rQbMSxyyv58R/md8vFvu3VGFgr3Y2Vtg
kTDrqnrsieF8GxSrbPeoAFlwjEV+U+8yZASpQYy9B8mdnB8ezlhJrGUN4A1afxhi4WtKpdvxvBFF
tv8+ewCi+ilGHlxk/gIH76+ETnrfuGrcLuS4T7T/Hgt6pLoFJ+fuF3aih8LfDwqvR93FqEz+h8Uz
+X0R5PG51Pq95tel2bqHp/uMnwxlGT+IuUr6iVc7YEN9saV6GdPxJ0pLTEPxHhuGTMDkAi2PXmvl
YENsgBDUjwAAAINXnzJ2f6RJ1rXIBMAlRGC52Qc/1MY7WwPErHUKNql/LCGgfW3+KE4vvSc83tkr
AKvddhrpaPPM5muK0TCJbYle3SVm8YSe7WpiDK7PTEcdOJvrzi6WAiRF13tzoD3qrTe9YWBLFRZt
t09VMiPE5cPluRg5vrJAkl9n4z4GYxKypaRzVjMP0KHUxOfMzNWMg1b1UVKAMeHqyr76hiRHzFZ+
Pf49VhHxitrlweVrXalxZZfQaYII4CYvTTGGCBKadjgMGMWbNhL67h5w2+SRp37G73spaafDDmfT
pkUpQTtx+1jcalyDiVdGiFT8+bpZoezmPgZZzoCw9TqfO3t2Dgz0oamDROvOveekd9nfsCbnOWDo
oDaB2I9rnw3JTrsX5bGnQElGuoZ15h0a6VrSMe0uKytu18o6n/phRU6WNi9ucSvGaki28tvbPy47
St+jMNAf067dYJYhWsLu8AS1iIhde/w0YJoOJ6cHFMkvJ2ZyZoXVWHIJeOFHLTjyAtyjXluiQpOe
phCB6b6fGthCMFliXs7KjQ1o+/3FW8tTWIHvzZFMzROnQE7aIboZI0jPnz5BX1XG3AOEF9h9Ay9q
6Dbt/odyl3qTMTSsNxXjgXmItQZu4RutYiNeUXuFZNM7TJWOEcjWMAG682SKfyJWsQhI+ZfKIZMP
+M4LtGeSSqRS+Bc+mucB6JLrMzXfA++qNp8MuYqBsDkEhr4xIj6YJwRa/SiahodozW2zd1qGEOMB
H4+vwzigEzaJsCvhP2VrDaReQx6IEDWDY8OTeaHdkNPOq2Pbz8j24n+XVJWOS8vg2SQUJlGk7cLW
KcxFRhRu37fu3uMyMqYn3oMtFjdUTG+zASO6bTjU2X/JDJjP13h9v3hqayclACCvtcRuAahFoK8f
wOQvQSWnStSlSl7+s0Z7Qf6U1qKizcxXsTv05mNmcOLPa24v9lyp9gpJ9ODg5B+hac21uBm+HqLq
IypLdTPXXX5Z/n0yUGCXSSOAKyKfQcMqiGoQ7L8HOl+NB4HEOSSM8Nehv9MVcVXpr5fog7ceaDh7
UEokT+CJbA9vJvhY/SVXNo6IOMDap8IOxvJlRblsWKSwdFsmXA27nwljLaeHlA4VI5gBqVniwuI7
vhVpUW5uP/g6m5OWPodZgi6qiUf5uINLHkJ2P/LKPrnkNwtmfyh7fUgAjiXD0oM+xQnoPs8aoy/e
xlqk1npxLbkr6AASH8eXoXJzM16NqjGcCY1Le+kWVkUTHDaBErc5HSfdCkTVXQiUIUTGPCyEb2G9
w0rDCtTHTUINgHtLnHm6XTF+xrXwu/cYRF+otVKli8SRYpARPZ5nk6L4MHU/BGyv9qx6sXQaIJ/r
Gj51EC4J0rBrLS5j2lXU+FoZG4PgtMIQ8LcLxzfnFJainlGiW5SG6I8hkgoi3qxi9jsXN1vTYQLk
W3zPfmritb7YpuPPVmp3ShgYmWOc3j0DAJadjlm8qvUKLWZaHy/Rh8KHVudj/v7VsTcRmux34swJ
snhp+IeX6bDP3jDB7v0wk2dkjR2V2cFkOO+NsjBRC8ZERKMzKxfx2UJsD9ePx5KoCsaHg8CGxQ38
aGmdwwBV2e6Xz8fobba9xf2d5D57tmDaY05XkMVEDJs3gh1p2Hhq3KvgH1v/HuJZGNkWSadQv82f
l4/ID8NzJr6ye2+QH1TBtQwoSonIVv7SjKiUfEn1eqRdnfM4BO9w1tc/cWXx1tMsKPypyM21JKok
A4wYfQkBX0a6IeVGZNtJIEfqFCKoSMzdmGStCuwqB88Jxsp7l+TEr0FuzMNZ2pV0vv5PGS7+weZ9
1XFiMOScFcCzR1wA6It97kXiUk656QMUY4JHJzHgbA0zKjoHfXGP15v7306gyx+Hzg/H+cfeAyL2
y/SBrDXfK0XfLKIxtPH/bMqNluJddJw6iOvEOqmJhDqwkWGVh3VbsNwCUPRDwRybDn3zmDRp7++W
UPLDk4RwgvuGvIN7s/DO32HTA43nGG6QBcu2G2xsyf06yCL/ryBLcg3Tg4TkHdmobJYI6I03WjUG
ckgmzLJsaLiK8Up3YWxwKZsM9JvRj4SOEVlAqhCMfJxudJb/GFJVhY1lP07JnsvwGGjy69icKTnP
jNAGSwyejoMmNuPVKNALCEVM8YRZUMjz738WfbjrTs6A7t2d02NcgPuIiydBwS+4W72wY9EI8vmc
AZ/07y/Phdl9RrLccEk973kEzaIAf8xKD13Cf08SMs2rwtB1er2HO9fNIBjtQHIO09Frf9QxKnud
PVMLZMJKyzV3CSGDSs38UkYY0O0OK7r5/SsAWzo0Cgdf4ls06LPpBAwCLD4TTbJ1/5vSCFaYsQkB
7gT0rHZaxSX5t7df1c5XqraiRYtaXvPiqFeNbYA1I2yzAj0EydjevPF84IqB1ypjEJoIWex0gNoF
HJ8KKgFKUin+3fsZuR0txl9hPhsvBS6io9vkXr0zIvCm0F1Ma8p2Q/Hl1xOSoeH6Wi+bFUbFjubp
aX6FwJUyYDl38uEUHNoiHVDemGyDD9VItF8rqtxUtFSamLFgKL7d92msxYLkjrGSmz4lQ82CQXoR
IXI5E0XWeZjmdu1uhQHxf75MMT3/zb/7WWjB0OwVlo5r4l/6ZCbYEfNEu3FERya3ClOr0vWce/XE
eQKTCcNXJDf7Jy80nLsuB/mjN8uHt2+60vn1CqCtVD2gtlYu6Gl6baHwYBkATMS1JZ+aV/gcZrne
cJebtifYyEYqEH1VNgLU7IQYTNl67jgF3Dk2blLQM8oC7SYpIR5U+ONXvE7Y76Y84Dr1cxJw8Fcr
/DoYMUaFBGmPCRzImdPGaCHrU86aa49Qf2hDnNHE4aGHiNUllXSk/xVu+FTZ33Yyxa2PO3EsVI7F
a5MjozVbnB2chFUAzzN4ikmyzEZGtHuToCS8fKOPvDYFayp0cSKvdcMR9J/uDS/T7cncVAAeFU7e
NsocZGg6gTN2fI2OVkakBg0pUmxDeAHaHeXLm/+x2t/7g4awNzPtctq+fXR6BrOvb37O1WRxGHhb
VVQj66NduFOxzvgFnWeI/ealFcFKJ+woFWvZjIhGhzibHoq85S22i61sVD17p6A0V4qhQlgM7NhA
F2n0tagfzeP2rgrdZERJErPMTI6DK6m1Y0vNUHzZ/2t7iyFaXh3GkGXnL0xVcpnJVOWyh0QlyreZ
Bj4ZDmTkpCB9Lhn3/qFFZWqwwbca4+0H7bTb71olKrIkXLkxPbkWQbHVVJjkjTuLqhaW6NCCVUuC
HXjWQkjlJlPBYYaJcay7aE6t5AaerUJkdnbdOukybscRxJIdqRn1+qCUVZEWn6ffRkmnRVOEbVg8
2sGQMMplsffOh3D3LcWjbXswEvSBz/aHdRtSO0lOVSD+uSXL18kdsl2GPBJ0Snvs+rlDa8NS/2yN
8fNZfmGZkGMOfARnSBXwmD9xDO8aCcw4y2zBRHtWFhKuvqcKZr05M4762yv0HbJ8d65KtEblHEwf
qwf4PHEFoFvnjHIrRFVMQby2GHaVFK18ZH7yccq1Hd4e9csoZ9isRT5BFpG5yJziSfDkGOFv1Z5C
eLhHE2zK3yb0XJCCs736+8QTpoFB06sT+rard82Np361yL3jhgrYGDT3VtFmYWk4bVNct0V8PzZa
PZiMM2QO5cqJaImflRPxqh+KDG4/iIYifQwQc2gQXUufvkAs/sJj+Lfr+4BKzaLOrgclw8kuBjX5
QRNhn+7ZYuOVqa+2yYJIH6b+olSouwTt6qPBcL6PqqtMm5Z7MDaH/5REoq0ppGhOp0HSjyVj2/3q
MFpKBXr+xh/9bfPZ+4LUleaOBxa/VWeqKuhxIFdpm/5+wnFokY8/6VZ2zx8S+F+9hxz0f9SFCpBy
yBYvkW9Fog/l25/9xaktezrESZ5KotQCjbvt8jGuzzm+nU65CvOAfL+1FneldEjmlbTHkrZ6nQLW
d8ZGrc7VVuhDD07I+WguMRFB/O0oKxiRkGBMrfx8hV1s8mDIo4adzaBwyKmDATcFX+PG+1OsrFiw
RTBG8lc4XrO9u9bFaCnVpErPaUL+JxOhrfYoS0oCBDldCBB3kEcp7uDFZFJHGguAmj9AKqY+SVYM
lxt0h1YCcx81Ng==
`pragma protect end_protected
