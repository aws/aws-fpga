./../../../cl_dram_hbm_dma/verif/tests/test_null.sv