`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
lwWLYpurGDQUNKI3KULuP+Qv8KUTy5fTGlHxW+X6JAfYer3mvPIm4RfkKv4gDQAuUTzf8sW+c7hr
OJiOAtmHq7yO1mWPk2ZKZlBWdSejlGzTaeU8+cn8lofIC2C4W7v1dzTw6hnHD6/zUIwbIEtFe/Y4
eOxlQfjORdQx0Zpx2rwiHiDrgiKpOyt8AIqpxewvgbBImjG1SbWeufCEQkwBtewyGEIxz6mdFUpd
cH3GQFxPQmJ6iMIlhj5NP6dBek2daJ8YManMwXtUHW4Qsphievok+GT7P+epjojlET+CcLtn3Rlv
jpDh6uwP5V3Y04tIBbCKa5rMcB0u7QRrgzh1Mg==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
ysTh04afus9RAuqaP9XbioRKSBJH3K8g5XzJWWauwZ9v0dJwUS+2jV5KWVfd1Wj7Mqt9pDTxU2gJ
s2ZTRqhHaCpBeaw51R+t54zaqmhhfJuowQpNDTLLAoEbLRkVInOjDi2T0OlGq/M7Shi776KvEARo
NPhNmaGJU01OTUk+7mI=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
MOCuwjUMuaGaYhvKzwDqJZnHUBohjJ8ilo9tDoIijIfcCL5y4r6wpfVDz9+UAqLGtmyZhQK6IS9e
XFe2S70BVmgW8WGAaDvxqaIgoSWeC39oiikNGIiCjAcT2BjyMz9sPvIhnRZL8qbqeZJebpztxNoO
z7xIc9W4cqr+Grm7f7w=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3248)
`pragma protect data_block
0FEKyu9+D5E41iMtiZdHKdRkjs6t2zX4pXmmITIeJ2+jqS7tiVnD2DshEjCjiGY/LJjj9jMntz8B
dLGyuodHRF8lG7aJKo0ae8I7idtMH8vs8uoTve4e0ubdrHYDrnswjLYVi+G1npx3ZN1JEECbaWXI
ixmZjiV+WrgjMtViYVPC8o0QbnQ4vBpvuWTgS1n5N3WuDXFrzqqWf9T3inAInsN+whN11OJIQtUG
y4M/WwW7d8ff5Bo7e3bAFDmLdnPTwDef+C8a1GiSZqW/GSx/Dz+Tz35/LQhgrEektbFdMV25/s2f
7kogB90K2nu6lDKZi/+GnhBp40CyjXqLOzX9g1S8uxzOp0OddQ103cCCHv3dxD/0VTrEgydWko1+
wXpE/GFO/vDzjavUUTj06sUaeTw/uZKjS8Wibm9jcpY7482CKMv/bBzsP2YhPW9bNlMWwOdejENA
cnxJfhzecywvqwPcsIMfIiSUew+0+p9hl4txwKVbWREMOpZt6dCbTYnZz9PAFCGK/hqIuTfw9OmQ
vB7z09HL722lSRM6whm+NBa+hHhBHta04n9dE+ffgEbXc45aEtXWePo9KRX3PbeWG5a2WFz9Teno
xValeje2XLc3PUIoo0z2rf1+GR7AsrVBBn20Bd/e7P3eOjPUddN0i/o+xAALLRE3UVUqpzNPTz9C
CCfjh+ViTlmqtOq75IvmKD/I3pe/n4SHbPzTHIRfsBMxCYSRaLmJSvBBdLJVRuEDblBNTqqzgBOY
KIC2Xd3L5u++zllWl3lOaaiJ7+QNT0qS9lMBa6WA7R2TVuYu+1M3xIvF0Nq+f9qDdmxqjqH6XRLF
vrtmXgDakmeNI2WOG+lXSj5ZWBm46jzS0C35U8C+3V33s7LQl1h8vi1/hQtgskUEgOj993pwZ3+r
dbjes6bnl/itXd+Ktepf39qXGTVXVd7ON1FUnpSvpIu97De7QFIXCitvTcpxzD0HfrgKdhRcUC1j
rxi/Q+bRbZAn1dBhmivlQtJfn0A0FJTyjDBJptB3OpZO0/MTRapnzZTlXBJ5X7Ftc9KYZWoA7prM
9yC0eOrVh2c+7+QG1/hmW/dexrOur1KPNMqvSZn+4CDUffzAh1v9itoseXYOxppCNRlkaHS/kr8Z
L/MgUQv0pc1OsHI7q7wwkxzy2g+Skxn+J1n1zRkM1d1goXCncd7xqDAxF8zDJugIU+GsKvN178gB
M0zJyxOjqzJC60gvfKgMbXZvefc9V3sKhkfP4bTU0X7FoRXjqqZVY772+51g/xaWMgX3mcLzwtw5
+bed62haIf6PJ4IipV2CZYR4diRZ9eHqdLmPaLmHWDuYI/YlQK5lEEPYfViX//IsId4LkMT6VK+z
HzKsTRs18Q6kFpluqaMNqpOyxCDkCLaps+IVUMNQmyxRPpOUyw38uJCbPu7r8UJmjZhg5+6POSR1
xQt+tV+NrWt/nXa+QF02Ydrdf0H/sXOxAVOE8rkWCrgqa1p9qaJMI8zR7I3O/XLONbNmNmSo1VV+
216pnx/bDXaWQ4MwinsdlKdlEM1vNOBjphYzifnkV2jDWvUEgktDHWgQjyrKlN72JVhRD6uIdwhe
hbvaB8fcyfY92jD+IA08y4itlSc1SIyONzQFuqQTVSQhGLZAKBe8OI2oDOp0NXKUTFpoFWzCBfpd
juPhHMlR0mqSnljmQnJrrR5uRP+kQAjT4779lwTpo2FcRKi3kYNvDTt07oU7yRpQ7XYyeTMawZbl
wT2SC7l1BQPTEWJ4XtnYiPhr/S7bkozPvEIsL7IELSb9dvtcK/eUIs6cZDPXagXQA7uRe+qJutQ5
+KXfDbjOSOeV1BkAg9HlfV2foWcBzh7G51ibPLHhE/vScd0VSN8ibTxzwmC7qVZBNkQrToyixGi0
AOmd07hgke2XxB+EYHecs/P8mRWtKgdiPoyutwedjIXSLjiG/LtVZBLDiiSketUdsK0whq98MAwn
Wc/AZgz87Kx4c9IDQCSbMiFaqvEEwcSxWGKDsHsjn4kukX199bmeNVgTd7ht2S39INtBY3HCRECt
0yBbUGTaVZm67zuatbYki7siH8hDGg9yPXNfcaFqq/rGc0/o81/4BcvbmLEt/9fr2eVr9ZsQaT4p
fUYHKEBBx1pBFwWpnuZgenHOTqmnRJY5UTC6nquZkQVBRqC7g07PoctLDOpstIvk3SA9PaEV+SZU
bcZapSsJOVF4CByawsuN48fwbhDdb++VoIqmWu/LuWXjyqH3/U1G7pF3cyoj+vfyRwIvXPsQ+Tlj
EXXNROmkgnZofUbA+D6F2IIqARNJNdIB8tf8PWOipfyMAiCobJF5KpkvRvqYh1LXI4esT+FqbXnU
mdu1xp+Esnsvb2ti0R4BW+oGzPL/npNcMf7Gdo0RiQ/pftKR7c1fopGq0vVOFoquauGKyJQuqLFv
HEvopKcb+/a3z0BKYVGFG6m+qdst43AvqtplwfINrGDB050t882P6ZZNxcpBcbCQ7VWpQ8prwHTo
NfL8/6IpWkFh/58/C/eTE5uauDBhwQOzzQih6PTI7G8pz01aQmpGMYdtxvp309ovuxMBVCuqnUM+
Oza9rFU6N5LFlf9KLKt9lfYyon1EY2NVC67pN4kI1qhWzoCCRY8M1fk0fabydSrbDP999Q5eQKcg
zz+tsXwi93tlHi9cCKA3znwI08RQyju20LHsIJ654GguVYBdYNq9hTpCxgsmahJhGc7wxQ31zXNj
xSNqQEyLHWCGGUTEgeGnDr3sVy1oNT9H178+zj6wucqVJ+3jmtjNlHHQRDsTFKw3sYB1vDA3ik/7
2WMqQ+7RINrNYRMYB1S/Al3c0kLdjhZrIrKaSefn/zaCfaxMPD+PBXu6SLSyil1SnRSEUPVAQLB6
h9oydUgFl8KVgtlL/RvCjDpzLOgP0I9tbhgloiaX8BvlBlb87vt4Jfk/ujwWazha/b/OWymRrU1a
faGo+TiuczH++saVAfWCBxH7T9IzY8TkmeBz8l9nj/7f8EQDRWWlpQ5e4eyw3dptPzdBXlcSSajQ
n+85Os29BAFfnnY6t2IF/RP18JMNOQh83NAVFkAQjMhgEeUfZDgA5YeBl81QO5V3pQMOG/CJH74J
5+8GWzd3UN13cfjth2r+beNGtlVa/4qmsPDYjFOaMPPvZYDRpYMfsSzln26fjFj2CqVzQ817D4sG
CJgtuA3NrRCmZ7JAQmDE+SOQoXK0w9WuFHo1AHLJER1lm/auniu+wMYCGysN2aiOok4xP+jnDlYM
tGQDXxWyV/2qYNW2i1ingXvRslFvtOb4NXZII8Dm7I8kGXtUvAfHydmqTfmrsIzlk+3GlKZA/afD
V2jZv/fnhGJS98k/zwq01KgVT8uRFNMp1XRcme1Ojvog5U0bEEWZaSwJH9GPZ4yIkfK444yAco8e
kZWNrPfxDFrtW728M0N4rr5ElrU2RNhjfx2NZBBhNOQtZY+nQERfQrj1zk+PBGNj3VNzn5QhF8og
mZCzNAaGP0fQl0Ohw+9JgncxyTFWxZAIcsPzF9Sq5UGvHCvPuz3I2OkKxgVcdBUQ18I+nv2p80lJ
KFLld3u3RzWldMu28AV3UHeULzPR7/UTJbfEN4UgEEsIlQ9229Wxy+j/CezW9UwO9BBAxbwTwqPG
c+ZOe5dfquEeeMBGuQ8Uqle52qDY8OgIYdHfA1JJ67tJmWZSqRsO57W7EBTwn/AugbLTo7Spmmu0
90San6eeqleJbwSCP/5Zt0d/bEKOIAcC7tTbJ/GfuXqD4iE4wLIHqeump8GT95N+LZC9CVUNmJ2g
xX2Zd6g9qx1fnJd9XzO7SbGoNoksliIZSDS59xxV4dBHhwjr2tvAUAELJaBvdasm+r1jEJpaSI6d
CHTyF7wDJuRSpYsxWKGhdCERsTi4VK/17UZzr184tyB5rwsvdeLtjMR0quAocD0y51gMPPJAgSh4
j0thhNtAwx9UAnIXhuWZo0eGspBWCCjamPfGwrdnAyWhOLJuz6vyWgoW5uhaSaGx7Y3iS5rBH6pA
vZ36qLmnwy+9J5K0ch2kOeoY/Gky8Yrx8Zw+noD6oskjLhg5oI6aWGWSdADoNC396zBKAzCU45wD
7rjT8TGFEFzJ4blFNugBp/V6X77yGbn2XOt+m+NMMb3PcM1AFa5tqG9G+fWQJjPeMpdIITe7THn0
FwqafNaBrXJU1lsvpL6uU12lK3A9KSoS2EUbPcTYOWG7t+1hZ97jDFeUMMxdeaWkiGLmKl9WQrJ8
xYYTafVO7qI2vjbHTSaLeLQFfbsdofSl1+UMS64E/7oNxSrkZqsw+tSh9JzuSeQRvvsg/8RQ/+o=
`pragma protect end_protected
