`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
OYNKDjOdz4rbT3ynkhZ7ubi26zW6kfdgQelR0zpVWqGJTXNU3fAGQ1+TJRzFnrxInV6jDCZJF/dS
yCEDrx2cQpHLppDOVpFL2pNlC3jsWwtvCbz1iweQW8NKsOIja86S9euGMdh8th6zxt6Xr9qv8oaC
A2K+Z7AlzHkXJQuQjLhg5dcD71gLOBpSrdeJa8m3gc53mohLvFggdXeCnE6SGHWiqRhCUzsyTuIT
3bAjqv5t+2omZMfxuGfaqeZfZ0CVF/tlGc+EeqLY7hFgx4xmi9/1+qvtOMq/v+HXhJlreHkPpoBL
fQbNaTP0Za5U6QGkzY8Tt7AAV0uuvdsAZxASlg==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
nFXgtHwvm+Mfwh7nLEFNPXbHcq/z3CxUE5fVKGx3RKn9c6X0JnTYyD1GIljXAYAfyXSv0EfjbTr5
KTTVGTD56okOlgTrWLP9OWWqOofkGOr1NYJGOMA4/+hdyAFftsQW19Kx/C25Pve3gOrX1jM6kmE3
lEu5xlB4U4Fueb+h6e0=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
Mc9g//lAa6IwQnM5UXWpfuilOs+IdRZqhRvHiuRYioMIH5VzdgjzZ0YWUkK8rxi7WDgUp0/N1RWY
oBpU/2wnuoCFwt55IpDFfD6UpBKXTV5OM2Gf3eR/8Sq1FJoa/EaQxbZ2Qgqf4ZNJUfSjU91mmpK0
Z9VW0j/ioGsEPJjQz1A=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 17568)
`pragma protect data_block
7s235GpQV+6IR9ovjq43jOxOfI/v6/a2tvtuxBuAQNDio8NUfGtOikreP0PWk1GIn/BRv2rlXwnn
xPyCHrECaVmZP7fpu6csx36Ytiha6sdhpYnaMJKMUreSKe4qvO/DfnohymxWmDt0yZ2EsBzKsfF1
/kX/jJXvoYb24NHzYaRoI6OrVrst26fqQoSvmcQf8WoIYpYv89nKmDN9kbEVH8YJO+z9StXkNvAT
WtJ3x+HMg4ze6UeA7dGBw7hH30DRBs8rYn2ZjWiuJFxq8LATgwJDY99On86b9NXOgGcjEcxjxh/s
aA1rM1ezAdFRJ+3xVNMlVZFX/lXwjSGMs5apP3MLvSWxaEuNHbUnUsHn9uz1OGTp83QVPldOCQex
kPxZdD/y2JbMQM6qy7x5E/zSi1kegqtBwMUHgRuMYrrXWwu4MXQl+LBgq0c1ZkVPwTbg65N023za
F+0rY2F2buOl81ktGomQISZy6I7a8aW8e0nW94OIQ19UtWIYaPEl0RDBa7Ymt780by9sIN9A3Uw2
RmfjKRWp0FJgZHEjlYm2cn6lrdt+wsX8B4RYFcU2R8eEcLpk9RzOhPHvSFyAosbTt7XsNDemaGNr
uHWRaTlFRy98lXKDMzgIyObpAiWHrOc7HVeYqkxG1GvJ70xGuglS/KffKrb1OvM2Nx8fIhW16aYP
3iQpVeat5QDUoTd0A4RZkBtxhpYMgprdvJzz6/Yhb8DPERPxV2bso0YdjKfX6p6/NRSv4nTnPz1H
mB6gQpPU+qjkm06pYdM9GvwBQ9qfPGLns3Tcnns3gyENxqcmN8Xca2oXwnR2XDGSf4qW+SzBRntM
XWnSaDBKiIC9+USZAFgZUTjTSrs9jprfDPEzfSYpS0HIHbsoWkOoRb0NA4z27QgdaJyNeo98j1fG
Frg0jkloEPQxzkt7aDNGaq8zw+HNmcdt1bV/bXTTwOfsJaf0Xazuuk7UjI7+Yj/FTQVrYCskZ88J
pHuGv3wK5Q+Wl0Qz/Eo4FBPolt/DmEIoZqiROa+PSrBlDlodKaTOobeltvLGRqJON7Arg+ldgFpt
5pT/SdZXM7HJZWlDWEjtK+0cnBDa5rNT92Ewj/PKv9YdBIQKPDFQKhyLmdfVIKk5FZYogF9X4/1F
8/pAM1/bcqu4Nwaof2F/N79tmDUGc5nN0vEh8DUEkYy0nPuw5uySRQnNHvLtub+Uu/x9hl7ERUTo
A//6e3nFynMolW0AF0ihjdwMb1uyZ6IubqTBHx7BCBrR70YBzaPhmIEwlSWkndVJdHaNFmaKEtKc
t+pA0FrCAtMMjxFXnRFwMQCZqMP1bUunNs8Dt5Aid5c/zoiSXgQcPBpwwGsfBIP2aLaHrvlC4K1j
Hc/5zAgZJKeE3OUyrHyTYoxKTGSH/RhmpMf8O97UXjLx5ngLdXETdJnUcT//SZ46y0jh+HngIR2k
zb1LWwUEit6eQ1Qvei7OJVIdmjpuO3TkZk60cxm3qbOI/dmpTu5ElOBeuHEe3fTMFvRqr6wvmNo/
b1pzKVHxmJ83r74GfurRO5chZcApEGc7xe8WugIkkqQV5pBnQpzurWCXyGiNTYj+ZdM9wrZd2lRI
G3biacsj9wHqJo0MgEsuZn9im6myVSIl3lkwuvpqPpiW8j0VVVwP30fv5ydAbk0v5aNLr2HYtnCX
rePnTrBft5p2YZXPv9+qE+mkIiwAK1lXEwO2oCfZdEitkW5SdU5qqRW97QGU+fqUuCTkmBaHBT7E
nAuRZKOKaBUR2+y5hiEysRr77GOvDPiZMA7tZSrQzqwKjD4Nqi7DV5p43IwrKETriYWgRxhWla2X
0Rq4uqa4xef2aN/d3TpxaIpQvrR5s9MJs8eIBbTlPvDzaV1MT2s1AjBMroxROFhvmQ5JR1nOI8Aa
/Li2ESCrfaaTnQDWRVrVMXdvZN9YcKU//89gmIHAw2FbGsDWTz0LA2GN9o4OA2xYiWQhbf9ypbAy
3nstsk7r7VeA7jqOiOfAHlCMgL/qUSm+VgXMaewjUf7RRWSNvMD1f5vnZ7LuKwig2k+L7EjVP4KH
6rfXKKZ/yHKdfudMaKBwQ3cPmoF3Qx8xdhNzIjQ4BGFn2ezYI7rfkxt99xaqF/0Y8NH1NRfIQHZ0
DTu9hoEvNCAHMOL+baYPi71bBphf6TEyCWOm9uWwjjq0ZxF4hLPVp1qFW6MRqVzCrsVgRXFZDPbx
15rpppAgPwKjmuVMGn2lpwj10sXsrtX5z9Az2ES6kND2AMEa6Wy+ZaPE6rVT5AO8ME/q+EdJENM+
cj3MaXfSLang3dq3lHTArMH3Jg2Mahn0Q2VXtcwo3DNEwtK+L4kFC5kzQrU7Zcy/E/Nthcts5fU0
dS2JHPdhPGM6TbFQY/M+Q6y4V3xZpDZDnRsz/CsfynTRQK2jIjnUFZ1pR8ki8+Hdd62sCCFKWX7h
9KumxnKp9gFG4IOntOXh5AlYoQTGGBeUj21ur6DtdGhU/WvIre7dNAvN4EjfQ74Yz6hB20fTao5/
iLfEjpK+EUt56+aAua2qRCwKppeZwyQYTs/OMp82a914EUwMb6X69XvCdl2LFf3VCL4oS8Ww+OzE
TrbeA0TdWahOXP0ZsHVtLJ6mwpteiuvVtOyGhQ45frVucfkg5nwSaLXAQziX+SI3PI94TDBTTqHU
dbj8/jMT8Bgzkf4B9bdeSU6pp/539qoiyNTkwHrSlUSDIa7piivyiHU1j1Z3XraR25PyAZTxiuo7
7tSFf5HHDYZNHhji1j2VOa4aX7XNiIjZ8/WayE0+tAfzspmaP+wAhG92wQGoj5597ORH7VrIR1n6
LvtbiVkiC0kajoACERZl9R6csNFGNGTllMXki6whA4RzI2orlId/mc2FyoFrs0Sg39pKC5qWGOA4
FM9041ZQSH6hYvK8TeTTeIkEY08sLkJW83OPYtIxqmzvHqLd2nr3x6EkKPcFvgE9cC1+E+9TmZNR
PVSjfbXmo1hjW6we4BPauRWj11dmA4Y6vwrp2g8bdm2sM3iQ0r0v/XYYSgUebOQjXZXUd+TZuOMu
2OK9rOIIkoT9hEkqD755bEVCEHSF1VpRTyAHn5RrnHlzYxo2gE0r3hNFIqRCGt7lPLBdWWgTDT7i
kWctUD4AX3aAKRr506kL5orj3CU0ogSgTqeTdrssPiAuNPbIpD/5A8LWBkJJJyzzYtSnSrKEF5J0
M/Mki6w0o42xe1ATgxmua0+yuuVygghJj2SSNGQTEjizyKbiGkNAnmZr5ukNPq9mRczVIud2uqf3
W+IjpWryBVb483WNvrLKusqLLcodFyJAJ/MAXeHpgG7sIN1emov8wuqjwX1kwG7elogcvHPnpvwn
BnmcHp+/0iOn/db3P6IRe7Off/vz2PK+07B4Y8As2ea84yoPO45u3AWxXRVCw//EHnrPtU+7v/Cr
OHPfqPvPtGte6ZRxR48x7Ys1kJhUWxsKbVQRBKCUWVYmni5ngXbI74o43SmnnWTXCl2Qg6vfFQPB
/3uTJm3cg7BSAu2//hwse7DeFnxgX/bwfvmAIKptt2hNPJV1T6u7uNQsEwRwRA1iTuMaYwKWffyq
qmvW9yRFRV7n9xbcNB4sQqyWPqu6g7hqspGU5WSSd7g0PLEsC1SuqewdnGMfMZQl4aZYmw6ShsLW
ax0QXGJeDeVMP87n6F196CLPYmjidJ5FkS/FGn867g5qn3BXMTd1rGvhi5Y8jg40scPt/E7qksg8
rWzW7aMPxo9/i9C+KeW67MBh8Vu3NyEcHTolDa93968eXYJ2Od5oMVkSlFOzU8nnqMxN4mfTSNY4
VIDwNpBw6Fi51X26o75SCyLpiceSBEuLyFgW7WWycsTYDnUwXMNPcuZc0EQemCAATqiw4gB5qQNp
GAVo7QXti8njSiSapLmEl2YbdmyK7ZTTcKYAhqaRo1fEbvFkLjrOW2UGtU8rrnz61vBbifMu0AUt
gaHkbBwAyv0+7QY7odlI1W1vEnvio17Vn8jj0ketDkSTfyBAUDInquXMNPCs68thyTpgyRgOzwXG
cYKMo3G5A4dt+dtPfI4wm5lywGBIk0Ysq+IXAzxuLgsqblC54Z6aQ+9s2DbM8TTdQCJzUePeT8Oj
yEICm3n7crgeAxnSr2i+9aRiR60JeLeTkiH6ZXPxvKYKhoKVT0RoAXIHmFfQOvb1tMSguF2+Jplg
LplkhaaRfXD86XRmgLkgzUf+6YvMxU1XMoNNNL26xRpOi6YV+GdfzrCujzoyjA5iGGdxzTp/8sGx
66oQxKI2K8Vk7QIDfR/hJxIA3vZmWHw8FrGL8MMmVd7ep+hP/Mb4XogG8/T1ffSrnWIuRGgt+Q25
skOmKuZJq/0RGiW4gEGca5GeOUjfyWNPcSgshFWLD3IEJ4ReCPaMg41hQYXKGCaGg4ERYzkqQBv/
+1kA6Y6qzoWcB0rfK/0jj4nJ2AVrgzfIk6uToNfHZJr6LtJHOFB6bLDFKbf6YzhDJYa3am3o7YjT
7PDLdvp3WrU2obs3mI6d5g8z4yK4RiTwczA1d79X/Srfz/S11RiLd0VnWYsyrdWe0NmIPGULwtED
xrN/mloNx6MOlaJIqvUm/RfSZ4/pfu+ynt5x9WjvHilNE6TpeB3u4mrEo8eV3Y6rCS9opmxncOG+
eg240s/L3Q67sj0o1Pgb97ed/6ziycJrifrbmVHtO2Knju3O2HT4xZC4GlPbEymRD0VsIape5PW8
lB0ALDQBkw2nr4G51rXVLtwZBLsG8IAF9DL6e/tjtZGbcxYi2qgdDxxW1dDoYA2Y3+LAfBv10h5n
tfSG0zNlwdU5CwIDeZwmPVqI9vJxB9yuyz3+yhQ2u5+sR5NnCHs2yE72mJLus+0v41IAKvFsytVi
n5KPhD+990mUERdjkHxta0IypG1sK8bFai6t7B2nVmmhDPVS6tq5JuFbTtlHwOkN95RIJ9cQ4Olb
BM5nyap53Yka2eneBvYxpX+nVZZ1V5U5aEp+38rya1jgUIGlu9HwkljSrsKIqgd4OSqL39T4cLyq
/nikTk9/ti5X3VmaqYVg06cgBXwP+wJnTsCjNBmzWYonjmCthtwNflEfbjUTNV9QhNW0od62rALe
A+YKwmxiGEpEWEO1nh/MlUD7MbONDQfDYIB9w+aQXM8FskuccF/0U4auIYUv6dcvSLlc3Vm/rB6D
Kt8h4X/yw0kHYYXUGy999jAfRKSAn3XtXivqaa2STbzPLHuBy2hYBTxV+5Xg041gx5zU4AwuUVH7
O+mjwf9OYK1OCpfOPbj0t6Euoc4bleqsgcd0V9xHGHUffiSaQEB39ktaM7/VvImMKWEHLBP1Fcy/
Bbd//qwBg0QqMkJ+li9f3oanDAH6u7Vc82EIBDjvQMuVyYwc0ySkcuN3CIo+d8bzJBGx2S8L7GI+
7iSU2D376Xd0W7uEyLMObZQBGMvhQguxFva8vQKLGbbgIgaGXlMJmaHU1bqUxbYsvxcXBIcBYvN1
RrT28UNFfsyx+7jK9RFAC8ChayX5f/WjkZWNL3ZAoEOCszIkUz2FTY6eNmMWc9TKHnxYbHxoDVH+
fgUcAtVB0kYi0YFG7wfXU4ZC5EVBN8yWfMzQSAhoTZ0OT97qt/3x9ymJ3PSCMwlqazglz8IuANuj
ZUEmkWyKybTH14GyHgmEoR7FMZP8N9Z0Q/9yakF1DXhMeKakvDrCMmFlI3paFiNl/4dCtYcYuHEb
6xHKqnziWb1NyFsMCPECAK6eWBoen2gDqLS/+gBTwa5oql2qndW3ONhsMowa5eLHcp42dQDlrh7f
KYEqITZL5DGQ6yxCic5eqYajaI621BiiH6dySs8Vy3175ewF0G7+NV2K7y8jjlGP3JKLtUFQS3Rc
CrFhU4fkla0wiaNhdcK6cqxXFblFmSp9ZqwHSRU3F9ACFz9ZkwVY5Q2UxRD0ZjA+Nwd6pGn/oOzI
ZE1Q+ZPxKT6mf7P9rWtiA791uTZTjqeFuMClZkkI7P+P+gmanmdaVZOxmM2C7WZUlPI1jpa1SK2K
cM+a7icTF8E9FJi2C3BPpi2uMP6Iw9A5XlgjgJ9V36oA7w0rYCKx0oz5jVcruWceyr1FxEuxpUG8
L1G75/haKXM2zCkdXam9jCwusCVLglRfHiGOPGrZmRXfUIWJ71fdG+XnlFcOYH3YqYyRJ/Jge8WX
mSq3Sx1rwiW+pjvu3fg57J1UGxYlW8eCjh/+sX0Gbx1ER5ALWBgHLZAkAtslMclfSoksalRbBiqr
M8FqcsV6tlCHw+zWnnWq6J5zosyakqw2s36WDAmM30NTy4n0tdZrpS3qd7nhaegeYJFHrTCgrfYg
lhwODNyYCuCHwXrzna6bK5pebTPf+xe5XXcZKMBl+5dQjZsUccAqED/APFnFEw0xYrqo2U0j4v5d
TiwmUxzrEIiS/4hoj6GG/69d7z0YEZPMJ+gSDQxvmptCv+iyFHuy2LPINxXBc9pT1TXFZ2Yuz8Rj
+x1sTYokk5MXdCTaxQUXS7pSAicwC0SAsHQPReL1rQ33YdxH3OC1tyau6w6m1l0IC8V2SXimhvtq
sX8zbVsNpXxuRKSP9QE8g/YjVjHG/mLMw4uj5rpbMnGBI1LVOHZgIixt+a1dTDpV0/L/8Fjd4APy
dk8HTo8NDkemiAi6SvV9GWMjY2WkCugkYcyKDgRTP/YFKIxYL3hQ8nsr5Jgt6bhkQYtOtxCIPR2S
WTdFFmDQYnsYu7Baifm0/k4Psl2pOyLyVLrq4a6lOtkD7EhYQIsdhQnfdAhSJnDoMIUli+JbvZQr
3Gs9N4f4PHm/Uy8p7XxPZj8jZfzGhvHmh9gcXbRg2Jocpk2SVPK3pSTssrpNWnR/VnJdB7gnpHH/
OAvhxlsbyKwlpkUSO9mnkLHAgmCSJwec4b6asHosHv02d/+QvwinDt8MSVA4j7YzW0yl1Ze4W/0E
iuEIUiZtSFS5yIHh/Q87e/46qn/vFW8qr/JNvp7B3W6mguSc82NzUWxJzEf9Y8IkjT8G5ZhSS/5z
xGQqEPOPxlfVDBgroOsWiacU04SIdVnSnd6QOzy+j0T+AR6gxtOd9U21/RU1PH3gTDlUa4LPzxy5
UxbDmpV61G4Vh2D02XUXdjwYYm74G3d3J1DQwP6azJdmLt/n4uVYzlVg7iPJJRX939aJaiVkMLDa
ovni9ZKBgLkTeuZFrBGXFj/6SInVWFrEkpVl0Aza9U2RBpWuyQbAP2jbqgf3klHrJpFSW35LmPTy
XviBdHcONeNEAtSEifex7FvHw7C1qMtY+9IIN4G1cld4o76ojq6MT2UQju7cyxJMtjRATlv7h22v
wUJH12nDUZIeG6paeCKzu/8rfk4VNUCbBKve6aBZ/thcGh2w/D55vwPnL3gtBn6PZHr0h+aATM6d
sE7xndmL0WSq8kuSIapzxQcY8qesdfAJR24NL956BE4T+xxXRwGHz6vrMnpeIgdpx0aEYeJMxjF2
psEEVZv7WpOy5sbTK4/HEczKJofQozHfFrfo/nrzIjSZZBvMB45sJT6b6MbOQzbJnCUlCfLxJyqU
ZRkgz7rjWCCtquieGZLQeXk4G3WrrvPFVTOMgLFFKwIXdcB+6bmqfuon99xSwhlGpQrJUxMrF8pY
jKRwf4BHCAVyqJa2Xn8JK4SQd4LjBly4khf0NZ6KmjNtv7mTqRAQih/y7cH4DEE3hJ+YmlFEm8VF
cNIKfySHpofywfBi8sJ2YWAjjrS52tESDgIpjfv/XQABHVxc58946wQOv9Zsw6/sY6HzAYD1EDZO
uGjBQjZTmyeeXk4wS7OMj6QOCkE/sIl3MnDUhM5iN0oPqN0VMPt3MhDAN2NVwGwb9hA1WkpsA40v
94cJTgV7LvbgX5Ym7fEnJMuaMdXHaUjiPFSHHLwKXfdw6n9snTQteMOAuZMlsdQ3mcktd5MHEG34
Eur+Wc8mPqx2bGpBLah2JzRp0AHqWhP0aB48e0D/xlZ7prFr7J0o+U2Q73+RRECsYIDnBrrcOJoB
Mrm7gpZGdmhY5TE0BMbMV7yJOa6meJLowCCA2PBUc+l2GqvcVRoDvJIfodJ6rOKmgnMU1cJz0RF3
9WrUugx3Cg5Q6B43wkGCmq8zvHd3daiFOH+VYYyr3N7kkQ97z/q4suFdioSetio8mv+0YY+amdJu
Fpc/KbNxUbjA8ySL1Ig78OFyAdPELAgdee2+h7XDJbcxXI0/NLL8twXAmtVkaEvtH1U5T5Y7RG9Q
UONM10RPkDJ4LhMxsTqn63D8olzDiVCnprYIXCDjExIM/6ruHKTRSeN6NVNSNWpaQL94qYVnjer3
NO+2aVzKGXLkcHajiDVUs7uRZ9LDE8Z43SGQGXv6tH21io4xg6g33EImRJKfO+CtpGzeMMZG8WaC
NCrzSjOKqRdmUjxs/ELUW4e2NaO8QvSpZzDxnjyMRrs6w9eEoRgGgkZde+rVuWEeqMxKzDrPz245
j+wmWvGRld6nGyvTCR77l6tfc8CTON87kW0wNrXcVxStjxImC+KSVIV/53Qh/tukpwEwLVccErVG
eQvoBobmv6PO2AfaWaT6cuLg2ibo5iRdZUbTT8dOnNkBl90dxDbClqG2SkK3GxFXa5/oIOnFKch3
1yM2X6bhKucjiGC1S4Xn99v3ZblUAn0ukoA0Kh/EckhCJcMvqyUxeKIp1QAY5ZnuM6R/u0xAtsWH
GkWJC/KwpyjDFsTn7S18UPz53R2sG7Hdc0tabxF+pfXOkJgwZMihyUeWj96MaaxTbpIKTgZF4jgp
omCm6Z8Zs1eaHSuRfB05wN4+JTLRjCui+qc+aJQWkLIVxcH0u8oq7XuzMyhZFoCYQJUxv8YxcJYo
/kaYYaeUsyfu1jXyhSR3E+y9LQj5RziTmSPhkpGKHhVYq4Wo6iNXF9YOQR/49lTABIhS0+dMF5/w
PlB8emjdcMI8r84ZTaO6OmrGWll65W512zyroXV82Lr6thyWN24Q47knkdZ9Vh+2iuZ5KfkOLcGb
8+KHN01CltaW/bPAXEemtQp1A7RVWsJWeqVXD37CgunV6Rc6R37mlJpENyK8RuV6ZtQfBC/r9IF1
ESpSVIxp0pfXbb+2F6nr4cqb+X9D0i3m/E34XBNrJ6lIZnTFtcnvGi4oq0jI5O+aluVFJMvvHjNy
zwgb4PL7iY+TbwcAawjcwjIdyvK8xLypZFp0GEiTWbobLlu9xNzW5ua9V6eUfmzdQac3ZzJHNu4B
Nqu6q9TlYx1gziRyy1EWO81sbFdSe3eVAF4PfjLjjdpk7pyQfwgESzi4VxMJx06KymWEaRIFlhac
S81OnYhTTJn7PfsARGmS0tjIxKxMyi/B+YvKNf5Q94zpFiFzJslanWK5LdbYAZFokSxEHaz6AaKf
urTiZ7+IE6zGCK5ziQ72LVjfS5mZtevrr+9uRYJlxcQ6dmdTcceOYKV+lqE0dvEXtFLR+l04P9nI
0d0jhd120TQsdHiCzwgHuztEfLK+kysLuazY9d269RLA5jlZlKsBDBGCY0ROnhhXK9yaGFhtwHWX
DIActyk8zvpjzT7GpAsx8rdagQs2CEvP2upejfUQuKxCs6dwX866D53BN6v0cEibDxeTswdiH9Go
UtbnMnTNfNLbggNTXzUgzYly/IOynZdZQfQqjaTPjM1+UhspGQXL+estGvrFsjC7HP+iFkMibAT8
9hVt5O621+H8onCEx9O8TQ4Hv/s6QEC+3MY8JsOK7nMWxrG0zAWz6CsdJKICgtj9oBcLJfz1bb7P
9RfjIvaJIfZPZHNWUgos/ekvhsPj1kzMleNdi0ttWXnMnzIs52htMkIzt560zmjW4/P+32qRbGfO
6LzPewVCFO2q7zHS5whgyBFaSVsQ47qonFU8jGf6PFfOluEJdPfq1l7OsSkPI8QgQuvpl8SQlLUe
b9UBZVzDY3DsTsZwHvIWlSZQ387X4MXdXiOEfkp+JnyctFXgntNhTrviogv53sPj7OX4gcJHKE4I
ZT36e8Yg9Nmg1KgplBKrDRqq9w+mnKPYIQVEK/+0P6RxFQyCx1IQICixq7PBorQtdRL8voHLut1P
1H5CodivN8zPV+5NyoZp6KGBse3/tfrkmI9qapK0xTf4lciGONSuE89MwX7wGi35wt862G3HmbOS
zk5+AK4VkVoBOz+o9vIN1FtGqTccAm3OtBgf6U2IE4CflhLIPkMXlcA3o6j0QfwC0V8VQbgvY0sF
UbWh57sb9NL2qFYKz4vwYUiOssnYVkj9svCyL95Siv7EGoXlQv8NvtMW09IP1SgHJNr+bxANDrel
XfXjSPiirESHYqqfuNdrKY6NL+fygZW7eGB0m2IvTa7/EFKUKAniUviqjWpiJDj45rb/ftnGw29s
AvKjvOtm3v3McunM8HHpMo7WL08MeI/XiiDVv920JBOID1Jv4hOrZN38etnagYijdJFqLgiT4nJm
Y+jsfQ091HCKcjnW1mUsc0/laJcYGXAywVaD8KOVuhI6p+JuipACoWqmspv/2OKcNaBJJDp2zkEo
Tl8c2ncY76cTrYJVfcKmkbtV+sb56aNTUVXASTcqgsEivW5ynwhOgurhSqru8OaLhCtthuqTkjLk
K/46wLeLSIhenIA2HJuhfvbHtDJC62Qpa23HOnaquCx7JoSbVyEeVvQ+/9u4zuuUCv9xuCbvnvXj
w6L0yQ6b3G+eIZdMgfqF0qWoRwETwiYEMuQkoYUbelMztFVqUgS4rfDWFY9DRxCbqRvTf6H0TIBH
X3QhPXheQinfv6Kg5e7K6cF9b1Qgq/YApe+0wbkComzMM1hjid2EkBagAyd7ffkUQUoX/MgjHK5A
+Rf/79GIBX0p7ffMjHonTZWKKv2PiDK/rXNVWB+yzxQIi0bLYOOU0uqPXI0Umste0egUa96W+OMJ
EDIUxnNHcJ3WzhEe6gm4DABgguLSmlLSygpG2cOvNgp5uswTb6sEMApY0uxC19h4L+2CkOPDUpyC
3rOCtJrirYanUN1AN2wssheWYDs43Ai/URLXLQN5PmDBib/0/yyCcEMLX4LzhJiAhx+E/OhXTIVm
aqzeIEzBk5WmPwM/jkfcEpSwK3oHr62zWUOtVhVc1ErgNnXKC6OvTT8CekredQ2bvqVcyCLkOVLA
edJmirLmkMBErye7JY6Zvxd+QocNW+jZI0j4RzkHuqaK3lBLsQ2Vh7A2Mv1O1RfTy7rq2scXLcZK
waSJ9y8feJ+TGtGPoZ1S+v8UTE+SaGSZFP9ca9UwNGfLgJ7BKnImbQm2Bhn7QclJxfw5DQ8henOg
So2n/2kK1S35uxfPpPAT3nw9lZi9rHLuli+cKxKvFeIzv6kYxlgzT6R2Ld5NtEdPfuhm3s6nqQhD
uG5mkqiQLHUX3bfI+IqzZ5t2u2WxYAEHirwc4JVLxC5J80w6ESnKrgoSttWNhzFBzKDkzo8n3+s8
UaZDwDISWZ/YqA7kvIXWDMKx+7uj/SKZk+f96Lz9+xa9eesWI7TvesbNfI8EeCYQ6L8CVmNrMmLR
jN0FVRWRebjfoozkG8QoeMkG+PY59pLXDwcxPcvzVe3eOD6z9tGwp583yzDTgFLJE93jzX4ZLxtE
l9FD4K1zAypizu6Dwg+twcaQ8P5JSxCVN+JNO7oh7fLETEB8twkkPy5HwaQ3LdFtC3IW01wHWx7l
m0VotwNihfHhZYKcX3GwLahs5ZYWgelz+mpBMtW+vskn99Zb/GjsTc3e3VmZo1u5GHfWIoq2Hyt4
UygNuZpmSbobfuBp6V0WwrznNUYJGEZ2gZoQOK5OiThso34K4o+vdwaZRAiHrHftgI9OSGQFqCiy
j0REN/1aW2ctuyu082knxf8Kmi14vt8FxxU8BaLqSuVpWpJZ+Fd6SlXT61c3GZ0MO/zejabQNPRg
cAPYSq2dJhPxDrEn93Jv2FcQH9XpPJPx1T0KanRvCJEyMmrOnBPx5+KHClorWy1YBMcAtQiJw+VN
+p53qqo+Fhq4Eoz0gY5vGqyCH+XSzMfTdyK130469AMrX107QqlkbLcwv8yXhdwnm1QCfgp5Chg5
BQDJLw4ZHtUME6ymF6/bDsf2eQTaIyrIUtlCO1hBM01Gfj7+eVxr/vDdU3rK4pbt0BaUZxeXLCjY
9YwPdRzlMWko8zz13cpJikLss6TMFqkE2sSBXMl1UzaYQiJs2vGZym46y+IXm+8wVEyT+sI42PJg
bUgJZu6t0vRM6E9ydP7uVdOANqIDF/tutDArlHmymMes3djFLpQ3lQNs3a345KbJrx/OGVGjvbKp
a4rnyUoDMgivD5lYRF8o6U4A4aTvSD8/Tna6u7Asv7RTZNZuTw4RyCzs7ulEcUtwwa7ZI0iBUpyi
T5ao22qD5GTqA/kpdMAjZmrS1SEi2yMrk0+CElK4KODUF+/p29RnUOEWEEQFApZRtawOqZET78zz
NxMUmm5TyOG93MHmpqMOgWSfIezD3Et0ID6QuIAVcbrw3QDiZbdKs8VYAD5tLTxsLFzZv6rSeBbb
7U7PvIqao3LtDBQHGfyU5tzCDGoXkPwuvCcHbxwEOu5i2D/MHtHqupo2VuuneLQllTi22HkhcSqX
7Gh8pxgpya3H1Byd0o5L0i0X7PwOfocU0dnDsT9qvkk81347Du4Q0UX7TgunuaC/MHV+th22bNDs
m+/mQJuxzyQMDtoE2b8JEFwPKB9iRGOvWipdJSWpCbuogzj0E3Sy8XtuaxtN8NHc1JuN3YXx+wFg
N9iw9qTFDoGUwVlMItPjZN5uEk6brtMmHTVntqXo7Y7RT0mtg1368ERYTeb0ZDVymKYqw1q9TJm2
0ag+zFB0tyr45a/7OqH3AwbCi8pulYwuC9/9tS+IJAjluSS6S9E5tmT9xzD4URSf4sV1xCTrKWSo
/O9xenE3RkvDN1W0W9sAKm37n1tGSIlcN2vgGCF727DssYXbuyQTS57bdjbE5JSQ6XYmH3TvwdkL
7g5XML0fp7YN5Xgo1kmZcRIo7C9sl4nwl2Id/iWbLrge6dtjJA/zYRAX1nqD1ys9u1g8FGySvlXM
XH7+8kHvJRNwg1710uZptxYLAd2L5xr1kDLXkPwsVSvCzetI8/EVKfdPkuTAaCVpcv2e8I5GhV7Z
u70MWbuqqWLGJmKyJxRkZWuKOvRtENamY7dRZ79v3sLBZItjXzUktgt8q4rYIMvTp338KoZ79KVP
F2trs/NVPQN7ErtpRAAdW6S685zJbH8HMkFJ1Np3839kcLn+TyFUWMK7heRVGC99GnPF+SnQrwG1
Qr9v9zTG6K1CElY2/e4F8e2OZxc1e7dbDhsu/teMnCEVA1rimyEfy0tchxlwd+4XhM4YVVnZmLnY
gId0i0NpcE5jqZQ7zljdjtLHxCmysnzPBn3eOFO+MQx38uxrkx56r8yEvSdqyeUCQH0sk46khMt2
odtHuz5TJ/eE4rkA8sQ/IhATRYMxgFdfTwVqnCfP6aRywtDQJr83ZJnBGR+bLGlhhD4Y9Um6VRHA
9Pew/O1P4hV6Hh7RRTOjrKmVwpo8VNT2uLWo4JjrZM9PAjscf+Un9aqs3fuXKCsm/2o4iUb/l+Sm
D96quyXzXvAIlamh++kU12uN/3p2XAYzUsfgITICd0umx+CJ1xb6olzjxHaaYbOgyryTG+jbuN9H
WoTzTYRGEjVuzcoCZIh5nHMeuXm3OlAIY+GN+Hyj+YHt19c3pb5I+KEiz2EOPTId/6dPj77On+ln
S9YCommLIBIzDVqubiUX+ttyqNVCwZKkRFvL7tspGfgewlnJUMbX6QcGKtLHU5DPTyVd+71w0q+b
jIO7i9QfJaRXWDD+ccaHuKUUdDv5JKo2bir/bzjAhHioIZuJqmAPA8h8LimqToL92GFQr/0ofHeE
+Eh3pMCuDaqE+HQ1gyyhjKite8euXe80djnwbku7Ok5XZq936BPZ4u1EZJH1Z7FF/HvZfIs2N+0y
57WkANmVtiYmPKnlUm1tCw1WUrDjgastzRZSjSppO9Rsblkug6uiAzj+TJanD577/pnAGDa+FIFj
clgCMfCJVx/ytaawh7NHRSx9dxH0PhteaJMoaxHzIKCw1N4FMTpe9sl6hvgj3x9px4fjAQb0XQD1
puZVM5WdSWh85yGStbbhRlxEjZyOaWOQG6+COmnFIPxKISVJcfwXPhf5TYCW8j/dZ/wpFWvT3/MW
5xP/Voy+R1ZGK5ezD/o2MonFsFiHba12ad54YM6KKZaNjad25qCnkKKC7hgxmN0L/vej9zHhx3BY
zio6+7QIFTP9Lr5EgT+vbUS5ajrDo71dYyExW5FnW9vFX2rNuUMg4YOHX9zE/X1jBSj190rC5q48
jTvHJEUT+1hm2YXZdauFNQlU/IyLP5KNHHYCXo6Sd+ZiIq1mw78iOvFy3xy3ppsf/ZW2PyAvnowA
U9A1/ndDqAq136dZ1SU++TArG3X5FRcSmKfMSnNTl38PEEsb0dn7wZ/ldsvjEw2m9Qqb6VpDehQP
OZMVBsnnPzTdrtFzzqVPBV/vSfLBT/dycFme6bu7LhAaaYM6nf3M5NJmp3mVnhXpLP1z0bI8FM9l
r1ZI9G6XkLMz2Q3Y4CbIG8sbSooocHS7nXCg9bwR+c728GsxlGUJaq4yDo/HnHZN1cbfQkkCT4U1
QVA31XsIi/4sUDSHgQei+wIXHX27IGanZclec6FP5G5ZnfejHljwu2Yv+7vcMyDZpl9tsTHIt/yX
rb1z+K6UzAY5YgaYw7HArxVgcs6QYX8dpZGfcisjeXIhSC/qpN5eC8DHFTWzVHfoD2Sv3hh0FXXV
6Pncw3wNhhodrGX05EqfZf0p8MAHJEF4G7j2JWnNlxIsJFd3leoq/akarsgYmZp8X+mWKPhO8L83
+3Lg+Qyw4gpLH/+XEEGzDrRQ/+ZTt8lvRE3Ba/0V2Vg9EilwEMHqbpDArXPeOKVffF42S7F5Ia9m
ZAc5aCkJhuCtlpxd7kLBLPpN0xDzscbUlmHpv8zywz4mLd1UyrgTRF78bvTc3aI5awZO+HqcrRjr
3Xoet4joEYM1hT0lk5rSUzdVHkiHB2jDmmiaFRazahtA7aVy9cUIuc22i9QMjlO46YU9BqpavUxX
z4Uub4sCGlMI+rhmQdUoDeo/8iqdicTnEZT0+Vr8mvHUutPkSnmL+7aKliwgGbTJluXxCZFi7gAV
zJTwe8nugeXPrNTZEL/pVBgSq2nXZYLx+pnJEPULzXtitTVgkmfurch6gPUaqkubUNDnGAGQwFX5
TwYRYUY3eqHtvg0Pqnuqr7ZGGhUTbSCmfL4IYNtd8VG6qLPY7/5IQRs7jR/MEjt0xpwSrBKer7iE
z7++jxmWMallVsisMkRyOgG53E7TKCZgFYVWG9l4phyAfE1ixR9eT5Ua4QpNRfvlBaDze2Tx5fPb
hDUDCdlgrpP83gDrS0gQCJHAodF9pIvuscfwzJoAp6zlaxGls8MTGTIqgReHnV2GaWJKBhnytPGy
M24a3ciuHdqzHUhrOsYzF4lFMD/Je+u17OcoE2KhyI2A8rIthkpfvDMOINifiXTVT0H2cQ37hjFG
LpIBq/T+kLGx9n/bZZpIsWKVqGUKo/QIMPmNjygzF7tZzRlAW/TLrYXiq0ompYZsWto6kfHNl2ZD
83At/P+dw0EgUIjbhmQCQis+iX/FaRX1+QOOqo6naCkd7GM+xFBurR9CRAAlewdhWd9CbEB0QZDl
PKGaHfnz7cy6jqcKJ08nopHauLggI7dmoKkwKELBwncXW0IUDi3wl+bua8TrCZKXMXAuaBAmEq5t
PO5e1uUE1psH5HywULRwzQqETrzHnEYVSgvjqB/NdKZhBGAfWP5QhH1qeoR/lgNod94c1DnEPhTO
mMKHnWBgk5tf3L4dMRQzXoCXiiGdAK4H7zgTxJKsDTp7/5oT1rjGHYGngaOkQo2Wq68hsE2pnFsS
fsO/fO7gV9Pec1EFAq5Qp3Nz6v1WW2tMuoECr1e8oxDeQcDpqzxKoxCeXbwYFXcyuePU4j7M//Fh
Syw/JkeovhhIesj7te7InlteKLBGCJnaKQrTxtZoFBUzteRXFKIKuzpyH/l2rr3oLXREaKQn6/Sj
nh4IpZwhnMUXsWtt9egUj2Sv1RtSrCaOUz4i7Oyj4QCpC14zYGStsST+e2eA5mpa96oHYmyV2Dpu
FPnFok/mTp35THnUtiPMq+QjvQL9TWvq6FCIGYLcEOwRassoxjAfShUklPynQxXRRugTUtQiGfRu
d/Fq/kdb9batxocPvloW1XDU4ItsHyB/tV1F43tJankey1xhzORNYZbfYpyy+fWvSxd63DBSCbHz
cS0qm/Wud6vcaABIcfjta64lwNzqrrzsi+h/9drwZOe6siJGFNflsdXaQR44n7m6JBQhbeL98oLF
VTLpZtzNcUj3eDRPtlyVAfPH5mL+ZqZmp7GL+NyJm2vhqPKF49iQgPuYiad6pLbQCp6hz78JAgh4
umNwhAF0EtTVm7MXWOywvlpBOsgfhgrqUEIqxILw4O0k8jI3PZWxhlaupMjV7L1K8jec22Zo7bPP
HCkEYv3hINzRsO8dAFAgbLrWLU3MTuDXR6DcAuAnIzwbBjwudnGQt3lEGkh/uUUoHMmcI41yxgZ8
4aKD/Tf7j+t/tfJnqGwXFSJXApooyq7mr2QpigcmthVUSBW2hhEQkMpKPn+elrb0mGLykCfdcpTd
ZNCb0sGSxzdissP7TK0G9jx6CMUc0aSi6vrza+auTkcLPdoVSiz0l3KmOcuLOOaBJwDsMnUMiDZt
WqKBRSWGbX9Q9hkYpYJkwR7qAmf4queDU4FtaFKZMlC1JGfF30kOtjQhIwi9umydWro1dhFi5qkn
ZDB2VZIvDvEJoD6TZp2c4jXxS2R4Y6QsL5z8FS5F5dl0tWaCSddSZTiafdN0UOrYVf5P9vdpNHSh
um0VoM6Rp5xU/m+i8IIwVyFc+OKLF34Y+81nAF6hW3VPRTgCNZVEDAEvVnf6euiJRnhP+VdCz+LI
6Ec7E2sqHUWKtKF3lPtKixYiBFRWyI321y/5rj3RXXqtnlwETg5iHHAVN7tOTMuzopvCus4wYurv
+gpKfY4nQqwrEjVBk/4WRct8t0aO3ytZF1jHyR+GgLUeRTlpOY2d17ow+lCMXeTowosAq/vNNN7Z
8oo8P+x4qm3C8hAJIAqXOvZrBHZSxnBiJeYKY3prQUMzWl4X7Uwhgby0ixDXXxRwxE0/mRq9F06+
053QT295NlUk3AQOcX9hNIC2g3t/W6TfMpwnMNHk0wl3/uh7YVaGm25ZhpgD58S20TAwR9vGJfq9
n0C3mAkYvyIDf4bpHp7sLZwRWi37hZYcwuwnPr6YCJNt6HO5I2RUDWLC0idyHMFzhTtelrdmMMCh
+gz7S/yUdfWRlJBUbUlb9ZvZfxivgNDh+xSHYIYBP9T5hrPHvf9rSr8p4YxD1YBxJWVdpnrQhtMJ
0W6L6xG0m5ijxcteUtT2kcoKdgelC/vfFui6n25y26whwYVbBJHO2mfU4fQ9WczrOCCngVHm0T9B
7Z4u39aWG/Qu30QWngXvB+bO1cpueclKRlGFKrHOlimiQyUHYAAHV5l9ffCW4H0aGRm+c3ENLUwt
uEpOvuD9qOAH1j0ctK6NM9iRzewzkLd9SArGeTViwiYYSElC3YrhpePfaLqojhb4FpR8WvAnHFwG
mq67zteIFGMqfjZVIvoL53WxyvmDwQvsia9+cqpA0FR8pYZbanOPKmrYCiBbHxhCatnXFwrUtlLN
Y7Fz2+6udDRNNS3/Vs130cmZUv5J56RsAVKKs5MI4VppsbogN0YFPnWsIenE4N0vpB2+PCQBCn4Y
Ke/JErJgEdoNkiyBpylhzAv96INzskKQ3irHGy/AZn4BAA0BX0cRquKZZZCOk6AQVdP3X96RYJt4
8YOFHdhDL50GxU3d9g9jrtpuC7z4Z1tPZ/eP1s9/jAZk2/RNBu3uU46DpkccNAjHGkmqoAwE3qqP
5NMb6AftOHU8N3azZZm2PATPg8HJYk1VEV342gcmTFc1wbbi+cuMh8LYkaZMA/x8PTC4fas3YJWy
NZ74OMevft7LKRsqrywnLGZwIZFdCPEXvVJzfmrQ0wHsXMUZ98hf4/NJyXOoXJZaXSdpAkLAGyvN
mxwC8eMBQfy4MfOPFzpfdPYZsh+vrwLG/UH0eYdZ3wceRNDETiRzryp1ndczg8EtbZKRJwVPXtLj
yTQ8GZdBtN4jw6CV6FZMnSy5kftHvVOUxtxeCwzpX9TLqvUHYIXX+Wp0VmbkX/7Y9RWyHQzSkkZ1
xa+FtUPgT9fcxgh53uoRReAZ11hH4zb/RXUz5EvamHFWeOfEk5MtMUH11MsIj3dJ2V+A5XlzAi6u
NDD4xud6OZ8tUtdDkWIqQ9NEbKQblo7VQmI4u+zqIqmjzbd8P6niqaNo7A/STnxal9UdJ4Ejd92k
DTRxm8EkdgGs6nINf/IAOKqGcesg2hnj05zPq5h/VoAuwNqa7ji9d3BQ3kjlIZBLXX3u6hYUYx7b
kWB/62Kppi++B5q3+aJBqfhm3u2UDmW+czYBbSbuDgyPKSrgTIbiRZIhlH4iOwcTrMwsGjB5UGZU
rpn+DU/yGf8muXjMJ3y6pcg+YLtlsNAPsE7nObHilytm0W/GSX8cVUtjbuTbJ25HVCVH1XxuOcpM
COKj2Kd9NtJ9hJ1R6XZW8NS9BUZXNTwHLTbzihn2eXHdNGAJ2G7zoOJHwZwdYpaqb52TYsyV+no2
pCYbQFhbW8bhRobLeqo/uXXMN0gBue+LKfKTCcFA+Gy/XKAu5YOuHc7lyUrPgJi8rFHGSvm7DEUN
hBv9gp0gW+H7yp4K8kJl9oNwCvkO/2JHVIPy+8SKnD84A6ofcv4EakJ/xtGEuVD9g/6PmDd6SB53
znyIUcL8yQkDY+Ax336g6Xxy3IjIO4YkXUnGhtgY4u7tZ6JYeVbh4+UnVJygfFGYjvme1KjTjHfI
2I6F/WtQA9amuh5lcad2r8+k58sr2dP9snFE7f/RPvETLzBk2eRbWjOS0mMk8yfdPUl8YxrQ9igi
b7bIwXZ75ZAq2hR+wuJZiJPZgUZHmfymArslU/s8hrWV+O2IwrFD2pzBWe4/RZvR4tkT6ufe/jBu
MP7IVe9PENA/MXHlZrYFxxT8yB5xcixYIE6LH8tqFN5TxIZ9rmVHotKiXPY5PuIaXrswQufPVZM+
NOF2yOeiNSOYrsY1OfRVYAlFG9fcstDZ4/s/z8k6PcyB7Ka08khVLHR4ql30XtC6ucyuDyqhwF/f
erR8YxdTmhMGNaAy5EkmgSudmPDXkTCvtwo3SFylvmU0S6HjuNdEwan1H7q73EjxfSLbeP3fsvEo
2zlFyvIBe9saHDRkIGMzBJywYCFxYMm11JDN8fgbG4w4fOm9kIOm2oP/pLyZ09YDdTPQzaGXtXVV
DOe6efsSfyL2KhwUBtg/9PfL68StG9K7PIpoKvOM+BG82PAKJvArDAvqXTl4D2i58T3ZwtWyW9dW
IcF+GS3nJSz1jXys8UIVqHxYj1Gqu/CkUMOpzJ+OmqLu/BZ0dVpyLBSp55dcdPMqGxfKRAAAhxM7
womSV8cQ9AaGJsZa9Oc7Ouko5Odn2449hgdgdMTcOszrpfx2HAsFd5XtjnMK6LPO3hfZftgCP1UO
F8d+fnqBOCKC1AelRKjNOEe2X6lz4ZSHAzzRy3FSfvH1KjD87tF1DwCyYM/6jm7Pjl8tx/fOfmTb
tUXy5Atl5yGc/1Id+owt1hefcN526sYarJCVZHIoaS5eYmGXA+m+Q+FwD1d8DYg31aSddN2y20Iv
cTinjXL1T0uHkshv9Sx8CJFoLqde15DSpaZFDvogzaOx6YEAeA25p7fcaQBcKRMDdIjwCF/l7o/i
iP3o0D31V6qm+EuKlVyJKKGdaqwwyuVpyp6tVlWQSeXTlf9bgceoDF2yF1edoOPrvCxXlaDbWuxb
pW8NVVobDBwn110llWA3ugc4pZD0PCoPIOY3EoW+q8V3Uxb+IEkiNAgiMWl3BVlDGc0SZVdA7Tpd
HQ0MtS0BPt3l8FLMqMr3GcJeh/olrcmgKnBY9+S39NGLp6Kfm085EWDQ3wG8xvoQyTLS0KsOwFqW
3BUYl51zj20vo27xP5FOZKwl9GOwLpxQvMzRtY1ewf0VEq8/lvgDdHpmTsAlRzz/woSdyjBSXoRA
sUCY+Ni/mVQrt2aFy5iTeNCemsUrC6qL7KsVHHIpsLabHa8HUlHvyZP3/EaNK1IJFDttLzS6eJwi
cOqNeQ448eI6HuK/GqSQVcSvjRXOEol1x9phqImK8LciApxpGw4LQRs2AVbTV7tse6vaaGA8lec9
D+1NMQXNLgyQ6KFxF4aOQ4bFbMcDtuCly0aBF4Xtgoj4kCZ92h6w9N9tkktOqq0pYRnt8ll0kikV
i83mMCVeLbbM7jkBvhpvTNyXQqKaehlVcS1qePJJxmAclkSjc07CDx54AM0RpWpPevrN2FfpGoK/
FyMTwZTMvkbhDYuIM9hOG9mMHu1BC0lh0uferJ+z532u8PUXFQRr3jUtCYqVqyT25hdscMq26hzv
htPD0BqNAmshbtfShoNI0VkVD9MdjefeJ+yj/VfH7NjzcMx8kDNewm/X1/Nt0yA0pgIIe0OtYRSW
39C50eW4yENSRLk0li+43/cKeCwa1DYS61J7RYLdeQphgQa9T7ymLP2G6Gb0/qIEeKSoip0F1Yfo
REwVZEfPFvMURlE2xp94JN+Eni1SjG8fV1WSvCNRCdGLYmxvMMndR8n/igVNzE1E2s2MAONmRk3j
j89tmPvExbRqa1R7D6ozsM3KzfppTrifrCQHnkztSECC9fjECtFNFinpUb1kEXTNo1VXSwaYzzpe
lhEflhtgopXbLkpfNEFJt/m+GjGDUTq4TSgEojHGnbVBL2JtIbm61vW1+cPgxNl1zYHxT/MNahu1
CGwo6dOQy/oux6cCzWPH2eRxmaXmB252A4BUX/KyMjeFefViWjiy+655pvComqlQa2Ik5ulZtWj7
CDBuFZWU056ZUVeRFrmcMl6rRzEVm528iMeTSai7Z7yCRDTeSjWI6PHWmYJxc2lcC4MFccLGhSFH
vOIwyaPjxcrmamfs+M/Tn90czpOvl2sLfoDJuvWrVNk97Da45hPSOO6XjaXVq+e//FbWXGwyZPkj
Mb+w14Wx1YMs+rFrcQm6BP1u/gerv58mMlZmDTy/EenZ41s2z+cy1c3W9jtasWBnJzvVEKwXPj/d
loNWJ5CM9MsgvC/TM882Sxix4DSFYKZl5PoTK3f8lbH+yB/TTolRS84DKVyajp85aXelqA0P4WI4
v1eDZUFtlhmQmTZ/WHlqEVqak1RBymizcKbdM59C9e3FFmte5Ez0WiBESrVi3dnYdMtliNcOpDlH
qQKpbKboiUGJhBBRCDxmClqJ2/CbgcqRJ1D8OTzZ7NXhPoKVlDds313i4YJ/tYvfb8pERxX9U6Ix
Zp1ClLMgJryahz5aiiy0sb3ew5pSqnKCwT/5x9gHtxpQZ9O1ldhIQZIr2g6gGfHCeRcdHIiFwXDc
F8UYAzpG845/6neBn9CymZZM7d3ZJ8neBv/1N/utNNjUeDN2SfIB2Ic6IXyF40TCep9uvGgKwJDm
I++7sYTf1vb/5vLpDKd+BYk2OgPaNhQKo8UXRXzcY2zHta+wQ/amHT+0H3m3/AJoYFh43V2EYNc0
LFRSyX1MdeyD1kCU2DffKsXB1Tml3TPuYnN2Oqx+cAjAIZvLeZSxPtemFVjaE7dqeZpJ4eYqYZ3i
sT5w7fhWGRSRlBz82oBgOrO2mWqoiJP412pYhzJhqsF9UHn4/31xfixvtComq0C6clRQ7/FLHFgR
+OvncEhAWvPzanvfvPQqovq6O9ftz5+XRugrsZVe/yGAh1zHqOfvQ4rwCIxOdgvyRpHjKVzw++Cw
ot2wH8k9tRdHw6SuhFTjS3+qjuRgGY5xR3p1uKn8mk4BCX0FkbxEUaXnGynFapE9eXcJI4k45439
V4uCdKoPOwYX2u1qWsMSYrzZlv3GTQo92JeNuB78BhGfB354MH5hGxdJ5Mal7W8FqoaGfLBUzw3W
8iGSXac1UJlbACzQwrQ5f0AbdM9N4o21zuYWq1DPOE759h01QY3H0uMOKusHKGm45JeLgh/BBR1I
wP38kFZ0X/NvgXW2gtUo8gFfPZ0LkFtqS9HjiKTubrevAbwGGQjEVfjB+81bIIZeCuwkUJRebn10
j8w0/DiW1gyCUqtC+hM/F0YaItHdyolXr+6s1QpOHd32XMEgGRwDQtyvaelM+48qthU6V1+uUL+U
9o46gxwZ6P41vuZsrkQbdqh1DAhGBMMjDEnSiUeSr4XKg7nsVqIsn7Dvdih1Fp/SAiRFuwnlvM00
qytr5mhzS3yZWpJdKfOfHZvk40J7aoxKIaEZpQhMLtRCDyE2KaVCf2OrL4CN5bXgW7DrKh5upEwg
4Om2sPkySgHozltSdVxdFDsFXQesUNoT4KRKVEg0MiibldUX5CSEiKNLNq1CVzEGFXDNhuLnZoYY
V83ymMRr2R5yzvlQN3n/y+yHGDQoA6gxGQDbi5+lgQnU1IcroUGItkxiNuv2Gp5mG6XHioKdiJJU
/yc+NPtapVScDXQBzT+lUm7/Fs08Tp83PmAwvZjm4B6tEamXDlmotcVMpcCfGujlXN7p0eJBuvyn
Dbqo2BkS1dGfWdWzwoibh+EbPKEcK5hKPqllDxKniNiQzt8ct/ocCHBEjvsBoT/OqobjaPau/J7L
urwH0kZ/q83V1XsGtJsdUcOwkfN/lkiwXR0171MQHlitm+T6RQ7AWoK8fzQeLRynAj1042P10n1J
ZO7mpZDCQWej4EqFXclHOfLx/uS4h6rmfIRH2FvWvdr/sZaNRpcFuUH8Tucg8lh6SyHWwdCte7Ii
YXk0T5bERdA6IKPZwLXgDkjndTohKcZckB/nprP9u6g8xYIygCYYsB/bBHrEcVSCKEhRF+t9IYHo
+wEgg9lijFGjwzwzHVjp6zlF3W4ZrPb0z9wPqKX2FbhhTOdrmpvd4VL2GmBMQwoF99NTRKjEdLc4
bxRqabjLf8Z+Xh5zZxFDB0i6mNKsAUXVT1+V+63GtpRn83bOS33XWMpZffXen/bG8C5xb4M31Vdv
Ymh9VpoY/WR64pqttdHg0n+U4UDSLAxlkw42m+471LuiG55YCk2OBMEil/wDwER2wdtEDLZAvkHa
G+l/UkaMg8dnouTSayvSzlLWtL6oWUlutFjdvAC+7f4Nt7LN02LlFQLRRnEDelqvNYIBH7ZSBfPf
hOShHbsCennLC4AI3X1gldxVYrpDlxIzi/hg48zOeLSTlg+ni9Y7cMjggPz3P3pl1Zqa2pOamtuR
l/vi4yA6kCLhA9hQ3ySOSm4E4FlMKVj5ZrYxIJ6FF6l23Qs4d8UkchdkKGreMgMPEWD1EF691gVB
+MVKNwcb+VfGM0KW
`pragma protect end_protected
