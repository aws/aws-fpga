// (c) Copyright 2023 Advanced Micro Devices, Inc. All rights reserved.
//
// This file contains confidential and proprietary information
// of AMD and is protected under U.S. and international copyright
// and other intellectual property laws.
//
// DISCLAIMER
// This disclaimer is not a license and does not grant any
// rights to the materials distributed herewith. Except as
// otherwise provided in a valid license issued to you by
// AMD, and to the maximum extent permitted by applicable
// law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
// WITH ALL FAULTS, AND AMD HEREBY DISCLAIMS ALL WARRANTIES
// AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
// BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
// INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
// (2) AMD shall not be liable (whether in contract or tort,
// including negligence, or under any other theory of
// liability) for any loss or damage of any kind or nature
// related to, arising under or in connection with these
// materials, including for any direct, or any indirect,
// special, incidental, or consequential loss or damage
// (including loss of data, profits, goodwill, or any type of
// loss or damage suffered as a result of any action brought
// by a third party) even if such damage or loss was
// reasonably foreseeable or AMD had been advised of the
// possibility of the same.
//
// CRITICAL APPLICATIONS
// AMD products are not designed or intended to be fail-
// safe, or for use in any application requiring fail-safe
// performance, such as life-support or safety devices or
// systems, Class III medical devices, nuclear facilities,
// applications related to the deployment of airbags, or any
// other applications that could lead to death, personal
// injury, or severe property or environmental damage
// (individually and collectively, "Critical
// Applications"). Customer assumes the sole risk and
// liability of any use of AMD products in Critical
// Applications, subject only to applicable laws and
// regulations governing limitations on product liability.
//
// THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
// PART OF THIS FILE AT ALL TIMES.
////////////////////////////////////////////////////////////
`timescale 1ps/1ps

module dir_detect(
 input MC_DQS_t,
 input MC_DQS_c,

 input Mem_DQS_t,
 input Mem_DQS_c,
 
 output wr_drive,
 output rd_drive );

 logic is_wr;
 logic is_rd;
 logic idle_state;

 always @(*) 
 begin
	if((MC_DQS_t === MC_DQS_c)  && (Mem_DQS_t === Mem_DQS_c))
	begin
		// idle state No one driving the DQ bus
		is_wr = 1'b0;
		is_rd = 1'b0;
		idle_state = 1'b1;
	end
	else if ((idle_state == 1'b1) && (MC_DQS_t !== MC_DQS_c) && (Mem_DQS_t === Mem_DQS_c))
	begin
		// DQS is driven from MC side => write_path.
		is_wr = 1'b1;
		is_rd = 1'b0;
		idle_state = 1'b0;
	end
	else if ((idle_state == 1'b1) && (MC_DQS_t === MC_DQS_c) && (Mem_DQS_t !== Mem_DQS_c))
	begin
		// DQS is driven from Mem side => read_path.
		is_wr = 1'b0;
		is_rd = 1'b1;
		idle_state = 1'b0;
	end
 end

 assign wr_drive = is_wr;
 assign rd_drive = is_rd;
endmodule
