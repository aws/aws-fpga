// Amazon FPGA Hardware Development Kit
//
// Copyright 2016 Amazon.com, Inc. or its affiliates. All Rights Reserved.
//
// Licensed under the Amazon Software License (the "License"). You may not use
// this file except in compliance with the License. A copy of the License is
// located at
//
//    http://aws.amazon.com/asl/
//
// or in the "license" file accompanying this file. This file is distributed on
// an "AS IS" BASIS, WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, express or
// implied. See the License for the specific language governing permissions and
// limitations under the License.

// SHA: f463fc25b8464dd6c1672ff28a603eec67bfcb40
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2016_05", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
WGl49kaxDgNkt4OFNMWNPEcSt2smeI862k4q1FRyKfWHCOhexDtbCMxxQk0MCUGapFpr6YS/2vpm
LpEO+OwItNaTovAdnKh2KkxWxVSXGbUvapkmldLb6mfnIotc95dCrRWc8jt2rKBrk+lvfDiAGWHz
zbtJEvINfSX1DpwU77DwR38LeX1+qSFhPjE1T5H1Y4rTnly9Kc1gP6Q/sQJOUxEEfhiHIOKuUKlI
R2A9dae7I+46g132QCoW094/bIzyM3AfPsO6cTy7HOZKok/BDL+UiCRNdNBnOigWmA07n3VvtmHs
HUYbvX2nmb2zW0xABljlpj4MaVZmNEsUtpnfYQ==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
NtSwoAPJik2TWyH6ABkJxVVZ4CgiMieyB7Q473CKmj0rY0QeG3MvnSZFexHBQJmBl+7JELTdS0lM
gaCGLAg6JtKJXAjfHjDJy6ED/9RZmh4beerLq2DvMaNFmFT2kBITL5oYk/buVVvUNr8VSPzub8VI
H6rHKdxOki6zr9Kto5E=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
FNxRaFczabsV6xctNaPwi22whoxhUm4wDoL3B9QB8OPvqUQ6OvKodfNnDyPcawgdqaxUxa4VgNsC
JDIYQ5GRLCwh+jn5M9743RxtFmXmZ1ZWXobfuH6PZ9II/2G61Ntm7sHwUrdbNF+sF9cJJJvV1jjF
Fkc1PKacxAdIO4/zRXw=

`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
EFYHv+o8HrcnxSbNONNUW/7kswWa6BVXERAPwK2Ghn05ljkbi6YENaYE24t2QJYTWq/PtZw1cCIv
bZkW0dD7Aw==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5824)
`pragma protect data_block
0xF7BsekOgGyQch76n7vq1X8vUrPZrL5+WqOT6b/TY3O4ldMTchXOpyeZgZ9URK+GoML7evIQBE3
KBQHCzFLuiKCtPIj2AZ01yAVZFWRmrtrUn5enYyIaMIuVD2ieMWsUcLXcCIhmoUbWnFt/Et50X3j
V7lT3LGvD0pkacjHFNhHFC+sbB2vpPT4Ph31QmlgnU/7/TmqPQGlgWoYMsBC1SdQxKs0FIjiolD3
nr4A/UImKypDyGx7KhgvzdJy3U15A/fMmR4foiFAndl4KCf13FRQoAC/3sxeoggdEIFL13VbRxaD
zuISNrHXKiwMl9Y0L1+LEHYeaR0HYpp4NMs68FVPwdf+uXzYqZz7zcigs3Ywp4H9q1yAo75Ic1Zz
w70GWANOFZJ0MJneB0pDpOxwuYzQmVaKc9mIBN8FcBS+BwCfd92pNiZoQjJJG3oyz+Y2qHoWmikL
6YmErJMyhQkdWI6onosieAn3N7A+hShTUtmk7Bw70cdNJenICdr87NQFNqyF2xL+xlyRePm4qmIp
yQgVgRI9Ktq06n7sj4nrqmvD2l0+JfwDmKMLJe6eBCgiFHiNfPadVB6b2dfcXxAnZSzi9NzKllm/
l+37F93oihK1gNmRQUX/PohkSaKs3IIppaQ7DRkyKqfizVB+V+zfMcydN46WdV+I4qymLu0o15D9
Pewe5CIkldlSeTOg7qR6eBcB94u4d0zYKnbhyDFurhOZeDo4Pq6f7eS1HjsSdgSc3OQeOQFbm0yi
0RH/HCy+0iyKv3H+K3wR78wWI+AT1uTFRMqYvrztqzyeYSTIVDeFwZPo9z1kI4WomBfh6DU2Gk9g
94+3pys4ihyXUbh0FN7ZOfkc5IzfJk/Sqr18eufQeEL41uHBkXqTjnaCWI/IwrZeQFOvlE3m/kiR
g3uC3Lh4zb/ke4zq76Xqjp9EzBLYlmIPnGRZzzuVYkjJFhPrYQVFWEkwUy/8Z84vUohDqQlnbZO5
dVKF3//mINNYOy86UHNJlyzdE1CKRKaj3xuQu0MdlX8SQ+VfYDExoq/m1BuNXW6XMe+iORhQbsC2
9cNLdntNa+M50nOZ01p8pnoJ4EZztdYtOOmBXKI8wEIZZqBvmoRQqV79370q75VEwcajJH+zRzdn
ew+tHkGzIU10JG/vAnIoH1goBlcnoNoCOlj9ye+lBhHGQaNhYcPbuQdKpoVercloRX8gmdHahgCI
8/Rh9C+JsJs3siRlbZwy6Q85+9ROUf/kute6U2qGMS74lDodS8iPwB/daOjV4rhnVKPBpUNDfhot
XfDAr7mCz5LM3pDbJGFZnQf7Uuq8XVisy3cqCmyNQ00tSRFSXCDxAc/rlRa/oGaRiZj3e+/pgzZj
9RrTFGPsCsIr0ugcw1cPGm7ADb/joi+bFJUssD4DNVYbWLt0hwZe6SUz177yJ5sxTpZ3kWEzKQRY
a0ZL7Kd+zhsob6Db6fKP/mCbfs/BaoLK1C3n0a+98UpDw9poc0shVzovrAV+jADNbpIQVbWlb6qw
MGZU9syTRSnfOgi9JA15AX38K35vh/RFPAj76J7uojwxarODIntJXPTY4payYNHXcj9tsujTPUfx
wixPLTFW+xb2Uh1oWJwobfsPcxbdkuHlLgbNUZYzs5TUzWssDbskuOSDgCRR65CNqng7u1gHPrs9
JGHSY/6YIrkjnCE05OZQS5pyYlbNCr6B5t5w/4/UW9Ob4KQDgGwRQsuW6IlKjkn+9nnEUFmyN+dw
OCngqkDsBT2XstOyepwaaZ4qY83B5kb5u04MwkT+H3DqAPTPtVVti61kHV4tju7q/aH/o83CwZy0
6fFoM1+U9juAaNxanC5LnWHoMTe/IY7mEY60+7nb9KrCT/R8MYGVL+aowk0taZGOy0hMyhQttdyg
aQWrXGN/jsUHKjK7VFau3Wblggr7IXdoEIpBjECT4Tb8+TPH6Cb2wGS1kOkTrp//UcTHjOpoUpuZ
Gop/aUUGnpQVDTXksjhm9NR3l8B8UI7jfsaZ5yq8cZiWkaxaZlyUWMexLIK0D822K50vOx+LJTGk
f40cC61c+aO8g9fzd4Y1rrj2RN8rz66ODhvr2Casu7gJ47f8IlIBgU9SNJAGAvRuZSdFllnLQ9lm
aThg2FRj0oyA3rOGH2WOqdJoMEOgj6Ozi9iWr/OCJoubHhbH95+V08nSYLtDgXpz/FqNUMAxrLZx
teYGWCF2JfCQzvRZItgaf3EKn4a5fWK4HKqcay7KDC8S3YGoTvJTpHMLd+XiJSomNUFjsKo1kFXZ
48Y5ktAWPOlAro8kUhTElq3dTW+QuukVF/PXOFGLDZY0ThKO/43t3jTatoHcM97iBvlYbjT5j4Gk
l9a5MkrC0g/u1lRO1jc0hHymjF5ENHEhosV0kJ0FHI1OY7SHTVir9kzuft3SJ46tlEGAXOS0TNjV
TGTWrYMRIvOLxhAwb5dWnZmQ6eDoKZIYg3/tytZteCgvoCfiW5cD9AXstjq4Xy3f/9NKe2LNXh+f
X8UPD0kdoJFf6hyopbTTjF5xhAdYsLCI7KGFGxSk3OmzvbAvNfLUk2ufghwKy83CASGJFYTOrJdS
DyNtDRXTlOnmvCwbTeFcqS/lIb2yKkc5XVknInvnoPXmwnTu/3yeYOnkjrhyFZvQECySCIBxv5eb
wwXuHFFOIkyCjvysvH9yBIxgZpBNzOxYYW9LwksSfmbCCN0ImZIuYNl9PJYWGzI4pAwuBt0JW7ej
6PJOBgmHSzGgLJjoehlI7pEPpZbasF3iY8gIxqbHSn9hspyLSXJu7HwctTkmrvmUCdnTx8xUbzHn
dAl9pYH9H8wxXDGCp8SqLjee5m3Iw8nrS4QeEl/XWpxV7hoOyfC/G5t93+1I22zpewdgWk4R7I9t
DHiyqgPEcFGKV04M7a6lHsamCpZwCuW1mLZGUiUWi4VenO1HdGU23FQH0p0Yr/S4TyHwfIt/fuZF
bFH6e1MQQa0PLQOnnIUv72tAKBesCJ4Q3zJIEfkzOzywGxbl0Tmdthc0cu/FzNbgY55IUkxOPYQe
UwuYDIFNN3cnG6crauLHBNdvQKVZTC8h8qXU/LgMUhMbhMoDiLLBTCHrFLxAtTlLe0BLqrLZld3D
rzg/deQ+4iMs2zuEHYKb4GCYyMxu2EVV4cy0lq2bNE/qBdMBxH6kwWY6y29bfgB2L4hLaZa3DRwD
WXHkvc1SObNeDH2KIKGKTqOQHUex77+ropSvGGTkDKaVg50RsIxFfrxTVovSdDXwjxxSIwBULyow
ljULdgfkFQbPOd4QfDjunPoC6AHlHDuoL2a5P5Lbx4pGG450/5kM79efuK/YTkNzNupZJliSmDj6
k24zXJWw/exPqj5a8U7J3Tc4VNbXz076xWDjxnSbTq+UyfNNd3DHBFE4qFgMYK/MsZW6NnDDKnR8
mhivKSLdL1fN7MH0U3hNt20hHRQW2xWSKdFjaDdQKjm2SsyJMIM/E3k3v9AeAS8aTgP5s9GPULRM
gW6U6FurRr/hjO0YjSiUIWFXsrwwYbz4RO0s/580NZnH2LKkGYUhyNjxT8Jd+3KzVhMtOfFpj1iK
mWEYZAHRDBZJkObHUk3gTv8XKkxwqnNT3SevopdqdnH1U1ZOQ1nz+sPJ0rwdsc6D4008PeW+ayk7
Ogip/ZrXIAhRgutEU1YGTgTUc9Loa8NemjZNa+nVV5KH/HfxL3DGmQjJAL/5bM1tYo3dv7rtH2Uk
XtldkJAvyKXGqHXMIT0cHHZDQOFNwI1iiOu1GuE+jvmZFYc8tiDH1f/HY6eCx/XEEri88nEs2VhX
LxBV/tyQkRiXkatnTSs23DsmLOTB+Fz50aGXGdlWTgwfgiR2BL5G9Y/qip4BhhTO5bg63ghziqP4
fvwZPdRrj8orPPjFj04jTnSqQTnkZUBMd1ZJvmI82P0FFCGstI/4ISC1tqQ/oy1j0TBRCOp00Csw
OjwzmuI8UNp3S7G/Sc1N8ojr3Xhcxmq+s8XfwwZRvzOf6ND8Bvy8PONdHiEvyYahKEwz0AvdVmKO
VvD095WR7Bo53XkdRNNr7rhoLGvgYq0wmLHtXMJO4mCpwZRRFr/veBHQJgyKN9af/ulZ3cjL++EP
fSxN9hxiuHKluyLi5XMVF3qTMdM7GoNDw+BuZcNotfKHijymw7GhRVaMv/OXf+gHmcnVRxwy93Rh
NP7PqaYpTcpdHJV2j8oa8i+fHP8mgj/dmJfD10wNj6+ftntHuPekpoAZ+VLZe+TEqslN0P6isn+G
gprO47oQh0aqfHw+wNejFInlSa/GLElPwbWTHTqdCpApQOUlxfIBVlySLnQGtDyLas1JRjLfpmeA
Dxm/KqVApjyO53dZt+Q785AY0G0DubkYUiHZcReQ6Xrkk2uWrpAZ0v4Sy+x9vIkrAeJDrzJVuQSz
nqCh0dJP3dzeQU6Cqug4jrTOMqjmnH55AK51TNk9GJ49IonvTM+jmAekGhl1q4SLWtLC3NVtIuom
R+roY2n9J6O8AmOs+0p8Z3nE9qNqPU8C4bWHqRiyPuse2CbkRZ7vcWtMeVM2sHIISFDYTBWJOWRO
7yG0+pS3HUE8Ubd2TpRwQ0p1LQT6iE2ya4W7GmsSx6OFRLSHMhF7OiyWfO+UGF2dWtKKeeOKcR5c
6tiyhi/d1rJU/SadsdguTsEFALhGncNhZa90b2lRxIG1APeFcOgZGlaCyDtBeSfGtLOsXcgQ+G2U
rk1p3SnSqJH21LSCu8x4Q1J+0Xdtc7BMql/RJUpl9bTqx++pkUPcPiE7kOztncWGay6MF62yGxGu
nedSGbGoe3LauzchOlI9bultjCb5nrDil+0VVnZB81tIQSr/YQjME3MXLW42dRudIIVbbEvH1YWN
LGtNFo/qIcCNbOHltEunorshJDUE3yPDkqGQx7hSl4zRykbGkbTrkDCBA32j98sTTboiT7Sp/gy+
D4pX9bXw0dSZQskUuouI5bZ0Fw+CtyFGKPiaFNq7/k0TbhK0aDBy70jKEst+Jr57MyfDN4fzxBsH
vQF1AVYcgG/kAGrc4aVIv3UcpsFk9vD5Feohj9L5ZYN5q2QDpiUANFlEW+iWGWQ+Uk0zjY3pzNei
M9QCsNNF4Wc1bR3RVJM7iflstPYk0gO906qBz4xK84FWjEYFpsXV42VaNaprkLVVuBfW4ZMSrFoJ
ZcJZclgIfYpsaap17/fDteUmF9S8Y1Vxke8IY+8WVQnQLJJPA1ltZRveinlmSsBK1mHyRZltpqgN
f7ubTbnGYgpvB7OaC1h264ZZ3jzu9apiBFJGseAbiz5DoiasMKUd0fp1FJKUXa1Drbcu8aSzbjfU
63610K5JN3fXUvTDLUCM9k55bjaEHUJP39GSbNFXZPOnXMebroNrOPEGMPgtTvB60/bOCMkuy3tR
slhoQLSRwGeoWwdTXDgsm6acgH8nLAyIG8JLS2tc4+onVL5RNspwE7X5uGuCDFnqJt8vI8Ybure4
NYDQIBIkI7742k+U2b6CL3+bRVXQ0yN4txtY9dMMKqhJLMSekcFORH5Q4fWIjA+2Pq/rpU7OjS0R
qIOGl8++Otq+O7dvwK8uEhLuAOIVqrh8Q8QTtEIsLVjveAIam3HTngPfQck+/DrJv5rTNyqjPYKp
tYX6scxNNkQJ5FHumttrk13awdIOalCF3gbx/luDQCwRqwe4rChPUVvrdBoIoEjqchRmbLm8lRt5
xZBq8b1/q3ajK6f7giBMfw5p/brs0yXxsGvw6lq+UpTteL0gy3lnF/GpF1KntWto5LqNfSqVNOlD
5awy1itMdXlPympnx+5z1bE5sk9wLgnXSn3n+mV05wP4Y0gI08K5XK47QUC9gj0zCEJzZPgHPNio
msAt/Kr+rgY76gWDp6juqYRYEXbHrlWHTIcD2UNEq0c+CvliYLrGhFKzp/XxvuUsPKvX3+0kaJ+9
He+agClrVdjyN3hCaXkouwMRup1P2bKqXcFEbPk9NbqAJQ1rifUDLRfOTr4zLcUwn7e2Y42doVS8
60WRrohCLc9hBIusacJcfasp4kFd4ZEURYan9LHLYj/+r6pMSCJ2UhhsD17xrCkUn70zeBk7pZ7v
pJtnabsJsTGcF8LcAtLvCKW6l3HFLUaxTuY3McmOonhJEZwJNiCWfwHBsu52m9AxsIWwdthi+d56
vi5gE5ie0ilF01IThV/GTKOWK6MtOyeCr2S0xMtaOdeLjJCvtANFJ0erwYfEhfuyOVjgh7zERdmO
F1qXvDNcjK4Jh0IvTYI9QlEvbunbwfVxfbLANK6+UbkBvjruathxrhLwSyerH1BJtHlLNT5DAM25
U7jvlinMLv5mFWf7a516emJV9uS0RlpMlr8jzYSWpLwJyTc6culwiA76rVgh8WIdOPIroRHISVOm
T65MKzZLduaT+RT5cHpl+xejW7vPE/gw8U8kstFkiB99qKfSGYUBl01GHddUmS8LEW0CiDVZwEpY
2eAu7J8bye+VAaoDK/DT4kjdTpRSQVlqhRsGmY8KfjdGasEyCnr0dRfqLqV3ThD01NsOU9T80sue
83O3ce6UcZvvu9JRIbisJEIuS5L+m5vCUlOJTK5YnGyVWEVFQmGIh5h697ImQnSD0dP0ULW3cTgZ
g9872eNpRbfJuNbtaiddPtR6RN0o0fGISp199mWOBH/yr415i41q8u++k5LbE0fdr5kmBpfCmA6A
+PsfCnHazcZJWZFPYvj/0QYQsrtop/GL6t7PMOZwGZbTSl7fe408awyJ3pMOvXU9O0pzdVJ6rbsB
LlPS+wbEHKW8TYX87mXuPQmh9dLQcLMiPImcXEwHJhoMJ9sLUsQmq/ox0e2MsIDiBQtwWu/v5Tje
lOv25D5isIfatwKArwLbSPAxZGNgGuco7+7Q3CP6wVBVvdpTx8FDvalgKgrM7fHRaYDZwQvWhNcg
5++YEl7wXUrCq1d9lhLThad3GiGO8p1Am6WwbC2KJYLbZlqi3jnzBojsi1MvAcQJd8kdm86j/5BG
SaShYtP6GNvrXxP0Kx9OxyPhhvLkxALjowHCB408dj9OLoJfXkuAJ2N6Qhf+uqJpDjEfnYN+0ycP
jqPrUIjHcFlml77YAW8Zsb9uadKVTSxJpXu7uig8A7A9rmIAZX6GHAadl711YmlrFhqjkUqnICRg
r9NxMbrAbCQOTbxsrodttEvQC8E9TmIxHnUQlJpU3BQGgM5zIF53ker3V1hE9MXqtoi28Wcje2mG
rM06geWcPLZyIf1GjFH6wyRiZNI/kj31ukMkF/EWjsn7y7Ui1JKNqAgZH+LlR6MZDp371sjPYS7P
Y81mWoueKQi01pgppVOMty4YMrCU7c87lh+8RWtQX9oj2r5IKdSaw9QdNFN0Y2IjC88ybRv9f4Ur
GEo6d2lVDw7FevhR7VlyjdjZUfM1qHgrewayDukh58CqG4/bG/RrHqx19Mrk1y+Pwp2RBDQcE9ne
kYAvjL/1IGkCL9gNZ6amaQ1T1XROL6QmmaB6CVFhwBIFJzLub2lfpCkz7wzHOnyUrs0KXWeFRoul
Q+3AH9mnVA7JNqRQk0hlENk98avI4M84IVuIC3HpYt3Lt94YrbVH9gEudbPiHLQdM40RNrWzbHeq
uOWaYtk3oAaCWWdHAXWGlGCT8xP4+s/FUdXXHX3qNlWDuZFvWprHeO3R0OdVSuRApauxb4c6xSXT
d2cAFY9Qa0idHyAetUYCZqnEOfvmKYGrZfNKcFEJiJNghCbTK1aWus6g82y0XzfBJzkhQfYY70oX
GonrIHvR41fw+w==
`pragma protect end_protected
