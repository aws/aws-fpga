`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
cdZKdDFlAHQ2xnKQ1kC+QNPPDthSJJXO30g8GOiv8GMLH5x2hFjlS/D0ULXoJDg4N2LNRLgeVY/V
h7QEizdaczfnvH3niSp1bGSOCs5mfeQ2lnCSNk18Kts2Zq8nAhffZY/TBvldIEVNzr4hx0SU1ovF
gviOH4LWHUMEAW0SUxqINqjD++heBQ/RZ36QdTMiT5SrJsk1jmU4df0C3IWxIH4sxnFPwa857OAK
GqV2jrIzeFiaqDuJ25kkbOkOytKHIfAITXflqmflaqMiTIW4vum1F6j4SuEqki14tv/AhCEB5C1w
8W4WH61WxGenFwpaVkX10eD1Ox8+Hqlq//HtJQ==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
BFBRCn+tsKw5bSopq2sUlJBnveulK5xCFsriIMXYZkb8z9wo74Y5mvAbj3EZi78Q7uby2sWmjGjU
DmPOz7FfyuyKYOjvNezfj/A+CKqK5sHqXYTtaDOHxDkKQ+bIK+rEngAKr6Z7tidNacjzBrm7WAzX
UYkL6sTGOYDVDFOjS2c=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
XxX6W2a3x4LXHfaDG53BarGw6ZfgSKx12CDEixWPsoJAcflo7MYNIFa61oTyzznsZ5ZjQv6N9psw
5A64oGYSurW7B1L+gZuPpn0o9PhvmsKmRtx+bK+xIJ3WOk+zFB2tsgcsaNZ+kea3aeTlUSUAgVRD
H4X7AG2MJP40Gd4RiWg=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2720)
`pragma protect data_block
znpEoZ8mJOMkOCnh8ikZlN5icByzhcMD6IqkmXES7Dcfb+KrQB0CxB5ZvMHHjweBs2zxnTKeC3bG
qpWYzf7plyw/bz3cj+PP9Vw0Zm289jaJw+N0rC8FMWt/C05L27Izrnt+sMtaQA9c2I0DHe0D+730
Z/5KOmPE8TbV5xhB9Z9omSk4Ar7lavrXBAYgihtubelsP8OCCK2aMBqyPhuv8rwN7q71ae7ZkPoH
GpLnUFeCa2EQeoGYdAdZx6S+Zy7MO7MWOScMW1RsyguwTfdRddq4tXWqj8dUXZ/XAMHERQSgJUIm
6QrwIbRAr8TL04doyfkMM/5P7ArF1ZzNR3PQuiD6Fe3Sm+hxB/LDqGxtgSC8imcIGPw7TkSNSwR6
TPw3IhdxwnSHsYiiBnDX1BvP8KU050bXA/2ziebDyvul4ZUXTwUJcqIzCUDaE+0FF7KBVfHyyz2t
aPIPpvW2vsM6z1iN0/dXD1FIm9XUYxKclvvzazbds3Cb5GVGG7sAiQDgz5/0CBqWeMKADLOmiOR+
QdsFa5IyQ0arENPl8y7BNghHIPurkhk5aEYN58HgFOJa5rulfNuxHU1p+oQBmRyT6wOgcxtFiMZC
nfUidfCKlnCwf80xqyu/q9AcQLyamr9kqW8izkq/BEkInXIoYv/vTi9OBZz1ci+pYfPshIe3dxRh
OWf4b/poqWQI1tKJz+RGNoE4qa9MCLqn5kzDuYd3rwEQoDXjapjhQqEdAfWMoCjCO0vDW/th6KuV
sRPE1u+qy/iuYGhli5mWQq8NFYjZvNnBuuqieIK3y8kCwnABCeS5BcIzEkPGz4xdlIdGTnGqdXzx
iWcnnbDhZ0DS+OC55lEGZsliPc4S82N5HVWuu/syla0AQMYx9kcTVx3K8tvcQinWtl7J6EK1sEBk
4XOJj7+lWFlDFkaCpjz5ePuQVIFUt3yoB0qmm8mBznP0VXV0bn7Yd8GmcPyVFA9Gbo02a0/pufUj
rHkRfCNc0tshTqBhdEniFWg0l2DCXrrFttDVJDZQabG7a97RvIGJEYEdOPsvFVirgE7hnXEm3Pdo
Al4fgrRKlR670OAd+3RTU+rN8d9c7s4+kFwIEPFTFljZ6yYws1TYX4r1sfY/8HNfFyBLhuoIiFwo
Q7exQHrYi+aZ7CKB5dAbMk+za14twanhG5EshO/gixLTJgCvAg4WMMF9PhYozYc1ok1Lw4vc3wP5
fGgO1jP4AHH7/QxtLI412z26vsChERBNXeFGZzoknKyIfEHqwByvFczV/SQUswONCU4jJG76oabU
etVasxtxVMkH0QtRWjF6z50zRyz7wzdvm8RHZUEAWJyGFqTw++ufs2ZEuKZYuzNoQhgZRljHj1/m
2/FUk/G39dQENZfTC1f2FBszqa6vNiGYfQVXybZ9yy944F3pwfKTKsiYiEHCneOgau4+E3pdvHJY
Gj19w2MIhqAsBmL6Ar4q1IOUwglZ1GzX97kAQLrAoQcwzihHM3UbsrktP8FOdKW1YapxZBVfgrIU
hBsJzjBsSK4WA3KZJJP9zwbDjXUDh050jmvQMgbdVnUkn242RNma3cxSyzVoMhMCHSLL7WaqPigC
Pi1njeToZi/Oq0g6RmCQQnu0DQ44KN0XNIQ2fFszablre2WHo9JsqFnWCtyR0ZgStikDH0QhtLqK
2oqSWgL5LD9sQPZo39ipyHP0FhQf2+4rWVgD9qCYVktNcSXzU9ZgmYRiGDcni/bx+p/vUiqs5kW7
dHcyw68PVTIprY7C2xI/cvADUwKf6VDQle/VZl1clxosKgVzAuwN8bDWtxZ/Kv+cOvzlYsb4xuiM
lu16HTrSPbcV7aYmiLv3TSq5Hf2uUX5blQ7ZsYUudCeYaP0i90nFc00m3/ExkJrmz5xiQuwyeM9W
qncRMRm6w6X4Pq7ThNNlLRlh5k19LECLr5UlWKA66oUibbyLMIB97k5l7E3XrfXUYVVF5Veox2me
SkGN+f2VEFmOuLfd/0XLhDHPqRWUkEsOMbFK+44KdGMqIEkZ6Nsi3Gdrf5asb8vLg9bpM6iD5GOi
e5kQpeGc3Zv9J1q2+pOFJK5emKxRr2EEToQUJyKMv4kPOB/UJllThZk7A4o4i2JmsZZr6qIu094B
yZG7ZaB30RqTrrn/jDvPmahPgjVUe3GrJHdZ0UrKk88/+SWXheU0oS9toyJknAYv0s3Qw2a3TWgN
ozH7/pZTqVNETmcBwZX0oUUoc2JO3/NscMgTs3K1mzGdVH8oTOHj/fcDIWbZhjGuQYIgQXRshNIU
I3uTUVk0KCKS/ewzzblOAmin1FJ+e5d7+/YRct+uIcRhvxIe83Vy498cSZfJlH8uS+4ocdd3scjw
xMrcnj+mZljA5rF8AjH6rnhIWlokIqM3gAWDogn1nWhLbcjE+sj9ulEej9+9mSHO2WFulRq4E4Pj
vMkuovTir5Q0ifAlakCNLoElq9BaI2RmC4+8/ZwkoL+0CU8XcxYslTAPuKC7gqiAwbGcjjK4Haft
5jKk2ofvflYCm9s/VFNPwqMZTP8ZBn2GihB9Z7IFnc3qAUG1TyUXX2AMiTcAWJR7tqX7JDmwnGrm
Oq/Mamwp5JCdb94vcmTWDSiijBDK0Dsuba8+eQySPrDLISxiuS2Y7ICu5EasrNnwFgUfbseJACyQ
Y763/rLHa28PIj5bCcDNPRfwSBDHQEwHMMQFp/XNuyWvfoSgh9SXMuaOzzG63ivKep2+K2bahTma
N90oPLMEuCiCXYzbffeTJV7VmD8PctPky9sly0WkcxQqM8iDrtKU/F8hWgxjgujTGq92EW3QiGEQ
2UbsdcveI5jfHpJOz8g4WnIDA6CA7yrCMS74SbMd+4z26hOe2D7yrkX4yO6PlSysjZQSw69DZjK+
RhBotZ0lTkq64kqgok068zZuE2aB+OpOIpE5J8mkmLaof5d2g/1E2RaJABmenAKY+rXUGHDkV7DR
1pJenb93fZez2tUJh2ar0TqGkELHfpy9ui7F/4NGyRRa+bMlO3Z+w0pZ0nE0dp4zZ6hjjH0oEEgs
em3Q0SDm8PVlC7qzTv50yI2RIhJ5ROq7loJQ5DYg/oeBmgiKrpxrwwC5SNOUxK7v50s1Kcqe9l11
qYpz3wK22TVIiv4SyMxYq2Q9xZiOFimOfdrficr9711AVOI3JlT9bJuty6h92L372NUefDPIvPlI
75z7Ebu/A0s/3ZPHe0ik+Vdo+JYSR8KFwrWTiUqnI59dqFhRzW5nSGszEjx1CorKCeRjCZb+Q7fD
kkG4+FIDYrVRFYUXFeNi97hPtakY8pKR27xpYlh+PC43WRlCR90KfpYHfXep/3vtUQ21PnxgmMQ/
0JZsaDTeThQIm9N3ylJUmodby9KD0JoRFn8VZ9BOC5Qv2LK3t5bTh8kLtZLhrTdqU9r6zScGfVm2
XzTjrTMMcgFw4YHuBeCjHaS39ESwgPwKCIWOSg+SbC2O18SvRrIyTUR3akXvrQ4TGUwUz8ajKbbM
2VlTPQ6BuBf9UVm4TGOMUWrB7TBqAkeoz6qnSpTaQ2SxCdcTIqNTf6Sa3BYWNQu0Doadq+18rfk7
syOPEpDOEuIURQkCdaK2PUdjC39HCKScoE4+WrutFo1AqW3U5U4s9ns=
`pragma protect end_protected
