// =============================================================================
// Copyright 2016 Amazon.com, Inc. or its affiliates.
// All Rights Reserved Worldwide.
// Amazon Confidential information
// Restricted NDA Material
// =============================================================================

 `define HMC_WRAPPER_PATH tb.TOP.CL.HMC_WRAPPER
 `define SH_PATH tb.TOP.SH
 `define CL_PATH tb.TOP.CL

  `define VENOM_CL
