// Amazon FPGA Hardware Development Kit
//
// Copyright 2016 Amazon.com, Inc. or its affiliates. All Rights Reserved.
//
// Licensed under the Amazon Software License (the "License"). You may not use
// this file except in compliance with the License. A copy of the License is
// located at
//
//    http://aws.amazon.com/asl/
//
// or in the "license" file accompanying this file. This file is distributed on
// an "AS IS" BASIS, WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, express or
// implied. See the License for the specific language governing permissions and
// limitations under the License.

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
j4deEXB1unuMV67pG+eByfxC+XiTdK6k7PVyZqPyZqK6acS0TvCkznD0OfH+j44uUz+pAjIZO68p
RicM2mkK8iKbep2IgOOySnRZ8WhTwYjMKLHlLupeQyM0dpHs6iw7y+7FGHducaj/E/POxAmnIPD9
XdIWOnqEpDL/BWCGqB38TaKllZxsFhB4zBM3MgHBXWD1PZ/nSJYKF97aa8CfNvM4MOIxkOJLnUfs
Cm4dODKjDazPHrcg1yWuPv8AHDXx/OLT/u9n87gZybdqYRkyiKpnEAbvkh/ugTdtd0DPUEc8EIWn
wRB/mp0mLtXP0af3XlHX36zZg7ycrINt/y/WJA==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
vxYeEGkzJyfN4+hABIdZixYwX00PYdtXtUm3uNzGPD+KD79vZO0Ujt8RwF3EgBx211yXNShu7DO4
tAwCf1I01ZmF40uFQIXQDiEDbTaDm/Gc0WmqJWdOMGOiXz9BV803ez7fsSXhRKV7uWMnowCauoQT
hZbYsRtIDNFlfm0BIHs=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
DQgWrj4d0aZ69TSIX7BE4p67WrosiKIGYGOIklCIcYDalEscTco/sFb8NUtzVYvn0PGU5Pd0B1ni
9rQUu+UMzO6MtZB8zj2gLPQB1UTXrFgjiFCCv4dFIXilOG3eHCMPbKSzZXU2DxmTARbiQE683hsX
hNy5hDkj25othAApHPQ=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5760)
`pragma protect data_block
8McTlzhdmq5+45QvryH5NETd8bwcJi3sLZdrWZ/ecVDt1jUgABYNsReKWmtTfmtfvxOHLmsvcS01
lZfnfxiOMdWgcV4i+Y/0YmorFzgixEC3Cyxw8sNeC79aLdc+j/Log1yMN2rgEM0zUVVMqRLCTc4W
AoXEm9K8g6kF7f73QdVRA9b4jmpjY1AETaV6DhkXa94eFqithNcWg0Ko1TD/+K9VtlODMGAYoPdA
uE3aKdSF5Z50CbCgvdZBnh3t0iK2QKskvAvWTv4jDRXP6fyr1GCK8SkNE50IENymGDL1DJWKThPM
LGDzX4EV3ALMI1JyMt+Epv0ymOn+rooAG9r47A352SS2I8rqdG8moW558JNIWx70xYP3qPZSNwQi
gPavh+RFym6sc3NBPX6IimrxOwcE2zvkpFSBHoYq0Z3nhpbhRq4QgXNGsVnNWJItsz6xHK6rhKB/
+usKJx6QtyRK2W3p7ApQVXzsv/8ptscB2nmwf1dI6lV8oBALHo+uCOsIpkFnfcBd2uEfRHeaHiKK
u0QAjeIMhvyBqkW7XFeyKooxrT9vcBrHH6qlc82bkf5+ssahNImezqfHi9Hw99Bu172Ao18VVKTr
aeKJq5JhhGs07m0etHnVQIVvlJAhGYD8K1ulrEylI7oCAoKn6APjPndClzURxpehR202pZgavq1q
iNVvZjo17hsujiYVOMGYBKLYm1zJMGOokIbUAqmr7uxkWQh0gigEiu3UCcWGA99CvYOYGg3lFpnR
IKrqBYZzaDkiNJ3ycouHbYj++noC+oLnCV4sieMzHKaoe50W1zEURVJpYdxt66b6jWRJS2ms6lol
/Z+nxaXgakVREMCgrLyER/+uvvHvlLoir/gaAYNmApsCodEwLTGbiZvNZt3JzrJt35olBILEXyqZ
gl+t+KzGaSNDSjQnxItOjfuPBhtl0/phyfLRzrlg+ExmezIB5hN3LjGtcjiMNKbE3RD5t7juynD1
TtzHqilqa9pXFSQmhnvctW6axL2B2+EAgyTxlyHbBH5+dKLh/BRmoZBz/lH4xSkTjHXDNkTvVDDZ
xbXgy5KB1p6buk2ZcqBLoOC6Hy4SEJOyjHCeQrHeUyHMl/9pQO8qnj62IJ2DOCWf23PvXWeoArXc
0vHJhSVM9GEcxQMvrLr3+MziQNN2UP2owMKf1XfM8LJ2Nmmvx+Ra7JzOpTxQCUxABzfNAa8HrUm3
TLQaXjIit1YJ2/v8Nuqd+ah7y6X3yPqlKM4KgCgn8kEYu/+4/rtu1JBSoymykQrsCp8hjLfVc8ll
I6dJpXKl9LaXJXRZOsFYRMVudsQCi7Q252wq9TSkS2j6Jv2CP1rtuAmjhToV9BMGGnxk+Ic7OxMA
yBva2FjfeVxh+ukT8D0PKoViHA/ZsWPj/RnV+AchictrHUlHNwCnSxX2RLsmZPVkJFBYngQLShDv
yL5HAImJEZCuZ2O8EU/Z6vD70HTgdTM+NdrX5qIBs9g3QP5wkeMzFe24wcS90ilB7uuQC9wUaOuS
r+JsDkSIu43T0Eer9iAZIil8Eux0uFCRZbnR9IFeBAo72luyeMxfCAcWwGblsC9taiFXOyxquwkw
ZeTUTkC0OLj017BKySDgJ+7lbvGZSRJTl7i9jkU7pnknmeVR+OoxedTC/AridrRRrLM9jVFHU31o
4tdq2E+pksB5d46Q8MLaUUVBwWzaH8nhGSDsOAWEIGVGbZxfU2fLx6f81VEz9gT/w6z5l5whAVXm
aG4kijBqDdBFP67YBVlz6MStqjkdY2YmTsA8gTHsCyzj6rJ7VK1Q86EoYCQOopElDVGMsrCwYVIw
0oBo6gHKJx/ZpFI+jqFRXcUIocKRp7dSqVuZDQlqDNWD0820QnBAVo5k5kwezUVADcwuj/MXSZDN
E/K4TNR51NxoCIlPY1QkEOFiNDWoavJ5pvidPIgypbFeWLi8KkdRUAMSajhlebD46HOFreUKR6cg
WRR4kU6Ya9xNcqapLQ6tlhOkJtEwtsmkm8/sTza+qUnToO0w9L9IEtZBtKgpxr2sknchsl/h+CTk
Wqi63Wp+56h4S57y3ZqD/zBYKIGOXH2Z7vJwH3cAvOcA/Z5SBldtAR8TZWpuzke4quKJbUupXm+b
6us6MYY++sKj+NLh+HEv3x4x6rmnHDcYngxJTKifqq/H55KTWx4OADSBSOz6fjMhBKum2n6u49b8
bHt6V+vxHj3rO8y+h0ifztA+mLykIuGflLRN76GQPzajg7SbPprf2k7tlmrUZGgY8HhRZF2IU7WB
qVEqK05Iw+71YmC+ShbJnd20fT7u0ITj2Z1X4KSH5OAVoZtxvMF56XWX5wNviWK8wwWk+eHuZ/FM
xwHVfuVB/SSVDh35HQ3yEGwe/iyLDUMDzQm1Pu+Mc6iWb/Dg9ISNQbJcT1eSm9QOQAVpowBxKSZJ
lHorGP/rNRE0QW+zCpH5vmvZxqItkk1PDkHgr4BpG/vmVV8lqLIG72GpQ22stQUw66Mx6rmEO4aM
A2IVThaZdZ8Q/qeS6aLSiehUtn/dQsAjoS17u04n+GguW34gtnfvtd6pe2Gja15Wps6cmUiILjxD
1/7mZslTg++gXdxm4If87it3pkA250tX2WG85QSWjCpnPkcvTugqidvVYFhH866kihtN1DiawwWi
L2m3cWBovpjHCOVpN9wdOIrUn4W0jQVX6y1xwKagOyH+ZadJaE86pc6jpiTpaIqjGzYNgbyR3i82
dP3gIMmVN3SA/+S6UZfTYWhKVGI4xRP1K4ugi3ZrawUy7/kEJQvsyZiU+ov107zPLdaxWaD6H5iT
uAftHxaNrict+JYRI2wC2IHCKOSgQfXQerIAx0KM+zpxC4W52FD9AELIkHzNFX4mWr+EEYGu/Sdt
Ara69r6Tz1KAowetDiTA9LtCEih/ZcIQg86HgzbCaxxUpw1N/o4uFW4LsHRDmZkiH5TOokZ5J6zT
G5r/h8fqbaQNxWjMH8HcbDVYWpLmygkSymrpZhgToD+KaY1w4LuaKe5C8j40qepsAvkZDjUN9wUn
Upb5gU0wX8MgdBn5liqZnmWzYRrkfiuLPVczRyDvQSp4Enz89Vwr1n6krGcAVGEXjxS/znyPgelj
YXz8apf4PF7xdwsirMnFxmVDmSGLHCK0Y+9Vxnu3XdC/ZSyfEVpq5Kr0CJU7LqhcIs3bLHaETqMB
SYDzvNJZd1X8CFslISKG6lXcO/ynm3cAvf7Fbk9Fbo/fzLoC/OeEBzdxpFqo0yJLVEpBtJ7EGsgL
vEfL9RSK2D+ox67AEPAKh+HBd9H1iHAL/iYyli1i/m+E6Cw7gp/GOqTomSjsqRBqZKn2gf4m9lQr
ai+DAiZtFZbdI+WIefYNrIA7xdf/ScIZNRIG98K+Y04od7FM3dYCAsv1VxYSBBrmZGD+6T7HO/7G
xVJu6Ve6BR+iWrRPo6Km0x5N+mD/j6Co3gBMzOGtRvVQ17ulLgEhsodr4dkYkcQFjkVrAbGAqqFv
5GhecuFMWH3jboCDUISIXhIjsDoXQ3m8yLnV8ARVmtbpmIBsEXnAyQ45IK5qRWm81jo+9rX1XQ5/
nrQu8pLNfh1qDtGqTpk6KGzDpNTVYV2S1JUjO4H614aq8ZGvoUPPAdKrIVN7gVCl/I6z9kOrgv9/
/2O74nlcuH2Heap+9+9jcu9PLU0a6S5IKmHuN2djKfaupcDlZl3rzpwl6+FhG02zAA0G0Ebsya4V
7vFbDDrgj1sA6xQ5dus/70fUzFSmipXQL/rsaUjYqTRI+Pe4cQdbO9NWEJ9iSJOqK8C7+nk3sq5t
ZrIv+c9iLPxMAzPfcIvB9FlTUzNvuQ1bIB5ZdAJfKDC8ED4wEh9nnZtoZbSWR/S7KcyZPZSkdBTU
rd4riAC7rXePob0J8WZarKcFRTHrERfOXls1lqaFrtKlTDCo7RUsnglLycvUZ3nO/PEYkFVVH68r
KuyTuefHA/hv3Wso2JnDa028TA1XjtKmqA/v00KmXbBGvagYcswr6tn9sA1sE++qZZhzMgZKE3fa
gBNTvpzHMpvv8wV9s9bt7kNabFtKS83+EjCR9Zwa6IB6waTqHe/nP00HM10htSdsQSYWcAFYUi92
iZsrFwHmLz7TTMKvVGH1FRuD65SLCOKHXKvles89hcf7M5w5AgzeqChv1lULR1rZ5Vlx82g+Q+wh
jq1q7kSv7VTUyP2LSTDywddM++7NEaRpjodNqzT4AGIrfezgRZrkPb+w+chOwh/4zZUyn7aJGmws
babyzomwOETe1C90pA9CFmgzGb4YH49P+WTcptTQ3+s1CFXu9cu5ZdOMnHAHbZUvisC20WdZev2W
SIHdNHItBrvTHblIyhqJYHofwc9S+mYMaWFIrS6gKR6Fy/RivJBHsYet1zOdUW7Y/D1ADMk9w60u
lyuQ7Wiac39XHfy9ZnKBMboIga9NFN82GHr1Yx7V5F/YKTp2Yn3HgrHjY0GGty+ww8qA9xCNNIs9
I0D3PFZJYInIAd9qBS58WRrzxWGvIXJkTMGZq05Qsyx5hMCg94H9QdflAjRHIXsg42pbBeClniNU
98x/1849axVnjzQ2S0Qnhldcf4YBR7EQHpE9qu0/iQvOR/70UYS3nibsQuwvIG+vYVvkIpxqdUea
0iiJAbd65E1CdD1HN9iQgQ0IZ8ztTXt44p524GiKwGwQxRR2eVTODQdiZa4Rfgk5tAjv9Y80FRQ1
goFxi7gXgwZ5bTaoudMuwS9VwR0hHEhI7Paet3Q8uhW6H490rlgKqkRnXjc+1Xqu5EkHaSplyhg2
h3zb+JLDZPDYLspRkM4dt7mG+s1Xfx+81ZkHf5y1vOn2NJ/KSTuzf2G4vzArh4B3LOdo7WbBa1mf
j7eCrA9cxS41xoLbiSUn/BgPqlGIFUTFLqoWOh2Tt2S096HZSGfy+QUm03vevrQczV5fI8y803Zb
Uzt4e2s+gLfnZebsgGklxqQZdIMdStq31oI8r7pKpiuy/3dE4+jJgj+4KZ5p9z7X63yoGJGqCR1s
vCAD7uHBfRMSTMRfYfiF5iDGjFhxtIx0+Ma5goSyQn+uMbM/+fnRsOWAgiHh48g/qKQ9fnnDQMQD
knT8u8NWSE7sGHaLZ8BBdnp7k9MSslpfyxPRgBGYHp872SxTKuWeQzHeoMucFvAXqpn1wZI2eFfZ
1XssAdYEtJQxbAat6Je/F+AfE+JAWksr8v0/JYYT1RNi46dD22wS3Q1Rnpp4HG4US+ZIbsIxqLzr
rNhJTIRvquDg0SeUjbjGg87kdEs6VnsEqpXT5mFfeLwfGpuqMnDJ1Xx/36U+wtaHF6LVSAeo0Yew
1SpoMHkk8ZWHXSSvG/x2XuLL9rftCIntBtIoGT1KjEpPRl2UtqJrtj4B+YtTAyDZpx7uT0qL1Evh
UiEKmSmepNJfeHuBMX3FxrpwNPFcqZoyLm0nvVIzvrXJNffJknt5beoJxMmNRx3RqXvVI39QM8uj
v+t7P8AGqh7PBPrvPqoNkAEf/xcn5Tgga2djcrTzdX78JsjuYCoWvNEY6VSwHFb+dpFTCNh4+9qQ
xop3eZpxz/AIPNWW1wqwspEMY/DAkU1jHchMbgw6gkykMUrGtABKnVByEhnOQzsLYYli0kOoZGNg
iMAegAAYdkfqZKY6+TRza0idZR/o2+5+JnJV1Fvd6O22xqWdojIGBLgm7w+phGz2ELqr1ADonMB6
Yt2C2ANZc8Uwr5Z90mhWx3lC7p/4F15FJqcDWd5SPv6Fc8GpsJqF7bfJzBsWuL5Is/wcy7J07wUE
jVpXWav0tO6Gspiwxwkei2tK5Ji1dvPjlWyWsMvagyyruKwydaa2zDJUkqrwxU2zR4vuE9rCOsaD
L5uhLLqZwj/nbaGq7cZHm+9VA1+9/zKSPsthzjogWCG4A7yaQKiS6IXS6vx206cxyjja1RrcCajt
LvevcvR06G5nCQ5nr9gDMx672mvaTKuxBBI6mLKMYiR4hOgdpy90B7NH5seCnncm2tYA7hAt92/i
NDF2RuY3z2YEFJMEF9dGeU3U31CzCA0gtzYBksRmmMsSLgRMo1EShHgtFg3pxufW/KheHfUzBMGv
agWfMDvb5azddxuIYBHzqIH4d+erJuRMqIkGJPEKm7lYo6Yo3tB412b4OghfEICFlVUT/OuIMbXf
fLNZa0yMhDaorJwZL+ltnPvtv8HlJ4L3Tix6tJiur6rMgjkPfvGzxjVQ47dN2jN2w0ae8BXjGMiw
gsgmLysQ0BoPyEWX0hlEV7IWfkCLhhPZyBPZM9833g9agkEeuiT1QxxqzoGmw5mYuerjhddz94Dj
xNOTVIGsR05mls7ckZvZdKJegUX0CS+ivhyDRTi+rCRncwDf7Qc9SJrVJeRxbwC8sJ4y6SOHVtvG
k7T6H4OPVUCTmFsFa2/X03wx8NMSXWpR7urXNFQTSeOJVYL6P2npika0G7BjcsCxxa2dv+k8fEzF
VF5UTXDQsHGSC3LtkAJOF2+8gIM3fQDxJVvX+RjHnW3/s5G023jal5B9ePYMS6sF5RDJbzV3ZTVu
KS+ZnE1iJiSx/TNFA3SrrihDYXxo55BuPuBT6T3EuHGW/Z/fDO/z04QG3rbx0z/+NdOWbSjHe2MJ
qigTWt45m0zwFaxRXJs+Qyy3pUnuuI+o0CBYKR0rVsZ6XIPWcm3zbPW85F1qek1Fnwp3x2IH9qyZ
APQQh8wTW5fKcala6J8ceWJ/RE0V9XwDRQ8Ag7GmXM85edWQw1bUC3fLlhk+EgGVkhHTHueYtw9j
VXO8RlqjVPZ3PlpaJgkibzj9Mrs7ruRwcLNlfRjn/DUv8gRfcruhpzDILRfvgRf9qpm38KrjoQTX
gAcgNwasQ9PmpJgUfHSl2+v3E3iusBAg8xzn/zZDwombdug5vjEZwkncmF+SO8xmc44y23O5h7sy
YEUJ63K9VAt4hrn4+R/N05lxIK3tjih+j97H3z2bPyXG4+/OPSf/eFC4tzCdq4zUcHhUNSrbUBbR
b8ALW5MlR6PuGuO3RHqEgcwuLTMxtD2U3ivlWMCbsCJSLpnw8TLh+pYPg9ahvxTf6E+0K6aZrAXa
W0XetQ5zmnc4DwreQ8kOQ4tCyCKVc1vERJfVebiL+mAKqnFt9JJNI2ry2ljnK77c3e/vYFfZcm1U
R06INk+W1ISjgBxZT2QQFAHoxyrgKWZI/vFQ/H4hx8/gcj19aMFw0jTIxsOOxvgEFr6wIOP6of1r
tm/WbQ99o7kOzJboNzkshb3kJ5JEymWWycyuyEhZa0ufW0g+as3Om4rR2oOq/xeRmgyrFPt7qyLi
DfooaCq8qRvK8z1puk4Jg+35t/3wiNxGSzaiViODOBo5hKD1kPzEZMPBr738jiREvjFfGuKoJeIK
BDxt8z/Jwi/m52UIg0p58bda0b8gxEBM//e+P5tLOi7aVGeTixLtwNvpdUG/8F4R+nwTKerYrBq+
7OeLrpi3WBpJn1o10xFwZwebTC/N4MoOulIXJbnykHB+ASf5Z4FPgppcwjF+ioUFGH7fE4ZjhnQT
lgBvKyiSI2uK6maKxcvQQNReIOcrYGsp3GYeESg0dDHThN59jJk0R4NtwQsBoW2JE2UbsTun4Z0A
XOYpXa2zfixbpZe1BKFqDbEygHvRFcCX8gIac+JTESk7nyVuOgIyoq6XwCvKifqdmzm9IfpOr3Pk
TYoL
`pragma protect end_protected
