`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
j0kD3nIUA+BXdwLRcBuUgK5scbmf6OQtrslQRRqsySceVUw4iFgSTaaom5wfb5aF10sMOEpsIlBx
Ntb3HhOIkvCUfxm57w0iQrJ0TXh7DYlE80I2SP4gkEkpe2jqm2JIsWzkSzRWmoTrqlusRBCyKKS3
iCMLvzZSyK+boxGE9bPJ0QNPYGSAhsSJTCFz7R6wv/Q8po+rFRC9n8DFB16se8zk3tbQt35Teg68
NfJfzhtleA0IcTYbTGfFRryy8obUjLVC2yxknvRFMXb3hQeir+zYn7HmeFs7Js05RV22SOhu7GvV
TcfojsplnXfIIQIDfYR052SuRH243rprq3M0Yg==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
k8cPnuhDeTlEBuTsgqhkF0wWXgDRI/PbT7soOzx4lJvrEx5gJGoJfmTMI/xQChmsIE60Iz4GLPuU
G/aWlkOJ2MbnptFQCBz+wRGjMKjqpA51DpiDS+VN/Mvj1MWQkn6UGMijtPon3MAnY8UpXG6FrRzw
whujcDXA7wR6aw2zDsA=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
DKccdOBjHwXgn7H4r3OTl+qWc3FghpCo6cQhglSZo9I2l+03vhlDOSC8UHYS0osl2eaxjZ16fpsC
5OQgmaWLT7cVxFFtox+gblKAy4/cXlPqG7RMSrROtRE7+rWykMfTdpvRLMiobmTg4jyDUG2nrRqN
ZCYWwBLPwVhyy/1TJG0=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 13120)
`pragma protect data_block
dwWNStEw5X+A8GObHWTtztJcO942waVTuQIwi4UBlZs0P63mZ0sEX7mN/pCwW+L8hpAMql3DZIwI
Yw9w6QxVCiuqKqGY0sLw3eMxvqNpboio6QnuGBRReYURpv60WG+2Gv+rveOJFHHHdDbjPwMfiT3A
yOIVqS2DLpV53yw+emmQgIqoF1gdWzvxLdOW0ey23itU+LWzjI18lA7LGlWJ4NKKV/R3IMk8XNgc
PbreBwJvEcHnJzCNe95PuYRy0xFTy91/oMQtL7/7UmWNt4GssOIJTJIdbIG+Gdpt7XWhXtn3mJag
wJKDQm2TW9Ftyr3vFSvqmNwxQ/b7vW4JDKT/nrzMJpDYszvt63GHrPai/Bz18GyhwuvJO8peeQke
gEMQ/WAAcPdN0LkumVIGO2Cf7lk24TOqoHOJRLnULxoky/bt+5Fr2bBHy2Y3/7XTIkUyOyRV6ipj
Ze4I0uXyC5hJvkaCc4tjF1KjG9ixNyspjQ6cRgRPfcJJd24dYVzqtIlWhEi8ZqF6vWhKOsjrYHYB
0GVe44bPT2jkndVb7ytcTZmO9ScY93T9RUIrkVmEkQTq5IjGLs0+oeMdRfIPhjRii2MQfVUuFG5m
qo/UkYZTCypb9UPWz7Ay8YvpMcPn/R6HmsCQG2T2nLYZgox4nUinS650T9K+HX7uTNY0mHOZ+KC5
c0iL3vrh3FcGhxufjDk77QPRwDNdDOrtBLMwh8a60DZfpEvYxunE1ve2zq1Hofe/ed3/1cujZdv9
wzD5vc7OlCGqQK/wgaRgB9mPyfSNUngRlnTeh1Gtp/7FSVivKlqMMDJOVPlZwITdNlMKD81ZkYGO
Pna2yzoZsNi5O5RD2iQlv3s9UVv6yMLbvdZtHfkRW3M/GCAoCTlrvJ+1uiFRwo3yk8+TCyRd4Jqk
chKczTkQaCyHMR9zeY5NWkAFe7skDhXzxm77w4Q0ZGWfd4z4aqVraDpLyER/IYfW0mcD+y2wkPTs
inhbOZYGHJdY+D4g5KtrlDE54bFTSvFHFgjony5mS6Nr6KrwCe9opTI+z3WLRUEqdXzWmrXD5udW
G86ARyZtX0ZjKDHCmzQkwWpbbXR/eyF+3Rf2XsvH+ksnaF8u6ts6mTdBAfCb6KN+n+/bWw/dEji2
Yo1FpT6dMuC+V3IhggZAiSqRCRwcXecmdCeGITeZJP/IrmzorfC9dbPR9WUmLBYeo1XBubx+7Wjc
3D225JEEa9VcJH5UaMOJG8EOlZ9LRxzyDIvU4b62FQg0+tP2kgIBWrAI/hCNSqgVnO2OHe3lV6Lj
W2SW+d52N35JT1Zi2tdlzTHwWijfrpAttO1Z+xdloMrHu6+MQlH0Z/hBgnxhuCpMmIOqqLq+lCVN
4ms/eDjQaSRLL+tNHHq3rcFBl0dqmvfaDeMWr/TXEF+Fkvl74zxUjq+ZEbgCELyaf7CmT+xZ9Zls
OiqZ7+2Co+FQ2HHB+6lArfk2GR6VR0/do/e1JsByt4NJiwgre/fObwqW4uhrTs9FhJAO0iLd0a3V
+pPG2Dyz7JSAYPNfgCJNX3EVKw/g+VNI/EG1SOpFFxRE90z4j6yLkiofGsopdLfS4clQD0iEhh5M
x3BjQVNVb7RJtB8KaBpfOIo8ZzYI9lEFmWGpL17sjvE7bT42/ArvqwoYDl/ydrcW4AyKC5QxToe0
OVFgrCyKbHIC+1f0679y+jwKB+QU0C9rf6539oVgjKJRiPJhRx1Bvc5X7kxum6aseFaeSQGDNH9/
FI/cj+CGmFaLAGj9fqAdbZlZCT85Elo7ypVsBwr38e/hN8QIfV98e5znKli/wRpOEqIjyAcCPrfF
ysejjjXBQH/dn7q1ME81jnFu47/nLIlJ0e7VSFsaftZ+z4LYlvywnEQag9yjOLM8Z1HJ+bsP6agH
+glZ/J7oovkRvDmtPJ92KKAs6iJGKeEoJ/+9wb5ZGiQallF28n4nGO35/2AR8/ChpIGiIxDtC0/i
QewZWu1wu1FClmXGQgh3YjYtNTxxHei27tJSu9XUg7x4U48IWGMWLSe2b77osQgb4Izt6Ui4v4oC
HupSRkGAq0aXcMU7NJ3YTgGErtVRDKjSK4BAaIDIWmd6Nb9CYi56hnZUsKoCLl/W09ErdclCC7nA
NBK2JeEXihfPgfjWwJkSvXwbOW65WKjEzMKG+n9oj3sAeHa38XzMDXEwAqaaWJPgYc0lBkQbIlOO
y+RE7Yqi3pUBuznweWAchkrwsUtT2gxR02Ou9qqnt5L1/E/wrF9k3SZJU38o1wfN/VL9pjE+9/sS
lsilqVfank+7GXFTnwc/+v+Op7ueNPl3CaaZTo6duk646CgGKYn2Ah5Xj9XPKAV/kSmsIN6n/DAs
+7hRRfzSJRlwYYCaDNXB2L03boRKWc2HPFc16ONuTUYQXBqvIloErd5GKGZew387ZtOVdKwZbM0p
gLOx19RiW30Wd4H94ssCxdmUTtdBW949PIrHPq2+2PfDkexRIvy80E6z0AUVVjNrSsUBxrVpY0Sc
98Js5xUye1YXLOgOoxWmhjfOj6dt07WxuVHUPOtV9jelQ4J7D9dhGwbZ7+IzRYTNQ8Txug6czpSF
1kvbBu4K+UPlhQuBhztiHZGucAceHtr4zPee6qIYlX3FDPLqg9Ei7l79tmaYHeU8qZ873HZv2kZq
tpO7T5x3FXVNpL0FR+L2Vmrj+aKfcks5L3v/2ythSpybVmZeajv+bacz5huR0Vjk6OjAvaoKNgBW
2tNmR+wCwnO8AgZ1hVUsmSUQmfGqSLNUyQwkhhTjstjzl3aKUSoAQZPY+NyNC2ZltnsEjdYM21So
lizUrP4HHmy4meNcKkmGxFkxbXpyfGnpnJX+QVF3D0oLPQGVDZQbPY8RnknhEdaSV2ProsxCGXDt
JRyoY/OzVyYlQG8sxf3E34zR0Gtf8rRaeFRoylEhXQfdf3GTBJy3ohtnKkqOtUXi1bordVmzf1GI
hCkRYlFTME/3yaxmgZPBCxfXQeV54GaNyTcktJxjEpniy9NIAocQmU6eFnLwb6zy2AdNna3cHj3t
x+SULYQqcOZPM/0Azbk403HwhDtvr2vo3MxxjKQqtoWle/KfIMJxkyR8QWB4l+Qc4yMmZJzLG5lX
EDWHvKf6xIwr0unL5Vfwitq6m6UrUA1o8UqpiMP8JW3x3puO1aUM7s/3+tMi1Ybw6HVSfZXLV/kt
beBTyl1ylYbBL0WN4VUD/wQvwwvdjktxkWd3Gl2lLOfo56zHzq1tseLxe/ei0RFRz4mo86S8SIGF
Ar+wvdknLzyTplKm6PqfjwvVTwDD9bw+cL3tDNCEXNv0JWjLEYqUQ6PyPO6CK5b1K5GL94/aI4cm
k+HdWHXR4e00gSWlhuLuM5Or4ZuhEeHsc8UQ37iIOEJENMa7iWyZa3J/XbWPdFK3fywJEFsy7Jd5
7vUbThF0Ly/WloJ7iZAlyK3K8vFC5vlznl94dMYcdUKgL6sKDUA2y+Dt07VxW6Sv5TpgaRqbayPo
B6iLii4Mxx1eAXHBWjkvO0IfPAHhjbxD+d+zPSSxoohKpnY616mIeWIovv8eiuIdtqeRPSBhVE6K
m/rqOUbI3AUUigAwu6chymnmeGdz4aIJIvw2J289TJM2JhHbHksibtLAvXKzJ1pv+Y9S3Qu+kq/Y
Jhq4Wk2Y19vDHYBvpBbDHosrvhx3M1+G/yOgToiTALL5WF/MYJpiJmMeFmCQ4f3HmDPIPdpS+Yk4
n2iLlSDAkOjoYxCz1ji0qJlPP/byH+9AoikT1p24irHzepz8mwcQaOv34SukccfYs8WiYZ4GDGYo
ViXU6ooqpoF4s6tiX67ttV2mVU3P8y+fiT0ACnfq9MZE7mIfJ6ba/PbeDxHhfwll7OchqBEyoEHO
GW+17XCzJkycjBKbIzQZpIFkbQsiTZspkJ3JhOZtGLM2CW97Q4QEAKSeLBtAyeZAn7mw5YI9kwt0
7Vzdlhu35oY+AIvrjyfRU7BWAnIseLlH6dlZR/Kh0F5GlXtKNZvf372hFFEfHPxFw02wGJ5+fayk
7J2rKiSmOXFCh/NbaL5kp5hQgKW8jXKe2HhcS5Wn7hR5Y7J4oi7t8ENmxLoDfyCIo4fpUWrngbqt
S4WJSP+Ap5emJ3NzyzDRp+4Nf6ZT8RzCJ97qc5dPfUsotEnaLgz9lrdqKFpG8W3OpwJ8Xur77ehZ
OKunvJn3+jcIHV8fMJ69Dkw644/uRKhrmthWxgzRPm1Cq4GtK7t1Y1AEmXhfJfajPQYqv+BUGycC
fd8aRpMIRqs2FirVmB1AIgBTj1TvplCY5XyTIfUZGo4XkZEDHEXXj/Zz+Pn5TpFug9lj7UT6OIqS
s4triK5bGLyMyBC440wL7vPd0rpdzmuF/fSoO8seaJUJCAoNWsTCm7G7lvvkUVjFJ68PW4krbU7s
V5n71Z537xhFeuc5Y5bcpTevoTm4x/Mr0ilrhloREFlNzZGJKxKaSUAoSvHNXClML80qndE7A3w1
Qjzt4JHQRxa3XvfKgh+O0Um5K1NSiGaOmYauEA052Jm8xSJdZADwrKvMaTaL3WfgcLuqj9I5wsZp
MGdtk3D7p5mc836W16YmyHxZGNVyZj+I5kA2F6G8LWG98XH+lNiVeFqg/O05ve9f/06ckRC8gKTZ
yrNZaC3r0jhkSWbV0wxflfPRqApcoZQ13BUqcT3LtOZcuYgEETgnsbibjmO1EHMqpfLLAQCJ8x/k
3//GXjY/OTrCFqmwuMGyHbvdILwWXpxshHdmyyzfqp6dx1uDzZ0OfOV7pg4njKHflhe8aqfNmYAg
xSdPj2UNkiEUFE9ABcyPC82nNmu35Cz293/yx7SLKik6RLBzb+TP04QyieTjBBWrBCa5aQ0ndgtn
h1V+uDLyH89SqYBb/EEGekeCLVB9eNZ6L40r5HA3VfzvpsUHmY5ZUN0hEk8SfS0dpolBEGxJ/ojl
aU9eGj17Qxkgk8NH7cP5fZ7VixqT2bzBfWQyNF1F5kckDt+/EhjrcOlkf/NvmfNG2J02v0KHaP7T
e0ROIXsgbK7ld+eTlVIyePZttvA/DN4mCN0ubvvhsm5bLdj2sPdV79SFtSrfRkMVqbotDddMiU3+
1ERjFDKCv7bajxZxTgZbsEUHzP5Li8pyb7vIR82ThneoNcvQEihOX68PkTgc0+wEXnSvdJmPIDJu
KwImgW1zdXSDZUgUtADdsxf5Ub3NOZGCscsec8bll9qfXHT8OjxYcpXx0iuHI+SvJhYwEGTSC9UP
3rGRTsh7d8RaefIeB/84XQm9oRN+GWewynFJzSl0YlAQACqkWXcvP4bGjH7/X+gqFFrfr+RzoiHb
QRxXNlYojr3lesslI5EPKzfE8lzgBynxblgjMzJcB7bsRN0FbJiOreYY+ZrTiX0/j4udThNXOCJq
Yu80/66aea1mg0yUAds92LS1DHmgBnZJlh1N+XrStCLl96PJJW0yMd4w9uTK1j4EP1sEuHnOomhd
6CQo3vhz9LsPZ5nZIXNXV4QogO+N+vdw7lsU5TJLdhSSngp934jy+BrZV5I0WFgzj+BN+gEdGHnJ
Wk29MRr1RhAO9Byu1LU4n5a4bjCGzMSd+jS87vixF2eIMwjxSeiASLgHcShUsHqEPYMYiitCtSAB
0NWVFRnkRUXEOf54BofYNYGuXeod5Hoha/6eiHDC3oiJJBGHw66qkeE7vOVb2+enCFmk6BuEzF1o
rj9z1FEydbjR5CtIYAkoQ0zLhIaoM6cOzpKgagHEL0etXJRJdTY0arf+Glad+fikYlV9tPtDtGE7
CVRsMQyF8+H88EMJTELiJdX2C6hm0zEa8VUwrsqaP6bEEo31kMStflWX5FEdICEAWHm7uhqnZInN
M7BAqVqN7G27+rLRNrA8n6XeDqAoBu6vrELv3kc6gsVb9+lwazCgURgsrrt+dMBRxK/AP0K4F+sV
GR4rhjPfskE9+5pTO4ZUBwovbDmvSflEljhDlixG4cLgXBKH8K2imn1OmmRNTZmsH+Zytb/h+/DT
g7bxLSTp6hEmndTN/BUL1zXUUVB3Jv/u0Faf+72NM5NNr20NHj80yETdJwqxVHaQQznhPX0RgQ0+
b/x9gDt6bUw7Nt1GDUBk30sBF4Fp+9shDElFGbNmZUkyxQ6MjRwvz1pKwmmwmht0E6tJ82ZZK1w2
qdosJcW8JmXQp3+cp5gIMSGpC5mLgcgKCqUqeT1/5pHsV9PvkKL4MVesjpV/CxZBPqH75PXGaDac
Pe8UgQ4PHtB6TmgxO7EkxJ9tfb1flQHCdTac9KA4b310zjGJR1zdxScqSuPlaK9PiWg/18+CHvZF
JuiHQeF9ME65qnoKivhOCg/iObysZUWOW1NsD1zPpvzjqGZQ5Kbcib87NpNVKYkIBfZ6r+8vnoMY
h/i3BtQVNlTaEtyfQM3e+snJEuBpxhXMtAL86kbxx0Yyk76EbijeOayrzFMDr5tg3VLh+hybYuYS
eOV3k2N5LAcv8OhcX7LMCjNctYEe9d3T2/3N0AbSgNy8uPhDkE2IHEvdT/7htwbsbV0NFWw2P28O
2aNQWAXzc/CSuF4olUTj3/VFGwGv6lY1m3ZPcrpHrSWGAcnOn0pCE4TCkLooCwb9N9ghAv/9WnJd
h/1HtBY/tCMe3NneMyC0ilwbH+tgviAnqofXvohFQLDhe28kNV2uZI8y1jMhnGpIz6wneFn0kC4T
Ujn1JbbPg7bCYWWGAaqoor6MVPSXl0oZkwBwI5655U7f3ALXfcTLLtaaC0hfU62FzIdRnw0iZDQA
PF0YjpAK7vb7PCm3MnDxxoZj/hMPstqfghqQWNo7Cq9Iol0xmY/vO7JX2BnK/oXWsDYVNcvrykYc
+Hko8qfgQRW+RDmARyKVlYoExDGfFZyeZ67nCpNYMuXpN8Ad3twJluWg0fYxcOuv5QCTbrqkzqZ1
0Ki/wQ1ON1VdPhEW/28g5/LT+uO8AIq2/KsTXPl1k8cJYHlbHlzDen0NuZ2xkAXCunvhbSGj7NK+
3FjR9tMar9WJb2THgaf9KSZfwTU1SgDaLQsuAoXBQbsSNoHJJVYc7jRp+5faSNq6I3s3HiOzi75G
lb3kffFrLXR7fuN2wyT02DasiLLezwSb+ourTwoHi+pWs5y/ZGLe0eS/sjLA8b0KZ4+SJ1GWIfKD
uyVhIlFq5HRE5MrpOqsSxDS40Fu3ELBA8AlsNsyVMKw3bSdhrWxaIriLMjS4JSqpsUHSaDkYzUEB
Fd3h3rK083INuev+WChIc+k6p0C0FlACVJu6kG0uMR2XYSWAdHASpON60MZ7yCkdMt3RfO9afmiG
VFmeJ4X3ZTyhON70CnVHKjtACvgA6WFmQB3ZWx594DD4ybWjHM6njoEDYpuEAOdb38BQgxtGSN9C
ZRzMEde5TfhH0ZbmLTx3OKApNflWrhTjsoXXkj0mcD44DQdmt4fh7kr5thXX6Lm1Fsg61mpzYfHq
iIUgeEY62X5e412oqgWnguuyOz0UM1MO1pWRZEWyh9n1+OTxAS6NHD+Rb+smwC/OWrOOc4KIw4la
ZCbgbgBW87LtS/spdsVKcd8ikHqwITrT+QtO6Bs2wa2ucVW0XXlujdfdF2LFqXUjMKpCrTM/U4F4
urT05RDFEOEyraKeWigMvqfcTcJm0L/5l9OHp5yr7XSPGDhLkPwrTGg80GhdRKz4IZTWbu4cPyn+
UI0O7rhs/Pne+vNOaPMWXzZkia8vBd2rbqa/k3OWq+q+8Hfo0QujrpKUrvYz9x1+H4UgeqdPXrIX
3HbSn1UT4/07B6t0l7y0BNDB3SyUYpp3oPpAvwYzR8ou4jbBVOEyMwMNfBps5kvh/AirgnNzQ2V2
wzbQHDDg+4SUFIfJFqYtm/7+o9hrQrAEyZAdIINfWeLZyvi/IINwn1wu8f0wWzMeNtH99OHj1j3r
cgoQoCqejlKv7Mx06XpraZNs93PTWKi1CXAINH3cYCU9DVIBJI0vQV0gpI9Ze+E9uL/7NLW3yL2G
0gmKMig2QUmUnJV33fsICv4ogPLzk2Wbc1CW9+CxB5jArB4v4mLub0ZLC7ApImcWBhsM1v2KH5aI
tzSiD+LAbpm84Pv6AGJiMy5KPwsVb/gYdP7hJOvYeiwltAIKqyBZ6eWXwCh6iDZIQ2wBMkDhrQCV
jMfrulfF8wcxP7X3q1vYH9KHSht+HON0+2H6MmlKeuPY0R1BLye3HO3tNpcst694KbERRZ4dfpzj
sRQm/ndNIkbMM9bKGgjA9o8OjMrNGquUGoGH8npDU0805u+CHOFwp4FhgAOBD4lOASosA+z1QEf5
UBECQDEA7nAke8P8ZGOyBeXjw9yrcrLLSXLFLgAjWHyQvs/Rcf+d7e8VFKV57c2osccmUrDOc+C/
qwJqCiocCR7KJuM7kHbkQuVQywB0gB3Kf2gjZg30NAvBfJpIY47mvJ9CFUhvGrfatwEgCyDplbiJ
32M4vrTzxpotmGftQu++o0c/95fuVeBbQGDOZm3fSzcJwY/P6DHhpeVJk84OgnFUTEr+O5Pqx7kT
W5caz44FkXaxpzucBZVmI7ia+YlfNqs6EERFeJQ3vpS65l9ejTzUv3Gof4vuaj5wc+/2LZYxEOkz
d/LiydXVGLYf8wx/PF5vivzYjZCnPptXGvT14JVNAbd7wfv6yTGWZnHuKR4Zl8hN6zAgrdcEk+9r
fchqOfgo3w2JBw0ZJl3Ul2QlXzTNCASsPJMcDrI7aDvP+h0wXnUK6AzQdWEVLMK/kMI4GaUQNRRY
m3/Noq2eKnB6kBEyTKBFKSsv/ewKkFUytJ8oC1lo1MBY0Zl30IoyakrpDOrHUtnJGmJapOOJnwUv
hU6JumcFt98LGAEPCNGlbXQj8/h+jXf8Qp2nITMV5t0Dpr2jjjkAoWuri8vg6lQMm/7PK7Ii5dun
MNcO6CA53af7M3LVrxdX//DYk7vh4G4H2LXfhsapda5W9V+Y0jC0dMmWA19UvslcpDmA1snDDFuM
sbs1H94FD2lRN2wUq2qhXm8P3wWGD7t4eB4DxYU/6uNg8N+shvkwEdJVp2e3pTn2wGjCg6ZVVV/G
CMr3OffhNYmKG4rJlX9eC9yKqT8OQnktO+SBPTw80ELiLY5MPf+8lHqoHN5GPeByDzhe4w3HUwMB
egWiizRn/tLaSJFvjZWL1Vl/1KQr/b7+4u1hLsgyzDKzmpd1YToD0EESWv7/jWixfd0ybY2+QqcJ
qSHnQlNL420lvjT9zFrzTpFLK1URSkrG2MVBlIrZSdbfOWFoeFKXUOJ5BFoqBf70+67+AkV2HlLE
+VraEbSkYOa1uSaZEdylBafPV7o6MJbpOjJlzi1cDn/wky/zHSc21MimyOR78X+SEKtSm0QbSfFk
XrMY6vyIsjnKoX60uWDs/DnOF62p5/aY8mr6JrUE3lbMaFgG0I8Ju8O3f8MEk1pGJJMvNUUM/LN9
W8673AqygpQ+2yx/xSy8hjbRzHREzuR3nW6V67Eqn2bysnLshGhRqGHnndx3yebg0lW3giamvtJh
h8JqbU/zjuVsdUAw7dy+XxB7UpzKFzhDk1hl1F5z1Sn/g0QsqXiGoDo7aG/1IAxNF4md7nTXVjLJ
rfnANZXHvDDdAlhnnt08vN2g/nw3UITE4YHgrtrZOxobDvt0GMGFNBq74noT1je1Wo7WeRpmCcTp
GnizA/xPfggqX5u/eMoLv/0t/yhy09KA2TJkd5abCa2LkUn30Hqx3pP9+VA55QxbqvFLHzsu/7Wu
4LAYGSCJMgIFahdNRLxCKdZJCvxGktfU5G6sfryQYA18iKcGenn99MqI5H7PXEQX7mxOipAhopv6
H/DRVK027I23BRaKX+xjuX54k7D4CijKyvq3YNj5nWjR9/KVPJwOWj8Ai8k+i5PG+cdsUxqh8Xjp
8BV6r/Nnodu3PpAA4qjHqgmTXxCO7Twk4NPTcRniy01xORIraIdjjc5X5UO8Gck37vWzMr85KPvo
I7MJyjiYT1ouZHcyphenGInC5IxO+iIx2fP9wCevb3cntzPwnKQCRa1It8sW8EM+g4WiTj9pvv84
jh4+84Byn9uqdF7/mx5cguTLv/y4vrMKCf6fxL5TZjZlWcLCfD5wSASCaVwcaD6zol1IouvY5RpR
XYAEoXrFO7QWHvktT974rnFkPIrxn1dBrw1WwZ9ziVTyaT5uWffH4PRGGPHtGmcJUe4tLuF27EVy
2D6PkjlOvC3Wpt2BToe8l9xkKv+4hpFYpf1FmowgabXPV5upw4Wf3LVkUr8Zen6A4Tt+5BlWYAH5
ZcAroo8jKYRYue9USjpbtUwuHCbycHxElDNLfC6uScraccBtMXnC71tHFJwLSo1JPGKsg7eKuCmL
+F+L794hI2eX1HQHp/7nf9L3dSQs1BNKlOCIupm8bHNHW6xYXVKuOREAnM1RjjLYjOlDdFWqt2Uy
UPIcvMOBspU4Zedr6MLYffaMH7vgcLeU/yaE8uZ1hKvaga3OemTnaMvC2wuxaOR8v9+F+XjlQ6DG
EFv2NltPNiKF0t1EAWEBMxDHxxJZMd/arMTnUYJN+NW4Y6hDDacbykp7xZM7Pn85Qmyf8xtGSODV
5UwPw1jezm6ZcH/77FdpBT7rxvHTSKEx95oCmWYNy4Yj4WByzhobVaPBxH4cU+/LiXea3aHUWBKw
uYvz6yyGvhw1Laou8lpqMi4o00S4dK/nPbsdijagdUjGUMoCKq/NR98W5Q2+Q8V5JX8ekj1ei/wF
UmGh8jkKwJlcTzGpROSPnt8KqaAbQ8AVHhgWVuHoW/GdPKOT48+/OJ16L4jUwlTi/K301iBQ19gO
K4+DGZE96UwZ6NjPhuXqD5J6/2RKhN6+n8JFueIgbrDXIrha5gTFarpyQL9hpHYvEeJ6Qv4p2++h
x3s4wCW093zSV8S8z8ibMELO8TezXcpMQVOrimJ/fL75GTMG6vY+GsOuDyqD+6SFddx4aQa9veL/
Ntfss5fvFvmzLE+pqiyOm01WbRrZ6yhW7+5yI570x1c3eqgSQSei9Nxg09ejCqH9/ZAEFJNUE8b2
iqZQl776R73mK/6VcZ510Oc2AtM8IqXb8FpNl2r2HIxRxUidFp+c9YEkLCfsr2sV8v1+Q4SE1bLg
3JJaBaPeJGjmc3s6jVxTntp3/BBYAPO7QE2qbdUSR8nYGH/Ehi10Rd91PmRH7mH2uSBNjPBAa3kC
COTHTo3Oh+9nZQGJCmDrz/S9yp8eVQMFQOiaCEj0tZFvLKJ4t8aakQhD1B/Jwz0Q8IknE/AeO6hf
Nj0whCzrO9G6GRJsf3FRTNPmHh6PcvJS7ncbNOcetP6cZXb5myXqWb0UjVBUaOg/ig8nkFCgHTbe
bIOYJ3CqTTLOhjezYrzQ4lwLbZwy0Svt+waeL1clu392SFbWXP7znxMjWR3X2a4E8SRg1KWzf+SK
pTZPUQmcwERgJ0/YnCHsBur22cpC+t3bFM7BUjnJ+Q/FlQ8LCyN1ti+g0UnDiV8xwsRPflPTTUp6
D+XiPjUAluf4bNgcwlAJ27W7XMMG8SLgDKVoTqb4O5zusgu4L5mjvMprpUILQQdqsfnsgFuPYhnr
olvOEMFzf82hVC/aIqoR8nW1jkTNt2MsFWqrPhrLgQjD2JhRssp633ASaOuJdqYCLDcppYjj8RoZ
lYJqZ2mrKiWsPKxZ91g9XIQc2E4pp6wxtC59TWme2qDq/dEkU6OLEXHe+NdYplyDhJ8ZKGoTmwKY
6iIo2nZHSZUOjSR3nf3m11V+8En7WoutKdV+3Zvp3ScG3AFc7PzT8zabolAGnVRmEbmBVxfbpkdl
gIKyZBiVODgvaEXFMBnuZHe87ZE11SmgooVuTv2Euefi+zOICQSG8uY0ILDOJCPtOm5unxHtB2nd
1M2vAWcL9ku7rJlDuoFRPaTYJvpD6vjp3mRG5QpgH2vj9oqK2cFBZdPEP0SnaoR8pdKBqAckkbkz
4We8DYSGaXcBwcfJCmCyxnznOMrPoKVklfvqBVGga0b1c/hGM4cv/7/ujpyy0NMe9QkiFkfjKtg3
1LJLTFtEH85BHD3jqBaAzJYLh5Y1zAO3MnhlnSeaw9xDOfQ22g6s3SXOvPAQ215PBSpzAiPop2+4
unZ4nKt3G6b4PRt7LaIxml7DqImvaigyqV1Qi+Gydiii/IFRN1aPTAovda91Mw+vCzh7+UW62lJN
Q87+TVByTThNycSvMJaMFiTZPsZFtCd+NPMs+sgIgDTd03gzGMDN9UV6Xc7FLsL3RoGhQ2fKcHNK
bwYqYgqDy2bUT84eWpP1WE1VeaYPoWTS3DnyGD11jkWeEjtbYS98mgE3/wm9uuDmFtd8rwcTB/kh
lWX6sHjYYAYvlQ5LWBq9AOIzEHNmQI0KbKicWItxRzjfFcR+PPdgG13DNUxSS13hlDubpxGDF/Qm
cJGPeE3yetL5Su1q9lkiOyjQqhROzxZxCnTPY61igZNQDNBG6CjkclTg3OwXSLb5tkXvDg11qgxD
Hyztwg5WeembY1PtE7/5LFkkmpen//ZDzBok9Hjym2q/0QuA3NmKTCw4zg9K7Q60UW8gXXdZzF1S
xxIt5rzoEviiS8nP8F2eV2K3TsHKgGyw4zQNeTTJ/gDZFaWY3uO2RLajjaxYMHkJv7b5EfMwEMyV
7+1NQcNooy7QPm7ADSbVtBPMxxMopMVLjhKqIRLqHFmcT6pJAiZjo5P/RcdtAzc7e07Vol5+7bg2
khJn1m6OwrSD2Zs5HjOc/KwkKh5F7nY9uRw3my3Z5UgbzKgtQ0ptSzxS7EUkc+97J0q30tGKjWQn
bEPi3KwQzK6+86UZff/ZKy4V0Ga2p0n9X1wpjZp028Jg6DbwGSQ2Tas4iO/C2BOerpxi3t1fVoE0
WZWHdQURSeDrEFbuuRlt3ztDn++0RMMkG3FEbj+3Pqkc/MQR7pywHIWmdPb2l/y4phJZZq10h3jM
ETiM+VUucMZEgH4nEIAnie9/kJQzaU5Em9gnQ6xLe3Dw6pbO+0ez/CtoY0dGT1Ht4/2noxPzSuVz
Rf2BjY0IQHukd8iP3fz/nFYBk7AR3lUEr53Il0KOkaP9GZZCSN7DjbgnvEYYBWmqG9Lvsbd40hg5
WtIaQCAyAhmWixzooAia6pa2YgqeKwGcAcoH99/SSfyiPlP6f9+tuM2mOSgtYygSDuPzLnIAlDyR
lUkYcs6DKZedHYL68N5NzEKfX/xVw9VUvZZrGboxy+pGNGWHtVgm8CvIJRdhSBJoWZD/jxOblpmr
nvjBKqLmRvxJh8395gRiRdecJOw/vlsoqM5DuOmIw6rgp1EAFE8QeDH/+vGplhuh2eMwigMiFDRc
4weP9ckTGISRRPxPzPFPFCduSKxFtld+4dUvO0HJ2TkrQo1oJxPJpyARcsUggoVOCnlpvwJbwoIN
/yoQgMwDdbF72rSKrmlybe7ZfBRvknb+5QQNd+aecL8TqN6unGu26CaWV48k6QN0Ejt3AoQFd9z2
8H3Ol83zYmc/iGenFrXXZ7ECgCP6BzoCthT83pZLfZjcnCP4wyjF6ZL6jdBPPIG3VkmwOKAiea2b
KRHQC676ckACcLFDP/QJLrnzlJ8/OmVkCLCqiinVG2WOVUH08Ku00A74Nsm52D3Cp+v/ejVV2Fsh
OXaOBtZrO646ITgteCzqwhNHC7+yijOEYaBZ37Qmej0VsgHi/3isSTZKDchoMyey4vIKVWR04FUA
KTf9ehv8WUMSr3b3mNeIiwZ4L6KDwj6HzD7vasIE/FLGXKaxmzncUd1qdV5MSvgyWf/LPVQkcmK+
rLA8Yt5d+K8nEJ4nzgulqS+pvym8pqf7t6F+HExaWTKBFYlCrBaQGGd0jX7A5zwOkAoPUl1uAHrU
aJ23gau71qTDODVuPZcTYmsgtRkKTYUEUDIK6HHaIBLycQVpEGr7AJ7D0VQViPgS9Tfzhd+wL3iT
Qq7oflFAYu285giBfZXk7hZucb62IdQ+hu6hVDxzqb9DGkmOzaX6dwgvJVtPob9PRX6UB6DJ4XZ2
owS1pLQXr9dDzcrzRDQ4TCUY+CX5wYOpB6SoH6hgtkhj1WafGq+5QQiVxe1o7HrT7wLa+T6GqZGw
i21tbrOan72UK07G2OEE6V4Ae2I+GNcz2TcL/59FrWSkE5H2MV4jFvQaOL29lVrKVTyCjG0Dnqui
PMeYin3t/2Ivq3z8ZucFCU9mRaQAZKXzMdxNhTdBHPV0QrCQY2rwzeN8Vj/EwmbX7VuE/bG/yuwL
62U/m5mqNZlEK/j7HyfHuZQkRelampUz970/g8HnrbdEZQ6DXf7SxNCk9SmzKKulT5HpXPrJTzQr
OSNFQ4OtPd8EttFxWAE1F3nFp3gIdKE/yUFAr1mDsz1AqqpFWEr+wjBeCvp3srnasuj3mmiXt2nb
v9cCLGmsLLlgs3eftLpXrlSDFmYeLoB2VdJPmEHF+UvtkBHLUY75sbixqdP9rN0BM7WxM4Xxac1A
XUj+N7CX0BT9XUkuRrGLizKGQTzwaH/jlGaAyfHmztB2SqwYFOolE0HoxD++6L5Q/Ie1XuKN2DIk
UMgzyDdcCJ0gcbV0xbWPVMmB95OyfbpvBD23xHfMPj6VbdUKw2IiV7xJ4NLsnFdvwZrgbal8TVii
znRsv1+mOpJPrphs5K4jDwo/tpxOravxhO67th8DTLUdwXV8+0qxvZXydgM3/iN94G1xk/pD+95K
iMUeXT6TIKazloZpk0a+JA071Q4hqe0ez4V3TGo41PQzy1rmtScyW1MN2j7Pkg9/CxdtvEi7cc7o
1X4QXhjxH3zn/+ahNyFpMr5fk8jXWfuWTVeppZRPXX8ZmjxfeO3SjbkeRQ4F/zbx+qRjGCkewa0u
acMATwwGVhXJ2ssjOBtDjvAtkIaeDv6dqqxeC4pkdDC5rZ0X0qsBrPfuWp/YUFtnyrzhah/M4f92
OyqyUUSnH/XFFWpfSsn7LLX66G1WdwnUdoZPk6W4c2EzHTuZQrCXj/PIqG9fSv2XH+hm/GYzgOCS
1bBlGeAaehSGoL8hECCr4iEDhHG5KtxrY921SZxprF8aB08Y7RlVoWofRiMyWkco+fcOI60n0KWU
Ci5B83ia8PSeTkxJNY8Nnw7TvdkRAP80kzciVb/5gASxTKAGeT2GrOcCuAzVHCPYtH94O388suRD
8DkJIcaIS/pEqJIU8ce9rH2eFm5njFM+tsl6peg6erpoYaZ1XhVlI//b/fmbTNIBkODWxTlXSRpp
rtdm5Fbe2dlTgovlIoeXfWbe0PYDN+lZt/gVtpyMYKV4H0mmtAaxqrHeXzZEYx6fh+FxfjlDf3s4
2t70RIMMD8A2ILS1xFrST3H71+KZXsA3MHzvjzHsJdBVsox/T7v2xK10rOcNRYfs7nyrYKcChBy9
F+cw46DYG2zpVap53ypZV3JWF8CHlGmcxFcK71iqzNr1MNDnRKZv+o7g5SRE9FPWuxMYj6EfcM6e
yBQgRYELNBH+UvW7n6BESoCxGlys2BRyCUsqEUIpUF79oA6YaC4kmfk6R9N7mEpyTW0JY0zt3vKe
2qiA2tz6QpLXK9kctJNzJ4hYuVTaU+zdbygwvqzODhr7HFOt5SHCho2scIzToZLmGUDtJk8loGzE
DWQFUkgKPQNjJz032UC/FPlMMhDy9qfEgDrhKTdZmQ95BLtovzXWz0CuVXIYeoew+HzE88mIwhDz
/u22ZK2t1ph2YhwLuREXc+RFZbbflYXXilywsqpMBfJW82RD6kOrLDDRjWYfBaWSSg7K23pR1kK7
qYoajTGcktVIcZ0sjzibkZPdLAEu68sJJdqVb9wPMXGJ3NHEtjnyOrfSO+QemaVOgJFnm1rYupmD
XWOsvLMkiIHDFEaNLZvDgg1WHiZdrEhopTQB/TGaWnjDZEpR11gnGNKWLx1uO5McWSBq1O9rFlQW
R0vHw3C1a2Aj9N21hZXp1WzniaxmOtB65wC2UXQbJEAAUMJcQ/VYviPjo337uiD49D4MwzuRE7SZ
jNH8usLHPnMyC9M99qx7Gzgk3p+RG0YbkTepUtbgjsGjT4sX3Ay0zdFpjG1038Pn1FHvjfwROBO4
ypbAx5OjD1ep3v78XzY+zi5jjgeYac1iwCo+37RDFLexc4OexohMBouU7kVS5VXkN83bM648wP1M
QJc7pWmkDCVs02UiHvD0MRmTJHr4WO8FJKLXpt7JKTfwFB3izAD1T8XoT9YjigUosSebyGvQ8LPR
Pc9X4rChRnwgk6lDCoUp2OBbf1x8WXJZZE+K8mX4uayHHXMU/Trey2zu1/cZt9M037O5y4+h/VBf
+FP4FHSzuQPsXxa1F20FHAjzOBUyMQEurun7f9WkpbUSiuwnMUIZKY9M+QEWzakFYwME7R3z5vON
kriFjxY91fh6KiziQutGru33G3GxwMtVXuBoG/9k5TI4nZq27CoNeiHbx4P17OXEgH7p2+YoOBSf
RDM1yaDM2qOt/Snd7/8F9aiwyoNAXEtYAdKhherXwsSlaMuEhvRVhWvL0hqMYplcu3cCfm1bleWR
qiSryJpfJaOlQhFD5Bq88NilKHmSQ2pwphq8Ret/p+S8ZMRxfpr18R+p6CilpgBO7nelPY/ipZcr
W4V0NB230eCRdngDUS/7aYUtZ6LijcXENdc/PSxaPL8p4ZhebZboYtqHruTUTUxn/xhRimsEpmJ3
LOw5sLvXiTKYtIng9LSZKRWS9KR2Jg16GAif1xIgcmHsq92ssI3IRq2efj31+r8OjLCyDvTw2EJM
DlgQBjJu8J/id7JHu+MJu0fpgrPUJjfSUPIp7P8j94cCYnFDu3kHHLEPaMaVa/fngI6M+nvZRSfd
O6hnkvn34KQdu+jzzvap/eehNbxrf0DO+BP7Eq7j4fHXv5Led+LBB1R6sdu1NEsVuvCp7pjbMp4I
gKvgg/MTzoU0npApihoPiYaj6S1AYXZglealTj8cVlnsgAEi93qeOpfwlQvaCF+k58cR2B6lHdUb
JOGEV4stWybKOweY9yLQYRTOzFErXV9/Aj4lIypXGtI803GkUVGv2CRNLLfxPImF1FhaoZgnEapK
NWqJgtbT90rK5oOIRUv6+heqIbM1X0vxa+CCd5gGUXSPBg0j3lf//hkp7yWlrWdic21u2Y2hF9FA
smWltkW0/oza1yU3FYrcoV/vZ51Zzso9wKGdK8Jv57/RSMiMQvqqoPBDReJ7tNnGaysR3Mc1c4ck
UokOtQZEahdTPJahu3gc4OUn2zRHDnDZA5HtFkW8IyO7LKkcAuD9ylrO49mq9u9HHtkKA077+iCX
Zh2ppAVVhPJGcng/kFzfs8L4Iqo6WiWW+nYyubW5km1TB1Qj/gP44TjR0QeOx1UmXD9P0Y3pooX/
QvR9nQTi/vuVA0xnQSG6Yd2DHtA3GhNIO+zejzS3Z4jP7bvdAsL4Kil78V3/EyYfwPKXr5FS/CEL
sqVJ1GlWZa5LYKZM4oJi2nQBToA5KnmeohtK5wM9BYCDDmxNsHSj8IhTW6TpxlvCZ+oEzA0tNg+B
KDAYabXtyu/Abg==
`pragma protect end_protected
