`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
ppgLQv0CJpVVr3Egw6p11wO+Q/Mp7RKu0NuFAXq+LGNj12wFjt5Suxu1owELCkn52e5LyMVM7rlw
qCAYboftgUlRAaE/ODgAccq7oKNKvGfdy9tXu3f0THwySO9oQ6JliR/x+3QTrewi3SGch1XUHDeV
XDZKpQJHk7XtIH+eTFVDcuPogeY1qzXMcscbVmGtwZGjTE1xP2mTHXT4EFJ+7RnhBakdFhF5f0ov
UNu5ZfpoEBJECfjYApI3RZmM4oDmB5LVx+bpLQq1HkNTAstDfRiZrlorQmW83cc7lQXbcq6HkBIL
uGrGF5kQbXQddTSQKxnVH/4FLFeyngpbL9qNFg==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
bDjlKjmNLYDzR0P+60wPTq1oNfdtKxn5S6Ma8tbEMigVcQRU98ZEdhpwT8xcS+oZGmn2EOF4Xvp+
NxLertRv+yPhbhQ/qeUKCpZ5gycHQp7sRdioSwK+18PvY3mBRvwfgKLP5iV5sk2dSlJtnVuvsLpN
IDZSZIiTrN5cITyVs7I=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
ox2fAYxA7cZjtuera3X4r62llIr0zD/9QGlvXaG3e7OsU94gmO0xEAJ+Nvk1XrWsjwI+CPFoLEOK
yZ4h6+Sp1Zw5BUhsDUNbh/1y/BTGYLAVqIZBKaT3S6wEqm1pbdUdNAODzzaZ2E0EFSf8N01jqXEM
tctpgON7M3O1bLYQVGs=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6048)
`pragma protect data_block
Svmp6DseoL2NVrGhbzzfuXBXAkZfCa0yUJ53Z0WIi4bFoYJ0I6rxcqIf9p22vlrhZL/T8i0w3Sc5
LwWaTOVqOsGLvAAHlBPXevy5Tux/MtDvpHDHnIiiR86MT/O/4ZzZ22YwaaVlEXgkZHqgZ/fgBfk/
C4AsYaycgrtirPs3+nch67Mn1kvyCrRXibBGaSVVZ+9AI0JOont1KHtsnJnGwDWVPyonnsAX9lbX
OBA4jv9vtGaDGNS/IhsAFXpw7L1Us+ce42n2D08Mqzafzg9d84wn7PB+9dfMXVmcfaTHAQMmbLL6
5Ld308vfcdKY81KT32GrPPHk6JKMIl7ZVlTVH4xy3WgZQQ3joBjHo4R8cl79CbN/o8QZyxQmuCbH
F8/PiJXYT7jp+DMF3AhyDdIQGkD1kdMyEGfzfCREbr6hX2MAQLgqs78C2xd0DYrZTz+Y8n/70coY
3q/N2qUwhLwZ1j+iGBgwy2JhPfEDL94C8dZd1u072U0UdGvbUEqbB2cL2g/3NWIacG4TzoR2DlCC
MQmVOCO45Y0AoLoWgI4U50R9k489b+5GAwsCSWkg/Mh2ITx5rM+Nx2vMq2D0UkKHM4B5T4V0bSiL
Xh3GpPfjc0/H6UcTsrg0KgeRxxmxd/qBL6Qk9STvSCeaehEGgt9IAKM/JGQetR6J8tiR+VtH8KkU
FzkriWDk5u3LpxfLBNx93E/8ffEMUHm4tJJxrqtkDz0oMh8++4TSI8dTWaQSmuU4rMiyyK70wLl6
jtxbJWhojylGL3L5TENkrCY24ceIUv88Z0vKgF82wcHUcq1Y1Caqjh23mVW8kG0SqVZpDQb9gS8A
oRyg7bbHKEtIUftHAHZSeQ9m79nH6EKRYFARk1WBcaoSSxLlZQokUdLon/Q+iweJ8EIOiIM4WIaF
zB0ZJAtSSHF46gDO2YCtViaODAs/ZQliIn9NmOYMqoYzr6clDcCkEVvl0Mqw17FTprevB8vJO8rn
P0HdTgdUPaOIkFIbPOeyFPXm9Zzx0K7K7GNrBd3oqJC/o9KlWI6oP/QgFhyZYQtpvqF3+uDAzxCX
NjQpRz2dSkCfTFxMqKK56U1e8gObcbrOcIZd/pUREUOdRFWfAuMooO2FbflcCebrMi+AjvHgsv7T
D0JKecqd1YLwDGx4xmrKHOzLKU0G6MoKzVtsTCZuFW9nuobVd2uHzSYU8HY/Lkm10yvPb/2WaKVP
5J3weODVriu0pfHewycqk/ZY5YAIxBRshv99rbEHTEyuB80FN6quZ56JNKUZViXxXVfjLgtvFrcG
kK6nmrK/z9rUwJY+khD3LN1u1321B7V0+j7eJImnAs1vLP3m6KzQGX/e5NgBCaO4oIAqrJo4ibmM
SQrg3wS7z5s77VNaExsiyvDw93aAsix9Z+Tt5bd1TW/ScR6Az6DViO1cZPHHCe5nNrIEhig8s2ib
sW4p1QiHCQEPIGqQRt0vG97zhe8VdXs/+oyOCACMPzKW/5LeaVCNvxGbFPaz60Kw2rF1z8Rdqu94
QpxL27hUd1OAEzjN2U84Dc/tfQ1s2yLE+Oa4QewJszyRk7zhtJAeZxXRGiZr4/766s/XJSD3RupD
Fga8lI1n0YJSk99zyfXSOR+7AGRIBQUcHI6gePeqX6ZNl83PfpNU1qQtIqdoR5wdFYNbGOF6GgIF
BLWojWyAEyCt0KcqtbH/ezRMcTukHd08n500B1Aut7VXIT6Pf1/5RA6b1TxRsYIrFJIQBBbOwB2n
oR8dJfGGZn6h6hSS68Diu+YDZ//82HiNho0ob9sZidCTgjueuNGTfpuBybOSa5AyixR2Y23XRMnS
XP5yVyOr2OlYNYURPrlmKDaWWL7Npuxl2Uxmoy/zTlqjTF7rWhKwSRaxNgioN4XMFHG1rkxvAedL
FqNxf/ZcI9eeRbqQSKVp0U/eU6j9C/mJ1n6Kza9Jje4o0WUKfD/HIoj3hg98agSGE965FTMO5y0S
FLhxn2aCpE03D+XAtzSo1sM9KhncX9gUyIAX6TbJa+NJZMBW1YVggn5ebHv0CG4iB0fRQakGOB1U
47YYgAcK1MIlP5mky033Bj2WYm6ANJD9evzAQmQdMB0dCwoe34DyCJ8Hk2hfWqqYiUrGDRoTP0q3
l4DvAr7qUrbG/dsjcHZiYAAByGvfyiRgCbUHCiRp9LJ2aVdJeGIpdcfdh5tDmSEaly5Ida3O2oU3
MoTy6d7KxKkFGDg9BKRHsW3hYNSsy4BFIcJShU3YJjPCD+GvjzYg5BR44VVYWkO3oPEtg1hjcSUC
mnZyCALAZxYz/EXG3TdTijmV3MFJZIcgRUB5ACb8K2HQnqc5MKHjL6GFS/7onfhlE7HDXWJ0ErDM
lYVVbKexQzXXDkHiaRe63zDlQjAzGaEoCHO8w8K/CyHccc9lW8VnqNs0B48zKw1dvhSUIm7YmEE4
b9U0SBCz+eDEEMFeEOM9wXoUA8gCruaautByJtxCpj6vmD6g+sslYOrv7vVRCusaJTJSOkA1lv5A
+CvI16PyK3tSk/edzgt8WyVh17WYCgHa4+gMoc1o8zS2zHGQYvUKQuXL72lUqZb8B287wbyglhvR
zIURphl1MvexXo8Ekry0+N0jhtcUl2ogdMDOB3RrG3MPLSUIt+xsaIZE4G5Uu9YS+S45gQdTon/B
J+3J/ZwbEoZEYqJ0P5S0FEUEzCkRWBAUPm4DeQKytl5oSaFM8mtf67uXJljDIGMQqCuD1NSomeZg
6vggspk7PJEaKe8CEKxHYnL9knEDGvN1vz1UiSD2rKu8qnKY1NHc2INgTBYjzYdEQQOqsVNEMt0n
ZGbUw9E5v4PEt2RwvVtG1t8G4sYYLVjxh1XrLLBGWEN/jGJCyv1XCc0g8o1nzoEzeNUuhrBwC9yR
sk5ql+JO4R4VcyHO9JKxCtp5ClAmTYUFgyPEAgZ/7JvyFpzKj+gDxLVjVIYVpTQp1O8XRSTBRENd
lIU+8sTbYGDWZAR8qv1CokW0VAtEA7PD1f2xz0AGqYGen0b1nED3wq6Ej+QAsYlu2aEhw20AysIo
LsOgfenQRJu7L21MCFVS7k9affrtnnY5sLbH0pA8hkHYlfc0JDRiDa5jlNPq1h/SV2f3kS+kfk7D
1ZMEVGbD9EBfQaPN+yeSNh78/FXWc3RrxAHW8Kq/wuq4/fvZwRBtldQiWysXvsBVLNykP2iXpHUf
VPj5Z2iDWCibGIjL2ifaqQ0TKjP2xo/A30TdOQVbj+wGgmPiZxk52EScVhIkHBOJJxvy9ZLS8wju
crtM/34T4IU3tWnKHap9CIM6Z93l+KhUs8sct0oNC54+QNQL4yl3H76W95Ou84kQx5K9drCg86NG
H7UPl9rU1/S1dyo+xz8UpCufYHOxRm0Og8pCXh0oBCleN+SaJngaoLz9HElpnu//xKV//twKS9z3
ufo/kGCeQvIxxTVNB8IvPKyWMJnGgSzPPmJus5MnM7GTs/+LZkGBFAphFfdz0a63WTAaLHdcQpeB
oa3c4CTAzLLj2vk9xlMhbTd8dEaHeNbjsmIOuK5QnmG7hU1tWAK0AuS2gfkNHnbO2AejYbP7DHCX
omZXSGQ3I0XUlB42n0rGqFoXTb48DzpUCEQsquNKZ5Qn6x0eXptsUU+C4YBN6FE2KscJPy5xwS2B
2H/aj47WpJjMKCqoS9p/pPMnOFqay8hQ9+pA++OfavbwHXCMKG7/Y688BizjC/b0dHyq28R3+Rbf
STt6HG2LXAsiD8vONr/q1X3nnBjFnXNa8E1HlBSDkS1yPkRoVDI+Kz7UXr91yAob5Uh+akPErxDW
Aznrq2vb0PbSxEBL8I/h0HVv/QyBxbv8N1TaFcmRk/0uPTYGPkpAHqkBCjbFqxMjHsgbVBlOpZsG
9GkxS4d86J52nidnNblZbrDaPFV7XR7c3d5ljvXvut4IWBgNOPm5BgUKsAcqsPmioIETmGeMiN1D
cHlaJU2nM9k7JC1z4Yu/eIjvtoe+SxbpO72uqxs40LavJIBiVcpk7iRAA/YrexEcoDQ4eP8O1W3Y
VdwC7mzFOOLorvx3unLJiHRQUuLAYR+miPyhQcdQkg8SQYc85Pa768gV2CMlTBS5eOpuiMABobtQ
wzTDN6Qt1Y/6NIBowdcI9whweMXedxNtBfeMEXjr3lq2aAppAyc7AUoF8jlsgKrXTVyIVEBBKaMR
GKsljQorp+aEnf2Vg8d/vQCOP+SouULbLJrFMn1s1l1bjwHM2Ewl8Gjz+0dtaWJjrsCpYYrSPNg9
jQfu/VDc5Aiz+JuHY04FTQxwTgrhXyDh4rijaRVJLSvEdNk4oqzHz2jMbIj6AQQ8TmYpCtpuhOpk
gBfBSe9b2c7QYhgba0ErxKLoanpwuIgfixcUWM9CQntCm3SSYwIeVGM6UUB9YY6qmHNG/i7jNgMN
C3U8G5MIGeUrJ1kwRNIOh+E4burvA98VYqNnmV5rXzN7H6TMR7611LHStvDeG3aek4PY2torRDEE
yU7Lr6w66fvXiXLhkAzmQEzDpUZ09vo5CVOSJyrFxm3tjbwaJkXTJOPGMOmka+fW3TYQhpipFOFg
d5ilJ9TeKzKg0j56L4p8rekwVW84D52rdUlwhVRlc+rX39b5fgz+H69jmbVNQPa2LjKuj+SVGZ2f
zmID/jnWhumiJQS4GasL+xMUTfQt8sXR5WJJ8tnfufZm9j4CD/YeHZaIh5mgPiVdmB0W27MrM0lm
smEeSpSRN8BsGngsIZ7fGE8/0TaE36Am8yzdSxgMH/kDvux7JSiy+FCTsZrlbrp6miAyVqucfGMN
TXVb4/E1qY28LE114qPkbaNiI/XoFh/8Rhi4zXSgCUIpJnEezcHJwgNdJ030URsQtVoyjXKcWhRJ
JGXql3WHvLYTxoxuSuHtqyLwUb606VBZaq4X+sA163A59JBNTcxjKB83FOw4/hzLIu8LECW+lSPf
pkgCZfinTplpy6OszDkNd3DlcEspvfv4B210hob/J8+8NvRMsnaHhy2a2+mifIaCMmtyDfhXiEel
3ICZfcCrRTTTJPrUTZBhadO8MmS0g0z0OsDO8DK8+JfDRaY7s/iDjKhw4ePQLxN4HHJf1fmVDOlS
IcYm3qNBg4OT+tKsLDeY3vgNpP7zuckkfVsCMdDth4lEzocWgnm5nq7vLhb1StQ2nKoMwX4ZbWv9
0qeaiXdxkadaPgVxTK4kHV1AGGV8ucwm4nvnV66b6Ru5lHSaiiuFCArWVI6twc5nKhMp4OIe8ppe
/IwDTYfWD7evNRBcrAwCYeWuXUIqZPL/z/bx/42HPzLKsN7lwoPFLaciMA0wE8juBbmbiD3h0TxV
oofAdV5q/Ce7Et39Ubpd1vsCNKzlTLk9YQ+Gbq6mHR+phhaQ6S82il9NHt6pTx4W9F/A3TZQcKmw
OvCbji1yDe9biSsrN/cuK4xYWH80bRLa9P9cUbIbYMkWohD9D2ZuyWFgPRj34WCKsJv29qGur7Z+
yQ9x7jj3nmdy51a6NXRLhRnG/gIJbUPlcgrAZ5/dl/j7VGM8Ik/Q/f/b5USbgDxN5+liDgMy9WGz
OMIZZtwM2USqVBcOjedOAZAEJ7s4UMwURaUk45QmD3evr4GML6dixOkWgnI1/0PenqpzQnvZUjUW
tRZXw0pPQ6gc77vxN5gJfr8jLQvgGGEpwdAh4sOJ9djiyHU6gYX1+guCOJYylQNvKpCzJynRYJHA
8QmseBBWNt4zlPDFx567KUBt0lJfMi9l8KRAvB1Y52pKvsW7V1Kvc9yDPnOrcYkU516tslTf/noo
s7M1xMbyWh2VOGAoBXWxGRHroZS2UJ25iut/l1PqqV/3aYI7o16dl9vumi6CnpqJbPvXp/GcX7PG
oEZefIjGuf/Y5rApZ2jJHYQHEK3D3bRc2JNY/iYiWl8N3cz2BICfL+01OyZe3xTLxkk45G6fy/Km
vqFFSiVHTsHC6XX63hV6+3bpO4BFJeTtSLnhfW7fNWlT4sTsyuiLaiMlGVkXdCBYmpfcCalLPP4a
TxRwhnQsFKvVbhRvXZI7JCEKF9hAO2X8iIxT9xuJWBm5E5lHuWlBmU5VRrC/PiauKmJw673+5YYk
mbvIPSEbgNu/CIIbh6yru7oIVJKnBxeNdOrPOyAIYvDefpGIgthG/892wX2gITLz1GW9ZEA/kHVo
i7DpuWTStnPTeBeO2vG7JNSWLLhsIrazZzrilcTqDQr3s3K/n7Z2H0/b1q4cknaG75BIJuWVUGNp
lgmBNPL6I2Zd2ICdnTYuIQVP4+PCwnnOo/DcDh3dePGRbf4XhvTKlLKio5enRGXMer5Ns/x/D9nF
B1lS7JuP+nDZxJp5bH7xOPf8kMl2GPIDPamu60tV8eOKsam/5HJsO1wNwIwDHW5fwtiaeAnLIzYx
GCT1ZcQyj19B4T8KhPW3N0Jw+hpgdM5lKf8tJ/n5fFdTnZ9HSJ3m/hMj3+hSoJ7NQAq9oPsz/zOX
cqt83k9+cyExVQLAtcqmpcu2lSbPL2Qtak33ngJB6/Ome0H8ihzFeF3u3Q4KPk1wQIvUDNVN9hQA
uOLFH2Ja5uEUjJMKf4I7WVz+72egPrPknHKGqHwL6HKN/f98O3dXrn8Ri/s87Fq05BLVkgcqRfzU
9pbzSpyqfuDVgU1w8Ox5+lR0gZOGmyZ22xsImgee60AI9ABlpdEOUCCSYsqIGahGfu8Kt9O3aa41
ZAdUaLs2hdMIyQXlyl7/S9d1M9PMZ+9lp4RJEISBepHNJ1Gv5Jj4VxevYp5Cr98j3cV9FfuVYGBi
v7fIklhwPuJXyCKVgiqkJ4iewusO78CKPBCR/P6nHV6YW0Z1QOoiitQEP9JQ7Wwagzf0XSjjltye
bp/OOGUx70AA2mFs3uetNL5zP48VZf7VBaVY7uaFCsIcyZvpYY6sji5MLGQgQha6bnso8KvjZ3jz
x9l7Z9eBe5FmahOUCdnRXUuuUEgtXWxzcuU+w0V405c7ov1Jbr2z4T8gzr4jfmnIZTRTdz9o5oWD
eaoVZUy3MCozeV3Q7+VxqTCdaPWlmvojoBxd9EM7VmTbVYeMdYYvDTTqqdbbF+WrmZW26y1tcafq
pF/MBAFtnOv4nP5lmrIBAU07gX9olRNDPKj6yRji1/k9CXWYcCXyJx4eERzUjpcFUinpai3Sd9Dc
bKYAvJFILHUP2ryFPOz12eMO4S0ShAFAFbCEvQV4lYbBIoXBEZTgUnCIH+kTF+Yn1zxwkispppxb
3lMIocTaiWJ2nBRjb6Em1IL/64QuA2SNH3/6bdWZSxgVpdIyYzltZhLWWV+B6ZDOtHJIxtk/Vd64
Nt8ojuyQ+vgEGUqfgKbtuKt5kL2bvaSIUkqOKBq9vyBwUcrqmdO5LHbSS1BHAJxb7mXF3sRPMcsP
iJnwjdUSQthKPJkJA8oycEQdo0YUmeCSF9mPgZGrU64TT6cNfNB1ZeGr/l+QTwTqVFBbUjcytUEr
Tz4n4MWftXQT2rR4pJnHymaJ8yMjWnGYGQYRebmSbnNGYEF+0tZqgp2TkPk4RmiMetuBg4aqxKI+
iiEpmGBc2M4LkHITooW1uQvE0MG8qQsmOC5X73uKSEiMtVBtCooi1w12zGJonpkwxaCUPdHZkQDS
ktxA+QQib9ttrj2IdIUet5yttDTGs1KLKRFf5B+E7UGoFcDTalvOnKDX5wOAFuPNCFughP9VbCjg
0d8QwzB5O2jSZP6uuVAROfEY57FJBPFcaXuZjwM+KKpk3ShSaDsWHjaNTAvVHv9IXtPR6h91uiuQ
gsVFoQqIj6pl1zpyZ8zQb7sJZUoD9d1Hq8vwWiFnLciv9bWmip0UgvJjeDNISXnH5gxT9bvnwt6h
+g1cAhkrkvhR3O/B+SNqk3A6CPQTgpAhiR6/zK1I03lf391JeNEEa53a0j7jFfO3zVlJQ/7+X2LU
FyVNSmToCXvKTG+YS4MOy8AULqET7YsxLzaqc43bU9EAUJ2LRRccQNT17TPX9u7j0jGWtcaxGrSO
9SL0fw/hxwgb4eJMRXU3H430npFfvRr+uGA/lozuUPrqnW0+FJ5WtslLR1otiwiNeM18Tbjqxa2U
nkAtAUuV
`pragma protect end_protected
