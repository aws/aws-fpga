// Amazon FPGA Hardware Development Kit
//
// Copyright 2016 Amazon.com, Inc. or its affiliates. All Rights Reserved.
//
// Licensed under the Amazon Software License (the "License"). You may not use
// this file except in compliance with the License. A copy of the License is
// located at
//
//    http://aws.amazon.com/asl/
//
// or in the "license" file accompanying this file. This file is distributed on
// an "AS IS" BASIS, WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, express or
// implied. See the License for the specific language governing permissions and
// limitations under the License.

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
WD4cqsLxwd9r3EcBmWj21J7u3pfLl5ix1hxKOsX+8Fly2CiJuzxhcP0puwAvLCi7J3A6vbrwH+lx
DIdplgDKgtrRVcbBYEV91vEOACTWkhg11bzvOTb9rcERUlHt/nrP6BkrObDPtJ2gZPQbg/oF+Brc
H0kkulccaiAKljWw0sZjTXe8kp2eZY5rHL0QVt6Vq1YVW/Hv2z3ioHvD1jjQtUJGWRQIaW26N947
BtE9Yo55M3A+PuVaBnjKU7qx4N0c/U1xg6LFRUVdUKa41mPnIKbxdj4Ar9bBC3e+pRvHCMnFRuY4
Sua1C20HW9ps6+y3L8nvzwnrtGO1Tj2iy+1R1w==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
q5mnN4O1tyMZHoRCfmWS1SEL+rMhXnaektgZHRWjyU0Wu/MmfWiAaJAit7S5WvJQ7//tgukt+OTv
DPVBSrjpT0AC6p001aGCeo7iGnDmFEh8PMo6DFzW+8xNjpqx9OwzMx4XnaSRLV2Hfmv4ZyH2iNTt
O7NaDpoDT8wgCeSSB+w=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
MJa5wVAQIqAMogSSQmdrxDbK1RCpHEJjgAc7dXDQYX0xB8ZfMj51gc08VBVa6xJ1aOdWIQMvhk/o
L1EzTqLZnxkvXyRCltgR9di5CL161IeltHB+0FJta3SYrj4T3d1mDdLFAB6xhdXGgOgSVTRdwLMF
ExyN+EQ2j1lHInVtYLs=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3056)
`pragma protect data_block
fNVIapDv2eqbYuziazGRhpkUYihsc5akhGbU/+mopaxa13bFnUGRTbkUXemZ22nSS/ZZWSJ0bPDj
yfZIFFr08WuMKus0viH0y2JF1npEDiFAkz1rLvROMHUQ9BZcDVyzeTZJ9fpF6cCMJDPvpYBALfq5
FStnsz7GExcLZrGovGPphfYZq37GvccONu38gEEl/AsDnVYpy1m/Eu4gYbrVZCbJ0xVuSuN9W8xK
hCF04nhV54Ipmup+RHU9Jbn8py4yza6ErUC/SeZxtXcLTRzMxZLeTYWBZAlg2fgbH4F44HRYkm4f
1+kJmiCi7M7GlUfFmXIfA2t1ZFPSjGl2nr8lmJ6zmH1QArYCkzb0TKru1ZoUvsRE/+9UGQd1eZHK
cdWFIPEJvI42nkiuVvqk1LDp1TPvmmrGkX9DDi/gmJZWRIP26jfRGx8W4AlCnFt/u4ii+ZJsQvmh
d9JyUP5vFHCOK5McBzkUGiMDl/iENOeBSqURCAlSg3l/HglUlx8YiwWmSnRaEZcqe6tInA0uG9G5
EX90LS9aAmum9CnhyWBWNtdZmosMvN7FZP5KenOXtuMm6dDhB6/V4N7a8e1YHIYA82XBIQwPRLqf
SS0RRMf2RdPY/Jw2QB07Y/1mkVm7xvt2l96uRcErtsUBzzu/o2us6D0n6w5L3rtQGe3jh8z249k9
EPV8aa0VHy+iiYITmXZk3+w2traYVjZOzatWwqXJ44e+nipsKiqJbEJbDCfMFFPsKWxE98s0bYGw
0nIn1H7o81wDe1UmWQ2LY97RP8h9rkJ+luUdRguIlHJBOAheWyWOB1Kgc12d0ixt5rniGClPJFxd
0G90WThLuCMZ+7yU6r/jqX0CqrsIphliJojz7F2yX8zzRwQos/LA506eXQa064xJEOIck12BCJ6K
JK3p6/dmw6fHQe1Dnntm1qb9cuC6ZNIjrNWu82Dy2hYtJpfT7i4mWU/TNwtbc0tMTTvFiIrZEzkz
CsB56vnrHOtF75/V4qQXEv5ygl6tLxKplyo8JQSrMXbydGh621+WtLdndX6zV3STOqjm/hXvM5Ah
UeRkr4GwoIHnhxSvEBIvG3VCFWlfX3WGjZtwSV9OIscV2VfGutNJObWIJr9Q7OYPK39A0odnWTwW
pzu5gxcjIbo31ihDZ+S0FgvWCWNK4UJboYO42lyQJvybsepxtu6EUiUJqrBkn1dxiBORnoFgX3OE
cMrGf/xNlGb1jfKgqnaqvSMUSTfZ7gC5p9EnYsmV9heI/gzHwoKtjs0CorESuQfXCzVwqUAKY3Ei
hVC/5/RnlC3pTNkapbzfrO20yWqOFIh/6RxDMPGHAnX3ShGJ0hhgdITMVYfnD6p9gVNbnAKc3CQb
Hpz+zku0W8GP0/+tve07lB6y5R2ysn6kod/ZC88qWiMvGE/l7oFYKfRB4WuYnR3K0z4fq/nFVGFN
4fD20CSqkLwdZYCC94JazM0fIvfB27eLbwwY7ljz9HjHe9Ozd9of6Se2+8yaJMk9uZQh/+58C/uG
6p38DFGtOqTt0QCTX5iTZhRdXYfJBF1msO4ip8Lgzlc8EKx9qJlDH6gGsJ8PE5w8RYlhpp1glaSN
b44W1Xp7aPEun0Np10iQCMr0fMBo4e4c/6hVTwmd6UWneqFoOB1to3U3LJiXqlRv2zEdoEtrIztI
0vNRY02W6mWEaJqHYyMqHYy8qNAoHD+Gucz/vJds7vQrtM4BQ3pjvauClwFLkjDvgNFMndBusnPk
+3AI9v9BZxfxnNrqpkmQDL//ViN4TyfYMZ9GQsmfvhFNj8hyXAQdLN6sdMT4IrJ2gk7XFmNiuPsS
ibaDOJt/P6jUrbiibyArI5X7gymzX7MrW0VlTwhSSpXKilIP9/GSRNYBos0BYXQwN0PCFBC8IIKr
KbzYtxKEnhzIrWd1QXyPNbwmfIHRuA/BFxBLAj51Bq1D28LO1ZvZd/wggLmEQNxUYZff20877lQZ
xSH+slojYn+mfOB0D+iqzVIZ4yYwXAqzKgvBrSZyRW5o3YMZlfqTftYsbiwm0oEx72ctemNtzyOg
+0dEL9fKWnrmqAa3kACs/+AZJ1WMQS4IoExpgrD42Uf1Uug/esaA5SdDFlqNTot3NtwgYSyr2A32
fbj9QRmwDnXXYsdpAyHT863iA40LyhsxxtojIlgoYYL7eh/kRBwIbuB2IwvUWonVuJTJJcMmx8IO
CkczaKFMZi0/s1wO3d9OC+pzbzVG3QiZSxhKMnzOdnnbOZYNEpH8lROBZFFhi3GvIxfk8TuZlaRu
GHjWPYwsoBzY8RourCI2ix62fwqB8Nb4nxVwXJetNsrGRH+bsHBgiaHVKBog91sr8i9YllNpaThP
CIRaLecWP5V1jxcBS3t6sBCESOZ/rG/udg44Ywbmgg3fBBB/JVA2tHmq934oJBBytSFsKAPiVyHz
fbuNSR9oY2CVwkEL6VkxOG/TFSlfSqIL2GtGbC8gHlt3pDGrdpe35Lwkd2cBX/LX5TZr+EtBIQ8p
UHnRYOxDEj2zXzZO0RvsQcTJP/boldoSdikLXD/tHG8smnOuFHSaSfaHjqfQsA+IYe4OMS3Ms1Xp
Kp+wyZQFgVc5Vy+si/lqGGuCBWSoMLN2Ht6xzSBR15mUPsdgUvcq9H4aRpd4G9waD/Xmr8OdEUEm
jsYe/NwhCvLIuyk6m/Pz3Mlvi3AcZMlpU5j/qYebiM2Y0DdW39QwUwjUWWACyt9V6V07/06hW29O
jInej2fnK1ZXdoEhLnxTTIQdBGeVRksh/XHJgpTNhYGRAixpNMz/2gVxAJqFO1p0zcrXV0BUm3Cq
/3QRaw+UqTNnYLevryd1pb/xygNwgU1m44/ol6uHmDvapAQMk2SyT+G6aUbwu66tHa5cTU+W5be4
hqx2ux9yxsPBF48JwtH4xXPTQ4bCXdA0qwIVZJHfljIKZlmRPB08CDvKuxZcWwAfvXDNv8fbbQIO
ExAuovavi6RbBnDxZsIax6SQH5ziZq9ZmripHM/jef94+hca8xLroSd1kPB5N8on09eQB9zHscCi
uZP7mByzYEMMO3fL99YwjCviEqrRxqJ3k9R7czx1xuulWbqTeeVB98Ag0U6/rmRsB5wHIx+7aR06
Qn1wj5yg58n40+VKReANdRFIfBtMvmw9+C0jukvN4PS69w3qsZsxnI3c9GgWTVESXAZ/2MBMPfeV
VOymW4wD+jrGMdQMZfKEDf2NJF7QDRB4suIHsb7jx2rcT8S1INYAA43r956JINXeXg8gQaPcWDGl
orr0OZEeSac9pE+D8eDwuyffoIJjOcSchlD9HDi9rPROfipqeig7NmuwjBQiY+N8wIun8BzQwaTd
M1R7BkR2tQPknjTtsn3dv14oC/SqIBU4eEvSvv7FRy0Z1UOsF0P/vNKE1GMhwOPf8AX2uAb1Ff98
qsqyZnvhuIPg+q7K+KtCluTuhThDPPw9jhZtvYEQZEwjC3TL3rAR7Qauxbs216AS86DN1GYJ0wdf
cv2FPS7tL6xWfMDsgTUbGVQ5xsM0jxoC3TI0lGaOEBBXlIosdOlvaxBWcrD8hbsJQVJ1bpK/Z0DB
mUHmZkgDGs/ryUApgkva8gDTW3qhQnqFN+sebHHDuULLCbH7i/1s3TDzpZomSUUa23ZfoXeXQcUg
cqrg32v0Y2jvxIxaSYo38eTj/QuDig8qW9+x2lkt2MV8L39U7Pu0tDFhh6LsYPprktZMYrCV4p25
u6u99TMCh/vOkaiMfxTDdNziTRS7fEX1xNj6wAHIymGpmn50gpC4FmBPOgm/O9Yuk/o9VEjORGie
RXYRBquRdye+6w7NaOxnhqj3NxDVtFa/gOJDmjqRB6q0jA8SgVqIFcCnBVFRAiBFZojB+0+B+mg+
Ip/7wyWYx4mRWSjuVRTaBza4PD+moklpGhheWdUXTprA18VXooYfWqRSMQgTJQojk/V3w9RYfsvU
DPvucIakDh13YqG+GjdWsbdT6Er240TYregLfgcLDW8IH2BqAcHChy7VZHOQ2vWp7+b7wUAaMVxm
UhQK3QUqGSFNH2vnF6EnZYSEz93JbMgz5BmNazv/Zi/luyY=
`pragma protect end_protected
