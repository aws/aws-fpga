`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
o75dNfPUT7VVszdAv0/QqFM07Ag+zem9aPNYQhfDkRp+Bq4LgASdY4z9kNYxN/0Frl8wgCUI0/0D
PBo3zmeJqpSqMn7gHXbjc9WRyaEpK9gIoC0CT1UkcFlP8ZMLOPIPkQK8XriA/gFvnkE4k7n5zab+
14Apy9xYXGcbV07HW8bLm1ySfwDThU2DJO1JziU+dDOtt0qqf46FmpoTcG4njECfKpeacEJv+gY5
6mcG4QBR9SKvC9fFf3vnsaK0LvukcuAdYAuAE5qS2tbNLBopJ11VAqWzR0NBI1I65wlmeNfmKAzV
ifG6JVy1nZYRuVidbARfe+4aa1HUPTFj+bF00Q==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
cIHMttxe9nkhQREZxq/vMJToxhosF8JGfOXxyeYOsMuuJ6TmYl/sodr2gj0h5XOKKH2kuVf2ISpo
3QeiYGISi70ZpWr7VKQc+efVWsjqiM/As2NLZ1w4klkgqQwSpURWRZwUcd9o1c6ojuILOFe5FhZE
Savg6yuuXXJ3tTVOsbk=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
HLJqJcsqo2gn+xgTyoD8G+SeMEFSFoEBU0G/0U3JwOyaijfRPY9YXOAPIm5GIx40zGz8aA8zGRXd
7WJokTsJreuRNfVfEH/DbY61ogqCHder3Z5ofJrntOsHwcT0xoU/rgDSDB37dID5oIQY3VFdHKNI
6me6daI2uPhu5Z1IuIo=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4208)
`pragma protect data_block
UNmX+ZFuqrwIRIQH1PNqZ8hLj7te9tsudVGzGiw7WskV4pjU5vrFbdveybX9KbQcgiz2x7rQGdX1
SiW+wPOrtyoYzh7ebfI2tWpfnDi/j9tZW41FXab2k/PUKqmzGh648j3NYi1VVOnXHjW6VvNaxIIb
29Lbmo95MyMs4Znc1r87NvPPDUfYPXivtQ5C/MtCCc7r0xtIUbAIIJPebyaqIJ2SihPwxbr9AJ00
nvYVTQT0ZIIrf39UQCqupSx8DFzlbwKeFo10gPrlTk2FP/Uq6jbV6ybKNAPZ9o9pNS156SXx7g0K
fXNCIjjaEPoZ82N+a3/j6cfJMdX/JfaGyygdF0wHGMPSVpEkt1Z6L0keGYC8SDUynTh2Pf/AglIB
BKvGluwmQr1uo6Dfncq2faunYIbf9d1BjGdBppWXkiEMmDM7ym1SuGiQDkBm0eWgOlTqj7pn2fOg
8c7Kdc7nZRNf20SYnoIg8VN7KMkIFCM78MxIMuq6OfwfIzGnPHdIi+EuJvaV2Q0l29chXjHiinRQ
vGiFWkrmpEQYwVFWrcqvEIeNjxCVMkcnnfQSDWZmvO/RbaUyRtajz/UM/3H7D0E4uInj/LBN+F64
AqMY3443AXft4mRAoPzRp1RoqOtsCtN73rQY2wtUYYG2/nKDPA4hGA7/840yh9ji2V4H4kd9ULhU
BXLVJOxoYIgRS+6ExiA3YXa7WoFUskAZtARM20LvPKifw8LzP7BcYNC7v5wkAjU4pYOtqoJ2z+Za
ocaW3SffvG6c24i0t7fqdkMxXadd1yr+k8v9quuPQ3iLZL9s3rBHAy/Wxd0mjtoKxhwEVvkvUcn4
HXvgt0KfWM25kcUxHJc9qGIRrdDHL+3m3xnH3KuQRcby4ZzLhuzr0XKMfJFvT+3S0nC8b8fv6JAu
7paSjR0MSEE07S/o8WfF5ZGiPOyFUyHdwSd5LHwlVgHxpFc7ud45O2EgG38Eve/d6QOmMW4Pyl0q
oIS21aEEtQOpXP3+cxAsXaXMqCJPdoPuGrRh/3iywaLXAdpxSqgsLEz8kiyWoE61n+a4mMe0rGtC
7O6RvAk2TxABEIeF9bedWKnzciritMk87145uGnSclTBn5MVTAu+cH3WAoR8YSFtljwIRv5V9BDx
FK3VsEBaPJ4325JuR0BKoDC6lf8hxSSnmXUWVpIOEozuFL621phMVQhSR4Cx+bar7Fqm03ng9auA
vsFkcmRMWTgbhCSNyEhFO46wE4fWNPXNLMUgAl1RlTewmWxp/2TRvicG7W+nedVHjGYYRHeksOzr
lMOcji4sPxFdGFCIc8/EXVEqU03UkHtZs3QG9aCqKly8ql+WZMDhOCNMabjDgoKDdACFwhZk7Khh
DmuyAxnpSSpjLe4ecXsEEDej+/vdoySSnCzCXgLtF0sPBl/KH+65INwQplWuoJoiHN4fqGICOcLO
hwB+15/XyCRo37Bd76KX78iP0OmebyZ1wDr3n5N+aLcxoO8uT7fhQZl/wqhhswbAkt4byquqErXF
T1jfqr9TzlHTPChQVPSfItuL5YPEooMFWvuvUVtcW96DY64Qq6bemvIvdluMxPZJ/bk6XBMgFE8S
BF1AY+/vTtwArqVkEpfIW/xxbmCtV4ydke8+qTecq7qCG+QiKVGp1PkEuowUDDagG7PjDTTxCwYs
taXnZF2jM22ajt/d8lie9r+1jFB6agdDtKJU3/eqoKohfYmTMjM9Xo+iBFcEqQXqyXB3VO78YqiW
SvNfZSXQbcnwzs52DJKks/Myclx6sGnaay9SPtX6eUjKbmT8CCNi+cLx3jZcHvzd+S5hESvc2zUB
vCJbsJbxAbF+RBstFOk5bpD7QIbk8SegpAOKeUIwwHD+8oe9FXcEpipvj6cQTa8yJt8WVrzYkc9V
xkkA7LihqRgIL6viIVYRns4n0IhSzcwy8GXC4+5WjW0nNoYjtAPyKmZaspF5GmR++reOuzzqH+db
kBFDCVjQEW7Je4s2z8zcHQSHeYXrNQ1+iIQrY/8Z8jNNM6uraYX1g24ndTZvSQUNKN8dADIah7lI
nBOwq5N8KdSYmrwfxfmNyD79ZQs+SST7WKlvLvkg8rY3cS0PXDKH7nyvcmB9UTmQbPxoAYVs5iBC
0nYGr6e6nycs5MWaaTeeeaMwDUQSy9ZsPqXgWgD9Nk3VOOzLmxVSF+84hbUMcXeCQFg02bNl5MmO
LlEsiu3wECEnDgnh+vXWzAcOYJPjxDS9DiaU8ZKhEf6USlNXNTRq+E3QCS3CpkDtA+tNjVdPlupk
snfqnWa2evAlVGPLnAI1fduxC5Uf4ixrufYjs9ZyYgYnXj5aLhQBuw3Qkc1PBJ21evK31bzUui2p
OlBwJtggS8dJ36EXdvKRDWYHzeR9ypTXw1T6ntkRJn6/Bmjp3xT44fWD5rSaCQXA5xS3danzdCtu
5ePbD+go8fdbX+LamFPNVhL4N0o9xeF4VQNHVOrd90Z0RA7kcoypdS3jbMlYHw2tgh+F0ErBtVQr
2Tj4VMRMr8yA9bNQhyo+kww2jsh0vMvPJjFe+klhi7VcyeEfibG7lrTzis9AKEkEah7+qkH0HB/R
U8IOu+xFGKyKvhbIqpxBK2RcDkW9jVmvIq0U9g2HloqOX9DrTV9eV2BkgGpbx9s4U/RZhbMFaGPQ
WTe46Jxtt0fdAf6wXygs6pKRG0GMd3OpspzGpSRoncZcD7fpfx411a1ZJIIdzXbhLbJKT5fkSyC4
tNuLHdTqZg35cXTWomyqUgnzhgxLS/V8pUrZAxasOKAKMCm/70sncHjYaCItsrkV/kBwYkkYPPSH
aOMcvIt8BPvBMFeALP0yx7n56lKIMCZIOSlsL8yXRXL2dONF1KRqshwS/vkaT1zpdc2g0ow7V8s3
szg/qHYR8yI4IEb3j9f0demTc7YVBgYiqwNrE0AB/eMpXhtSpvVCF/qo/zSRj1Dl7XJN2SxXzNAX
5IyfgHw3+7QGZ0X8clUdiLgHvbXUfIPlP1fOwBpWP8Bgw5PzsgWxLCPDD+jGumccrpWC4bqqffxi
TdmpLruP2KdHhAT1i4V8dOnmbKM+aDiFX4pi/Xj9PX7JAf7NKMocAZc979SL581ilzUHngr8pb2V
YY24mOoUfGQf9viSJXt2zn8Cjj9ZW5DscaQuy4IDjZsiCnrv0pzp1LKzfoE4YtqnYmnVHPhqdRb2
cv9iMbKzXx19BKZGxFDHFKCfKN20jq+crUuiiGQ7U3WI8jKDLnG6ghaaveVzdFdgKijILypO8pdO
w+LsOYbgrAykhF0QORMEDOcguk7qSHHiGvKv3wM6JxzODN8FxXGyD8kI5+QhPTvDzGi1WF84nERU
WBziErteU7KZ+pQ5VyyfnViCEjmxJRoe2grq04q4hkX4hSlQBdoj16oqiXqTDPudRqXcfQj6rgVz
QY2d2dYWp4fl0Ccr7+6Pk0HWPW41iFqlYdvkXHvquagZrfFAIcBHzGtu6uOSLPmTPjAx8M/bZaNF
3i4i15OMd2m+Wgpn5nY4BDPezqGcl1k0FR1jd/ij8ciF4z9Dz0jjDZPRHs21to5xG5Zmbz63Z55N
U9oSv3Hm7oOelMOrwp3j7sFtRxuur73Q9H3RhOC+5ewxTd2qSTU9B5t24VXKUIsVGBIMeBxS5bhZ
6I+UWwkWaPDUS1rlHSDETQTJ7tMcU3oiPQw6qs6KpLVhhQWTG0MoC8cMnwFKeMaMBk6f6WfGN6pw
i34hoeb/hK3U8DruRvvIvqNKY4CScOi2qiSTRLrCH10vdiC9U+DtAxUefkc6ik1F0btVDimE2wWg
UnI2onjW/MgRz8oA9jepgQo91ah5Jw8HMZ5SyirXk4qMiRDZZrlEzS0r5F+OheT+GT1gnrUUUzJ1
h+GbVkQ7ZhX1Y9OojUGnL84H3Y4WvluQquty538KmGcpr5rnh8XK+sqVpjb2E9XKC8q2A2LNGuUV
lr+bR6SHiBk+NtbmJYZvPaXJbmR94M6qq2DFl4Xzl3ZVFDYGqk6X2XoYIZmW/vnARjq4ZSoSK4XB
I9yOYxN0t0/4ZlQQFFJUrk7/W8XYvwX3mHN29UgGy2wAdsRoOcVJwEbYwtymwEBNKZjPa+GwLJ9n
gsnzGVOeDB9bSofkw5RgJoogiMORZQBODi2xjgbamFK65szgP5wvtw1DONBdbM8sgW1hBYIZv1aQ
hi3LG8g3nChFEyQC5RPvQdzPM1QOPtpHCuD6c6j+VN3HDSB4SUIg9iG5fDgBG7Aa2gZkUYKXjee6
XVbf0DJmuxG+CaiaIMf/K/tCHu+oMm2mYRFM1TqXrXj3UQmL5sNAYrYyH8GwMM0TxkAv5W18m98e
yxpUvHRPWE4ZUhaEZFG/a81173bOirLjZUFR05JwMohWIpWHQyf2ix7lmO8HihHAG0wd1hgqz0P8
OxNmvYxjiQ80gRoPKvQOCP/FBynFqKciKI/GOCYRP3nlL4rT4betkEFwd1TgAdydr0SVzXHkfLop
wP4tsz0A0Nz2XOZ47lqSrpBJiNRLdV9AM0M7y1rVuQvnZh6HVaVyfCCM/ncuZL2RlIahENO5f0qb
FnjQzmWZFZi3m1h2AoyH/JpubnbeJHoMlCbYFgTKAOoLgGXSxJjD8ZXtXCYfhz1MyhJcpUQajPMP
O68t4b9V0KbnuCtFVjPk2rEfypZbkM10IToGAOIucroYuiVrMQs+01DT+9Bt475u+70atwiAaBkZ
PYmO/4jiaxxMNXTghhOxkNlLDXx+AZg+UHDWp+lgqJfd835kqJrzkg0Lf/QKEP5m/2ouFgC8rVb+
Yused+Wf6BtZ0kAgYjixp/eUhUbICZmCI0fv+5hEThpZUH2IeEa+QNQL6rmoytTnGtkJkxwpwa1g
p7kw8cz4nHjLrnfToN8qv304QeH7vtRmY4DqGeUGgMKddQY/fN/YR3qyNC+O1rYW2IfOOCxx96ft
XtNhpyOgRJfthoKNtz2qkqrxiTu9AX+IfAAIP9oDaeZ2YzYdKo2D9aCFRO3UNr8Q8jSIWwEFqEY9
5DjiQyMPCqfNM5C/TBmyqCn6waEtyLBtMFA1DReYe/RqJ94w2p80G7rVunOAHHVm25Kz+JZTm6HS
t+A6WIn/AuJzKht6nJT4pBX7mU3amKqSrCXqtykCdAX/qbk0ttYqFZ5geBLWLR9BSZs8YU1jWjo/
smGSDdUd6ifjRReFhezE9OaI4RqE51+d0PiS/MvhxL2OCoyba6qNV6TDvTPDwbmBH/Gz6COqE8hR
H75tcUcNmK2touDpHnaH85469Ng+eaekSR6zT1NB3RVQHD7F5jVBqvSMyzE32rxcGaJtg4Ji5Y4R
3nSGo/isOueiYvH3bzxyYzzty6pL98Fgh1wf9Kl84RFIDgNiv502TRVAzKIG1Uz1g8ITuWVS3TqM
XXffaLRwPr1rS5ak13JaSjZz1argT3N8lzOoRjaDBgffzFRUpaoDyWk0+UkVzZz/B0b7u26KYbF0
VaHePlw9YkjPW+IZSfjjNuX6aMBZp+nYWhJU+/kzGJR9Sq1pQb8XUZDKjBu8HAuR7mcZXwL8U1Iw
PX+hm5ni55YOuDJ2eX9AOGpVJ8dYlmAXzSUH518KnoW0MIRIBxpxnkfhwHF3gFA=
`pragma protect end_protected
