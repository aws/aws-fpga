`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
JSkKVWRpHf3ntDjy3iVx21OgsA3lb33jQqR8cALPi45MRFbhME5iASao4ihDr0+9N721Xbk+WwiI
0owy1gdbXtMRKi2Lzi2Jbnk/EDNSmh14Vn6wJe4F+LYgGsSZOEY88VqqOZBp1jgrmTIZiujaqTD/
KWtVCtzlkUGCO2sK77Ccz8pQPVsBgXrym3hrTeKzH13bxD8MEp+b/3XhSgJIvo6lli9LcivCmAUq
z38UOLfDM9ZcpePBpKFn32ZZu/PK2rGdvLMAtiymetJATj6ki/HozPj7WQ7YvO5u6hOnZFFRCrhH
RfzKqkmE0Kfo+JL1hJLg2h1mXUV7ehd1dqsXTw==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
Ek0mADiNpb1/sFVJLrwMFnJf+fn/q5RGJ/+eCBCr8EFLnfm17Mm0tRmXgwaJafrF3ffh+KKP13/7
3+7IbGhuM0QqM6gYLILEsCaS+tzCwxYtn/CdopDCcOsvfrvHXY7PDeHZq6V4KGeiH+6Abzi+VvbF
TGbavIdXRDAPEE0TnIY=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
kLG1AV5VPq3/AVc7+0+zwmrcg9P7+Az8BLLlYlXEgTaFrGuFLupxw38eBn+GOZvLsg/2b5m1xF6P
x2aVALPsyNkTYkY/9eMWbGOpppFtG7wTmZKhOCi1DnGGXZSeC+m0lf6F/g3g6RU0vGaz6YqyGTls
gtJ/UcJHGjMFylGeX7Q=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3504)
`pragma protect data_block
axysK5j6P9etuFktvLJjdqUCKvjTc//rciOa7vsM3ZvLmebUMcO0eC8/amgJMVLVy+3cWvm0N3r5
eChMjjjtwY3gyDU2Za5UN5RJLwMpA+mMnvt1q6U4IbPq47EiKeKRK5nWN50Xri1FgIh+yFUTUJJT
eY1aXk2wjTvhNgNbNg5YtTrm8MWvONshUpB0M0AuaerkBrvVeMt0Ew3dEQ9vqKDx8aNdktFCKefw
NxK+6myzOntj9dBlbUOS81FqOHStnKX1knok6h23X+Sr2pdYimNgNPZl83/b6Iw55q/+j0FdkfZV
pt8X4O5JVLZya7jS3nXaYgChmAlLMLkERnS1kQZU2nYfi3yWkQFIoWIS6J4SM9UElK7XvARozCSY
hecfUKkpkNY5STnE7g4CLVzGLVkKKuMENu+xECe7CPxz0xDh7X8teIJg5OGBzXdbNmDfoeVT/fPB
ayhOWSO1iczaSngf0osONGANHptCR1q+QTZwlZj2gdhHzl2qMOG/tZ3QiCLuB5+jodwUHNCQelVX
3+fPQ0G6ejnBVrcKXXO24FtOr7xuZSoBMa1x2BOljZF78HZJTfWU11fY+FA8OTCbGXG2svNAJsJR
HpLfvoOEgyyafDD3mxUvzJQ4zr9vUpD6128/Tq9vqATBF3cH9Q5cs+empHGbDfO81miEmx1AvdhN
giMNJXWxzXJx34Pv57raU3iQMEV39O/gh/UAI1O1eZT2vqrNXs6AytwsIhoFXO5F2U5OQ/1dEjOv
69hxEG9aR1+6NFJGpdtkidTXAn5sNia5j8Kgs7/8zho6p/8hcam9kKnBfDIBx9VSgSIUhK7Wu/da
VfiaqXZgHr3OFfXOVK/bwJgFg/HtHNlBrUss1zhq3kNEfGP1F05y496bLQq5bc7GHcYPzXHlC8Ze
WLqTVxwgJaFyc5XXpmJCnNFfcwktmNw1ov+nxCuOhtetfJSoj2cuQ/H7sE5oJLQFFe/Y7dGcyAcp
N+3iFgsL5QC781aTdLbZxjX9vVryTPu+XWlv//vi4aaEAM+qn5yQ8kSLYP6lkr6NDMgal0JnoK2M
rV8r4TEMokA8YvD9VUN+avpn7FZrJ+Le1jdwzuLevQztEgEpfn22jhFbMNtozoHjIRagyxoYZIf0
2+dXpC8RYZ9/Zm2LwgNkJjGZ8vSrcxU2BRMCvVDZb8QA1EvapXQFCe3npUxZ+hUd9tBvaHxc2Gf1
4Udpv4dUv2WagoJc1sEvym7f95+965BScoPA49fysrI/N9CNTbRWNTJNckNf1uyVKnr7VFo1E5Ts
SfqtKUGEj+BcL2oQWLc1Kl0uouwBuVDSJElJepbHCa/bnBC16F7c66026blgNKsiaiLwt/zeoY5Z
vJRFjAlyMvh6R73z+Rn/MvKVM3GDw3C3FtzLqm7k0e20vYb88Ru/aefyjj9f6CXyTaJrNbrTnywW
VmrvJDmkQKsvVEjAI49FAbARBYqQEyJfWb31pw8WieyiPS5fTOlSz0C2WKT1A9Uz5d7ZRq3s+6ZX
61bE+HwN2jiKG6+qYZ5ARYgQl9G9YTqHfVWvkiUOa/ilLxwV6wRDQmTvK6OKADxqS6jFdeLctlpP
UubpefdwCiw7MiEVll53+8VpBIo0DMssmNf2Xx2TiBXhH3sng++tg55z/5iaNJ5j8V8ldjiSdf+E
S9BzCfH1ZOpmpROSmMmmflBYlJQWKbI35+t+AdGDak8HRwcNRLJqJTmVO+hBGTItoLdyZEnA1jAD
eytEhBi+JLtB1pHkOl0anYshs8b8vAczg1jq6bB9rFda1J6kxvFl70+bvXUfG0o9aIfJrmMQ1a6S
rb9Mlm/hN4gzlaRJYRN3rtOlFhMaCi8w+wlBIndESYOwLeUuAmwL06Fy+C7dyZaY3UUD83CTECW3
h+le65bvlse397A4F78k8rPc0KjPfEqx763iZk+PVCbzRG7G9hnFS3K+FWjcRVBCZ48l5h7YF7P9
rhq0MC1AO2SVWuNW52e+KeID9RCx7AGtANzDk1InsvHH8WRjPiAmq2m4WVlpklqFnUYrLHsV5iFh
pvxu5LbEsSfFyw3r2j51UzQwjB/6mhoOOjqUK0tHPpkA3k/sMoOGBa+qzWLdMRFJsVV+qK/lyKTQ
zpGxgdRkBDS8IYDE/DCYnHMKO4D0KR6cNybox7TUdzHc23DQC2xmkHio0FfI0rWZ4ViIk93XXaJw
YVMQxw/SQBkPj46bPUMKJ1SNKAh3Y20QdvWw/I31a8reYSzSLdTaB4613iJz6UDLqezhsx39pSes
HvgSuhvKaF1Wx6LBAUK/6OUgd8sqfkvI1THicq+t9bFmua566FlgdfcgGkSzFKFVZChLLmNpRkRm
kEC1GCIo2PBRzkVwnoth7ugWU8Appup6k4Mp7g2yqV1PvfUIKkdo2lLEwBuwtvaIg2y0QnCN6iKK
sgAVfVh3iJwAxR43BKfYBMJoGlunzocmP7dsNOPi9TWjwGmAdkmgacXZ/BfbAFSiASl1PAy6xcV9
8e0koDP3ily0cWh1SHEP2XgrAFQJV9vx/h9mh0Gu2ZgcMKpw559wN2ETVW+dpFVPCvlOGnmcL1T9
Dde7keHEbmSF6HKRvVjAWQAWbMlUt03oYakVHk1Bt0/l4P3rTaPSD4yqaTj0HN5WylFWKM2dwlDe
jYmpn+TkQaFvBKjW0zqDAo9H0DjbIsudQdpKDa+XHlCJEq7XzKWA9mouH3+jbGH4Sd+gl2DPcH5I
UrGRjqsZmspXoqK7R/9AA36nzSKY2HSmZaNcfSgvcHdpMNYb8dXG1QIUaSinAJB5XA4uEEMLbJ74
j8v+OC/Hb3UI05Ut3jcl7y7u/JdtBYH1YRyZGNp6u3+WdW3bg/0ktaC7HtkeF6J6BAKAX7YBqXkk
0OVTyCfHQbNuiLvDWzkbO6zzMi/wT6BOCChsARyuU8KQ5ydhF37pjZz65g2bTnrYNMzZfGqvU6En
Z43xzn0T+xOT70C/a5g0Tmwb9EIsioSo8AnI0iwns8l8ZqrywbWSbEH3vlcupVlcSW+X1SYzRD6X
TC3v9r1FXTH0DzhP2tzVPdWFmAmZpJAcXvpVcRHRHAFsL67wdvRS6e+5PsgUsjMOnAB4I3zPBOjc
ZN/tZXDizMFQ9bdCiJQG/hcRqeUqUjS8CD/45d09awEGtgvQSVbNJ9nDrZQLdwgfp/Witr5WDo2z
caSOXyZxKdcJbX5J/uapPcVzNQpZ0r7e4RjkLUtxyplV1ZjnXjYzEww958UlegmI/f1CmFWNYtc/
O70gqUYbAQutFiuWYhLCMwuldAoeiMxR2XLypWLQ+PKe5LwaM+TJRrDMt2h0/DH2ap8VuHhHoRMz
79neediNCl/VDg6QhMJFN3Z+8eJhvYOoXI865ShggHy1TGKnaDKuxpiqhSXad0VvDvo7Cd/24FKC
R5knvphzSHcN8Wv4IPUKTvMt8m4uzjjKs5S3FdeZdgyrjBEVJ2euky8HiHL/TXypiWHuWzM+chZJ
53ba1sUgdI868lxzgZYflNYzcRfAj/xiOLymIMfhZPN5Ol+27lLuq7UHrG8n9ykPStdfUoT9A05J
J2vLCfwH49nh+y1kMWohb3a3n9BCXjmsUFnne/zRhlVmHSlIAa65nt11ZlsBoLVTKwp+KIA/AHna
w0A7E70r2++J4u+pa+WJVPQgaFG/naRlZj1xwVykR0G5wug9p1ALOQexZ7dw3PXnTN/bw/6t6g5K
BanznWKnUN2HUypCaV87JCWwsw8gr4s+90OAhQBwLPk4bj/8u1cYcyyUX/hgU4EZd1+D0/GFMEaa
d1/P/hgYHc53Ld/focCcinOgI5BxVXuhMLAAQOJnoc0dfAMFk5kXjOZ4qMChBJQmFblK23EsaQmZ
C/r2hFK2BsCYtdxqZrbcQxO9rFdSLd03eNUkraP2+vgEU43No+gLcp+0KRxJ3A9VOCpO797sUves
bfuynLzu6C39lfjxw+bRMYE7bHbnifH6l0UHBLMKghTWGqFajdcScyVqEYxnYHmrGoXToN/Z5KSR
zsg3/26pPZRpRHW1acZDGv0hrK+wcId/i+2SS8CQhU4bg/r9yLg6fW3lBSrdv+TWQkROXK98jMGs
5xinBkh0SxK+9cRC86jKJgDrM6dBv6OdLErUFGlzT2rDl+3ZHsyAOpnW3+SayzQigXDdF9upc0Mn
OCejzzAxutC/P7pRE2aB5JTmMhDslaSnz5UCO1A9ptbjK8Jn18Tw+7Ve63Z0pa2dEXW32oudx7ci
7bFnN+TW8IgMSVd5MeIbLiDwG3RZpLr+x4oDYfQyAgoiSxkzRJkeJUDC4+uD8ExLuttpBLl9xTxT
DQXoXPJ4iNfPcKlS2u7BRJg2txROHOAMxOXSPXnnbUGJ9rdAf0HdNUBoaV1MhOEYcl7Y/9o6/VR6
KlUPa2wJtX+x9SvkObxIRzKoBwvwSlh/t0Ke1cLOEjSgiwnMaVqlsWfmWJASgrirTQuA4ekqlz6w
Vnw2XnZEpVQzZqzca2v1sWglczoG4flgK7fDeGS+stEarcqXwwoee6t348NTfU1r7nP3mEuPweId
onl0iDcQF4tlxZ2Z1XMRm9QeV6KVzN82Gf5DIrpEUke6YsD/D7SrFPxd8p+VxJ/onfoI4TmHFuh0
2PMvog+ZlbnLDwb/cvlLvTmACI6H0mfCS5sZ
`pragma protect end_protected
