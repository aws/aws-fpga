`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect begin_commonblock
`pragma protect control error_handling="delegated"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa", key_block
XOSV9Zyuh5CgCA1eUygl/ZPxm53IXEGUuKhkjzO12LeYWxifAMVlUCedjWchJETRlBnZKb7rSTfN
EV5c2Y5h/QYKxGQ3lhGTFLQCKfyG/SF5NhR+jebgrCXOJY1DFiznjEMs1Yv+LBLkPzlurUI5reVR
IFVGXQNT9ATuOM4OgTwTpvQCl4dsRgO4VXXd4OGlfOUkBOJJ53V1BVB5y0dwpCyE1zajbTgi7US9
3K0JauCxjoXn8fLHk6yyzcATX8IuM5Bs4cHWQTtWYZMdVv0wHZpGnofqIIENwtN75Rl97KkcdQLR
W1jGpdPBpmTQM77ZLIEE2mWOkgMGK81EI3eAuQ==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect end_toolblock="Fg/4nE7Y6AGTmyh0ZvJpehhGsi8nKfEmuTLRQjwj3Ds="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3488)
`pragma protect data_block
kVJ8A3pS+ok+ycgnexS4nr6WZC6fVOoG5MVgP0IvIeg9WFXFLBymjIan9phGiC7FU8Kd5YzWOH8I
ghpJ6hcA3dem58zTXRUGz3EOaM9mBH3aomoEf+lz4PZJaJeHmMkOKBl2ryyW2aESilJP5JXpuzOo
h/ivHXUFg+TbYA8hQ2cFP0r7inut4RSEaBdAPUOtB6qrF3z7L5lHNps1xhqwbVKPLwxow5q6Vky0
Szxkz2YbyNJw9MeDs9AdG0jJvPtqp+OVwgBNy4Zlb46gSfKw24URzdYChmqlSAfttiU8q1+gXu1z
kCs2fYcCdBuDl/Z+fGduTVrbs6zf7BLpQGXPiA3lAUsHixSwUQLG8Zi/s+evo9xtzcTOTrW+mG4A
ikEbt2FENtwsFc4vfP6Qub8IF9nF9ShBdYX/i19eSyCf+y3r2tbJnRLOHVnJa22yGTuMgrPMTyce
92FOadQCIETKdPJQCsWTvNobvP1WwmeWP+ocUoGh4Son+I0ZjmFPII2uwzgfi86PWe8Ak9tGukHo
jDuA/hg9Y8Xpss5sz95S1At6Io3X4S8tOYlgMp/ypf+X+qTBm3un1Umh+bfCkTk2rt/Ur5VGplRi
c238hQtYh6tkpox1itcLwdkLTkWJWINBGaHQN/fTpMnAOGGhtCllG9wyGFWNNNp7zl1dsQuyK+DS
4EFRjlxBhe7diyfv2WQN5WIhekWjD5ieKve7TrOsZGitwML4ZPUEAieuCFRdedPSzIqcO8kOFfxh
XdOZKjkUZzQBKHoyJxa3wpQMlo+mr9VnxaOaIBW4orXVh0uZ7/mAgcNlFRxh1S09ngEJhqYUUU2W
rhsd6iDojR/+sP4twNTRkI7A/R/qNyBmNCR+uZy7/9QIYOctKozbG0NbVmHx0zyt12uy7fiViTii
YEPp8ol9SvAVnfDgiy1ojPQn1DobGn5a9IROa28UIvZnUvX2gEPe0dtLrrGCppylDOn+XMyv4X2j
UN6TZ7IZd1eLPuU1PfgmdRw4KhRBzMBTCdD2tGTac4wF9TQo1gfQCSC/tkxHvrIPQtfdc7jukclj
RZmDbDpjc8qTw10gpI3p9vXiPJGizaq/fEcKowVVayfz9NzWIuUWwSDGV9SISjQGKxAWO61u7DbR
hv1MNdihZPscWiw7WOUDySttS+Nt8u2cbhy8AWjNkGzCJxi52MGaA48ug30VhCLHcR7IvEe6yhIU
WF2gnn1MjkghXovzkcXqGphuCNvwVo3Gy+BupLvCnx8nFKJs6ZHIKdpwwrxfXHNLvRRLEyQY8dHu
Rv96skzibxI4WWfpHaTwSaH05s/3lW6u1GHaNAct42tULeY3JmanwX1A12Eq6b8PPM5lXPlY/Z90
kqarOWp9d5cJ5TOuoUY+sd5MR9SgZBYVh2b03bFsAPXyTtD5kvNm+EYGOKSekVkpKjOj4WyhAl+X
eacIEAX8KMcehSRGjc8FgWI6hXywUxEaXvkI9VHO329OEuO51ZYFpNPb+J7yaBq/3e8ykEXd4wfO
Ypvxek1R1OwcFmX4v2GIri3j2Z7clwPyl4dxb+3XTuX1fMB1AhWtkM69B+BHLnxGYR/yenUqm5bz
LIV7eMdArC+/f6RpaTRi49D4tXDcID/S9Cwa+KTOquM8U+E2S2/V8VwHyoOXqz0+49G6XWxAnWeu
5/Owwvkse4+6xikJwI5zLbA9RVAMUpwDeao2KOq3tH8aeJJOmrO+3fwRibyNQ16VZtBpXhylQWO3
UXi4rj16uILliEwyNJf/0QGCT6A+rSOLVbUTGOM/g7lv3gOCjpWJmftu9MhnXSzfvE1JDI63N12G
T3zpEwRLvNIMLxjj0VIuuit6ElAjyCYmvVrOP0WqETqyr+T4rXwve9mPvnPrc50p0DE5/0KB2A+l
cu6/ExJc+cseZJCXJMTOmv5qE0JG1nIMSoNLe0xXLaZ2jvGpHnkwQFMLR0Io51scbqYwki/m64zn
9eMMg37yadd8K7P5iqughqQbCtkJ2n5iwq8/2nYZ6gnZcerb4y9SMhfPtYzn/Nl7o70j3Yzw6dB4
R2uhHl9b7jpoavs41ieQldw/iRgeOJ23bqV1tDcsUDKHyh+aXleGOGQv6HVN14be/D948GbY/i8M
K9fFs5H3QRB6k4BGEwCnBLrq0hjNsMZ+g+muFZ7pI1DutKQN1EAz6QdzeAwr0owGMBKR19D6UhNn
8gRkoEBVK1lPua9XAeBtdtnUyy1qf8dLA4o/qlDzBwQQDC+Wb1QJEI9yPicQUVuxdeF/onl6JTRX
DNIOEE7A7ORQYGOHraLHAoCcAcnXhBBUSd7mWf0ov2e6jPlav06Jc+2tk+MynFcOn9yzsCcMClBO
wWnzG7yFl2UMzV/jdkpGRzWK3KCHhcbE9Sh/m4Aq2eQQ4xbGwojPBeMLg0XnT0X2BHVpXVwo1Zmy
o9YzUxsjxrwAGjYsScBId3RRRBnIYRNutT5Ou4bIBA3c190TY/S8LPwrjEubzb7f6BSMBBWCrX/c
7LbLQqrsIhKrZYbfqgH1jjxgiW0Jj3sX5poMM8hizExA7xD8U6sHOvU1NgPm0Ikx5FtlOoFiPl8G
FMpKJwBdJVa7EPWX21FgJyzzVpT8YShLt2xOMx3jLu+sf8d5GoIvbaHYL1jSLauxqC965UNejI9a
0XYnUz0zB2SjpqIzvLyoNFk0don6CoOBve/r93mX2X8xc/WpVh1Ym5UQHgQyDOfDwY5Kz04kPML/
ljbe5kCLAGbSt3O0JCWEpDajYXYuoNN5dmp2TVWnCrHwU+99YeGwSbf6uqnb8n7gWGZdqio5XNac
Cu30/j1jlyE9RiPUSNALYaxkeUMAuR+3bVWf47x/TDTIZT+cx6yUZM2/zrkzWF+r7awUKSw8BzSj
od6a1EC1gWVpxekZWEK97gfvARQT7Li1TzX/XBbpF4/XroPhGRLgBwc7MAFdnWQcI0GCZg4AtU59
xtzC1d7n9QuG0XfMsbo/DixU+XF7t92tRKAS68CR5IecwQf6EktEgILbJbGgyL42g0NoI1EdOkB7
IkH1kR0BfQhTEodSPt1KVqOBXAy71i6QuMLHkxcchwdksWmTtl22iziwCKNZGiekJSY5UKaANx/q
pqD5ZprQp4gvLcPAhzJByiRx1kh06OQJgvx97VG0bwnBtoet49b0Z8NF1iRWVXtn4/hkkNZa73Ms
UDP42YAZgkMQgXLI/d1Ca6lWLaNDJK01jtOaZdUUtYLHVf+5L0MgdyuhZ1emafnXuZbKcP3kHvFC
CoR3tbFqJzHPheRE5UcVxFqg6TP9gl6AK2IrncRGDQryEJRPNgnayif8+jKox45H64U14Ipxc0G4
ZrNGAOSpyWr7gJqo0ZGNUBgTOVxC0/zOCtVK5mfwMb9CPUJIQjRFHp1syPzcH7oSoCxXJAc+szkF
QdoJns4qjKZqZLggHAzeBmeEAXlcz+MJCOhhaXU7147cHBO245rPf/3f2wJH1+8mNQAlTMlUvKhk
eoKkrDFRJBBbuptDL5OHtahBzJB0izWTq8B9e1QPiqkqRkNko7069rkFhX8vDqel9ofXx9BP02gH
XnyJcZkxEfMiPIy5OQf+sC1lpVfRiFJE91GG5YhSfOEdv9L73KR1uCIpsdQlAYdoAP0mC7u1LMqo
GXYL5HGxtbHsww0hPMitAazkbGmmqM1QY6pLsZnnHTEezhInLzwEKl1n9+M1KkNElr6qBbVXgrL2
SKbeljdzj3tRiLQv7r/GpBU0cqYr4gDdnvKcDSOgYulIgfv8HwQSe4KZhvYQ0T6pgJZG8meYXIo9
HRjNmAmagFMvx9rIimtiLohoHCI47erktOISMOYe9LKgg3HkC+2EeevIEhdN/fkEjY7waPJzSGlG
dOnGS7jFaSqCMHelVvbY/3dN5K9LY9pHNMa8GQ2U7rX+Ki4fMaCcXhVV68Eyqsli/haSi7pg1Il5
r5tW2uA5VrRGXkk7phSsuQo3Ws1jrenVdWtEv3tyQEvOSsHlxSjYkj1TXKQBLpkU7CI9IP5v38uK
mJ9lbzz8DHBFHqR21zwDMawYCU7zcsCrbbeI2l/xhzlqDAutuyRGb5X1Kfh/xv9t57Z8dMvsgd2W
/fZ2eLFw9ChWpZ8FnUYp9e+itbOJg+3T1f6oD92Em18wf5+vRv14kMEgNp9ixGLoRElc9WRvoCI4
52nvBVfMJv7pEW5JMICZUB/v41VyiN90bv0WYStxi4XxGdGRcydtyCAXeGg+YPlbA2zIofEaKodG
+D6ni5lZ+9FB2Y0aOsEXg4z18Ve3bT8lWgVUAqqKu2QKR1JHbQcI/T2FEB+ypY2ZgkD4WG1EPN+y
XIzIvhyPFvfPnPATX/EpbFDNzrZz2wqiA8tAh/hy7Us0dY1Di6IJi76C/5ZCtf5jQCPrCX0nc11p
12K4J/e/mgSDzjovzX423JSMSay81jO8emCPZTEBV15tNYI5YPHgdS4Vz7/HVkcMNgcGuwD+Tujx
MA6lAanqkXIDevx1gY+aSBRsDcJYeDmTAk0o/3+6tE5wmz4sByHJ0sp85huv+Y45j9SKhvGya1Cz
6zLiXF11WvNBo4G+QqqHDlRG3L7P03f1DlTBOieQT6+tVffAYHieInzIn6Z8edRWNP+3iQHVd637
xN5M7eSe/tXM0dE=
`pragma protect end_protected
