// Amazon FPGA Hardware Development Kit
//
// Copyright 2016 Amazon.com, Inc. or its affiliates. All Rights Reserved.
//
// Licensed under the Amazon Software License (the "License"). You may not use
// this file except in compliance with the License. A copy of the License is
// located at
//
// http://aws.amazon.com/asl/
//
// or in the "license" file accompanying this file. This file is distributed on
// an "AS IS" BASIS, WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, express or
// implied. See the License for the specific language governing permissions and
// limitations under the License.

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Wk+TXwj5EV/WssyuiUdklCfjGwgwlctZK7+eXb+Zomx92GBj14YwpMs3Ja3FNZquTm+e9HFiqJMR
JjfkRGWbjvXS39siyJrhjZ/mI60lWKQT92v6joY9xq8M7g02W1eaXy0sMrmuHYLzfWNKm34NPydw
m2je/zJSIAXNtG8u2HxnyvDq0HuhEEl5sRC/gcOnoucGuuq3idcHJ8GEe1RxnxyxlyA3kbaZX/5k
3M6S82ZK51HilfDnOw0/fA3uW1gmz8y6iEfB80ny40sPh8uATgWAqO5tfWrwZo7SXB23VpHEYd+c
0w/Qpq46nu4KPnlJgBMUuhGB7whCZtZ0SCuLag==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
wa4UU3lttpDAy8/C2U4p/rmSp+gMtVirTLBZY7avb0XBtm7gDjFBBWy56ZbEE0u+5LYxVlax2gRK
lzLd5hmfYnXBOA1jycaN6h32b1EXoyXPgRtU09J0ogCeuw09iXGojnieqCNirbbXue+FhrO60guW
3mbGLSWZrS9pV/fF7WQ=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
fCGhkObbgItruJPZ+8H/HNyXVfMuAKb9t3G6/P3gcCoA4dFGnRdUWId9sSpQqfP39vVg7IBWmQO6
2qwoQzHe8menskfo3PXY/Zm9XiC19ZYZC2zx8QSZmWybgPZUn9/hi04HkLbdmrshotL+woypwFNU
1Z8IfeU7DdWIXRcAiaU=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4208)
`pragma protect data_block
W2fYtfRJpK3r0sAA3xmahQsBwxW+9uhdtGnMs5UYbJMkPhL0EfmiNM7hfpGVEPngvE5aYshNXKbQ
ew3uvf39WXpv5fzPPrs/zEAhbfyRATWB2iK9SR19r5EHlBUSmQW0UtbzOayO2DMH2Nut+mXpG4bC
pt54YAbjEBBJ3ySO8ga5jukUsJbLmmUc4UDRBu7kfRdVGGS+R8kbiGj0OXTtElQHseZRzkru41jo
bJBZHPJz71YBISvY/Q3fvAGdYUJdnSWInoL4l2KDfZEKpQ6qAiqGy5bILZ4kT+kgdrXVhJwYb8Ft
YJ9IaOStG6ix29vOniQPVrikm+CKasCrEqqTF00yRcwJ+Dw3s0XD/xtQT5aJt85jeixosHFmGGnf
4oYIOrRgdx+psJ5SozDpndCNXOIVbeQTMLP+eM7JDrqjbHUEtOUdu6VAOU+0mHt5nC1m0UMtjWlj
h30i4aFYJ6agrg/kEgQZC2bNcIxnfAKXCDwVXYOBY7+R27OR/xqmZPpV1z7KCuAjmHbQUhPcsoK0
2nfWtZEyOAEZ+IFPvfrtpvpj5gSTpHDVOW39hQWtpTC9ReFFYSzRjrubcj8PmDJtfJzr+csHX6Tm
xq3YmipxIck1lUBs/AUU7yqXSnZip7TIq08+fOLHT4hpK/RWKH5VOB3fxing03EZ12ebYp9uNKtq
HMHLar342xddATYrlnm+L3nqGsbHUfvJTFw+KkxMrtjR/CMg6W9v52WLT4KpUvckuYEZBHi29urh
XMT7ETTwiXF4LTOFVeI0aeJXlMBWTiXQzCN6cdMlOvH00dUP1OrXHKqUi2sOmvs9/L6XvpYAAmzN
dzSMX4mMNWFCDCKIcyY7JczQbtnZgdAKF/NbslbgIZGAUz/nZddLwDWvaNbEjZX+SYS5gNJusO6b
V07WzUowI8UPzsFpE8Xp0/1SSb7+hnTv1bDpySRaAmRqBOOZaWEjLhWtpAVMmq2prAku18zVrVZt
rTsG7MCzw9q+yWOc7vYEuk70NF9/blrktwmlq8w2iMUhFoTwZB7aVK0mEhp90XSDmlRmipj86hja
0ngWKOEU2EvHCZH0/jWs5Vy5ufyR7zSkknUVynFyyCIf1WSyYg4x2B6LmMIrbQGx++kchGXUw+7M
R+YWjd8C9Gmq5UJhG5TYkw02TAMH0DIJHzfB84pTMsU70uVLM9fcv/fH0UngBFAxA1zRW95lkcJA
v8myNL3jyHeoUSa7/o/F5QXc7RvezV0fCvlTcjaS0uBv3cKGUuFUmjTG4R1zc4e3bs1zF5n010vQ
8qIrp6Sc2LZ7fH8y1svgxHlnLGNHiZYr91nQPStRSuVRgms8xL0we9hFIf6Qa7bllJjWoi3hnD8v
cJhd7f715X06bBjSi8tpSHHJtFZxqYRrMUOfTCqSMkJW+5tLlscnfchYEOr0AQhEr8CAJEFaRtvY
nmU0GH6U3ZI0zc1DxqQZAVwVb/JcEDmQ5k1kOfttudUQ5jNVfW7QbEG4P2rhyaf4cAH6GSAU5KAC
aTI05AnMO9ydbEp7ctbyFbEUxxnDug4mu4mMS10neOIIYINLanewHVAcOx5bGMwFU+xbxwz+janI
SXJQ85pnXB0dnfpnD9CpIcFRXINCZ4a6w5TTNdLiGj5Ey/ygKrAahiUccoP7iEhFTltkKpeadaJq
ExH0IiQo0GoxMa2G8LHJ0jJrGT/IF4ah1tC+/nBtB1Auzinz+fVoOqFHuj7BrxIGjwvQNQA4gcYG
BNUDKENUGbihXHZYQw0b8Agw+Im8tAhj2+mActS3fWmt5RFMGPqLeEYkjs9YeGsZuBhxhWOkCr8k
LAwzO0lcgQFDtV1KK5zD9o1sjE50Lv1CA+xEBEswXIrI5P36YeFQzh8lUTyS/VVl/UlPnTG7CObo
lEVCWhyaRN1Ofgs6THchMwOclt5Z4h6isGi8NEi+iNsJAaxtlxI/dUw24ugxO6tmg9VsvWfRKQi2
7k+TpCCLEOyK+euC/mKm5sWpIfFOvuyFIwSoZRAWE95htdbCq4zYhiS7nXkMoc7EuP7KA/Uxuv2y
HRvW5R2jFLDtabIPL2HUqjFSXUSwqzOIYmLoVwnoRaXNOoriAz0fb/+L+uSZTYcB3J/AzGFdgemx
8yfru7T+gxxI2drOQG2FCLFxmDY0t0NnLTSOInK6f0jZrdt6ViHJRG62PEh2DjC/HDJMqrDBuzLG
119wZ/86DLCMIF4zWBcebGvYNUXv5KGtZ70oWxqurHQ+NbjWlg+lEXY0+5k0aPgg/lHvD4Uhc7Kb
iuBkiELxcvXOUBOe9E+Vlgj7RuHbMSfCtMalmyTNcT8FrOm5CQPQQL68ViVXloGNXWY65vAvx/Af
0oOQrlShjChOJxty6r6NSmHHEhuun3OehiXWNJ9Vu3a2ryrrCtu0yVNrK8JZZIEZVRWPB+VZazKI
mM3rO8RXQSdQLGI1YoiU/z3HbcbYh/wKhz/qf3FLGz21+R5nlJful94NwgWfSBLxBWidN3ds0OUU
HG4P4z8A8EM4iUdBMIRtkCWQYM3m097rOO0vusWCuaWhpOv6fahxF6mZEkjidReIyvE06WKp3fmF
TIJF0G3nMSEY3ZX1zlXmoNgZaU2DfCjfiDccBj+f1w8amqyYAv3koNy0/sb+Dlyhh9B8RStIVizq
giDJ6fU6tc4nO0qusj+Wn6bcrZTysSdHgVzDT7XDWqNFauItPHd3qk3vwgw+848zCD5gfadE1gf1
07Sro61fTd4kjhe9ml2QaeAx+zKLPejA+ZU6IB6ptYB0Oye4gbn1AW5z6MWC2sNBZhwn+DR4Rbzo
cMzj6eIMFGdguRQTIn1cqMKNyb6kNdXYlEO4qn9CU0gL5tmzRWb28RPymIdL52xOCDxqXMhJc2Tx
nriQGtoysyfqWtPE5hEUD5/jbFAIU9/LtolxZjsgBIMQJySWWfREKaa4vcLGGZNKu7Chu+9hnN3v
z6x9KCTYOhEFz6Jg5sBm+BzrzNIZDuDO/9tPhVcXYbq/L+xzbLHzRyLfqGeUzpkfWIUHF8LQSQNQ
nevuQqg3Zw60w1o9ae+HdG9D5eRi0RW4e5SGJKSr4y40sUA2t9fYOY+cHm6uFHJtVpcoDLL4QS2G
1sccxO3ZUiX8qFPu/Pvgi/rVD7oEmy4DrUtKn1fhJRJZOvussjDN3EbUxt69gqPrJLfgO+VMd9F7
DQkwd0z+hCs/KCu+lzD+BZMjDMfPSWNjCuuc7ceVvpFBNFW5iKH0lLLv1TXMxNugF1vgmEIs+09z
x8BAhTz83O0NgOSD1IWHXH8LZhz0ND94ExsdwGEP+n4VuGwOxj98GkAA7DqRokk5VjCQW1+9OtcI
w8QJUx0GJ88c71XfU8vVOen4r8qS9NipRGBioHttUNjjERGwC8Ie7UIwP12q0PUYdZTZpRHZgXoh
lpbKjpM0UbNxbxojYKeFiTqGQBBCDWfeet7lwZ30ie3h8vEycs6Ge4zcYECaR3T1PQAXYFeO5XX7
b1HcXqQew78INwj8xF8ejrR5QutcSiL8PAOdKc0IDTb1MZTqNH9QfTV1yfi4v8YX6hoZTF4k5cfN
r7lbixvBXJvb+7XS7MWAU2WTdduZABP64nQqZ90vxxLCzXv1zvpyvDtl5QYktNYmnJSlfFLVdbAr
Y8VnMeeTOlMTWzdaHz40LVMW+j3Bb0+QlWlT+2r3MYbOdeY0i3TjCwx7z9F7MeAbT/HeziqAgReA
43cg8A4qt84He+3VR1sXtocrmlq4QcuaoU/8XzZnhUqYS1XBO30wGnx+uPhiMKvQuON8ha9Gxjn9
ARQW14ORjfR3Hu53DhPOVHoCqFg5K7PiUl6sc1ByntI7vYEYFiWz19U0Km0dPGebguzgFT8Qhul/
jWX+eAzdw4Xmvc4sLTJ1ijVpeGZpf3aRxQDZCo51O+IVdAS4spsM43ZLni5YSdAa9Y0hJ4/yS6YA
3GM2Ot2l3arC+UB8dYgrUtjCIGMlKBJCP44kXpld5ZVCZwE+2iAm0GpODocOzbCDqWHwUqu7p4y1
CVk/sTxNeyqGhQEuSrMSpcJ6sCYs+hLH84B0iG+FGFv99ftA98cAmdllx3gpWXq5/AtbtkB9DKMF
ORmOIM0TChJ2X0RT7OyAijuxoC5Il4RpvOC8N3GFnsstNHxjUFxfqiipWHZzKjUytP1igk+J8o2k
Aj5UhW86oz4heT2yopoAdFG1B8MMyFPb9onfX/yJLKMcu0mJp5nocjAkt01KPUzgGnGSPW1fJ1o3
P7wgx6HOLSe417Ru6zrJGWgfO43XPD0fAdKpF4ZfFIFc0+8FU3QefLCVoiSO8QtyHJF+q8Gg9Hr2
P7XbNtD06/Rd5F/vP99ALE6hLs3ULn5jKsPqZ65KmMHgTqJ0HF3pNL6BXUMEWQeTtxjXy5w7q0xf
MKN/O/nYbyjwfJEtdKwIArRYL2Fnc6HoaaeDFmAn2FKtbnrB2F97OGGr0Jikob8mftrcibbI/Ykj
qebkWWTvvihABFedthRjlbFBExeD2oxtnIEr6b2nI6jFoUvv9D4HjB3Wkr8tup63S/nQZVguKGho
CzGkDxH4jCGZ6vtP8ebQVur2R/fEN2ki62ip8N93b8Qds9maDuJ9vPrfHetdkeAp0oTyvS+puLOz
YM/AZH1H2bSpNh1z7vUGf27qiYiQy87jojsWuxESwXjMM76PbDbAFngIE0k20OhTvVx4QG/wV4J9
+lauUEqesw76+yUVurUUSaJKOpxvFBKL2zf/JgdjfR89iLHNIJH3lBrfBmjMc07vDNVZCRvSrit0
pmuwCdYcz3uAvVWCwjgrTbngM2LhGgbOIM5LfULWstXFjgnIQwPIve8KF3OTGsk96BBgU0P8J7fg
s8mOJomhI0wJd6Ka+BiNH0F4v1JaYetJda66WWdsijD/7yQxveotkhgymNQTeyZfU7uhizwxVQn3
AivvP6p4h0Ql9F7ymveDqsXH2aai/7YJ9mOlP5TFFIl9CUjugWgRyqSleevCLCh0MPTL8z1+Y3y8
sbgGgXozkHDYqgZpHK6/eV/ZqZi73HlsxExLT8TsNmTwrJkojpHv2VamfcuK+2tbty79BFZ43w05
9VOnZ5fG3GJdA9UdX4jPlmvbE0eFMkmbOyd0uAvDSqd+XmpucTIlZ6PuR9dzMKt/UhrZA4MmZr1e
Z7FJmSMPOX50qmLVjJ5w4NN3sBayDiTXGq7kq5NsSb67q0Z4kmtlXEh1m2852TBgg3Cb9/rOlty9
ycklRwqafIt0UucG6/8pv7lc/5sz4q1ARAABJnOEa7qtiplR6aycLbDfAsoZ8ZkzA8Rd/i38gVWr
Rzn/JheQxDxLjqVrZbyFo21g7vy6am+Q7Pxw4qcG6FKwpkUMsdpowuw7xisQRRr7pfWVMgkVW9fg
4D9+jOQytDT5aUXuOI3d23w84yMcERREKmmOUlJy0GU3OUWrFVnkML9kCoKrnWCDMDZ8JymW6iDM
mLgjBn8ST5RLfUW43ZI025U0M/5QW/qjjGpFpNYnqbPWmSRwO1zCWoHdMW6Pgfw1pJFSMBBXaTL0
QKFO/rDJYxXB4YT+tdmtwgtsGeMcBCkXGm2XMOgHI3pJj3qZo8McC77zt5wsa6k=
`pragma protect end_protected
