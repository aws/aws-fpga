`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
hpNJhWywMnWMisa+Mh3Hk1r5BXHMdVSh0OYE6eIJpLagjYqnktoIQVlqAyndjEp9deLoVyncf+xV
o+AzIxoNgI4RgnghmR4yeIp4IUbGAOGE7B7XGIIXiAL8iE6yLsPKtMka5pkTNK0GvvOaKCAbxk67
r+jIfOinbp2CpTJzUpJjnkw51dguI4EUV/i3uUTd7aDZp7EpmVPUES/WB49/aj/LiMflJ13g9kDS
7oGAYQEhXjNocfvKcT7az6BSXgcDjK6N/q3fY2peF7S+OA2TKR0CpwxtAK4BWoGvExxFP/lOejaj
V7nW/6mQEcR4YW6UCJbtheLRoMrz81GXU2A9xQ==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
AkA5EVZUWdOB15aWBFJCf4gQ12UIbcIT/EzOILNvmVM4SaUkPUz+llhMHUEanzg5713pp+h4jfve
lBA0c92MulMUKd5lFj/HgZM2REX+152sIgH7SHVVBGlqtTVT8n3OcQe66UN5ImuEn7qvdORZLDkH
jnUwMZ0+g31BjSgsmVw=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
BDfapU7EbOF+ouX1ZRJIUd57zfynMx7OC5V6GdRBJWBBDRGaTDO2G+JEo9wCKmY3S9+8b2PqcD76
PimDUWaspIBi7bMx+w3fWkTnn0A0/N499t/ErhFZ8NZ4MCzkZDHa8MiW9NsIAtGNK4fb3HPlhlEQ
Y2S/EKaN1Clgbdc6MUI=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 136816)
`pragma protect data_block
gACvrv76guV3D39jdREh4BSfCTfVX1JmBpP6r2b1ZKYkyow3WiBkvME5AM3HDIa3RjHnqdjY095N
zVCMRcZEZ8PjTQl6Pt68KA1mtf9HEIUtY6KnV/ZkJb55AS3XxHGWpdRDQe4WtCVADS9RiRfLTUrM
hni5IFm3M8ZSPv1VTb1Bbd7X64TprUXOmvxsR9bDyXy7GvAqj/CEjEeqa/gbrWlhha0dQxVxFdB/
RqvIsUz02hkPg/E7jwu8OrEsAdEQVas8eJnEjsdcaq2/W55lITXJpGch2gj6jeYkr71k9t7i2VBi
CliFBF4ltK8E65eWTEMosWT0xmR/U1k9mdH+ASENmgw+kib5kYG5ZHjV5vJzOxcg5Mlx+30l8akf
1ZeChY3wqeAVp7d2pRN3YSIS9gMY66o86G5BBl93XYQrcgYLI9ulM9brF/BiauNkW9IfWei3OFTM
UZKe6GaaEvJmYjfGpILFhOLX56pGVQBaxBY1yp03N0OyxchcP1fRWlT0kKiFYF/EBqKDjOq47S5d
bTaCBieXsZoVCkWb0nYQDV8MnloW6ndvhpUvJhpKok8M9zlg84LN7RAt9O7qXB297VbCjuHC1XTy
dNps1q+WDpG6ZRER7YSUhFJ76YK9CtkbEdxc/TTlkI/yMsI5EK18+xlRAbH6Btxe5pNynMyiWjJD
CIsEhp3a6fGjAuXmf3wOReU/l5sUi/UN3dLA/PvvtLln5VN+tJX3VMzGWEAGBa1u5gG3Tvv3mLBP
co1+jo+1byzfjGPqkdVE2Ko1GF/FEn+ye1tVvDZWyaSRxesq+bTG1vnmd64qZJzVDNzHT+OGTfrw
pNtK7j0ajsnyE3KSYdIegnqZNKLoRcSWqd9oIjfqZ6nEmzZjFMinlgN3ck4iMui1xehKm81dP+8U
y9ZqzAvtKQTLV8cAG0rlneawam50Ll/u6AwKRZiRbITXUW/SsquNspjIuaSe93f/bvQS0MB1dJ5r
tX0/bVok/d+0oswKAcW7UPAn1et0pFbGJz/XJLFExCgzt9icZir0+0j2ivCNmeBcvXussAYFg9gU
QFgJiYgWzXM/T8ObFQP8fTYfN8lDBWoh2TesIjLawZLW3nQW/jCNR6ESxwpivdbbA6jzXnPqsv/z
/ZVPX4NBX7Zu9D/Vn2Qiknrk0YPgk/pWUTikxNteYb2YEgi4Yf7zgzi2P0ge79kKy/tvpna4JT8g
sDcpz+PVbqcP8inBBVFpZXHAs2DENvFl35m6MRUQl2vlexUx40a4O9P/JLeboZJ0h4vouUMu/7op
R9fBy1ybjBPXa3N7UCgfbexqD4gvj/L8BKbNfeyedWswkN6qmzeQ6Z6/XJKaqbg4aa7/GY6yTFfJ
DRjkHb6kv2dkYZMwylQoZCfz6tNhtmLCxs5raQP987TX0oFevc+wM/swThKHMR6PMtu/3hy1L2JT
LQQ6iuyOW1PSCqXdQ1/xKsPB3+1UwwQ/aNJ9q6lqcr0ITEQNubeIJPIt1ocjVONVHx+lZAfHk54J
X69CrGFhI+dNj3YR0698/y4OMiMXwXUQzfjFvzHpZ15GWneFsy4QG77XgwlDu6BhdAyW7R/TO83i
TMqm2TPpRNF6vIxUATnUSUtu32SqpnfzxcTkaJAzWhewO+IQG0dcMxKg6TdBwHo7IT7ZJxryVsNl
xSZfM9h0oYkOp1HHgpOdYKcMBpuRfRUonfVwaVVyAgzNsWmPG4xMHs91F5yooRoqwDXSVw6nSWy9
k+lhLCtDowr3wZSRx8LEHLU/VCKMR0HO2tiyEEnBBAnyYc7StmCGegO83fwG8VKKGbRda90Z9u8r
ELzgz64G7D71PLGBQOXY84mqpPwZ6+YJN/9rPmKEGfiU38P3/WZ99RuV0RhBtg+GqIK6OLcQPBur
XKRAyrZ5NvVv2snEwR8kOkluBrUiX4yZIISmak7uFYRRlCQd6rOFIO38nqh222EEH7hT8WTz0Mwm
ouq3poBFWotwPYQc4ohD5cal1wtQEERZxRCgxYLYw/Z1LRzhhei6QLlr8bc2oxUgmOoXvtqFs3i0
nNxiElBJsmuwjTXa8oFLXR7MCqLnM83ukBoSoiIDUJVa3w+YNfrxyiUndXsoVfvNeOGsS3SyBzM1
Iadm2Eh2F831tXWeaiKEkRGiWrVccXTClfZuimZ74Q15+Dk4y9K/ifIUoO3GQ7NrTnMd3/p8q09V
KgJmYwVspJd71hfIOMYbLhVo1ggFH2lyzm+0zw1DA0abqsq8IKlex7/ecx/CADddduhkx5USzxwX
9IlN7PytKAQGka8f30FVR+3ZmQqkqqwPdPBR5KrhISC6HX5BJjSYXLTSP+BN3nzWoZcgoQl0zlT1
5exTMOnSXp2L+eGI21uk6kg+mMQDYVWSmDP8MWdzqYTtwO96e8eAR6Ak6lqxCvaMabhhcxujiKrE
Y4LEBgENuH0rk4yw7nLIQ81FFw/5RUnq57VUjhi0c/x/biJH5SRsjQqSlfx9Xkcs39Ceq1wq9EPK
U2ypGktUdgi2vbCc0U9E0UxWZvsL8bX3i3OaGcpY6fovBUeeG+YV9+KSJZcgzxuRojGFfH79Xhv2
0JiGl8YQieaZ9LkyVReO0A7n9N7dYxJOTYC+PFxuNee9cqCgzMaJdjHuw25HVJkGaBwC8QpObdlB
CoTfn26V2dLBHqrlu1ClxwN7JxipK7rwXfVxOEX8b5M5iNjlLmiop3pjD/3J+MuQkEJuZeKbeBrp
JLpYZmjJq5ov1DxGgOOmm8mPx4zVwZ3323HGTX5XNioHrVr+D0mS/x1YTwTHWLTWqVOccays+cgk
XC9uyWZuXZYFEz1CvZXYjoViUYQn8inhB5uk1t8kGAAsje6IzG6RgUx+sc62fjo1UCm05dLPl7EB
rJveFnmJyJrZSpQuyfo9wDnXZYqRHAbTSY/U4BcazKsnICrzkoZ4HTod3pKdnJ/7eBj2hnYxA+Fn
3onQAOvdBoEdd9bGJ2J9yjPXXnI6sMUNvwCLKPURqV59fqNsaRrhbXDYgsurOWhuQPL0hchMqKM5
rDnRIKQ3TBiltWCBlr6V0O6KIKDxnRqDSWCU/0oBSxvCDkjq0mixGSpv1M5CbQWxW4f3nfGFbpOF
cp946DynK4A7+gzWblvW9F6PMDT5xcl9nyvOgqK4um1A4C1j0l/+kYi65Zink+2gwDKxsmas/fRr
Ot+c0cL2UVtUZe8aR8o0bvSFmgmL9vRujq+5S7SLbdU97acWZ1eRs3lLMXfGSS0wYbDrFR/Z+c2r
jcU1SJiBzu2KsiP+82Bx7V0rV0l518UIcTtG7BMBYH5uPDQz8AUuYdSihqQ53cd9QMsZ8nDoapxe
ge6XCuTcO8txYJFJPSmI0nmKDbX8V7lLyrNk01l1XF1XmA2KQ0BVNssU6i5WeymLl0w3HRrikacu
J2ZmSAoF1viQ76EQ0CvmKQklKe6olwdbUr7NolMvv51HR0PYN18kJYFJjLi+F2xDGMCIWW44YYji
1hI65ASoEA2gY3eyAR8EDUit1KxQvp9KUPOuvGdbtG/xuFPFVAgFgXZJW+dQ2IkJDRWMxRHVuug7
0P1hJ/zMr+z83CVWrm7cZIUMCE281RMFNlz49Jj/xHqk3yyQqE0+HpzSSbkCDODS2mlL7QUsOdSY
4looiQ/DDKmxVzGZRJTiAgsnMXLDpSGbd/cA4rr13Mxn8t6g4gah19J+0h8ghdiIbq7PJSA3bUJb
1KL+XRDquxR6lxATaHDhPuTmqYnbKJSYBIcZ9mdeLfPvoU72pHcvRq9H5o/Lev+5ovJVKnYWpAnF
tXXyMR+kea3EE/8OTVriO7Ert9KClV+oLnIjxbmrsjWqTKt418l2PCjPj0CcO54xurkKgNaeXitc
z8OmMaTUle6ApfEIlCBlRrHyowfojsn/V7hKq1tP8PMwCHW5dH6Gvxtv3JH3t4RlVnClSu6nH/xA
V4UzVcFKY6BirOIHLMtxcB2HRe1iOUL8dRMO/Y8y1GzYtccJ2DauR0MlnrqqReyLSyzrolARsuaY
4tuYz6jIznDwz+yL/Wp5cHwsBkRQJnCyx3G4IPZEtgGRVdxbG34SVFlySmjqBAf+6+0jiISw1GaF
ElQzb73ua73u2XWK0IhsyYybhQsrCdxo65pNDSfN/CTWCnbO+0mDGfJGaidaT74pxNUidAQSMnxt
jDP6MAn9QPzB/Nx0Rw5kmfQJCIG0axKayv+K90VHGhzHWQpxkdFSE+9VWNLoXGeCSqptk/2FiXMS
+1sPkQlgJUqy3W/nGzMZ0qTBL14Z9nl+j0VtazkyQLOmNZGmtDeB9LFET3aiPq6OWKGiE74G2YjW
LYIsi0orfG5T5xIUplgjxIDRnM+V1RJpPX13E6/5n2c+cEXggPg/gOUfDgovhaGXqPXWhZ9eWuEf
1LgKuBGTj8uMlYK6hb/ZWlwE/8g2+7cv8NT7RUTPmwZjF3uCggtFeANziTQHnCqKpDDiMpOVYZHB
SFPdifZYAfCC7nh/rI1tKvJvCP325R+z9d+VNQ1JZ22o9JfpUUlZ4ozyW0IKlnIXIWAwM2WIWmT5
4Q5XOUpjAgr1Pdp2LThhJ1HXunfPZC8n+4jhM3Bz4uiO6rboDOcSQdPgMsqkzm+XcKSJwN6E3OYY
RC/gPfS6c/ASJyKdldgdam20GM1694BBj0GQFlToEOKS7OefucCgr+feV6rGcnLpe5trOoLxCBvH
waqI2bVtxqiEveRCwuf4WcXNw4+8abkdSHy2nLomMpUirSocHfpE2E6CIgC2l02xaWwNDIEEhEo3
9/o4suw6YxohMuo3J47DbYYvI8bM6J/cqZMkMrxfAV5OGN5s/LiLXSetzZsx3NGFgiDAQxtSxKCi
Zv81iTgwS5gwgmZQmAle1naDs2GXW3szU9c1DhfDUderbxBzxGedFudad22AMQH0r0Uqbmn/9YJ6
57oL+UGCw4Wq9R3aYG7AwzCDRFn/IUb36d5CzGFWJ6V4vXs6nP54nFX4uB8DEo+yEIzNcL8jlcTi
Dk0IUBNtyX0nf0aNHy9BDbVpH+KrANPg8EInV30eKDFxS4C+4LGy+YAakdUstj9gkka2lovvGJ20
AiSA6/c3RJQmQF3HDrU/fw4dw4dFPyEJMBmmCr/ajO5DE7QJNJGGj0g9NOF8NOGZHkckP+7FGlIR
4EeRxeOzgnoHNjsv+rv/G9Ksauj/CGvtIBqDJNyGTRTfk57vTaVhsSRDKf3Eduwi9WnwVYwHXOgL
lt7lwwnP553IKDTtUfRGDgnMDAk4qSPi6z3NgNdPSCVlG6XdUXrar85iTyY/5XJDdZfsxyMOmkKw
Kh8cr/WYJOiloImlGPNlmQ0wvR41jq1if6SXixN7Vc1Ohwumfh20svLwuG+v+IpcQSD28lsASw3+
MlagAOAjHlxdCcKLkjl9WQUjhc+h4FgZ+VVZn9Q53U487BCZ8zjws5GyocHPqJQhgddtjCP7eL7v
Kv6V1g0dzt16e25oH348c7s5EjydpTls94AKhH0jVlGDZsJjfuWf6wtOpkNsPGxQ2YLzzlyYkShS
dlR8zmUgWDdGzf5ayryzl+ww3rVe6y97u++2oJTOSVbz0qvazvDVfBClVwLnI9MqtTpj2fO1lQfY
YbPwQkKspsjeNmkUZgT67UJac+sVMGUC6vRrty/dFxwx9m2XmDFC7A4Ad1tbJ3keaZGHdg2vJ/Ld
YAT8REJg+H6jDgqOTkufPgngVdQcadKP2Ajr9gmWuJuetYK16hirul7GliY+/c7zZ1IekLPYKes0
rUBbj0nHmzzA+ZR4RfCnNE03UurgzS+v5k0+mLMDX2K3/FqQcX7UjaT4l+UAbn6dEOculn8fPEKO
OO2uZ7GxtlKSpeLyjztA0vRZZl/JjITLmXqaodDHmXIf4pMertIkVua/IqsmpFNSDM3bN1kDCBZn
5tTUkKjnXi9k48HO8+QzEy5wV1TZ50qYTfnqmb80l0+E6MSkGfAskHXzmaecAvztqjC2f+UH0w41
eMP7z2y85s5QkjorGC7UQNuo5Yo3SlQLMa5uDSdcRENOjfuXDk6l9F2svVKKMvc85QoQ/8T6yFPi
sAlG+7UJR5CUPy7XwNslydpPuiJoU5BzppQLWxivcbQpLNiWys1x9tJTFXAyeNvFJthPlnRlo8hD
yhp9e6aRhP2xgrx/E2/M8Wy2HbDPODIhUgMu0jjzBr50D4oxrTCM8623SChd44WLH/JVbMgdfC61
OQgtWXu/mh4Z3fH2VoJwWHCnHxfGrK7TkMK7L01CDBiRmBdwCsPl7HuCwMo/5ti67QjE5ZFrYD1Q
e7qwOPqrKykfthmEW3wGMiBcgW1ewHkb3yJNMApZFUbS8xoP00b1x5DrC9ewSgPNcfYnp4eGrrf9
S1TKpv3AEslw5mZUwIMnPMQKLnjfm6uR1DwAeXVZQC64QMQFWJ5nQPioP/YkE/wLDeQE657AL0FF
qS8Gw2/6h+aJOgxzJNiKiwqaK96GTkVSabtTjVfih/8Q8hVn7ddX+oTIX1otXOJlBYNxJq6V9WT3
lKwauYEt121r5i7DiRuSVDQgT8T+gNk3AaRrhUt9BkEHbx6U949Z84qln8AY06LlNPvB5ja4sTIC
J2jjsRZMpnU3SOa+ds+YYXYy14d0sW9kNHgi5XmR5Xz3FcWS6Td7XrpHqTzUghOVLp1DQDY0C5EP
Cc2f2nZ1AB2eeqj77qPvGEpzICZ1IqOdmOwGF9JjZCRs6Ez+IvjzVJlqVJuBASxc/qq7fWpxvDpH
gXteiUtJOaYvGRBLBjY5M/16E3amk3HEnIBb78+IJoj2+YXVDMk3jme56zFFMG/l6+aiOIokGT65
DCRUyZIMHhnOg78odLLLlrSJVbCJVLCmFPJ6GO319rg7jgnM3eQ4X7tv4Q2v7ODjWBry9PEhzCRH
+V8+0h0RBPaGwegkpCN+CJeViO5S+WJec+Zbb9XcUnCJCZ4JOVVIstKMQUTvbWlAANSeQRFZNaG6
8t0R2dN3T+WmlHb/jIEvTlIA89Jv8CDiS2qYecQc9/nfWQC5t7aDv4Ll0T6/MLNboIIih9aaqWgv
dmMwTonfVMjQogGhiRYYRCdJVhjOSp4DJPgBHZK+6minjw1CncqsC+Bzjq8drY7//IZkv6EUJoCt
SSi2BzJpAcnmQEfJyjJtVfaBCeZRwRUJ5C/7KTZQ5Sw6jHFO6n+rbOVgVZjpzn2MArZf0Ibc440g
c4E515uAwrsjjEwuw6k9bStbDA88qeJgf/WgY30hQmF4inC1ffWCAv9BOV2t3hXjHC3m9lBiSm07
HQEA5DFuwbBQ5qn1RIpEDnzqGx2cDB7Vm/NXdv8ZVdVvPSCEgjBp5jgTm428EDfwvfRxbStygPGF
n7jxW9Vkj+dYhrqcN9xm2nlNXerRJyHx9IkWkdXhLIPZ6taSWMlVsYUOwEZUmyiJH9QJFGRb7J9I
YcFaFOYHKVgRe1HRCkVZBIBH108nBZjI7BCK3Cq3gSc319yGIEIcNuWoINQ7ev/3Iv26eOYaQC1x
SLGiKdkhWL3Zqp2ty1GXlwgKJYIM9e5EDpa6ZBNjH9SXkAtAIljR3cLb4M1VQjVVVJkNHK6WAX3q
nOVQ3YCXbryAV0LZeGVv2PHMKFaRXRn5YEsRwkMyOeMoZ8n6ZRT/aje6j73/7zaYZkyEi0j1/2Ou
oV0oVQpPfgFLspm1izTgJqipvmnf9wLBU1v+jqBZ93xoEUze8tZfdtPuFiFitWh0WyS+UXXprS9R
+O9UUnwQf0NcdNIE42Iya8uvn9DTtrdU6rRn0K+ynLJvsaUq6NFXflo4jmt/gKq2apSjOtYOGdvY
Ndw3V/17XPPVr/1uVzsZRyCIE91vr93BctSfbnlEHGk9zjYkvB6IUwUUF2GuimKB8eGYdUfroIKc
qtUIaxddMY5CyP6rZE4BM4cV6WfaLBx9d4pbNibArVI5ADh2yNJC5qXqPSNR2JiiCB5NiS7arhg1
6cBV0mo9RdJqg6CIMw5EtpZpfVDtN0wj/pklrIDgOWiTjuiLP3l+BtCVgiqmPr6sJpUcBMe2jS/L
ZF1hmLXNWxv3zNpq50Oekj3U76seeiS6Unw0b/qgfr8ceKhTMniszUXW1sUt61vp06Q2i6+ruV8t
HXM6YGi6OMVB9PokQtFYqKzWiwG6Y0zRoL5RCOV5nlnis3qAxje6WP4cpkRaHan0VeKKJXmxOwNH
iZbPWL8o/IDUNGmW05GDRhFKyl6n5rmn2lPA/5daN0dFUTns7Nvlk/JKg5DGGVyAf6uq2nvPhHPR
i62CCSyI8OpAMr/SdbRaF36b4Y5b4wLowXFKkw63VfmW0gMTz6og6Wwx3lHedFwAYZMCPjN7GKMV
qJdlHXOcJ2iJ6z71d5eCNFvv4+Bad/Cxu/BHCfE7/gwVTGMTRjfwtL7JdFvBUu3V+PO6dJu44gu3
j00w71hPSsRPuDg6hf8K7jAJ9V1DwcRdFJjJQF868lTyjId6fnw8G/EwrsroBW/y+4cJjQM+eFyl
ZCLJthqQih/faPqCryhK2cSzxAGiOG22uPqAWm4bFuMNShRngPpkIbkJwxBRsPcrPN3tVA3hqc1H
vT7wZmottK+R4j2lReVh4rvfKd3nCYlw08QgrAg7MyqeefTEKNd4CPLa1LJcKE6RqeOoByvfKAut
aQUksI+cKzD8HGmrCPtbhpeJv4EdVbbK0zAgY/ZsDtbj2lIuZrati97h+bOkBONX883iehZYOdDG
SzzpTmWrT6fH4T+95t1JsB6pp46bvPiINA49TWHlB/lK66YebbYQgjbNqS2t37OZ6BBLbioCCNHZ
zYJ8GFv5FOHIJwJtccmsasKTANPQjiihwbPL6EQVjjxXKSgqz8QqyH+YUBXnWKZda1T/tq3j5c+D
91p5f/0hcKbc2H13Db6+mpTeLK+ndBI/BZwFNKLp87zNro9rQGcNYnqIUSfFSlMxj2+TXGwHAeVu
SaHFSnqrEKnBLY/SJG+BEBpF4xjHeJHxhF/PSSu88qOruzoGgmdiHS8WbZvsBxWdHEPu1u4oKyAF
XmjlT34udpbSqbPYAICgP4eRJZi9Ip+oUm/pUAOtFx5xfYJXFzD32LPuzeRBad/iXqr2ld1Tm6qD
tV3goJlbZvdV6d8GS1eoofCZwqXVZMb75OWSRlRwKmvBxeOhQsy+zdGr0Y3uxZMAFsAPdBsx78er
pF2nzNU9mId1ZHoJb668/NUGTuCwQQEnGhun+jxZ5nmq1fCvY8yA89Qofo/75dO/CoNxlQ5euzOY
Z2d0OdKnaZgk0skRewpkol2Ywh+nwk53nm13yRHV+XZZyu5vFigC0f5VebEaEYcbIs3676pex9o/
7b0k16TjdPAcezOstts/F57Zi7YYryGYzaBzCLVzVC/b5+A0wbBWnyImTAbmOTK7RFVKFA3q3TQk
cvtYu5wnYFTAjje1klJBHSOSH9Zln5ofJyWmqbqkQnR+BoGmN7KPjfyIFMByKD94oQ6tT8Q9g9Of
6FA47k2Mkde63xVByisyHTMBf1r9EzmtdzEQGuUoakCq2eKx78fGWsj5iRi668Xdf2/kTO4E5iGi
kBK9BDaq9n/L8yDNGnuk0qe5UBOD031CGZySdBZMVcY/UENAN1aACQovY/MKRydlhnVa658uyNkF
B5keWAdvorxymZV+dFBiiEm8EsJ04yvV6j/FZrHVjABDvHPrnnsA+z5M0/FOJwdXCyIdM5ZJHHu+
9DmhaCK+34hhpEwASprw/G/J21ycL31s9MYE9KU8zjwOo18/CETI0IthXB+6SyGvkomdBQsbKZtx
wAce9jkAKTFfWAXOBUIH3VeA8+VyNXMBkC5FBM9kCIMjdNT3GS1hLTTJTSwks6tq2k91HCNWcEnk
eRTD44lCFHOP1p6p3LwM1xODjylQYdy6olyFeVYvqOzYGgph2MzvqEnMLMfHr5HFtEZqxuhJf5gM
GooRdBNQWMN8yJWgrCxx/W1BMJEqL+5Y6+5URyXCRGtkk220D7+4qLEP5bvl1xpERYzG64ES27i+
MwVDVC4MhnagfSy2WSiFtjOWpEUDKj0cSCZw3WNZYpD6nJPdDy1F3U5XWnho6lDpY+qhe81MRCvP
mqdi6LOC1boCQkV3OOpxUgCEv4gojDYatTIdrvQtU48lGhkGwOT5DdBW+YoXevyNofqcndsUddAo
B+eEn0H/jgS/0id85gACWxmXpFA6jS3VXWgXAP2vE8Y7U0Zpr1FE1ncovKfEMUj6PLc3kAi5BKa6
hoOGma5eF9lHO2fz03rLDNLZGgQ5V5llXrEQBtgBga2qMbnxRtVCBKY/XHUEdWEOQL+ltsIskgvU
9Pl/l7ffkKRR5LWP4sE0B2C1gMdyhvLsOxNziHrWbJROWo5eKQex+uhzXAQh+W3qVhmOTn5hfK7a
WtfKDgC8g8Cr9l/ljKDIqgfhDXjyPsnigzK8iN7DIueZKglsVrotwh5JPy+b/T0lTaPZMN+7IDFQ
9TBRcdwiuTZaCXWqRnL40FyOtk7rQ9NmcU3U5HcwT0qrEqZ21zgCJYV1AxOLcriuMfBAgJnjks2l
XAqfMavAZlOlJbRdsI3oU0yBInS6nleMBymsAyWnVe/a21EpVfCLRyVoeVgQ3cmfYGNgLGHtS7Km
VDFJjJ74p1xJy/aK9o96cdaERWq4nunLbqmxbkfXFBmPxoz5pQ3vzQ+T6DstGJdi/c9MIimN99yb
9ZyTrvgcmd9qb+aj0a5X/WovuV5mtI8WAs/bAFrm6Gkbmrc2ZNfxpN4GEDEm0aVFL4/ZiLQskocv
0bo4knCqaPG5zgdP74zhTaITyHjiYGpxma3+m3Phw8A3sQ195G5cucxogl4cR2BzF7IncOTnRzLQ
GPYGA3S01568NadpW4yv82kMRBa02NEw3nTr3xZ9U1D+B1Bc48GfNMqpSezOE8jRwUriREzxlzdl
+lm1I77os9PIy+4BuwnK7XS+APLQP48aGVDGA8L0/SNKYTeZ/TN6SCEpqDHhQm8TPts4tYgmaUSz
CA7feoh73MX0TDFfjo+9HYAgsYKklbFF4wk1Wb7NyH7qEvPH0SiEFwrRfkti0ajOt3YSqVZk56My
KaXeCCFGZa8oD0Gyo6TFTbJ5AExdO8OFrSmQ8Vml/yQOr1PeLGSNlzmYVX3xFxpLtHoemWLnjCRI
J+41j2dlNN7S5KlLvONVQ+SqY/jLsEu+NXsDzXW6ZOXM/Zv4tDiRVYm9Fg7tJ+DEgVV3Kh4KmKX8
rN6HvjYTos8XyfuvQZrgUv6m5vK9IXBT8wsok1FnA07YAwSQm0JP8NysEUSg9RI/coHSR74lQ0wx
b+sf1bjK0tJVqguBBjoRb+a4SzZTuSiZjGMVk9iAoHizc8ZDzq2+tJMd2/uYCQKlqRsRvqyL8EOz
Wx5RJrdTS8BPXgYGFVt6nCfxaOqO3G6ApS/dWu3ILzk7CIf3/uKxppipW6ie8klBJyF5awtvWOKH
RBmBp6LCdUHRPspDhNgjqzvtKI6gvPLhKMFBsh1cTIGjWjqw3Qnqp0bKtOQ0otZm46WG+h5JjWIw
jGL7DuThIOjkbNYcrre8aUj28FjJddXaW/dUm1+iH1yLgTKAWYlRfeIzQS/DjZ6SRZNFXSoXo3Tt
N8DCNw+S0fM74mYI3MUFgSJtnQ9MLQUZGT1SkanWqd4KqjhbgWd8knZaOTaDSzUTwWroTh+jPh4l
Xu84j3/kodYQfx69oIksK896oAxAvLa7wlRYOVYRupxdO5NGWr/J4R5xQd0FR+T6Jf16D6qZUntR
rHR2TMbVBkHGrdndKUWwZEZG6j+Xczdb0LctoUbxd67t04zUs+fEE6zOPr0t/c7WZ0wo3crCd5rG
tNw+vgRJPocJW5RXxt72NkTReC4n5NZ0PYjM8M6SbTglJNgiwDvmo3ivguSasmdGLPLz2o6JZp9q
k1y1B9hZp8oHn0lUSRH7FrEDM1kKlPxsWtKel0R96JcAsFQFCPIv0Q785zhbd3dlC9zy6qoR9cYB
KGyEEmoJ72BGyhFYUI1Kq0dFNwHdoO0wQPPHjiGAyq+NzdXnOp4z6uXnQ/Wn0JEP6b6X8v6PcBL0
C+BweOkKMd9sg3nHYKtBrrfWrjArOj5exVzHCyD9LgzBanXEu8A1P5vtPXL0sWb5RO099aiJK0o5
cHM6lJHVLpHjXJQQbJZ4a3I5lNrK6KJYirMcdT9LiFBK4CmPFMjHfw0uxgMiifsuikGL+fPLMIiH
/4Qxopj7OBbA5zop2gSxEq+8cHkwOHjtTt0RO/kpnIb0gJdNy3d1Ba3oPeLleHTZXQuvp95NoAqy
Tj2MenAb7hhh9jchSnm6siDgP5Mnu2wsXCeMlUQbSX83pEYkWVZgdPJMxhLdbdfXVyUtxfjPWYgR
76LiaNP5LCCavFlYpiNyQPCAbUZEz0aMGUXoUomQiGMmpFGyBPXh7ySMtcEO9DNf6+CpCRslWzS8
Vp4UpI9t9uLBNN8WJ4yLDsS2Cu2/vcjttQdfCEtOKg8bq9FZcaoqZjqy2K3TWApns1wSYCOEfFuA
h8aAsHDc+AdzT07f9YcOlHIhXVEI83mREw5p9NCulOAbAXQEAjgbRCVDF7UFpIRvqPM8nYX78Isq
AuzEhgNNEUQY+7aBED0w/aEi4/gtUFIIU+ljsCNLv0Lv41ZE5iWfpWkxh3WlcxBBE7ULwzoDYlQ5
ZcuiFUqdNrCw198WKBlq/fn0JppenSv8fprEmznsf47a0Uy6mZyUXZHaE9iCYGXQdDxOIBtOxH60
+WmsYFii8Fuoyn6JEstyXffC5Tfx9IvPI5IzqPk6qaDxm/b3aTYfHmFb8YxJk7G/jj40uqu+7bKA
3N6ETD8yTuNuCTksgUdb6wCQgGhV499UN/IYB3Zqk/gxZIOUsP/8WyPhnJVN2WI2j+4rldtOjjTn
Yn0CPHTyIQV+Ewezyd6c5he/Lhi0O8HsEDZCCPAifL5V3wVpWQgLFmDUAy2vwdPjKYw3B69EkWIx
ZMDIIc0uu1dKf6sDBbOixx0MmqFlWPPwhIgSH3mtfQtWpEV72KrvsDM5ALuQI7cV+vYDln4TbiJr
gIBhhr53WN81fHytN2P1dlq4ID1KZOcaApt/GyJ4dZZ2YAApMvFZb0C5g32Ym7g0zUKZSjlK83WE
R81GHCSLaVS1BjlX+DSXy+46kvQtSHwlMv6sjwfGlwxmLcYBWlqksnFrVzPMLyX5VlWd79aYjXO5
bgbi0HMWciI5Ethfrujv2+fxnEq5JoF9PrUw06GJXO7gA4IFWzzm8MPuMfn/Im6Uiku8UX2FOlqk
gqb2+xKraaK4DKn+oGqQS2ayICa+X7VhHSmzMkM/YtfdxU9mnEThJxQZaPvWsfVWQHqxOfCckj5e
Cu7qxotqlao0W3OwCDTSRB+kx92PXhOhHjVzijHEV8dumZa26yuDmim82ROH5XpS+6vvF+DI9ohA
F79jz21BUszEvDXctCOcX6B8K4uS/ibYLsCQ0GHmJdyr0dactP8ZrDzp9oIF/8od/CEe+X3gTp6G
u1l7JqYFcNwDu4/Eo/+ydEMmpEdc9BUskjRqfZ91OQqXI+3wknxnPeniRpAd/IBd/GhlywWW/fgu
Xei8pP0+bCxRzARDdHUIADr8FgnvLxBLGY/MqJqUnnRapDSS22WmtrWnuOe7cOk+NVvEB6/BNz4p
iGjdkLCKeWjDzgYGRYhpdYACwDnqf0x7VCLNJxCz7HObVonVJFDhtdKDVMtgCB99mE+lGs9UdS3D
9NODl5RgsKqSz71JTOFPBjPRcf0rayb/Vv0iclSa3jkupBZAM82Sp2BLvsnqP/Pssh5FHy+4yDqf
AruDNmwyGSh0ud27fOZZmzXGci7KTjA+DaNn6lDqvCrgmfSHInprgaWFOJmXrqj2fVsHrHEM7qHS
Fq1RJyESsvJpSwPSFfyNB/ZTGYl782piqvUt1KIMSiJr1ZAR+MuRmdfY0TWzFQMsI8DaikKgcfOI
uYHI+4ravcZGJoa3EVnS9xLrw7bSHL7TbEQFwwqjBLB/5DSSMRH2Ryo1DtRRt5lA+z+n5GM3p1Ne
th3GKHPfVjX/tfxjfqZkd+BwLxybrT0GOb2CRWJOs4AeDFPvKl8yIH+Ik/wbcW+yH6UoZhB33Oda
XRTf9Lb2hj0ud/SVRkemNbWhx3hAIxt6cMWDimUVJzVt/xCRyXF7oiRlvO5ek/3kHTUhFLoG87mH
LRIgNnae9DENCYp4e4IFtXbuiaw0K2EbBfCnpE/Hla7eRH36oj8qiHynqutGzx0IeM5hbd7XiEZH
m4dMpAqsKD8g8NR83lbAvyNnTSYrsrkQSqb9TmhEKYj05dIL8f0IAtoVW0QwQ4koL4J8J/b9quo/
kwnvAPUzvQEE7CaCQV68WympeSBWy8/OChdXt1ggPF7AyZZtNw28nXe8XvA33R2imYcO6aNiidBS
AFRf1GkCyyPQsDzEAaUG7AG0EX/tIdTX1S4FPCfbcZk6zuGyfw2aOL/PlEI2cVwV16mrvbZPXxGw
8QP88JS+mv0JJs+C/0BeoEMzK+EdHdpY59BQz9pUPJgKP9fvfpxIRFZ/cbyLQA3miUE9rDnSdGYX
cS0IjDQ+jp8ECsca9UVdKhYOjdse9JIgUWOwLr1+pihXQ2QSma8jrGQDvv8+FF28Pyy13RIDCeDi
SPM/pYBlaVCers2m6hxNPwQomunL8O9/Iz/C0Y6PiOVthCXyRgKCYqxb2DXUdWZAomebIFk+9gR0
CngBrGNw6HDk775bSKQ64qiCR8htIFU1g1iLbBfP/i0yPSoOniofL1sD/Vn0eyAUefmVp+FT1gm8
TPmSDCRIMuBCwfVCWBXpRZvfFU4gIenn8IQW3B0StHDAuBltK/y3KJ/POwQADqwdJir1CXztyCFG
ZgrgLpnrZVlL0FC0bpTE/TpG+xQpcF6NcMc34WoeW10l+YDte8pMTrecfP6AtaGA9RTWymWfGLXg
pc/H6yYLf6vwe8NA2LIHiTXOxA9PSX6nw1mUC4pojsn6lhqZzYvbLCDFrKODpQfdVVyhXu4uVoD1
Wm3fYE/E5V18OoOxpwclWTJRs/4kpvfFzXEYb/Y4svFo3WWaVUfpwBIb/HW6o66apqRZeZCmwEH2
jj5RQsOTmJremjs+qh6nNghw+DbeDPYSLWFHDro+URQy7S3RIv2LDqtCDVgELthWHe2kkXWCl7fJ
Gtb1XFzm8vYKvn0rjl1/zS9H0m/LlahBUqt9F+YqR5NtlSoE/3hHo28P4L8oKbDCCmcTT3cgt9fH
aMSG8frvVlo7qktYl0gVG75+UuIXJl6CMtMOvJLuU5HS3Fs/BVwook+XKFuEmew2uzZG8Fkp1cf+
Ks49NmMZ96BWyGa1CXTggDRSwPojBB//abZ0LcicDxLV5prIWG3qmLWZk2jWvKAyoEio1PVKlmCy
5Sgd1MBgtJy0WjzSeRPucl3ZyuvPA8yA0uaKcP/kKXrdneWmKI68rGL4NVyh8JbTumPamMN/l3v/
2Wpy3ttVB3k2qQTJv8K9MP8LHSUmnva6uM/08vW8GxNFo2IeAxets7enjlCrrpjHwP2A5siBUHSi
td/u1Bdme+msXaXuTY9tG0AibEtZIVEQiusAzB/jLLKjeCKQPkO0AMEr1pGSdEDP9oa6YZhTXkx0
rOwWEXLDtQ3+mo28DlbJHiw8dKbmI3C4gBXA9WH/EVfHSguxPVN/WrPcE7ghDPYa2bSIOMD0CcsF
uSYSUnHpigfXt6cJQx1Ea+B6vvrGWOMEglngqiOLl+9mChesIhw0blVc1Ux4T15ml3WSKY7EpK0D
U+Vyq8Z1vmt1AbMe86EM9fQ2Szzjiidb/AsQAw8b8wFpv9WLibT15VETmT7U0vVSm9dP9tK0yiAL
e8K+bAEB91pETlbJrdYHJ9ido5eduDSX0wz4s3WVz0NfwlxBx+J6FEgrP5hVXzicsBqVBmdXSMw0
J72i5UgcJfXlmn6rrV8oUi1YrqDZgTH6iHcDRoIhL0acvkKSoKKOyaTcffMZwlZEGCvr0y/YtToq
ubNyzA+TL4hbtYhq3WzKG8lgl2W8sW4MzyW9H6WCImhrpDqZgckqBjsx8+oqYWJhTsJfxX2DfL4f
dTfbNfJvvTbl75DY8oFYkgwZm8jlD6qoQOSxKPogXkNJtNFqthSHu9FRPflt2lERFxUjxmJ0CfXG
0EoSn4Xnt6Mydhf2fkjXrxWnpI7mZKsCzNQd5eQneSIMaimR7gVLigG9X8/mV+Wop12JcLqn4UJf
NKYtzaB1v87KSvzi8t9iC9KZn8vCdiaD4Ca2c2aGW1T8zyTGDGUzLpjmGbo11l+/tT+qyUsUXdmT
vyRYnzTyAH5rOTJ52+3QDEhIUAOICJMH2XhVZCqCZ8wfSxfA/iUjHULHrPQNwHLAn53M4dwTU0iv
AG1QpBKqOs8LHkTWxp5eE7ThYUDvg5pLeJy3lXNRj6+ghKVKOpMoAfw0vv/Lmv53MOp1Ws5lMZ/q
vpVE7LGbfnLpZFEcZnTZFyNgOAYkzoh/n2U1lPFlzGkbspsBAUymKkRDSVmIjk1h0uphsZcLHyEJ
826+9FqPggDzZN7La9Oyd1GOFIe3btmVRhfMn74SqsHJItJcxDKGKUQa5B8cePA+YXmq1OCK31ht
a9I4Zq/95mCuXOUAYTYl17d7AGmDOtFZur6ZAugCWVZTtXiyGer6lXTGy6rYgZcWYdvmk07LDQ/j
sczpgktbx4b60aGyisQ6+remTNuZJbRheKv9jmCiiSFBTUwri7PO7hh287TpNAFvtEkjK3sb5xrJ
/bwIBmtwzodbLHbVAyc7E3v5UjukQ9s/8fXUjf+7B6dCwJePA/qLl3lTfeahQuMx8shNkUBGTm4A
uTfGP6hqEh5ot6nIlbDqZbidlAfNy0YPozGgWCGigCWmn8HFQSBolHopdCiWzooA85Co28pVxsyW
DrE0man1jR0vrsM+1RJuyNl27Hx/vLlkQPaCC1qCsjuM6gdnzkmTlBEoPpmhueElLgGFXh1L2iDF
jwPUQJireII/rjcfFU6xrUS0LiZeiZbSvikmMLphbGAraVmrYzEYATTjgLYnub0sl3rvHmnk4yZl
ML1nPUDeZ/a743T3ONfLU/tjlqmTG44RP3K5Lm48XK7i0poYjvOJZqLceHo3zl2ypZY5l1S6VD93
fGZT5fbZjneEVjVeiXBLmL8QfOXs4UewO34uawlytdbDjKpLxvVyN1f9hFOGD5ZQymbxgNnKiZjb
Kjgq7acsdlTuDfGJsaVFFqPBQ959Xn7MypIiAVwlaQTdlLAWTuG928jMwCtZhgpD5LBXIb6j/CTw
mZjI2KBnTLeGz5ctP19Ur/e42kdxNpJB/t74hTx+Ch4fHVOK80uB/p+CQTE8X+kCXvrArQ9htiPP
UUBBXLVYUIsOOinUIaf57ln3JCv0gogievOcQglt4sjM/ZeB9j+ZCqS4nuWkLZEVh0ivAr39cCcc
2IAeiAiqLtnKvotPfO0gkFB8+pYCWQMMZhC/xHodoDNDhV6hbfTW0XLzBJVYPLZXCpHVUS1Lxshs
UZw7lQxK5+ev0GGumBVnaQjNsT2LNVfn6ZkHvh9uka11V8ObEgsPrMzS2/y4IV4Jt1zxfyxrZQQN
jARC3tGsytDF1BVneQtFCyXOrkdSZkbKPK3yGZBOvKcIuCyV2Qgmz54fiuyRT5AjHzQlu45kDksW
Gji/ZtcNSsPCQs4AR00o/D38Ne7waJOqIFjEXWytXcsJPb/XOWg3lGxqJMs4vthws5lv4Hb/nGBr
9GWcnT4bXWe5hPVKy1VAqFSWZ/PHZC6oAJtxa5oiwYDXYH0RMA2tUIqHnL/f1MBoJKhxd2owcFG6
u6jsxBSZDyP8OEkNaGPwUKOSxI3dvKdrK93wINZfu+K0OpKG54eKSO4dPYpUWKwd8WJ2guhp0NBz
yCi83zuspKzxUrLucewb6c58JjUr8axDYocnuLdEnFRESLA7rcfB1jFNhqSVtvqjJkrOEPNFvHzI
ocr9c9GLRr1VHe5mkD367Woy7m/WEpKqmc/m8z9h2uJKbSddb8c8l5JhQsiVwRgg1t7PQ1DO6c/Q
6Ex5bnA2uyun0ruv7yP5gcsIQTH7BZsity8UnQ1xZWzYI85tE5U0vBLiuXj1elK015FplAxacHX6
wKIus4jhv/V2aoqGiWszYt4H9zfo20IB0OfYfdKG0cX66sOCHzAUlNP+4cTwbOnoosgU3b8vfdKM
yiUz7G3Lt8bhoexZ0IRDdGLM4vUQi50/Iwt0TpVzd0Mf/b+eXc4Bn1SJ1C7wLX1g8pP0KCWtP1LD
sCzKhKlA+xdeMI1Xvm4Q/M7EMVkiTYJzKcm5naU8xSn8iy2fO6d9p8JwkrTpUW1KAuPvf0UMtprr
Nh4drb+HktF8JSMphIvYZLJJyOKWLcbtvl2dFzGtoih4Ym7TPM5gipxI6wZv2fZ+w0/dWrFWGsGy
MJu9HGWz/+8hjZ5zYp8PhDGPIy+NP8HQktWF4ENZJQdHbMgwTUyl5CHUp9TL/PTozPSnpjYqhU42
40hdvY+BYTZpXs7+/PxptyjT6vfwcLfPR585zBXnV+j21GRa7PVdKWAkolWNpwtELjSRC9mqJF2Q
wKzLgY/zFTK8LPyClsqy2F9ktTsGdqxaUcF/qlJySbO4uaCNBSTQb71a95ITcCaU+L/ldEE0PhkH
2FOYdHiGvW4yZpSWfrhxQ/xomclyg0O7hkxaX05dIE81OeIyt08gEAN2cFCo40MV0c7ull+a1tcg
0vxbaxk0wv6jOorQJ043n0kV2AkNSTEzyjTWBjnKSV6lQXXrv8kZSgiQbzGAZvqbqLctN2QYDtm7
HpNgpT9WCogiM63BadfWa4a85Mafa8Wv1iEzioGoXmAiPt5u5Q5NeRTU2kIgstVTRYlokeWLvLqh
yCoEWb1IJjlVrT5ORs2KYne+l3+mr4/xKsYoG1RizwCKnzSP021lO0AYwIj0+sDF0tdhWIrv0Raj
kb0Dq8T/YPhcFy5eJdLPlkh4pKe9QdYrrNRF7oSaIV/aFxqwfMCEwc93PqyJ3uyhdR/D67ePEss8
xArNN7Pg/Wi4e1W4SbM/QE0DN13qIbygJLpATHE3EJ9WU6neh5Hs4deJ+zbPgAqFMvsE1D0LXbNj
fSeTLoweEk2zK3NATwdO//Ze5Qs/jYcJcf+kVe5KJUjRSIlUd1gYgl9X6wYc1sIb0nxtWXS4Guo3
mnQehwDCW04gdBD4bbwrrV/XD5xYPMhgaiLaVaNYARvDfP483fbIAZOYH0RrofRQU/EoNIY9KF8I
qr4iNMWY3tWlleBzC1oUi7YrTmthpmzSYiYwbC0Ec9ZkT23959nTpLVE8txPW6zvkRV99MNPcosQ
KHIWR6pJnNto5NFF5EFYpSBAWWFTSFaXUX/2xzYDotW9TRn4k8Io9Spc1gtmhOWz9XduKacy0/3z
dhJGJHUFtlmsslM8uSLOgBqfBcH0PkgMZjSrRJuUbTcg+CW10zMWBQNodbH9TxEId6cOvB1671NO
E0NyC0On0y/GgkZoV9WlNdEEMZsmZd8wyGuscLwLaoIL94g90u0enx5/oidOPG+pq/tLW6NsCQsQ
GgeKzPpmPjyXcz1EQwdBDTTQ/3up00112EvxYQ9urFyLR+7p0ND4ehk6pQ7szWwj8cB1+A+xQua8
xGNO4fDPD9MvmvaJkV7S355gMjxmeqx3TXqNRiO16Ezbw+4uVQ33ng4wzHkY8tp9TvtDjTQ60CP5
kp2kJttMSgUQqAQIx63NBQQhN2aLNIhw9HljxSzll0gEqoA/sxPtNsZrgzzlVtjuvi+EIK/q2GeI
2IrfcdKvWkd8Bl8cadt9Rro0G/YKZVlK96dMs0Ip1SxFEUxuCcYJNthp9Sc1jsn4bOab6yiAmY8H
IiP7zh5xUyu1fBhFgnXJ0VQD57+RZbaifYn0xR0fMvHRNTH0rgMRPf14tC7ALuce1k+YgIDTSMua
wEe/RogCmeVeKgeea2Ka9S1/nTZ+EeniMKS909gOmqp4ctUFitFoRg9GKmak/lRIY4ipg1l+TlUW
xfdU6VpIGcV8em+/ybrDzlXLbOaHYa8CuveCZLTMLb9d+XyyLM6OmIQGRUbFAxAfyDapjk745FMD
ggzawb9PJBG992weg9qQF07eFi4d2z4ow/lbFwSvXHW+gXjf60JlAr5msw8MUL3VV3cDBLouMUIA
sw9YpU+TEvz8/ern/WfH+w+xZ1lWZDzmlpxqXtJbUAm68DtxmoETLtneyW5S1oCm8BVbuEEC8dnW
D1K5IZ2vZdmv9A5T+u06942pSErdxovIShcZIM/WgADcI+dT+jEixxZla1RJvoCUWIKAeHyw1YF8
rLqGB0Az4dhDWQJsa55OCzPZpSssKqTlUTfwc92092YfBik5GwTRHz75CToLNV+dMC/+bPJ7Y1km
DMH47oA7afiJ2nPS3+gWjrrPlO4KFonOwZ7xeCLQGzhiFVttBsbcUnNJ3m/XUowaOLGxyN98xhvq
0AiUWH5X9S5z/9p3+nfvTgx21riuxnrhOSVOiQ0q6cTUBbwoys5GySzaMkgqQjuBvMd5x27Xo0Jb
B4m1cQlD/9U1QUx0h4Q1vf91+FQupPPyQHnLfP1n8fZ63uQmxwveo+nexHdvrEFo3HHYKTbflU+J
s8KBDHWplJ9ojgNszrCxtH5jrZGjnj2f4sSqBDjDwitawLWS5A5TvVORbz7CxDgrC37WHkR18n6s
BtFoKgg09bkF2aVGd9VnTLXFRt+F531ddAqyj7EaNBdooMa1mdar2nR1xT36CURI/Cas54cVT62d
zJL2RHRGh5LRMxhc+yJvah80gDPgTHOjaWeW11wpvRj/ol18va8cKzWsQ/+9hK8mD7ghzIDWWhHU
4Y5hmSQke9n40q7u1/XwnOra+UPJO1DhIEYWtKBSu9I4FtzpMxqPPBzd3rS6y7t2hSFV9YaK3dq+
pz9n/OnSm9TEPqZ+15uhgFtofUpM7s7yLozyHp3JtoWroMtG4JcIQu3bNTWSmUzm/YRq561r+oNn
bJ+XgEvqZGaTFoRtn7H0UfyMCf2Rsm4SeKutFYpCTOZNlVE/3spfmcTL2n3u5uzqSsMAsndIviil
BmGP5QLhff0ms9e38Hi7OHe0dA4j8+t3a5L6pM4O8NkW09K50itZsdjcqOcj3iivY0sW1tcF1TsJ
uzaY4dSIpGdBMK3P/SlktvY/OoyJE4Gsdw5Qqh9wvVQ+7rcQrsb1v4nv7WVLzneCYfwSB4tsatiU
VX61gaTZMqgJ4KhdIvqzplPxkIdPf/NWAJQGqfZrle87R8u2JTMrmHRI5d8MSb5v6R60PorZssdY
8QmB+XJOosutXu1TM9+gwi1VPuApQOTYnJJJ3ZIJtAq2z04/Dwk2haf7kBJK/NA75vsV+RfHa5SM
1HcJWy93xHY4dKOUbJJODJ2IAmSNLr4TkqPoxfmH+e5ZM0sdUVz0UII6XzVPPyr3TVyslZ0pSIll
DHrFr5DRXhPmaLYK26Xda/pvRJi+x+VTxju7T8CBpgFixcp9WvrHcjlr8D0CjlKxVJ+Hz/ufW/6K
QZpzPAJQAjGghQ89qxNCdP3GZzfgIW9xAacWx7+MpXbF4pHz+M2KuwMKsUCoqGu9B9EO540nyXf5
eMvD0z5jdZtQTUXbHg14dxMxADkOOWSkJ0JEGLCMikV72o2U5KpBdlOUplM1aqPOqzupzGqJAJmj
ebdCxggM89JCAMMk2FxQvWAs1mP5P+lwP8rHACn7cxyTnCT768KkchKn4077cafh2YSuu8JY7FdQ
boeRYjCRUKiCN68pdB7wQ1N6yYtYhsSt+So6MZkrr7kmMZUSJOoiE7Y3XEZVA0L7DpNEhElrBMJT
sgAjujeuCReeVKj6aavzk6UROdegwx0zB7Y7EsNnaLvpNc+v+2wkLCkTQJcwHojdoJg9ZvtmMvPW
gUuGWOqQW/PI2REfkZeIdIrDwW/RRtATPgCmgY3nSXB61jtbqyIpXoM9KO7y+KCDOekx6Ikh70/E
yGRD4L4PauVffqbH8gcgAPUQzYv31dtfddF6XKH+el0crcalDZoygb0aCo8SqpWzaPBc0arLn2cV
Cze0UzyN9d51/yhKnnWviBc9pc4DLtYjqg9B853ThMRcaY6Pf9mUP5sS6hLJIVnV9ymYe3ajtxuO
vO6844UhiDpwky1tBDrJBnBM5rWOTEaZxuqMFG9ucKWImfrinntIpUGiZia88rlMSJHthZxIeqq6
5u4O4vcb8AqqQHQhtwDe5wj8Q0N3G9sAlN1IGyH00U5Yd5PhreTQXOw0Q8Hp2bdhsZCHw7MAEmoF
ZKyvyqQ+HxmMCDEQlIEvS6OwVaPCgHXWJG3CVljopNbUJTcuC8wPeaL3xOT1P9TLYsMNuH9J6195
bEShCpQUH3JtLn6sK7/EgiK+xdYcmqGTsugp0UWATU1OL7q3BKM588qVyfQA19FtchGNEa98yjI3
lqI9XoVI+iTKoJetE1ch5KQGBLFmhpfrPlWjXjHlfFU16pLJnVoGZ+3HDkxvLjvpOhAKz8uc6auB
y6oL6WFvuMu5iKB+EdNGquWqo6R/QoEPVD4SxhXJwFR1xDMN2LuLlqenlqi3D/WI/ZJjiadlZc0W
afaAjYZ6rM/o4ZGwteU/AVxYK2RpI6Srba0kt+iD2O3mGOkmWdUjMaEUcVbuwwC2PTkg/W0IrYzv
BWh4P8RiIcG/FIKfXApw+ka00buG3hEjV2ZDYpBpf/bAHXa82h8tEWBEhtyaLawa6vV1dwqDxQ3D
OR4HiJU/4UKPdAosiPR1M3J3/zl6rTR/fF84ulySh+8yC3doepK2jH3+BZWBgkfAIIO1NawXUmDs
CCCihNJEbHNmZRVyi7lyza2KfLw1dxt5hvm6rc94T+1TdZ5dbz4s2OEe4AI7k8M/tGjBoteIsOUA
+z9t6JDmVJX1Yd1mBhkb0ZezI5FvE7FqHGRxh068T0HkfPL4G3i2924sNur+zeXCkNHm3bLCmd1q
KVlqb4DE/TOqMaVpu+0ObjP9ueMgywmDU1OYR/arZ5PM9QtIxdIn7zOgMKLRT/FEHIDGFnTc4RU/
jSnn3xYEr9nNdKWVQoCSRgdZsQpsKv5C7dIZQmEU/wNQmcvhU+gyjl5U8ODS/NaiJnTZmL7Pql8S
rOmVVEi2kswnYAlyHnMK3BNnSQethOEcTW0xsUYHKVgJ8tHY2dvC2gFjOw60V74UTvS/u0Jo2LGz
pSdreaSSiaoUTekEkdjARhNM6+IloAMvyz1w9QlCxdFsdTPhUNEUwSQCUa3+eW46ibcmmIG7I24a
njuENl5+gnpmEh5VDQxbAHls2/0Unl4iD3xWBGish6sz2S+qhosqBqKXIrQnqzAHsS52FRm3I3os
xvXFjv+m57FjkKmhPHcaTJ4ReivOFSImUzaqRUD+863fVdmktTQu2cO8uiwBtjUvRufklvK/zfaz
Gaepg168ICgUMK+vNfQAA/N7pK3Oj4p/t/byiBe6iJ6FgAh2SfL+vwiTr7qeTCDFvVsE0enLnbjc
BZpySVPnn8FrAmfMbhGZJQmilh2J52SgpHDHv1Q25Oi9z4deTZo4fJcIv4vnt61VucVT0lefC44B
psZ6tjdWRPHbqmsL1iMRW6RoT0gkiAJgvd9Qsa/bXXu0VX7yqxZYbOHZUpX7pFE3IkaCojxQyhyQ
jp4C5T5NnKEHwWBJC/2YShEiCjN6Q+O43ma1oRAR6qD3erxAbqO0HDxatzh5AD+CIEL4VVfmwHCS
s4LdgtvSdhjouQnC8lJPA9z/60AUPRRof0mwhPnL8UPYUGE9HM6foqAnQDTX7KovXtZuz11FIZ9O
tn+/qjTGufWDORTqpoxkLO3c+xKYu/oDFCUJ2QMKEJzjFi8kEApNhv6EhtHvFJ6UrcF5TUYnQ607
HjrnT9TSLjk8pFgBEOhrZYznMHqVm0PgRbP8NXrhglnJ2P5dV6X1XKsiUTwBwGpBYPpzbcBxiL4A
or5bZyUkAAPXD+jy8f1ooXOvDygU4JLUCX3L/U7Qin4Kf+ZJej+fX4EaO8y5RGwO2siDfy5xVAF8
/F9TGNe7JBHLrdeDqaDcFY+kgL6EABlC/f0EBuNQ+B+geRx8aNVTDnojcYP/GBuZ9N5vXX3Xvltx
GXvTTLnYjp6MHmsgre5+i8obafwu5bpEtgcLg5Ls72JvR5s73L+Hu3Y4T+lGF+8QeUHw49ogGa9l
UNU7ilOcJCulVJzs2i+wtxwe2wrmR8j+tbalIoAEQXC0NpGpMPKgDX9vHZfUbJ8uYilzGlwx1Lxw
r9yog7exvWteQXj+ekqqPdi0Xh+CXuK/CDqwRVDBgYxNow1QG2E6QsKZFZpiQs7TijhWcDT+8+rX
X1M8hd3JDC1uYsFyobXx80Ab6lgcAez2zGlvNi1VC61+PU7K4D9Mb2ujFccuB8O9Jj6MWYgsXen9
TLSmO5w8QRmbemFMxsLROebqWmgkH7H+ZiI6QFw8BmXH92pIa9WMikXPlwnd2i7p2M36Mxe/H6MQ
3GOYXCRUWlKDZVy2TLAbqEN4t357Wc10G7S8F69jebKEaRsTRNb/ZmSyCKleHuPbJBOtgL+b6h1o
bv/yLrX6HX5DK9QLwenc9T7IVr9B8AHdAf8L+3ulHqSYl7dfTbpwvGrv2295vKMqHeGP22S5n5+J
gqlmlzvSMqKvzzopKimAD9RbpQnwUtKMOsEO4o/wRad+8lud27sIQ91h1A7wEOv98GC9mS9GmIKe
IaBAxiQdLEUNTyqsVwIqfOdLeTEFl5xxI7AbWZeieel9wxRrOwb3lvLXSm9mop3D9c1EDM7qzmPo
LQfyftt/fbxqmJkeFrbM5lzx3HAX0mCG0nuAUPsgWmycahc1OEAiwebtKMgrMuvp8axM6tDL4u3K
03TaDaS6hPWHUAbbt8xyxfIH0mczHf7Nbsi1zTpc9HXnxUecNg+qf70V+ndICqBE28G26jqyyywS
f/EYcqhdwbZR4a5koMbxuSth7ArGJH2ePr0itiP2PSRWu58oPUx/dd2Iv4tiee9NJu1eaMXWirIh
vetHgWmWnt0lywfFeV9bdUvA6VKvRObeYAFiEjTEhMDIh88JTt2tG1tpYlTEoUkam+1Gb+DhpQWp
VIz9sltqZ4JRKWjP9aSXqyEFBdSl/Uljj0iHG1kpdH125DN0Y6WbSLDyURuaTx+RpJ48zlV4mhO6
J+RGIKiaLNUDYv4FYSncehQeBDlMAg22KjUcbHwEpPoL4u2ujv1fRi9MozVRSzHMuDowOEJ8Bxa9
Ntmt4W3rBAmudUtrORb9D5kfkogsj6jJvNZSTvijr8S4pNYadDprUh10VDn4jBpg6TKHzr6havOg
2Gk2Wh4abAaE5gp5askI4A+2JQGrBGy4ov+GP2Ca+TNQT+af35oxM+wRxrBBm0wOd23mRlWRGA6+
lNSfBGg65G3ObacM447hUGHb6P5g0BDiIZQlCH5aXJ9J9m5Zz+rSbGM/pXgB7Br9Ck6fAoGq3RLA
p+iDFzM0vZ1M70+kK/IuUT9PN1S5UigyGUusjC8XgBO/9niPsFUXMnlwyQVVroZSR2k9kmOyV0pQ
TMraJ1aSH9r6OW0Daj0hqFHgMN7RtGONdls52h1qf4KHjyIVaaDNzXvij6X62c21DU06DpCrpz3T
I/oci2mkfTUWsQJYsu9XQbnDWsjnwem71SsXLuinZIvT2OiazIeASsMDfwm2sVPmo7eLzcdOd3db
7Zw6P0hGcVur3Es1eT9qHTU9i0BjAZTSSxW7zMNtIpMBj9oRRTjl90IpjB7AX0jCWswNuQEO0uKQ
mDy5y9C4DpqYLH/X2yQW7O0Sv8QacADOa+rPEaz0EE18+qWQ7WajbXsOkNNbHtMtPOiUKrSgjwRf
6I1bloemKGcQf34d6U/CmqYIFlN655EFnD5U1l6slV8R7PwzOF4bCBg4OeRSk6E1ZLjB7oKLHVpV
G2Uk/WdPkV96uVvSmbnDRhLHEugVMFF9Y7LlJVJBedg1vPsfQ7XFQqs0WSdKmbYrZoGGo4OHbimw
NJWSZJ64T4bC0AkEYI0HAAVi9pLhdWxTgcvezPJE0QjtfTIGGp0iKtK/jl2jVR2QVysFaefF5A5J
Bd2BBYsCQHP3XWPYkvduGvsu9cgoKz6tEey10k5ChMRr6ovFHgdHMSdEsnpDM8zhAJPwtGcIcBMM
a05RPEt/1kLpGaVo6nOjZDma8Hf310T0kMxRDdO2HAsvVhTR3O3WwTkWUWWwkMEAiXPl3BOSTAMl
soafnvBqNVr28cvucjxRWOWRwtpgHPzh/0vL3DesuTQlEPuPEdngDxsx6Vg7MMLkXA7Cjl1109Vk
ao+8Wc1oXdeK9jCTkrFV7RhCOS2hanji0zrzv80LgfcLsXwkSJXcXh6MZfrePUFDvTtKTGMBr+F7
yJPSsYyztI9LVKXrP6ptPDQgLl+rGqt2yfqHYYC+0bSrh82Rmqc4puxVKwW/+rGWNpOb7EAIbYfR
yoNOv6QSg50z0mkrLGsGuwmp2O3RtbAvsQGZaJ1Tov71N7McAHeGQosUJ08rnK6HPgdt2YBTMpBv
4l9tK3BavwfUmZN/DKGXaEvfdjIuaS4xXNm9SDQACBqkAE7LB2gws8Qz8u4w8yTHNoUO2pN9X3T3
IBwQQvdanWtglpYIPokueNIiuBYQoNAdb71uVuXQnmmNYi77EZLe4ms8E5hKVYR29FSZ6tCaD6y5
WpwnCmg4Pr4ZatzWVabgH7vco68hvndQU3WeO6bozd1/pog9SZMYwMQRJQU6Y+2KJAdeKHPS6vO6
kNWzIRERZiy15r/q3IjOS4v1VnEX+vAtNCIEXnsiRE5aRSPB77vhWbmcPAy9Z+nnk+Ma+ioCfUZD
J2BD46tKMPZO7fJOeZWTOMIuDiEiqN07dmyheVaQqE7URfC2yPnmCJpB6gezHDbi/wWzUYQDk+B/
0ecZ14cCG7rkQyfReI13J49ZodbDUZlR9aZy8l6e8dNuBbV0y1dcogDe0XDLtl/l6bslH3oOvxjj
dmZzzKD0NGBRhNBs6BPw3ViBlbk9prpUQsmXOunyB0jwwhdydHghfwNp+DHl73BxBng3DR3lnd3i
Trx7q2QsorD6FImmILkIbKCtPfTGKtGdstbFcgOfSdkoxOMr/fSPUyGMm6ptX+vFsC1A80oQvmPF
K+U2BbAKJiR4aEj/869l1WGYVC4g8aTbnIul3kUco4M1l2vQxGEpQsqMuQj0AHV1uX2GiYBELxPB
XtHn+TgX9/dqxkF6keATwFHDxvA1HRjmXe7p8x8hsaFRb6/2QFT3CcyFjcUVrTTUgLibTe7aIeoe
bMoZyyl2mBG5QETmevr62DBZ5SWpDjbhYSaa4t/tQSTh2w83uYF+T9qqHzAj+HiKqz3Q+GpSD3kO
nmUTnO5jrxnwcx5hhsfgNGbPJ8VldfoIuxgVxSa4TkhaD/QDjJrKHK7fEfxDhbO2JVtYpF7NrgVw
jXmURElpOYmbu5HL6YFtsYxkAu0IRHHdYzjvuNI1WtopClde2L5csyeIuUjAFHVXa4Dc3i7e1vFn
pTdUmWa+7IP7mfSKxKr3aGTGzxd0tdVt5rNwf4utcem21WrFlP9EONmMhW+hpmwgdspE+4eGCToQ
p0GgDEAYzRfz2eOSQ5HXXE3FfJosDx958PtoaGNJuymNTIr+gmESBcISzEYpkpm0zY+H7vXApk3G
07mMWOVIX78JIEpoFP+UJFyPLYuN5254QjHPM8JGGuMHNYf4gSuW5cCj6I0/wa1+vSDaaoxSvyrn
LOpQMPHCJkX6j63YLfyiWEo+9u1me2ncSChJZQp78RC6zEt7OeyEQw/ogXXVQzUlQ8gPCWufSbni
KmHSdZQ89UByRrw00uyJ86FGjmGD66YINwVfrcnUZEk7vtNf0EO3XewaJY1s0u3nTG4bpl+NYWtQ
5wfqHf9FgTHimsr4WA5WItmfYovz+JGyqJ8QTBf42oR2y8lgrbKtIj/cjH03miV1t3fdHfCl7OHW
f38/DWxh3C4Dv+ghNl/PIKzyT1EWBpb+VjLaZQnkrqWA78EXs8y3LVJLtAvOFnSfs62EaQLc3KLR
9Cy/y8oBMNHix+2l5GFK206VYwrIvn91Xd6wmV6EbELgGrb45zn05Hyt9rq597tRo+e5v+j2EZn1
FIaEE/xFBUy/veGLftHtgjQqFCEfobCdZ+uMljj2YLUTTqj6gFZgPAdf6clr3L65cCTbp8rvd+f8
0Srof+ZT77FBPZWTUepQsm50PAbpe0bwND9H2RUeAi5xQJHIMskPzEsYZg3XdatBbwlaaUBJoCBo
VEXQWndEo5hl7wj78PhhHkFqG6bMf2O6syCry/qERLi0ZUcfeF1n82LXMjWXOU0C5vAG1b5CrvnD
N+h3Ee1feoAriAoa1cuEaI2U1Lr/VeTCYcb3ZqbCdu8guayNpkX/N5HGgmwjI+rT6ihLM1Qh268i
fedk0kcDjcFQLOZUIAXTwB1iUngUCuxHN5JqChXmGu7KZ1B3PRWQxvoSPdClcKeybAOjTnzSR7lA
Hm0n0fXVnaJvYfqvxIi5JUf0z6pfnq+UFK9RPRdOIhyiN0VD9eyL1e9LueqWPmWB19oEO67uqS1b
BOwuo0lTXgu1pCQi867+IisPXYIP3Ioz2mBhI96EuZKcGZHCSv2MsscqNfgcIZAWcH1diXpt4dVU
zfMJ+/fWWIvRA3HUP2TDiYw8BJUOFPIxE8PCT3VRmbXx7aclnaSNXp23sKY1ZgmJM9n0lpYc5OJ9
p9ZAxugP/zHbz3gzawWJfrugOn0WRSSuc3J61Fn2Vh4cLyZFBbxg68yZCW5Lcp05Rilw1pW7bQkn
JPRmj3Mp6hom5L6eRMIqhexkn2j/kXSN87+wzLzKAMdlpe1ZwxBUbRgSp3YM1ID8ZdjUG2YtL0hh
UFRXzJaTrjgKoLTysE6fl65fGMktuzBT/tOmEYOHKL2pQ+mW8QQjUS0qFQNQ2CqcFXzz8BXYJ9sc
kg/bxDZS9tCUlXruyqC8fdSnsQrUlFd2PXrglE8u9oRjMIa2k/rqTh4hzxayQZ6oXkZcNUWh3lOa
QIETA45THTPb4s5iRclEq0XrNIl7Kcrsmqf7jEegtS5FbRyVEj5QNxtVY9XXbwnJEZjLxR7RbxLp
dtj+bLWUTQVDNjekmoz1HkMfAxBhLyXlUc8zWwoj3/Z1y95nGJC4a7yKlglC+iu/YikWqcYF39Wb
U2mL2OVMxs2gMDo79T0d+H9QZ/I50qpRhk//ripyEDSeqD3HHByc2mmoDlLLt4r3Sa433BoKpRlv
pOg4hClJ6o+P+Qkp/HT2Sn4ksZ9t6aia9xk8DzAE6GfnqgPET1QaQb+f5I8QUzFr+ZMCB1BQRZCL
Gue57gNF83RLq3MGU0eVFoqbBzsLUVa5Ov4QUDOov3iXQYmNMt+PfjBfzqEDxI/tzf7vH+o/QpQe
xOYQ15p9tlADT+cbvp1l3d0h7zFsLiWgRgcYmlhvCyJIOhIiYy/Ih2g4yk/a8aBNZqmIRiZsyTpU
i1GCQAbSJTQ+LDBwRmkegx2HsybRgFHCMncpPPQDLIdyUd+HQ5b+VYFU8a/jEtoWJxqktJnlovZC
LkbEwl92D9qqlvDQd72HPlBTh5P5qHdoRbkIzBbc0SX+lhVpQiW9NJBPQ8f39f5suYAmMkK9P5F1
+CJQQq0aDLX4A06tYozrymXxPk+3TjGtm+7CbUT39xch7ZaTx9Jax3dhYxCl4lOs0IV8Fp8glPvS
w62V42L2nTt0JGMmN+snIYmgccp2bM5+zS2E7SqbipCLYofjBc8nAU+m4JgGpcO+vpb0Dv8oas5z
MwTheazItz6mYxiaE6Pwfl8vp/6dYIE3TaXuaaPo9RyqXqOSWFy5NOh8KwL2N4d2Q+op9p/IXlfW
0C1/tKPKqdDV05iczyO2Pe5aNaW28T8QdLSK61JnnXuxTwugNlU5A8VzzioOjVudgYhMQFFG4ZNT
t/+Yn+SypAv+WbFWXWrS7/xjlLRbZ8Ntxuf6YoVGoyH+nxfvxnnSL8rZwSN1kOfhYENV4mVCX5X4
joX2qkUWeoq4RzL+BpFljC0AJsJbM+lw5wQnLKKeY0ZgT5IpSVHlrj0y/yIcBE5yJN87o42ODmIJ
Vd0+OlSqtzZWA9tSkveD6vBzctde+lc0kETbUYAVQo+egLhxDHz9OMieHE3WiKE7gAqQYrNgdUtk
NEenZKXwETyHdwANbIYC4ah6Rm6//i5i2zcIXzI9iWXdwQOIQMGSjXn27K++3/5aJyhLxyQGEHZS
5vkbqupWa4tGWB/ysganGpw/A1fO2zyu6mmoaYCQWJzdkUioknMP/xLIrZeJk34/CRZYIk11FHZ4
Sj2PyS6plTuj/LCJS8wgdzwZwmDYbHOGEqFdU9nLLfsy3UFVysYhupSkxtzrAgx61YOoFG5ThDYB
4XIt6xs7ClUNJo7Rgr6fA/6Kum+D+GlRTnWXGKk1Dx0ZlVNKw1oVCd3v/8c3+sVEDnz1y1fKFNUW
qoXk07OImiWeoz6beZ+8I9mnhZ2NHxufM+Pz6qwyUGIcVLsxIwhmTYbu4uBpS8TYVcr6NHj8+xwa
1ugvJovqlukW7SWtOubf5TGeEQigw2FUuhu2J9PXYIP5Ce2R0HKP4khYhW03UK0qAcExQJFF3IdI
DGDLp5gH9SQn+P31Go2sioCiIEeIilBbpycU8wrJNSk8XnU48D2yorjxOD5lgQZnuQ2KjefrOyOQ
hT9a8tJYH3suF7qlRan66Xx35LtJkPtvrqUnda72OsnfF5NrOqhNSNGvcUuAjBOro8JO76PA12TB
ElpSfpScRIjFLGLpcz7ZSEwdmrHzCbXDliF/idsE8ojVVW+mRKOCIAeRr/LMMJrGZcFtp0mJPxEX
BEQCwKJGC23CQDXbQUBq4BDaG/yJyOBOLbJhY98RCSeWOQ8umQOvH+hvYOsm2yx2+VuN/yhskYgg
S5Kpo1IGwiYEAbpJowCn3Ex7yTNq3ZPuiblGeai0fc13iHwNmcWHywyBvfNJKvDk5pLOmc9MWpg7
7LiaKLNoE/0NG6hQ676TPwppsgFt4MfWL6ciUnFNORd3GBLNQrm6lDcd1LKh6sdjaYsm3FRGqsO2
Dx7CslSoox83gaNPN8rtfX6r+gRrOSm4ppF1etTVMnyr6fzwyy2g2GiJlVb1+Bs+MMWMBsGEYqFl
L0NSWSkWxxzXRjRImBeukIqR+dTzzVlRtkiK+AHfDiPDqDUm7tlBR51/qIEEarLS0cW/RaD/4C5Z
1KEG8YcEgKJpDY/NQPNsrUbhCEZv2QVqhayWbBVGePSjeum/HbVNCnV/fDW0MYzsr1+yAir7kLdA
+yVeAvH13iaoMoqsxBXhyuHBApZScWjyLE24+DXRUZWPO32kz1S0mrrYbL4pnm9l1i4Hxsegbz83
0urb+PaG0SzNwX/VeG8BqEqo6i9sRnN8Q5P97jLDiHNhJXq0VF7t41QE42MrBvN2xR5UnOUe2CLz
ELA4klTaheFUTd59L31OWoVuLzE0xCQY3AJHsNIKEHTagwPn2kHfHLTX7MF41DK+VCghkplRtmF5
5oG5q+Knw6aOA4pthd/fiE+ptvrY8JeoY2W+tjgKyJcq2XBFriNOesb0ctB1Q+Poccgr3l2awAx3
Dr+paTniR5Tn6owDDqeqpZWLhZbyWIsvgL50vACVIw4iXe6TUaP6Jo1lVNR+CsCFwoq8Bu1YfKsM
pLr5i76HKxrWFydUNoIXcxjVAarhpdau2Pc6roKO3f3QeOTAP3hhae/NvRTNXiro9wdHMIUCIa/l
72RC3Ti3/eBbjjfglzVHPZoblZHod9o8huDv68tX2vHtZeyzqFUhRdMkhG9WDpX+/3PFLO/SFdnE
mpyf+y+8xoyWd25mxPZqjCpEP4CiHmy2oKzf3E6QQYei/TCIMoSLNbRdThAz7IdbiFXoo0k5iPsy
easWnHByISdkuLVgH7l5jp2HBb4BoW0Kk8H7n4pgK9yGqTy3TZ+E+BejwmLNV3F0D/qIM6gmQiQK
nP2m6W5OHX3RHhydxJqgM/nsYxBxk5qLEUK6RNjXzwPFYiX+fPQ+UPeOLFzVkEUN+j0Nz4E621nb
UxQhy+DSnLyVONOPOxLRNzc1L3VWDzC/06PUQhBhs42t/vSvrLTZJMz4jBm+yYA+oVvd+tZHn7tj
2H0WOvn6tVq8deBSKDdmReb6ppzaMfph5A7jc2slnaQ6hamDwPLUpeurncPPWkTHrGZIxW88OrhW
JwT0txptCX+nlDVTe3w33G9oawoF7uE8QXdkbGTe+I/PMBJVyOqv8u/mA0Ag57RPIUxUVNT45wxD
wSNetIA4wNLDX+CDZiZYvj/zw4M4lBqApvLWojHfRaud2bVLILiNHaztoZIudcpY3XT9Y7kxc+Ek
tlQMlO85ijRrlNMakp7aVPkaztv5un50NNNCFRuNrKFO55448mh1mhJKuQPjnY3Q7YTA38b7THgY
cW4/Yw61apM8mTW8HhgGJEG6ea8swIMqNeHy6pkLTVyqNQhBJXiIoisKDJfdCvazp4KxhAg4G5Ab
2TRlVTIXjulPa/EVyUdyPcRzRXqkE2WpgxbWObNux6QrbFsnadptcGIak1/Awuu3J13xXNg6WxXK
KXEGYUrD6XvO1fVYfYRZhnkiwTcw7GRyvqPucaPyoDIsX7afTP2JspubURq3yPxSSocMFwlrF8R2
W699QLdwgqDtudquecFbZL/ODLklebkXhxSXriJjjQXq0a3XbuV/TiggdV1YXWRtdnVCARUfAmOZ
YOfkhKE8gcyYvpA6NtymNxtwZX6AcQ4rU1QnTkZgK51gGTole7fehEzmogRnOUD0Sj6hEMilcOtV
gpjc7c18RMUDGsuL0wA411gyO60SS8aqbVluT/zH/zvAMxWVMkS33OhU2QEKXJD3efP6SaRmOZ5W
IDvuuDOz3wr+1nSzt4n73PZ0it5lPbDi+w/NlGlkQDcGGrZ9+wv8VXwH/gHv9jNoXo7LpO9F+v3M
VLD2lYOU6RdIFSHenBy3YGlJFe65FXFLd3xJ4WJqdvuvAL1/96u5gkAcbiW1ONWMp0vYJ9chcRUN
YWGe6FYMqmmqdyMrEB7oPXbEvbK/ivCl7HoXnUhXp//+wd59BS3MxSGqCZoiT2OFZH8895lAtahb
Z0sS6WvPopoKVVxIwiwo2b2G9nQzoZIJAvLRd+mbxzhLT4eroGP0oX+ju5VGXtLCNXi5Rvd5frC9
luryqxaT7uUOTBFFGUOd7F+iUolBiA0Sb+YP++X47L2Jae+gs/47liRfakNApwrkCNW7ir9fPG07
cWpKRWvasdwSONaKKs38Oo3dqUDguhEd+varDrXx1JGzHWaI4bulfS4+zZRMxF2LX7HcF/s+1ZB8
FUVR5QMxMd+8XLyPAtE9CkcJMeRFef45AgZkyxa3vscOmC+ffYmnEvCnbZLs32lWst16QsaFnbKr
PiBYlK+Pwg2WH4yjMybfRczDpQWaprW6AKxl/EaE5ye4vHnQIFM+pYkEFRC2WuOuMI+7gHbZ9LjV
TooTunklmH9j6KRrfUktV02JRHpP+t095n0EJz/RP9aV7xF5EYkjljvVIWYYyfIdbxBk02lFWHAQ
Eg/JyJmc6P55tLMhTrmgpaY1G/5CHOl1IR4Kt3U7pesTCc8xmxXsiJyrNNvIa44ZJRe+ow5MkXnd
f/Jh9aBEWC8kbE4x/Ew8OqoaKpfFc6jaDMyrV1DtQKbm55YvnDgkGkZDIVWP8zQtbPGLCi14hQm5
/hQqzdDfT4PSHxhmHLe3oCQRJ8pWFEAhv0GYoWKH9YhepCQuo5WDd9yy5Mh1+U4ayStKwOH7ieVl
rU905VHNN6DXLB7fmH4jUIO+dC2XjyWIdECzuKRVPTnE1Ho9FBnPnvndDTmOZcCBs7cC64WXFYDx
iM++0aUSzZtJVWQjnylxZ3MLjTwOM4O81wqoX1k2oh/Ot9HPCyVm4Ugl3QCAm96yJsBoYPNMJ4FU
DW7kRfR+1+u5jlq+xVDQ3AbuOK7vBiPrwtKccIn+B1EgHMPOMLBRsPnfP8pzbhfppQ90KPKIkrZT
TWUguc+a9pmmzTUZUJz8dFiXQ0SYMKjs47WFb+6AidOnf5aBJzqDuJBJ4TlqQj7iTtS++JGb1M0g
SFwA5gli8uit8KTIQMWU8n9h9Tj+ijappoWqQMTeM4FYptJujhVrISJtzTnWPO0Yq4mhqabBLvTH
ehw3UYKAYMIm3PxpIXUVMWDmksU40P346JcGUFT0b3DbnbZkiCElzMJOAeterKR4Rr6R4bVXcHuj
MEA2zJrcmKypP9HcuQ1L/0wk1KGvtkPRsfQUyTtXB0toWTiW8o18yXcV6o6kZZFbLXcGpYFkelIO
uDgTp1ZOkgIOSgeYAI6LQpqj9pM+E1IMhxoKoKGUEDVkNruJJSmZf+X2IeRa2NtBNVfLt+OsE04q
P7TG8CeC6Qqx8xzIu+55gjyli/a81Z6yoV5du/ZAmy2n5ldxIFeiQLpSsSfHV50ZOVw1p+HrMcBo
ttVXF6iLF1OEBMRKKdXe6X1OllsG3bCaSrHwiNXpfEwmxfm/kJraf9JA6nT9L7e96Kfs2e/NMFOf
mKAzEimEui3J+/6tb4pbYt73Zv7co8PHV03LlYfQjqB5a3ZgeHdEGCsOmFt/bHdoH3jwxwmreCQD
HfgUCrV9Mik2O8e1v2Kn4a389/0tc8WjwGC62UDxuDFbkx3LabnIP+KSdKlHs+NDcUJacCDsmQKg
Dxi69ZlrrMVvCzOj3FNaBZTLlhdHW+l3Bnk28vcXOJzMjW4HsLNczZAvvl5STWL2ra/QfgOeg4zx
TdRFqs91MZjwQWu96ocw1Wy9D/0H6W3mDoUHx3c/73gb/yWy1l07ODiu4cUtNnlKu7OmEVrPdM85
USRsfTnuoSNZkNZqBDKg7Sw6XrnjvUMr646hRhwu9MW2A1HlQBnFXSJ+Qw768ODlzUtsfef/Cpb0
+u5FnMtSPRO0tg3/U/D55lskGFMkJ26BzxO0ZDr/83uNmrOv2RvgA2178J+7k69QLNWwt42Im2Eu
VgyxWRgvzxlcO3KSt7N106Z3S6xrAPliouu+9folKCEq/dPrKrA97CtweLZbJWCsrNFL4Z0UEyqG
xsGRZQSvufYgNuTd1UkAa40/r2EF+Dhwqe+/t9DCTkMRRAwI5WcoGkOe0+SAwZ0jch4J0EjT7Vh9
ACSRMIW6d+Wn0ttGuVeXku22sH7kF63SK7SaFg65ZpdRsYFKiwOPpYbedWW+3Y0PsbyEXU3ZiWD3
4B+mfp1kEFySLcoe4kj1FEn4H9cQU3lK0/dSsn40NOroirS/bpERhkmMUUL8+aXekPTb6sA5jOI0
+QkIg6kOnaE+xZiCjdF5lgIXeh38BQx1tSLpCDm4I1vSkB23uE8g/COYV7JMs+VSXZtshQjhXx4P
eeheX0mKoUYU8BDP+c+oiPDkgcxUFwmUoXhue4NjU1UPYNn+idTc2nlZZVzBtXT3LmvUJNQlj2fF
6RomtQEGXPtUPSn1qA2EwOXnyLDZTkK/siDdUYPKDGkhYJk24dcKB4F3rDK6/gqfvw7Eq+v4wsGe
kPE9uWDd2WlBhMH7bJr3j2ySWHAUV1JnDiEj4i8KXyiiT78s8MTOZ2KgfWRCgJVIOxlVxgEuqEn6
kPkTWInisqHEZ1LANrxkLtgro/4SZ/LMYLxu2mY/otnZ2skjEifWbAV9N/Aei/tRX4wJPCOYL/cE
tqDKt2W/Nsv66oLJgoCVX5csH0gXfvohVZRIULI362toa2jyhjrx2S5nC8JTk4T4xcRYF2tKcsk1
512/CZaPZplsP8NFZi/HZXarziWDIYHlxOHrKNiCFvxcCojSlB6ufykUyJnrFYpC3G0cJtu4hClZ
69GmexDUIpIwy4YcbnMC8PYFwMkO+C76Z41w+4l82G2m58KlTyUX6KKU3ayH5TPVLVGW3zrazQhU
ZKg/V7oRzIY/o9qqjL7znPbaXFle8djy5gjLkUt6S71SLH+xz2h0dhzaLe4QeeKHxLmIUVGRPgOz
rm2H1lFT8ThqXGc2Q6FN4TZ5tf1p3IjJaikmyM05LLACa1BIjzHr4X2i8DuiPSP656LWnw3INUVo
v8SMYxf9TVuH637Qmplh2Mh9PRHBHNpvLEQnCSy7quhSnri9RVMXhYVdXSN3gPfT6WxzkCa8650d
UISy5kBeLGN+AAxhf8uL0fU2MVL9StML/FCxG8wNJYQhbB4OG19aGJey2rDZ2eoUWiX6PMIxUOhn
orT7H3MzVqfLKjLQCh2kOq4kDVkI8CpybjOoSNned86dFMwKAyCUm/OjGYEviELXb0TvzaiQ4kK8
obiN+A7XlYF/4+8bjn3OUxohP4GJKQmkslwmFoBisZHAg0FTY16YPd55GJUhnHpMW/lRWmom6/4L
I6Yk1EQGxFWuNnEtH0IZsVUZd8oHgEPaJV3iXrqk3KWcrkC2bjnsjw6CwcfXpjuhXped285fDB80
aREST3ukfFwHscIXNaFsLOYVVAlLSPjpbSHDwPQG0fCSyZukA560VnJU2Mb++AW8V+b2P3Q6vHoe
NwNPXCu0F7PpB7VSed1kIpo4cAhiCFahZzq6AivbG0vBPZO2AKT/XwtM2PGdHC4YP0Yo+M0GDjhc
P2DruMLG0OjLvLWPPsmMyoJ0/Pbx4NrWYgpwzsHgL5dnwWQUmtaswnX5kYaaNEor7c+4/fog3EZ/
b3hK/RMd4H/0WiwQK6VL2yKu2bSMOIpKAvXpy1cXt2qDlm5cO3rxzTq0LIjT68iStkl6QKCY5r39
RfYl6vKJBECtfntAfOGpXaA9jCeu97RLusNJo6FeGsE7nsmWRTsMNc56j3laLp0r41N9Tnvc2TZx
jAzgXNkwJyNI48y6+NW8kMDdyftshaBy78fF2taoJQbUe10v1k13CfjmHC2fzOagSL/SAZ5xBk+7
LtY3FQDLaZBoJFzbZM5nIOTNoorOe39rlnt7s4PeJGHYum22eifSLio7h7Y/IY3EL51mgJPU6ukc
aFVrLdrMEI07VXELho/rGs7RVxxf9QS3C00/xiQNObZeIyP5lZh8r+VUhe+5rQUtBXjmG34/aPnO
Ws+Tg1OTQAmvCfnOi+nhXigu53PPZ2jKJLvt1g6XhNstI5B6kjgbewBIH1bdJX3rW5/wFF760kaz
n18K+j7lDDfweSAp2F1Lv1g1PGb5DQd+SzvsrTi8UxMan3DlyfApGSfw/gbgqaz8lZaySOp+Srl6
MJTHu0z5gMEb2Mfrl/068PiyN1pjk3SoGdQhKH4/ZfbyUBWB4hCBwLvL5Lm1iKP0+FRGTDpeuk7B
lp1+LBuXybJ2kUbOnKuLRszazmALj9zWwKJgcNH092zTNrUrxZ6csKHpVRZ4lE4H4b2LRRcKslXf
DAwmn0s0qKjhsnD14vjTRnPkA+HePTFlDxAbn9SW+HKmH+EnTfDwOLrgtBx80V/guH9H3/5RQw30
ONDOzI7tMuMWxdXX2NKMRv1jP152hwFE9lVn3R/mPTRA7l082iRZPtPL5qKG12tKN14e0OG+hxzf
nJ4D4mz3Ba/mm47GStLvVJATlPdmh5OrWNdbZjwCk7vZxatkeS7aFxwtM4Ptxd9X6CTV09zPouZX
/9KjY88Qr+82PB7bZLrB1GFT8HTdiCnei3UvjDz3+cGba63K3eUKMu6S+7upZBAROVZ2Qgj0wIov
cJ6H9inf1oPmfrrebC7RBglui+xwh1NXuFj6fZClVFw0UXiwbZj8/oEL+u9H8yhjROa88tXaQ0XT
FcK4XkadxV8Qm16BqkseC/6k0s76xNgl4ap6GR6GjgrDKMGDxEX6ehm2woVr1eU4ComyPbhqfRXx
I0vk16ChV+jbx5GN4nplv/63OdsTxTG5JEVCwfjfzO9lkphwPiWlHlx+5b1MCWry2CRR44yo6jOB
wxx0pu1IqRmC5L/GYPbfPfzRInqVCQa9Qrbw7CNB0/k+WPN6k1fc/a7I9G1uTJGdq0hUvJZnXgNT
dudeDsocfaEI6uqS0TFfTIEOumHArVSPsmjMfeF1HZLOXHENAspYl5v2wRhtS3mRP2ctBHuw+BTa
pbm3cIiA7ZyhLCRyq6+LwoBCYr2gYM1MoNhuAGfzqcCEBoRyWBk7pwfFJjIPhF7jF/bP1cgL40j1
jWaDK07sVHl3nl4lew75x5YWKQVWaPsg1JbTjmZDfEt2yt9rGw3zV6vYvngkjeBq2CkAlJPxsdM9
Dr50dR6IQ8gYuIgiUyXQUmyl2WM2xDMvlOMXuS2vQhg03dYQJVYZl+3G+7LEZG/wswpr5WC6M3cC
v0FL7aJDvMvK+zgrm8yGplh/pG60oei9cSLZ6MQbZHqKrw4nlUU/To9fnlMdc1x9UxZJhkT7m37d
iNYWSEDyCXZLV5GWsdUaGi7PutCDURv8gZteh3rLf1rZ/3xNNkvbvkgtoYMUNmo+TneQ0rPlkCQs
tQIjf5eDFWsDOgmF0bFJoZo0Lu0JmXNalRCqW0/e6CY0x8FW9IXcMmM0jP0x1n9JTOAlZgKyVVJP
CXq6jrIZhO0tExzdzUFb40zuupsFYktS9Vrhf6nlrdJU3bD4QQZBUgxfmY5nOcUumHMvL83AXl5I
/z6jjcrS5oithrvrzD3lt9OEC0/PA7r/m/Ar6QoBx7NQEqzwr4eVyauNTV6K5K/UmlhpUsjQ3bZC
aatS+2fFucw9irjiTqVDQ8D6qq8X72RznD8C0FnM53XGCpKBIlrmWBPA7E8ekcOX3gj85iVEptK7
bam5JNP0ZveISCbWuncfnEtefSTP+VRKZH9fQP21L9+4jTiu3evCzuqXZA8Aq+tQFsRso0JjPQqU
IeUVY+VjkSaItVJR52t/y0kRDtsdWGu2T6sM3CJyM0kuOU4CgKuvfuGIhGA+y1Ru7W2D1WgktRBQ
9Bp4ggbZZd2jgLkEykVKQX+/CWEHG46RLAEUv4/VS1sYWp4/zCEOAHTBAdPGVPDoA+ZhAl/RQkhQ
HuoGmlp5E6QxFtDIPVrHkto/8g0tDaiANlYei+Q80NAEbSiUcN9QvLYXSeMSPuUS/+DHmqKGVGe+
2yYH5aP7LvWHPjlIflxMp8Cz+SZT9ddSA+jGBw8v/m20Bb3RPI49VyVrMV1PyY+WTyYsuuQOh391
kXH5nGWHSvopi7dAh4AdDYvp1nqPxJ2093fMbINww4b/eFxbiJK1nxe85JlwgwAFB1vXf9gTcI5b
JSQsNUHe6Fkvva8qLlq0H9CQ0HyhbWGqfZYKJ2N0Lnrk/qlaOIpcDUdVPK4wfz+dgW1g1kgJTAHW
7ldvDvqSTKtcXxs+rFgt+GIHSxQAwWJsjBRrfpN+Dj5ooCxRy0YWGW7qdSZa2GrF9AH6jiqOO2g+
TifVhC/tONmDXGXnj42hdugmpE+7Ppp9rV5WRqKKh3u+NClSP1QxlKy6ZUq0JgZZ3rOqH4RPnU/q
fWLJzvLURg+8vJjOhuhHfKCtxhgn5VxVUUwgR8CCIN5cxLgMkjUh4D6sCOnnb3dJiTfjwm+C+kjn
AUhvy0mw4qodqHVzirHMOgqRW8xZxovKxCGr+9+MqHfBmpe58XUMBnf5oNSIo2efUxqPYWme+qNs
xEkQ/ow2yujYbY84sZ0BgIXMUoH3CVUESTogsbpmxOTZOar8RC1ZN0W/dVeLhbpDdn0yFCAdQ3pp
jOCH7EJDVj5wfXOoB6kftzJAoDtixiaVUJP1+eQpfkVgwUYfl8wKzaAKuAkECK1EFYBADYqr2pB4
9RJRrKUGQ15sfJEIGixAy9EtthB5VmkjXZwUBj6yyCeOXJX0lSwcUlQ6Y3I9PVtoLDkdApq+xmZD
9JuN88NNBe3+b4XUJFED4bFdcLyPcyAWncc/GsnfMFGj+EBU0AAuVfGQ6QT0qCE0FkWz4qok281S
Rc39Ssozdmihkh6TnlFZnwNpLpouhWPYPl1zVd1CAlz571MTuMWZsjnpY+vX/hy98I/2jfZzkw4E
hAWT2AAdxjRq8Ton3PZPxsnjZbZ0TZafs5+oNHOC5DSyV06b6drBJZOoKs9HLVIgf7GQT/51YJI7
7mawgreae0LhENxiSoT9WSXBgV1TBbTuVkpSTgdZ/9qonmUTGp8SKTs+RqofpYc5x5VENhQw/v89
6b3Eq91fLija2OSf3dzRD4x4fDDxH2P8Ld20uZpfnx+sPKqoHdi1J+5aD5/5+kzNB54rMQ2cKeZJ
rJSDRcxTd4qS9t/AUKrzXC0n1j4SHaId9j9Ud5C/n0WIHQIJODcEVyBbW0HDa88NwMLg9hQhNrLC
RveyS/VVE/VFDX2vBt56AXpM16t7ToNxnkX7SRcBmEigMbof/R0hFfJgITXGgNSuZKTvZFd+8Zh2
EmbZvwhYfVoJoqlsLxiOjrA+X/bbghDRIgLQ17AEh34FEjmAm5LFsI/T/3kFBz8gbaa4Dxeq3x+a
hXiCqmjyD8tYEGTKn3w9Sx365frr4XwFLoFRCR3Fp/SlE7rCVVwGssNaXvx1napwcPK2uU0+I4e5
5emjtTyaUOI5Omnazsatu0ScOrFCmrORhQa3yHiOujGYe3kFOIdSQ8pRZpL7n61pwCRtjEEyHfKH
E75+xNTz7OeR1xB2ImBygxbF0hvLUlBUTzkb23QH4jMfMETk/1rGiZQr7Vzdl231XN7DpGYyfpOm
aTUMUmr+Bzkl4hX+GGAR5F2FN1xTPioVuTlc7p9eRfR28/Rviyw4ZbtqrzO2lacWWmrBuMF/l9vF
Te0FaolCVUUcR3Sq6U6uZz/jLq81NnkPoij1I8elvMeUUVgGoqqR6xr04wLKnopHfdwBGcUMkfS8
AZQSd5P8Mk82/MiXYOz75ePUqdvO0L72TM2u8RA5aPilz6GvDvb7je9Cxhoi0O6yyWKvNOMs5UVM
riIgyS3i9ckwH0fnESC6nJqjbN+h154T4wPKhmKlusGxOR+m7qCZTSTBK5NzzvfUHHfXk6m6KIwn
Tmn7ixnORmrUCGQ6+oeHdcD72WIx7zHp6qGU4l2bF3t+7bkUOT0ELOSvUGI3zyS3w2Q9sVE+JU5p
g9pKRk98owOktE6OdLPuo7qRlhHRl840AOsY+hwWnQXRJD6CHKSxBeHFyk23meR1gDNR68AEnB19
r24nVMVxP0xGCsNFqo+tB/YKy++rKEVqcoIwtYvtvM4fzK6rkLxkFQhceyvZcSi2wUcS9RPHimZ+
J8bBTmJo5QUGzeeVJhJ5KHK5Cf6swl0ekYiBfXYMPtFbhRitoPx8xAa8JPgfA6LKmM6he7mD69mM
270KxFC8GXd5vi2lAxHaHjwPbpcYrYL+hNTT+QvTbcl7yH7HsF7dZlbIjrFXFCPLhrhFhlTY6kRH
BNs3qB1TtNfuDjSMct1R3KYVfKnjH+gBJnFkckYUTuXlyRrwPvmYZXf5ub+NWUobliQh1HXrUrxM
m7zIUoXwquQvL1osfMOm40fywgbAJlzZ5dVqIOU0KXKLFt0LQfvtL9fJTq022lDLOumO64q++Nnd
q8+63lZE+XXiU63ZsrYZ/5Ylc3YoFUog7ZtnXs0bnofUoYRExNlh0JzWGYHRa9SRztLgO9RCzX3s
iH5HWhTCxJwVumQ94ph8cv2D76ulxl0KQXfKpGgmvJp5aLskkWWl8/fjiBKEBfFgSsXLbNC24WSi
KDchnZayFHCECvXNHBFiHTv9jr7MJH3/VQ6+TOUHh+KEnjCXYuJkhv2itHCZfNCxm1jP8ku/44ml
3W8PeNaj78QLVEmWHICDl+rN6a21ZjoZHBvLFpyi8hrsGmTO6OAbhH9mGgvGa7yNbfFdwHM06gH5
fiI5PSlsX2HpVjsoL+qit7vHAox9IQb+PgDuQdB3OWe4purW6W04RgoF1NMbsR7F4X/YpwuZr4Io
46ZS7wppttgzBfKqoZ6p4V09O3Rpz2CTzl4UDQMqXLFfhQlQpy6I05yi93u4i4Ge0hJeOAFbRPgG
W6J+OgQ8WFtZozXbedraFvdTdnznGT1Nwih05OB43p7qWIX7yiHXBO92udEOXaCTm40AAjUGFLhH
uuZCqwkdmruEI9T3IrdZoITTVtqYt/xqamr0A1oTGYYKSw/iwPN7BRqyxL5U5Kd7RHRmL/9vE2LM
hg5Y3Fh8rkAKZgEc+aHUadIVXuG4Ii54k+7LSsbLadrM6tBDKIqYrBA+a7nDwd4EZZPs8hvbbL9U
C0tuygjU9nK+ZqF7jNaEiNs7pNZ0lIoeDagGD+Shcgz99ndontWOQcKocAvaXrAE+Cb8LOaShj0T
XJ6fx8pW3ek1KkGgO5QrM8fBD2vC6Ygvw27kpyJQtRL/UkCvoygnJ8b1EgUvnC8gdlSwOiWb1jwr
w/JoHlVvSbsEXif0MqasVP2ajo7bgn+0FM1T8XGmdzW/M4ZjjhGycC/Vzp1eIJjQE+ydlP8w9L3D
xdlJsHNSR9ifaIjilePWY0DSeim35fokVCJspi5eziyS9wNBd+RYlaAGIp9Q3r7Hq6kJw20PjNNQ
I7DY1Pl6SuS+28MrqdyUJNeW+L3c3Pj8J1wI9o/tjxf3Qlrid7GDBqIGXmW1wJPBTNgiU6vX9o3Z
HnrjST2UE5gECDG5sycFJxYe098T6tIKdYtiGYtN4YDPhU+yeOVlosnskaK0BUq28yi0+1nL/L0t
rFjLVc8pAyq+OMwl3Ad09EvwOaOaF3YWFC9Z+0flKNh/YMbmmJPkBYXUc/usOEkjl0KqajpPxTSH
8uAFFeMP+mPKDM36dHP44/2AFJncv5zBZkjbArtHwWrbD3C7ZekESNl/VCPbadxayC5hZ/Cnzb9f
7pXsZuqMKFRWgcbu4OTYBZeRnfsok1u6D+XHHHPXQxPD9tb/NuSkA+kps1dz9YA4kirItJaijIaq
MO4EarpLa8X5ffJwpBbC0adXH02N882yAgCoOnliuPudQYOK2hk/RFM9EDsLH6JoZnwjSz5GZ4r8
E1pIhz4+0lxTLnY0Bj83li9h/NSVzgfVREkC7hNlsd55cf19wXtFIl0O7Klpop84fInm3VYNkSUW
9/HcOQx35sW0Vum/uWTY5o3pqkscHLbRBG+PTgf0NiszMuWi55nbP0tW3tageslkDO2I0rlngCtc
OXLDspBOSDSQEw+syQBDf2QWdkBqfWP1aLGG86xpOpNEkeqULUhRHN8NGLScMFt750xUbvauqJtT
oYJmG8ZyKi8kTM1I+qafNGnJ4FyP5Ip4UyMHR69j8IwGlhE/m1HCxtsNt8S+02M79CcPo+R0dsNU
i8OQ5WJIbjUXaDZpFe0ru1yIs/BAtySzMnq/ag8W9ZtbjQ1NaoWbJgVQPtbp22w37PKvQgjkn/pj
52/51ZQfcwfGxnPloWz3RlqiQfAFfZgJJ7yhpAxvNNXmQNeCt1jg+OxEGVL97RouoT781kJStBw1
2MHyAHMvbDif9kLlia1tCyOlH8oBgKo3MXNDZB2knEn1Fqy4QkwvyCHQnsFJ0XznrIm7BvBhjEeN
ow0kIRXozFK0h6Vci4MAJRQZbhnJU+VfLVFBnlMacOTd+PZnbtC5Iy9ZxuepfMcTW7B5pmIbSt+W
94jkYT5z6oB7DCwf091C2YsdqbsFSTSJCEEaIRDDrkkmdnVLe1CFV9v0b/Gv5jpJh/mZNttn6P81
N0+Xt7ZlNn+8R7JcJ7nkAn3Pt4I/8NdzlSyqFJXbNEK3hQOHZm+eFVSglOcok4VxW11dyC6VynC2
YTeAacxBAU8WH0JTHt6yl9GPAtJKne7mPVU289CNB91Qy/azpz5dIhrbMqfGVyqutEtr+Ya2W2B1
+RH6a7hi/j0TNbetVei5H42ShreXT6S/eVQmDahmZhqvUxEUXLmlAZLPEHa1CpeJIbrlPvw1eHgh
i6HPSqb4I+7NwlqcByZbYBLx/xLcOLr66kOizWBx/69/Z4Kq+Y1bpZ5NeF84wWCy1N16Adjsqg6W
ksRMg8vWtVPBH15VPVriSrE8T32kqvMQFUkLMYFFDbTaSOwHx66x5OkQRYLdL4I1ySOJMbuC1nOf
DGJ7IJlZ2/iUbocGff0WD/+iKbdI/+/LZcxiKtCUIms35Ni4VkDz2rkb2wlbxs1/DfieVf2oZ+mu
BzMpO90aRzbP5VLqtD68bRBQ9a77t0Ly2Vn0njbEVc3njEX5XIttp97RI4dQOYFmvIlnP5omJd1Y
Jc1GX9aB3FdgCTvCF9pAfMeLMGYtU/sucb75/ehd3XEfcUe1MU4H/aGRVjsNaa+0hgSbpkghYDS8
luZmxtKqXp/2oceqCN+59CtDHpm4NyeFBTGoX6UZSSMWW0VC/bGT2I35RmvBjhcQyeHur+BAYM5N
mKCF/XNJfuRhxfV+9eVNuI46M4cc87lB6VSg+oOJ7dKWh9RFMzggDvumQARwWOAGzmB9j3LnPDV3
lv51YVHB4MysJZgO+D36XJ6Fp5ZVPQ4IhogyUXpIUYgwedbA6VVVRotSHm3n9a/Q/Sa6ySSZ7pmA
ZMNB4r2GwD/CrlxLkNY5xcP69k+NLieAckrHvqcFjHedRYWQYJV0+PukO5mc4GxKyfPTITWF7GXn
cinkaIMkKEbfsULAhirDgVZ9Hu7PQVMeW4QdCaUtiul3Jt3HOTqJOf3+DZAr+ZStiKK5ebfg8OOC
9vh+oghELGy3dx6RcXKx2BhZLZR9OTCHtwLKuDnHQFEOlxWRCdxEi1Hv1+cbZaxugYJcZ+mHZaU+
cQa4Rej5qma6CFNXbhR1kz+5Em3BYWtsG2IcTqsABrC6+CSWfgCHIp8Gzgt8lgaq9LU5ffcqzj9W
mWhztHRBji5YIglAi8B4Dp4SDFTMEmWI3l7hs/saZFfiwSMIcGQ/asJ6dLiUcHuAw+iM4zpPjfTo
6ECbCbdgnCUN6aXPb5i84Ag5dvtk0sghtRj6MCS6RkZWxlQrDPWZwBqcFaEp+bHGip719OGd3flN
KuvKGjZsxI268fwfQPwFJqIO0ZcU/Ny4ng5nyWYB5dkqXHx8z8ZO2EAStt+aGtWTkFo+2MjL28nJ
pMKLIBf3oyhbOAIUhnk/Cqov6Yg4pjd5eojQFPqdoPV55xms72dBmYOJBlZMS5vM+vQn4T35TUWC
PoTSpbY9hN/pTUweIZVK4ap6YmC8NYWR8oVCl4dew0/sql419oimwELJkeDxQHQh8injtXMxaTNf
bCtvJoKo8hp+5CBoifw4KuRtCQNFiIXlgIF0mkb+AzAEGTesBuzKqYawWTJhfXZ6o/eG1uAyD1J5
4qQ4E4grOcaTv1apvV/T/7eNWVDpblWBSNrNlu0VLxlVkmjXaG1bqLiqv0Ntat6mRvn8ZYbBcBqV
5c8F6FM6D5YElIrSJV+r96dzM4bG81TZ61/KQXiAyRiKgJ+qQHKK746lJBUVy0WODFvZxZ6xSyeM
vltbN8Dj7MCtLN6YGOoPP198hWJ3LwjrYVBRAO+uXuagzKsrJX4OyUmVEl9be/Uj9S/9bqh0qoE0
y+2picgEWW//aOKdFi0XiB7zXBwX4NGEr+0/hgWx1NYHAPTCYdLYHB4lMt6pbT8y8v31/OVPwXnb
/uwX7xqpp+vM6WkpbOQ85uWEgvms59a0tSp590bW6ro3YRJIV+B0p9ZJM9Bihf1PjwjWFU+NIwFo
r2QH7HO+/Sg9WGAzf762gmqp4CdimEdtz/HJBE1GyEjnSm4P4G8275Y1QNJafGciIgy0lQKG4GaP
fDh82fSOSzoVswAkqkAXQUzkih4KT4xqj8yBXt1XxR0WddWNW9aFPBU43K4n7XcxhaMUuWvDYZy2
4D/3Cs60Uf3J1vunDxJyXlCsNtH4H6iD12JErCjKlWQB2Zwk2vaAbnVzqimQVKyYzmturwrK2BHa
CdnrwxYQx9tWWNpymQqg/QUEoM74jJiDTVve6RrYSacPObipkb3UbFLSzVZAZhrSJm4wNLOtj1nl
UBoXqUKxx2eU0l23hlNNHbmpTT6mzajBscQyNYiNIgJoYDH2ubrGjfpWip9x1z5HKbb+3wRB7LFn
Z7NY4d600l29bsyZ+widKYdA3idwyQr/XOM72T+gDfc239irhPAwA2xZIDLw5mHjIdpMx6W3H97w
YJZwwseYVMHh3iaDMI+o5I7p/rBFBSupBhgEpQOMTNvp3WcpnuL/GewM2goGmVBKxCUw8NvAY3Ks
ujCWp6hcrfrIf7+vqUTGT5K8DqXFYWmzrdOPnYvy+jfysrKsRqCO03ddkc0nMabxCTprCu0pVsaE
BrEackUSZ4pZn4TAqydb/6aVX9Ck5LDoG33q0/1N2mYfyKeVUYqxQTvhYGJARrvlcyLJ92TARZAZ
ewvG5OBL/5QKZyEIjlTHpWA93dzp49uyATzSdAhQWOpHm5S7ys8eN15rqLk4owFWBqUBHM/MbpoJ
4kFgAqPjfUjQVq4qa9th+9yCTVtlqXvC6wQozvYNLiaVIVM+9v6pEtzzXsHtfa7UXJbeCUZJRhVg
kj4T7QafExWmlFqw0pJkQLfm2EXLuhMPvz9uUtRXzOMB4c4ZVvZcLbufbgAFrjCbKEuhr5SnuekN
gW/ERwm/y1/oBkfagaXHzehYuI6OCOJgOPP2wqHtJWFpkADMoblvqRHmgB3zX09ePG737UYHiicw
bGIXWoxYwnJz9GydJE1Br3VD6WhF7R/2/b6ZGCYtqDVjSnAQEY/R8WsWqnPCeIg0g9WXm+ANuDmh
HzAvsHwcm9iKLHO3EwUYi6PTNyVQVG9PYshbjAD+xKp574r9LIsturTB+/AF+MqZVu9D4StlQJLP
0tUPmmvN7Q9maSiM3uvY6LuZOBD6zhow/pSB+xAJBPL3oPZKG8J+D0SjGU3c0+9yurVSYcb1K4MA
YvjmwKB9aUwtNmB6L3PkQQQ9h9WbS0Xiev6+KCG5x0ua90RIh7Yrw9T8Au53N71193bd77UTHwzl
D2ppJIDlLmxc/440/3wGac5bK0Ni07gPoHYd5rmVCQEt10KMJqaGs+zJ7Rhz33V6y4PB3xZ/A9H5
19daid0W8Vayzk+vh4cbErVcEoLpjhYYtR+OVgNxwTU4o2Grgcv6PSBgkf6UcZn1bH9rkARfiAEM
XtHYy3HvvyQ5QZci2ROJsppG/iqS1NPmIvKN6SYfg0w9nm8EEjgVGsxrHDo2HhxJjSlaYrf8swH2
2AuYomrODN8E9nGE80ekzEJ9HGhJtHRVBADFvi4/ai2JcxUy/BKRGXn8iCm8svX/lwZJQzoNzJkb
7fVpZWxMKD39BhLZt9KjNrt/rZYW81sQoZSX7Umkel+D/FVanoTJlM5+DbADW5wquMRRK2hSNfQV
TNnYjqQmAEa/RLjj33D7WSZDIDEa+t1A3BNCyBp9csZo6qfEBVozeSeDzy9LusCzm74O/Q8DYYv1
rQMa3naLV1F18y2AlgQYXLbFRcp9roHIeP6IoBVVje9I/bJu0fKWflB4TlrFmYk52W2SOwmiHBNa
m6SHEDu4MLuHquFqVYUhwE8ky87NcLVYsPGpcO+c1leu+bNHm8Rh6utAKK3o680PxRZVmI1LyfgA
FAjIlKziD+D6lMHU81+b8H2TpDTy37eG+vhi3gS+GBqD0yXXyLlvmWMSeK/+TbziZlVEmX6t6Epc
Yp95asvGqAX5ajjAPjhSPYe9rgHAXa4J2b6/sBTLt7ZQngNH8n7VvLlF8DD7ttFglYuHX5yTvM19
GVLXImCuoaYyHmlajxDSTIw33wi+ycDHR5ZmBATbuhMgm2EaidzrtaWJ3P7YEKeGkLtyLTMEIajU
cEeA0sZAZOd9x9GRScoIzyhSOQPXh5R/ZWoapIwor+slys+9/R7vammVpqwL60yDa+4fZr8x9PIU
kkTvWx0btdMuuynJrdS54YO3Nwzb4dBQuoZBYpqb1m+xHiBozkpWFEYDp+vnNRGVh6nR9QW1xpEQ
SaKArY1rwDyo6PFp+b/HUco1l5UyINxV0GxoGmQ0zLnS7MiM099kZu8oDAJdFNZLhzlTmmLZobNH
sL4rOSaAr9I+TW7lZx0FoPF1SEJ+MTE5kMO7tDr2CKJyxpwsJNdOGJxDJP4tJizOoHqJmkygB6Aq
p7Emlb/7UNXC/Mzsii2HHrrR5WnfyQE7ejPaNKnJtmJ0jhwpa96O0hO6zWJK8oV8VVB3whzK3e15
hBmBE4u6Dt+Yc5992BZtBx5sMIRbjlp3IWYYcKzK0Ci3pmnCEgc+RQ+bYWnOU+XyXJiRFMtTPcFy
VjnpdY5GPBY6J1p/vaQ21nDQcSBckQR6j7mbF4dBnHuedGV5PGbZ3IeYh7NFvq1CAfWRwp7ZiOmm
3TvPvwOT0DlTgmWPpKf2sGuIgyAInoxhqgo8AGJj6peJtfFfZuoqRyoUyGKpPaNuq2H125Oy7lcc
27RwlcqXucOlLwsvnAK+pLaiPxYV1nXrzefnVy6irjfZUK+V5dBwTx75enbgDrnF7TRt/cGaCEv2
bMlKxTcNwa1DLrW/2psJgF2H3yZkil0IAoW0ODVVPMSSB4mP9db0O8wVE+MJtMEsQ7QShGZOTUro
raNME616PAooxs7QDZ1WQz35zDsfhamFB8PdsZOY0/fWbsA18PLywHk6uUsoyEzWt8kViw+fD4nO
+T5rwzknIh7mdR9XDaA1ZtaHa9exuFYRP1vlMbb8ZohWaq7pMA64ezex4rurkdQl3PLIw8P8eJnI
TOMSlmYo940T6MaSZj0eQgO12Gx+mS1plEfb7HfXlEG+impoDs6WmWeEiYlaQ1lqWidg6Vjd6qmq
8xdmXm4QzO4AIWOt7avS3Ut0lGhvncYVpoS8BOgFKJh1batbxXtNN3L1vKNpHScv1yGvbSTUARM0
SYgRnysMf+a0vhrkSmKsriB+vcnjDIFvPOtBY9EEvhlZZH/rXAgzlPd9nMqld6StnZ8Cfpu7OtNK
qRXSTkpNv9UH/cWd5PBQ+mXWJQV3w0WWaODhVviKHQdinATouUUDMMH8sv4uHCRkJwqSOmA3JAZz
244vYBUj9JULKVTC0EwAYtV8Fdxcj9AUUTEZDgsCd8YaEjJf638Vw9I34+zj3egeJA8GzRCzXDOV
UU5S2msG9pnShxnURihjukXkhokZqFnt93jiVmYNmXlxweDoGYh2ej51Hz8nguOQn3tFfP8UjBC4
Zx4+KLiDjUHkN1tIgZNbBDuX6QPWJKS8JYT0UYmZTkD9BQ0MUaT2N/hSse93GJ+YaiNhnhDPI9Ou
7MPbAMLCc3hVfniey+rjSpWb9Svt5SJnuptCUamjiU4FKvmkAFlwq8bVUXrOjcebJgc9NgvSDUQA
0sBsZhWdiJxs6IcdmZqZhsxIRtKQS4mIe/mW5cYqbGv2RyRhjHKatPRqfQqFTuWchmI+/D4DN3jq
7SU6ECkMKLdo+cli3Q8xHPne2fnEKpTVVGpcJaZi3Ox+JkHAwAHjOUhrm5/Ae44EElS5yv6O5Z4Y
COigKdLrNZNCymQWj5KXHWT7C+H65fGiNzPODV5jjgUNOdPQ4cBaiF2d2tJe/2c5oRYcAI8KLbgG
lMteKGvgB6SVrsHAXqyOoW2r9iRELeY+iH07ByQm4GIP4PneqseeVSQkl3Khc0UN5b5cjGj+gpQL
zSUzD+MpPhm/nkklhZCqUnblMiHjSz0P0Rg7kOWOCMZwcZqsG5NuM15tsGLNBJza3pJxHPb7IFgG
SAL1Lg7N24kz7s2/cMiLaPlfthVHRTwniQ86xWD6GeKD0TdwAbQAX8GGk5vOf68rUeZcpnTqB/jS
o1qBKAd39s3DdfI4dal5SLVv2Cyx5rzfoY9XCrdpTGDf1Ulbvdkg+Hx8q+Ns+MW5PbEudoXZU5Mu
ZDUsNZJ+awx8qjE6gE8XCE+TLbaa7GK3LXJJX4E6IyXpLcbwXwlvn5oLoruvRJf7ZTchB9jhOKTM
U3zxv6i6AmlKnmvZJKh2GIYmAHqtodODEXSHG0cAsAs0mw/HeZ6naDf8O3cTcC+tjMgtzOllkPWM
GOAaGS+m2ozT8L7HJb5SBOGj+fCYExhjmHSAsyRsX+plkx2p0w0xXmhzC0qvUnkMYaQiBfXAr8sE
otWSOjnzPI0R58Ayb7ELNh3TBBbNX0LH9tOfaidBgjbB2ZRNwnzrrRl3E2Q+icoAnwtiFVVufMw5
SStdnfiIrpkel/satwqccTf5UYgMNoH/sB0Umviq0W5ZgUbujUB92yIkrtipGtICinWqSsGQ8a8u
1XqQKmOkTx0sjMQ/oPddXl/jlkiENoQ6VFP+htjJksEqhk+TY262XspyOKCOwvxMObq8eJNRpFeu
dby9qwHLl7VsjSv7oMyEr7cIIsrWxmIsytiZ4nS3EnwS5waxOCkDXIjeuYcUe67TG2XRn9SMyM00
vy+2Yo5+6ESGZu9yVWIAznykMYOAkaBbMCEoP1LJ6IZw3eDYR8wsmbSo16M+Bvk+iWBX0jCR4tbs
lIUYBIg2BQN+i2Uisixt3CNdbe6+yeaEK9DAXtxDYHJvfWJ02uDfxjC1sK60DTCVTmc4tA2NpZz5
VpfJ0IqI62SEtJo9TSf2woZhwe5UyiWbCfA5FZvR7/nM5w26uFty+RMx7U7ddTEiNI/Ec6Z9GOkc
LCAdhhswA5a0/pFecj3XPq2nnMc5mV71qjcciYqHZSee4kbjt81LUwjUa3M69t6kG9G8WttpNyJF
gsLC93WU5ZCaMtdqNilWnFeKWAQb7q0O9o5NZY3vzxgI5TWtLGqHhkoPrXgpTxlRs7KboQ1aB+Ny
A/+YoaI42e3utmtg/GILZZMALDIXoALPqdf8beQJVdPvTwp9TwtGOqO2T0l2V6aLYP1pB7BMepEm
sasCCRFAAAdwzC/UAO8qE6vI56vUARbdqHmxerVrrDr5t0dPAxw8K4KeTX+OSl8yrSxbDvgolRc3
u4dSLRsZbELnYAsmzbLefiquWS9+O/AR2I+bdF+taBWQmr9CJJFMlBJTa6R1n9vFxa1ud2zQnWo0
Zg4XBSv5VW4KUFDgOOsDB6zgSMWYSSh9kG4U1nb48JCJuMgMjAmmPTD+WtEPfSS4hiMJf+LcHigR
G38sq8jdQjIoJdVzCe7kKMJ5LKd999+vxRf5XcOBKkmmBq7ZN3QQv2aEG7ayxUXHGATlOdbbus3C
b+OaHkZPF0HDkInpCugCzGd0HoRuK/Fk523fj1LNpxFwZeKsMc/SDv+ca5jMUbHoKM0VAuugu8mw
utoBJ5KvwtV1lNlve3cI2XZPsNEgv4I/gV/flGtzNxqIO+Ama08RjMzeEb+tdzfkfF+83+8Ncflu
2UgvoXLIBc5idTLruwVK87cXoZTyZ1k0JhCvGHE0R1cTcgZi5n9KXb9EKiEbPJQyyrVFZEPub90A
jcFfo1aeMJA0/Vw+DX1ffn2sLLJcZm+RSSGobh5PI6XgO28NFb25EStL+q2uqReB8k2J+NybJhw2
B5CDdU2BnpObkUOJ3vERPtcw0lQbAgBB6RkJjJu5D4iFX3WT7DwFwKumXO5xJ9n44vFjnFxLDMVS
Iu5T2Ws2RgyxdqJulNxq9U7DrgJ1T73K+8aLKAag0nCOXFdc5iAbbLqNHKwCx4IbvvzR1DLZCl45
ve99N42mgz6YuEpbAefCUXbJuMUBCgQ3PMHa8tKOFLwYMCTuLcp9kQndFOeuhJ3229bURt35BaJP
N3Jv9VZawcp3e4hMZp6bLzXrvoP81tPQ7GxoHZ2j9BWmYPPjgc5k0QH5j0tzmn91F9HMhPUXmRF1
KpIEqwDhakG+5boeSg8Zfz+mRixmwzP4lxuUvsKP5kXfBfngtK1m1NqlAX+bzt73mYVGAhkgtFAo
iy59BKAlXm5G/gjXPVrAIXPdHnp9aCro0Js+LoWOrqUxyTONp8LeysMusZpmt2J/1RbO2eM39bVz
kC0xECOgjDEKszMNfCkYqCOnLLlo6PB5y10SnyrB/I/PJ1BHLMaKCQMgRdCLGCx80ZGIYTVvMgxF
FNqngOzl6KofV74T0vnjru41k6YuHiqgaZuAf1+AyAkWfipcJO5bYafoEGY7EK48Fr82X9wnH4DB
W+qoST3N/mZDEBeQIe7OlEuFMXMkUBMK+esaG4gNaKjLxglDTZAKCsmoeZEcNSuBy1/lOgexTKSy
cI7Zjrc98HLrJYrk5cS4+B9wBW9YaBc8oPV84I1ha+lyTunLnIWGMwt05su38cn0fjYqo/cj561h
s8PSquQsiF3WiiVPIh1ddlrBU89fHB6omu8bhwmvRZSBk6fYZhQrsRnHDmaQwVVBq1VIFYMJ3vUO
XCiSNwrgrPopz6bRbxt1ZNb79waZ4M8UQAl0heUaw9XZ5tF9SXGx0P1T4LU19/xT1WQX3ZcPwS0q
zcX8NwKoVFfgdluI1vSQJtjPUTiadsKcaXg5YuvA2sknZMyAswSh3a7uMOnjzFmCqvSx8nsuGSXq
H52Klw61bTh10o4+BYmnLzGSg0j1b6gib9frPuDEMYER3uazo7HFGWOy85gjUPy1nLZ6nKmmigjM
Q7N5fUdSwy7eZIUFU+RA4bbBQLLuYxfqhwZLyv7ZTojUeT/mKv1/S8UqRScsw6c+wdkYZ0ONP2sG
aRpFXiev1CDUjNpH32hIavLzq4tXh1Twf7o4aN5s8YTMCUqYQ9M3Vbg0jxAjOggZH4Kq3krGmGO0
dQFceyBivjpli+Pbc5Z8TB4cof+zcG/Ld6/vct3t3asb/3KLYivOAq/sqEsJWw/VBBWva1FnLv4X
ulYHhJG8AeB5CWAHxkPp5p7+dsLoiiOjQyhdD012or8LyYsb3PLZya/vCrCujlCxi4OZo78tgDmJ
L67FqgY9gPbyygGOz1qDIIz3D/nENQSCIgNwRrZZhtYrUuVAjzGq8RTUAJIQqr6ufAkfhnCTdtIU
ynt5xKMcMLIaFZ5NgSU5JjFZpeDBn+i3T3qP3yCELBqI3KkF4lmKFUveVDdIPZjqNHGCCGOzZ3fZ
vOfBp9FuhJC5s8SS+scpX0oORi7P+kqeCy4tAUofq8Byi+/C1ValbFmdty+/fKNiMo5WvoI5V+6D
LWJ7AvO8V3da5QtXYYoQLQquB9oSnKEoqFWYNLhsXsMQ6nRA/eRY9y0ATyfPUqsAABzEv7L0CWki
JdRY3CfVKyYBEPhaMoQ9YrwoPxh5p0H7NJML/I5E+uvgxurL7ruGSKxzOe1qmbG7BUhKuDZIqEya
q8roga9HvHIT/2zxQcIc3hbIcQx0SVm77kdQxN3jJa869PXBKNvbrDwdDVJM8IPnUwT4CGYxluKV
tcJBT+wlzF0pkkASQX/dZJmrZXPy1C06pMjSHxey2Z7ACyaiNUGsSQ7mqDuhIXiHIgIPFyIk8AnI
szc5u32RJ//eiJ9GNbOXMWnQOGY+Z1ui48N5BOPm2b7wMskGf9VS8He25tBkbzBS3SMduDADshVq
yeWE2cTIhkz+d6uEImVuEOSC+zyz0TZjj7Fw33v5os63fGtcMGJ1l9+cCBF0jeZZuu8pr68Fbsm2
SrKA7/VAOMTpOEDS2STG6du6HIgEfrCU+p+y8RLDdqpoo6Ccs+U/XLDhTAdNLtgdSXd2t95RpIhw
RohTBkh7OeNNq34qr3s40bGkkOILqSW68KbTcBzYioQeRg2nXx7myxXDKDu/984B/Aoafz7KmPpz
S8G6mvL/dqMdyUklcfrryIjhzJ4zYCIU9KnqzkxclQRK3pEVy5hPfwIGvXlTVV+IbaVFL68imFVP
Ho7fo3C3JYu5z1GhBgLrlaJ0+qvUnbLPVLZ4Gi8ppzbXNPAADQiHVIrSh7U0FxT+uuY0yL3KVfKc
Mdz3RVCYIKc0skV0zBIYr/q3xgX9iiObRriUsQ9Nh+b8tescGFYimCKDkyIWJGJ9Q6P9joX0YEAe
dv82yCswOK2v04cNS4O/SBpNBj7sREKQFmfbe9Ma02YgYV5KWLBRyApSk86v0xFMbk7To1CiwAP8
6hr7A4ZoE27CtvnNoDLX8qPtjVD7/K6msjY1tWJ2ItKeLZN+Y3DfOQ8tN/woVdTgwZa29F8VbxtS
TuXH4Wyl9kYM8uBEkoEwCbTl4i4upxcSvPq3cobnaN2sIaubRIi5tT4t+YruMI0+PknIujnq4Urt
oGPxLy1dY0xlZnoWNyYS0qibrDnfLTe1rW/MeF9wHVI+yV5GLNLRvEMqmTAgL9ajthB39GwDwdrU
NXkP8w7VJQ31kp9XTMGhMlplpvM82YfVHZ3BDkz7zm9tHZUqS7VuJDBfWeg9/dZHTxh4OkJnIDAO
6ivC5dfY76BugyckRAEL0W5EYnHOW/aM9vyho/9gyPTV1lpwqhlyDJ8/Bp8k9E9W9A1wV/SeONh2
1cA1IAKqvKlNSMDuMW9/0TXe70glajuqbtc91CrB9z0w/osgZAfH0wcS56dt0jOgr6k9BFl2CO9I
1wKLhr3GSuFPRqG3YwK1Lu/fqi5FwnzDf7tn7TMhZgYsN8JZMZD9rjz6PhO1adwo0FbSBcJiWYB0
ULNATIXf8WxfIZ/JaM9451w4EMX2321aXZLcVJLkYPL1GTtoPvkP7QTk2bxz3BHUG1tbSkz5eVvy
NT9Vw3jkMsGCsxbG5gKWbxgifAXqKbKzcsNzuVQvYcyiPQjdZtfEYTetX1myKKoqzG6NC14WxqJG
A95f8wv+M+dFYQXulq/JnCmiHnzSg8l5xzQ9350piAtZbsB7+/Iak7dqJxPjNPQZyOVdV8x64Mue
AlHpVwwI99HqLzjIW32TGOaLuJrvi5X9A+0iHN0800nm5H7rUhgzhZ33iXvLCIz+HYFG3vmp2MCh
JlLg6ZrmLfOlk0AKShDsgclz+kQvWfnjcA+B/apnH7YZ1eymEdYydlfr/mxSfkBt4TeQScv6yy0N
KkzVJcXNMCc5rvom4V5hPd5641NxTe/if6ofV8IwcMoO0dhXtP9vNQ37r8M2hdAuJ/LkrDsE84Qs
pCVtX98Ru/yLYax8tKwKkHZDaChAcdwcKvJlVWP7401kpvgd54veOxrLmf3SQCRfmyFy0h0LACCf
dAUTzZi2a+I1IzQDXxMy4tAEmrcHkPZmIoBvG7lpXe/5epkIfp++m9tc8Z769qehgusmvhmnnbIQ
DgZe33fcIUJr/BOdIsxls85oEuVfo2GMEnnUrLGOV/v5WAhV72LkRP8lflSs73ndcERQu53u2r+2
36LxzNvNU1Kr+xuwZN7vfwUZlEBN1NZLSQjUHwNd9/+Z7U0xuWK5y9CUv+i+L5cQJtDSMKPPrFWt
ru3lj0E+i0N2ZpnMXhFlK5llHzdLuVytB+OMmtiA8wwaIECEHYPmvfR/GRJd6dnC0T7BUfXTga0c
kq5Iq7KP70fgDmWPJ71quGTB3MId7WhoUKRm6u09Pj5KyXFYXoyTNwbNeUgIUuy1nJFtJyoYCrCP
6H2uJpKwsDEi7HT4rw3+vWptKRXzOVBRkLQkcf8WYujKpsRCnD7IAFpQMg99kW3vXC6FXZVnH6qS
ncUwmR6nIUYfk8a0RzN/lTTNjyg0P69CbW//67SvwTkHzNVTg0DNBHMNCT6uvau/GaaQaqxjCK+B
ql/0zRC9KhYEJiky9ymd9L6/1TBzithj8AB/1kErC19Dglw4TwNJR24rpYb9KO3Tp6UQDvGDlT1H
adXFDL9Xu7I7453h8Y8LKWzi6iYQ7D2VRFnSH1Crb8CJ/gT9qCQV0k15MtLS5JRruuWjwNfvzqYi
Chtnyv+LnDqB0pYj3hhYjueiJvUCJQWNfpBSZvAf+/1L+ENjAtRGo1pYs1Ma3g4ho7sstVjDmIMB
H/uetmakvdJLH9a9qL7lGLInELQKScgD5aa6ZU7blgz1jbC22acVp6raoDxTqbnsEnlHzXzM0rIz
3iQIkNDL1kbcvcSQSbzb1cP+6OXZwOd8a6J9BT/etxPIxuZYGi17if5zWEWa7/nyoWhxa8sdjLx/
9R+cogo0O9MMACm++0vMzygMIjxlCiliiMMrTngySFWb5QLh3+ZZyhvmx984cQcOc0kkRZrOP5pv
ZWYNNhuDpw6SBP/dl3ypYdBMO3Stledkl2JlIk7TJDiyUcJ4eqvo5g9A54v7ZpYYRMBrrzbCYm5e
tZE3kzyD9uUJ/aIUTiCX9KPlI6IFKbY9NGaJAgM7NyJPgnUMROvrj39QICR/LyTPK5hQileLOeE9
HaWiRonVXietCJd+qGDG2KYVbA5rU2oOPTFaAEpgRWlMZIUk+Y/kDmZjJa88bS3ZxEVOiRvitpqR
/uq1m82COgfDC0cHXu6vEwp+VWaPmo+Cr8m6kU3C9Bq54jWEEyyg/fWkxPGakopr5X17ngO92mgi
axCBaktwoNj1vk5/MqUcr3Y2o3lgyRnKCY9OHcJBXRXzp4CoML7mjmnPW5+3nbwSKeuV013t/4S+
+75AIIc8quNxXz3swYdMh7llLIu+c3CP+k9S8JK6iivlzhJK74lvowdJqZqcmB6tEVzp/nDsHz8y
5xCbVdIRcgQBMgOW4hrIQkD0/tYwyRSvGbzGsPp3FuW7dwbxAskmF2uPtQfPynbM4+81RuQL3t4c
ZgW+tl21YCWVLKqruA2xae5B5JQxAVbiVOYaaACZusERKW8RQRwo0ebZL8McQzZBsD6RSil3Voj4
sjb4iJtiEDJzOEu1M5h+b/F0Lu1lH6MsXn6mRlH052iw8cvL7FFtpL7Q3kygfOoauKV5174JJGHT
xKSYpXPy+bGvFKX1BdPzs/zayKKalm+9QciBTxPCiVaeVXVjbBfJOXKH2KAYfn/DmKqUfsPN3GgP
CXR3z1Rh3Bp+uqYGdLZzH1maQ6hA05r70Mx/AIlDVVhmLFVBb99cUJzXLHiQY4e78QW6sPeVP6yI
1GsjXdYUWEMoXpJdokXxumVQbRV7yNJiHAlA5a4M1UV1cc3gUb1LnX0PnussbX3KLg5LqK4Z0yJZ
s42Wzd0made27bpIgHSigk2oExwOFNZe3m5203UJP9Bex9QVcvdNumVA+Nl4VQhvjHvVeeftEj0Z
N6U1zPV5GTRvJ8ltDumHZh9utXWRAhN3XonzKxyN8r0b2Y5h+CgvCB3eLEMnAPX2ldvYFWk4fykj
gVOpXxrqLTqoeEqGqdGVThPmAnhrtuxaDe8UGXLlQIXN5O/PWVMiPTJEzzkPBPfB07hmKFLA38Dr
wG9nJgDq6ePS0XSskm2w2A2LcD2qqQLsTIJ3cTEuTW6fisV/5b8kDHi9wopjACXGDc4RSBg9vJdr
jJzaw0pQeiYJ5lWRcgIX7TpG3Bdu/4V0SmjohabyehXCTnYHH9dc7765KY9Au06zmasu+vqz1+l+
Dlq/XU4U/nP0+vzkguwCA/26Z4BKkDnydcdIynnkmGdS/EM3smI96AyIJpQtADQrEN7+fjYle6lo
BzBe8tUBRgR2j67UkxmyKVXh/6v0l8tERFX+0PZbhkHtGBUh3Us7YmJjWkqvmVBWgjjCqsRV+XVt
T8v9Irss7pJDd5oLWG9awVK+p2wiSjyaKuykgdleEoHxSTfrvCP+JJ6X19s0ZfSjbITlSPfutr9T
thY6swlvJTj/e/DC9PXdzr7BOuCy2pk1YSKINYhZpLjwvyA/5M66Piu/skGZTeFa72VSvEPBKeJ3
EU/WiapYzmQ1OAqoZ+EOCeUYmD8Y7z6QTpQYTtF4rMyD49NEtqmsPCI1mec7rdAvXOAEOZJHyqA9
nroy55EGjo5eizgW+tKNQkUuNJYafjzI/iq2sMmj72YjFJJShTi5cI7wdipNK/+pFWPHbMzvLW1r
sULA3bjOKKjPE+DJi9l1ISG2ejUIxEwraEmu2+Xw4jczzf0Ix5cMyayyeEao5G9+OD3K/i9YK+OB
7fB34/Sq9ZDHervct9qNPMPDBg13c9UZmFrKUJ0wsoNiorKt6BUj8Pa+19yfbyhPDZRsriEruVCu
Q5v9zPkRfgfRUMspViZxVzdaBmZKNUtOvy+guVHt59jFLGoNu8r3Bv5bBB4U2pHPqAIvsbJToZcb
FZ0eBy/MirJKxi1j3e+BdYpYN3KDqxq79i5HmMDHBdcoP7yXQEep+OXq8/WQGLQ2KUe5/gHBl7Cu
uqMG1J0Mh5ck8Dsz5J/L48i1FrlyBL2+nLeMIzsmDCm94dpDVwBiZIq2EnoqD9/gEtTyWXDUFomM
Pux50SFGy0gZiADt0c1jzkbRmWa+Qo0tsc2adaEbsyZ7Imo7NVj3Ucu9ex1PxoDvRh5ejJNDRyJZ
d4U+8Szn3CKULDJ7FMmWNBcRNunWTOrRFQ6mkLWOz0U8+kgIWRUsatJV4AjxV1vs3CLSObuCOL7P
gUocYJlHqFi+LfbdO0/iPlgAytmjEd0w/Rdk4ttPwa32204Z0CP0WdGjh574NfzFkK4osQtCwRIP
E8B7s8XL6E2jp0mfP2Qn9vZQcSLwoSkoRWLIlvkUJQyZI9YdLOVSXYV4L/6SfSPZoHt/w4wQzL7E
nbOUsBNsJj+zX4IiqfFu9QahMZahEaZ6OHo5vLrBYyWUIN2aNYRtVjaDncpr1jk88aWxl620kJof
owq25MdWE6L6bYxB2dH5OgVvZyZJ7EPweUabpytmB5yXV7/Y8UOoRJONjK2hTMpPRPkZ9BI3SA4l
9mGgW4gfmya0lbX1oPjiDKolPXr/3ZKJ+VDPhosCwRRooPTh+O2zOqDBzQgdylIqDwZV+2qIXwPx
RKjabN6L3PN8njcSus+Wty1fvbTXmkHNKw2BLJRgziPRo/quTuMuBAn0738sd8Y3QFAPJ4/xGzkm
FjOYxFT3pgJ3ddWL7ArQDrVSDPhNXAR3AOoVdOVbveabKBahfZ3q13W/LWLEAIp1vG3raQgUUch8
/Q6ziP2FDU6/bRfh6xdwu/MqgRbhI1/uQBU7hhJuKljsZX75LjmE2J6CX0UKnWr5F5XqKd4oGPdO
IvXj1NgMzEJ64kmhK0AYnKQSxVfMXmw7HFPM5ZdFcYehoH5TeiuWCfUof2CdCXg5G+yGOPmwfeeo
XgW/GP/qSrQVYgC9VIdJ/9BGFQNvv2tmHer+jE7n+4oJLeQyaDHNcoFJEBpvS+pMZ9xE5NQjtQEy
k9f9i9v3FWFgYdQ7a5FS6ubixBMna0LtgM28oo8juv+Jj73xdbw3ug6loOKZSf2AG6YD7CoMvw7h
EhLqREw/tZZQa/JDtyYmi6oDlRLvXztB0mDpbjZ2eP4bPpKQTupGTbBrFxDjf6ZM8BKwi2wSz8GM
nF///QHSLcg/vNScN6eT3pEUbcgRe5GzufkYzMmhMjfvF9QGRvD1ZCLrfUhEEBLjvYEO6hfTih72
vMDm2zXeoSyPAd8jh7rPnKT+0+5KPKX1Y+5uFcfZou8dSD3rXesP4yyqIeRd2sQRUo55dlxZM7eq
aKHM18Yxfd5I4vrrJIHzo9xMi9JoBbYSlxF7+7WNi6x4qNGlAu2oWyz7G4WMiJza+4nl2Dm8o4Ih
NYQMH9E46r81eCR1A59BhDedasqpJkwGi4Sd0S4m5FBwkTrnhvzwJkoKk+qu3HQU7FUsQTJSoESH
5HduuX//2urHpm28CeyZkUOolwxRKF4b1gICjJtG1CxkiMvyMss1SazKukyXVvtJ6ld2EMFAELRX
n2t6F5at3uN3pKiLGxpK3m/r+sUhyemEfjCDTyzegO6xEqr78oitfp6hpL4YImj2cVEXWHCTYJTw
5ZOa0zL30JZsE1b/gyJ0DSRfrq3KiUqWGM7ufvUhNxe6z8EZR9g9B1O6zO/Q1b2agKMrilFQ2BNX
YOzTZ14gEjUmmHDVqcE24JDEHPfjnugGP63UzgTqT/r37hvsN2Zv7vGuCu9eWduwLFkYMeiE0Z1N
3I98Fxy+OSc4fEP7czUR59Os0Odj+HoB6TXTUG+iZLwYbQHeAFi+4ODGAwW7uvEtjBzPow8MYMDJ
jFVxWX4/3l+2LE0GpOfjRHJhZDx08jB5lkhhjoy3x/wGgZupopL1vrfnebW1WR66k52POG6ER/aj
OV6nVVGp26GY9vh4rucvPEBvmXcbQRv0s8PN9lbdhTuzNansgtSpXnES7pmxHNJgiY1YbZox4JD0
itZePrf/Yt6enuj4HakOzX4Ljc+2+EIoRsV0bB2aCuvB6q26qmg5PYmwHUAzJLhJcLEI8434TjiS
vSBZVZs2oeDRBO+Jfy7YGf5cTErYjZCRWnf2znVMXodPsLdP2PvQOOIGCPVRDQ2Tkq/uHfgmrfA9
b7PkxL1WIp50hUg6BXS3OXkOsFFIcXxa7AyWq552fCQeE7tj/1zvGx+THBAE15PtDX7PG1WkbOhv
780cgJOctXlouw7JtZkpsWnOgDaCWEIjtBtUULss95pC274SCy3B5O0arWcBbu4XRonMI/T69emq
DpYu5W+iKetYIZweZ0LIzcyQ8b+OrdavJOV9JlxSQTVf6cH79jfyXTfIFseHTGyzaOv6361fzrQH
UXxaUQ7orsgAxUE5vGc0y3OQAwDBkVTJ1MKLyGXhLXP0E7lWJyaJLWH/R/HTwPxIMmwfQW/X08wI
kIns55340P4P0a/tZEX041fqqYs2oc3R19jKYLAvqaWSNHypMuHo8MzL/l60+eSgokoGOvRR6Tcd
Wgaqfit8V9mzAa5fI75jSm/0b247Qs8+21n6gsL7QaqyO5q7DC7obdd1P7XlfNtepjaa/wSXt/gs
ukaXvw2x6GNUjNXc+PaKkSIPaPwbRTAswwn7JqfupANHdcuuR+pWSKhFIyCyBo3/0fHL4zpc4qKI
jFlBk/fHgIcL2jgkBCaHh44aWWv4mVn32PGYbOypLfFdiv5tnFkvSkiHJ8U9uPAQCTn5VF0dRDzU
9MNA2MGu+q5ofr/N5L7+Q3oONkYLbk2vk+6RYx0UGdp6cHbun3e0rjlrU/51qADwzMc30sd5Os9l
UpXvT9Ij70ERyRzkJ29kuSV3AxFrg21ZjhQgTna9Aw+2gUptTNpz6MZnQTTIG7V6DHWq7EPbMJx+
JQNZeirf66jRvKXtuMCx6usjBtq/uTvJ/l2AQ9w7IcW+JuFZgYefQuYlNMneqWjKqUnWbmj0jS9f
kL2PD9bYuICuVRAQZffKWwwHeWYS1Z5H15zkd9s1anVUdMggkBm1BUtoZjd+1ZWSRYQrBHEYlt5y
z6xi215eavrU1B0JC29OlD7rIU0eaN234uEAJmZe56PbxpQqai3/gvstV32J69msHLvZ0vbMsrcI
saL95DfCAaQVKUdPuql65O9QbCZ4KVgA4v+NO49lfVaZub7AOFWr46Fy/7oamox5mpKp0fvPN9AV
z12GdU0gvNpMwG0Gghc8hucFPXqlWVSh/mmVVwR2O32OKZDzgC+Eo8IOXadz/yE/W04c9UOKDnJw
uZNb3G8QWjTA1m16c4amM1kX7x6ZdTZasWk2IJdb8p02FoHHsMiwneGUSXtuH8YR6P0BCHE+yc93
abikAESOLrkFv4Mhko+hQF/+W4DsmBiDuKZOfoKro0WoIgALzeWE2KqgY9I3MM+EjimPPfpfV/jM
2vJrXTMqgDQOTBl3niIBKW4YPOyLDHCJJaBsKbBtYrhlAQz0DZ/b+oQRUj+fBthsxEj2FakEHGXo
kgMiqk+DtgqdcZhzw8U4vEs8PdNvQEG+xbj8MqtklysR5NB8B24WtPIRE3yxnqnrpDri4Zhb/Jxp
kdVFomXHH0WLWmF2L9oGO6cNa11mtSUZoYgC4jww7i1wC707nPoUrUPNcJEKAr6ielQsuTL383Oj
hZwvFBVlebVQm8rUzBuGHHLJr59kzi90EQEANRsz/UB5c+ydrpO3K+2bzgJYYR6IJnXN1ZR+3yMp
+So856LcoXh4HYEYgwGgH6QGBYcYL8LwYx58WfFRHn3kmG5Od80tMUOwygp7qEGBN8qLxHK8KF6Y
f2XtI9C79uBVU1z2KnnE6M7XMgAGwb+l9u0BijA769MWHx1x60IoDJzFqfb9r6Dq9KYHjfpJMQdn
FznGtrN3d6kTrFZR6+MoQSjREfYvj97FYBpEZ3ppW8FhxkVd2im8e7HvvvpMjjYb5bl+B0bNuh3T
xFOcImQJLFjGUHls5Oa80dV418QHAVpvNssCf+ynz3rKpzFa0Qr8hxFILrhbC2L8YME5qJvr7R3X
euE7Gul2YOp4K2lR7KwbTekjrYw5UjD/XGzH0/fY/f6nrx3ldW/XENZrGiRuYe3a9167LlODPE5k
WgCMvPOSEneX4v2y0e6CZ+Mlrns0DP8QID0f9yLI8JkShZfzE0ft79qgqpS2E5V/GUEIZx8VA1U2
X5DpFCkSs7cz2Gr44ZlabXdu1QMr1Xf5ClGgYW+cfaHxVeyh0UOkpoxCuEqZ9eup4j3ydpu/4gwl
offamxd+9JFeoUumyS4XVqX3z/vcZcpyzlXyLTn3wzdw8KnKBhhF98JjEJPLcEjg5DH3q8Or/86f
/fr+Yvw/hkQZEufPRaF6je+1YqIqE0D2WZqT8sejgNlnen1w8yIOkXybxKqMmzT952YFSfT481Vz
cPaWqksXHOpThIJtuu21J9Hlrl51ZWxIAk56Ck3C68O1gf5UWTlnyrNxbLL48uDGHJ+ufRAKzdoZ
+Mi8fste5QVHWNTBS+n/gALjAyFAEYSQHO02ciInFBe5bkxKTs2Bm1wk6GYU3H34umebGwTBysde
hMWPAtoByiiKMmCQJlbqqFpTZEy8IfEUmEFWfJswlHqGI9n4MjwL1Wo9fo+JvkqekFajV4z6/drM
s8n4Mp5OtjMqjwsLIzXkBg9q9aFGiaEUys5LQ3Kk4SjyCIJ282eRd67uxN7vOOg2PEFQyWDaxL4r
T/nNwz93AH0xILg6C4fVxJtx0k6SogmyqXEyhmGFe7b2azE9fj/KdXphDaphsMZU8TkIDc51+Hs5
aKEhXtWYInDTlW3cuEM6feO8XxcADbRC7YhqyudAsUzXFyBHYO4UIcv4sG2oZh+RdnOQsoyA0l5L
0r9HSI+wc6zBPMwCxWr6I7o61DdYmJwUI2ejNi97meKo8r5jXI9bjCHWStyyqlRELtO3Q0iXoqvV
KW1Nq3AHckVnOKl7UAOk6Q+ipAwLbv3LKPvSsBsEm2xFKIjfPNssq2DhY2o/6t719wqclBHbvuTD
Nf2ADr7KYzmnfKbqU/ZP4WOUcpcsfrm4SSkzlv0Ic/PF2XVJXjRdnCVEpvGm2tR+b6PjcG+vX6b/
7je2hVtllFhK9GAPm8d1eXDBKBh30Nid+VK8Od9tzQAm4IXGv3BTQdVxo/+iHsLjrTuNnFZIiY/R
W3SbOi/p3ZZyptUpEcbta0esxXXyUEycgl1Ykolkng0IharC9txJMjBoeWONOiVZWgeuFfi9HBs/
5aF0/ywFi9RLrHcqikpHgv22TqhA+DzuSKVu/G5o1p+UpcF/gRcIUmLq63lQaHkl2mb2PpTTUxPj
zfSCTdXWPW0oWL90S3SEpZ426ykqZEE8/228JgiHxO4u57faT6MbePn46KBmMYMLGE9TmQJ9c5As
PBQF1eZyG1uBKokL1py9GwwsnNm3FaOziz1Hb4psQ6BgFE+ZylcKpw7HvbtUzmsjOewVQN4U7VpU
ojBn6uV11EjqdCfBJd28/quFjgXpUYNh/PtXHC92iQm3tEjjFtk9v3345c4NVqgsLxjZpn/3FyxB
6iKIR1wGuii/gDGivhE0PJAII6t26/UBZ9zDtw966bPWeWHvycsi6h3bORSAd+HTPU9z7vdRB3Vv
mDwjhxuoDdNLfoTw2odgYgvTd5SdbcXgESlGsCwuyfcNNYkRyth2IZ/mZKgVKU4GIeD9+PRcUgD3
7NKJpQyCUAijEhZoduRjaU0Y6TXrT8FuO+GXJlS0jgTplG+Q6i0EmUWRRANPNveNe6lEDqyzb1f0
TBVJ7Vp3/1I4CRounixI1UILrRCXuCktAtOtR7r/YszkqAWICwg0uTV1dK+00BtB2o1DrUY+/ANS
Hsl4l8ningaqCS7UdDc+4+AqVs3K2NOtJvpqCiSq17QVrE7zTCNYqqllH556agVng6SUzseCYSJN
BMQEi0HpXLTNA4CHnPNXyvmYet7zmJLnQ2+yH0MlU9tdsTEizag4GR8n8FmH8aHzkd/crv8WkrFu
RkI5e7HMZjZWk/lzA+rkH9ABRNMC/tiRWKMBwf1Jnk+LFMzQ7fIlR2pLOpwvDHWYJBjbnMj0nOWI
LWc7AZFDRk/OXMvx622mqzPSzxZr2dPB9Rje9yhwdpQXZsKLklpeq5m5uSxYKtMuTLWQeMQOsj9q
tQWEIcl0mdATh5SqJmpXLc9Q0/pQPBEMCTO3NDtByKgXa0pXWttg4vhTuWpKn5Er4lpQ9igOoPZJ
rJDJxI7WwKbS6wVQ46FksUrRmLpDXcKHtsFhp8EaF2ojvsX6E7KL5Q4SrPoc5GpMfO12PSRqOFZ3
YvzVabprUJsWTmXzGP+c47tO7AxzlY3IRiF+ULkPc2nQzPjNW/Bj1tjeexK6SMbiMh6TV72gI/lF
ZgPQQoqv0Ds2r8cdwe0Q53ahDkNXb3Q05JLjj5KjoFYDWyOSF3KMceIRJ5hXTNvv1KKUi08vR1/Q
e7dQi6fM9VnOxNUcTrGlpGmCJ1fr5T18teHdZU8Kne5H4te6aCObb9xoWNn7TfSOqHdyybGpxaQl
L3dnZV3PcAPU44n20hrvDN2YWjf9IN2O26hupHJEJDWgyfoIMG09wPiRm+vAAE6jmyXXQp81w60M
08yqEFg8TCYV9/d3qo5Z61XfYr7wK5Dgtg4awRgjIe4vM9WIBBKzLY3Yhz7Zxw5Lq0sGrCDXAJUt
wEGfqbaKmQIXaSWbMWYv+5XXcmdl+xWciwzOQUhv0iSnstLnatnS01U0ZbwjqBiEKQd8fEgP4TzV
pjKnp1Co5yEtDWVgXyEhj37l9WlYU8g0b0YRb+Nc4LtKjNL0niz0I4h+9Gf65bbDs5Hu28Itqeku
qfn7aySkguEUaRnjK0Qjfq/dANXzD3zC6pukheTPvQn+7gDEORxriI2FVSaHJK42jnvlTdFPSOAM
MJj0LkSWr8PBQt1r3Mr1G5P2aOh0/p/4CteiSJCKiGbe4fyo3Xy95qrMBCZCpKyja68yEu3Cv498
3yZwNNdzNBamy9qjpi3VFzbAooA/aIkGe/9H0bwEcQeBddAbfPNazWTb8PChRqEWgvevzXZ0l97Y
TmVyRQopX9GuIFsshHxCu8t0XeEWpfdDd0VHSYBjRY5Kvi1ZIPX6fbIr9zUFsSSn7vtmXmgIHOa9
UXmL0UuYgwGkt6/AZVRXEU78nn+mK9N3x8aZZs8ivQ3YYuY9JhTaab8exyu5d/XAbYUnmkk0XxBz
OFB2SPAcAtQd/xqU5MJHihXUDpKxy/xl4TVdMOlHxJbTKQOymsyGDhA/hJ4l2DV4OljYyZ4th97P
h978tgYYo5LhlELNZpWCO0TYobSa0/Lmt0JH6atmyQS3/AqLbtPrIY1liawHxRbk8SPGW91ZuIv6
DuU/jDZm5LREAfb0rW3vatxpI1XO+qYh5kFHiX7YNcpr2bYMUyUWnUwCFxBd0l3GcabJB2F1Asb8
U2au3hdOjPk3qfw8h+YZbPbKNVN+rRCvHTu4EKGvxS4Umqs0BmcrLUawx9WBTfMEFybSFnuK+o+A
zPa4Rdf+/jI1T6CfIYAyhdDIeeOtfUgPzz4kvDxx7yeRD9Nup03W7d3VRaxZbUqNQiiIBsowkhnK
nAdCXzFHZ9qt3JPPPNGRG7cmVg5EI4bXZtUgdlW3efyMFijVdHSYCoU6Ogj9WHluOQVRZ+hTzI1r
AIpbBIjD/P6NhIcGtMulA2OeQrTpWYwOVA8uczEBp1l0fh0zuQki26gAkJQFyFA8GWyGLW5k8qga
b90ADZyHvJ4P/0vN7tzu1Ty29XgpN9eh4AHRbfFBcYvrahdx3MM4atwgWbcBnvDmIvZ+b0zVKIrE
pS1O0kXU3hqZM8wQtIi6ddJBYMZjQa1lyP0WfcCrsJ+1DCz/PhS7URxm08UhtJTF/Ji6xVpYkKVE
FCyPlprdNPbbAPkLclgQAIhbVV1CGCXcqh7DhnEYRcbKY1wpOKyhuKuN+gOtcMaaq6EOGBDXm5pB
4hJVT/Al4vmI5tyc1ZFrFeww6m8lh5H9Z8k0gNlH3qWr7fBhgyJsIYI1tqxAG6E6X43PfcGSI5Ns
+RuQoWaCDnNREqh9sWuUOQRToHwZchYeUwmUeHB6qOH7mAl6oajF9x6UhsWToXGWwlcV8HqH+032
LpuCukeDT8osWN4ESjqKGprDh8CJHeZvHoEWAyKLx3g/fkWrSlBq+qh7o9LXWLXzcR/OJ5HrSley
H0ffdALuCmlg/eu2WYJVKsNjCvTUNILbl1omE0qwJVVtTHazzqq8BerVYW+0B+3LUSnS0fnAoVEZ
FnW4b5Gv7MtU++xARltjTaukX+CCzB7tHrG+BkeS1LPri9B6USkarG674DJCy/3vPZrmBBPcG/Ti
aKVXILRZlFbr2PHh4Chb8/l7Z1MOYSjCEL7LQ6e24yixLfdLL172RJJTSel00hkjQLW5lGRfu/Zd
aO0hPHq4nGjWbwkuKUInprrxOsyTxwAhb7R1koZjbCKIY+9i+T4qRp9k5ccd//7C+phhFzJSWZi3
P5zQ09OjtGFhoda7mB2bbAfFFHsiryQmWoR0u1MlDztMNi00P8Nbkt8yo125K+uTLURHNyrMqoQe
Shc1xBK+oLVVqP2q3wlkxFa3Ol25DC0M6qrbZ0ccClPhOv9g6Z4XbCOu3PfJUDulJZKExUbFnZnj
ec4exdUNyeZOcEiKmn49R4p5UP4JEt2rZdLvuXwRKlfxBf/WOTfkwxx0FPJlIASwKDXWSqjaTYRB
HnJ9mDuAYyHnNjef3pXRqxbzECzem5gyuzbKzxtToHoZhF2EEzdxTI/IivZLbQW1cqFeA2aDM3uT
twA9i5/I97zZHaoUPagEqSq/YUZr9m6vhOa7JLJKmPh8fVhCaoDUtLQFMYweasjEuTsGrnsTskmU
XaAAHDLF0Oa6ixxm2RQ/cOZm5o+7+4W+evONFqWNJibREsYgD4rNWN2sIin8NUTY8FOx9tOuMUYF
q+wrZ00br1dRAZmRpjoNP7/gvLAJKqlPOGxRT9rJReJP+pSVTrWXn5I82c+6f2FMI5Zk2QH0HIDn
1puMlSmfGyq+rJgC2Emw2h388BoUZGnLe1nRkVg7fT5ns9BvZoxMW0oJsqxXR3n3J2HqFAXI3DZE
QgUEyaKog/FKQ7vWbzcoEfqbjQKCGMfeJeozhiCW0FOAoJmfBhD+Gz5XuA7W6p6/Z/zxBD67EwLY
DtrBInvz90dSuNeEeyauJie7O9peFnd99cXxQKD4xelewp6WbqqQ686Q9hsmb/VuqTpTthNOzL0I
qGP/hN27wbm6w1ZqThZKc8PsO0PnIaIRhO+c6V0YEvaTaREmCgkwF5mfI1x/6a/YiNuEzGZemKx2
1lNWvafx34dzNbsE+r3+JxHh81AiHVoTUog4ZLHriRShLVMmqyoFsm2z08Fl7T0pg/BkQews9lU7
BSyi5XS7fqBaeJdL9OkHYmKWYs076BYaXGpRGAxa4tRB2wBaNmaxcPOwYXW5QgbXfHEyuSmwbeJ6
Jf7vAUUu2ugeKpG8XtMw/g0K7jESWAlG/UiRF9uObpjOXaHI+3YHUsslPO+asJSzF9Tpbu3ZmkNU
8L5/6EzZerB7wOdJhSPTwSBg6GIjvXBcT1HpvwRrzqxz4LPDAtzM63hCxE6SAtsmF1TkjdGj5G7U
iHDo1SA2lZvkvrMa2U1WZy7Z1puROxFU8TMW+8xPcVPxkGmrnnjZmyP1usbxHzsVBC1ZicL3e/0X
vdl95xRB0HNE8A0kSSYPxbjdYylJkbdyd6KCY3D2RN4n+PpL+iun9ErPOFX8xbtP1QbRDvno9a1B
+7wuJRhKnzFGyIkByETphs6RPLW0OAsWu7jAQfdRHCnTuySK45UeHbWYpH0/sQNwzmkutyTTWsf5
SARVevel/R0UvkC/GSMGv00wf9TNj05VGaFMlE5cNFljgRVzrlytN/SINdnUa8I2NeRJsRNss8di
tFe5xRms6FIWsfLDY6deJAnLdNPJLlAp+AxtEBP27oNm0VNnVl7ucIXxzOrZRkXVgL+Cx52sy2EM
+qfhlqxv9lAp/Ba+JEhHNeUnl87lWb8Q0GR9nTm0PQisSHJIzLTplJkpPKfuzQJERCHbnD2qGey4
JUZbzorPaDJyu3ow/2v531ZUuvmKJ9BwPWrDgX7VyIOgBvYQa6rUaADTbPMhzqdMfOMV6Sws+VTZ
5WwsPC75p6WbSqydml46kgKjoXhRV2xGlyfee6gEW8PFfY0xeJEYlRuxb0XlSUH8lzSDLR5C02Mn
JvoHyVm9qlWipihLlFZmJAYrS3EVXyGsoNVTDRIPhaIh204TwgoVNcEKFYmWnOMq44TYPfUaUA/u
/vM2QtQr5D7M/En5KFqKXD0g6D9d4OsAbzRc8cHxhqA4I1PQgxYQwfkB/zQMZBqm/8cG50PcpzyW
KEDpdMXGAg61wrhVvvA17/AAkT2iaSE2tgQKMW+xyL8hCjTvsbEwTB1SrgF6aWQnX7ep/P4S+I5Z
tPIqw3SVYtkcBxwgcHYhgInUYPfiyMoktdaSO4dNmaqzgNuSpX9Qk640A8yNKujnsFIGCzHwlP2H
bEEOG+evUUEYDX5DpQxNBY6GR7oAYIFMDVDLF6lqkeUwH9tB1bRK+n3N2htag8PdY6XQB052KK5c
lwKEtQbZ+OPSoGrv7CrDthbJWuCsJvILHE+FUtTqNel6UHQROdaV9f5qNDt25AbAwYeC6lbPfCPi
hB8hMUfg+hZiQEWbYiX7BrPItTmcEealtQISvJtl9cqm2MUI9bD12c1qvnVbWgbD62DJp3sIKYIt
xhCG6+gwbnSiSfW8Sh93TCQsfUO8wYdSiuCvWituXogIAVMqnMQ9JBQIk99Jpm0NL7m9yKtW3nQG
Kyyy0s8RBoRs7SYcrJXvEjwFpee6sSiZvDwTPi4R7jP257Hhpcw5dFCMzdiIXDfptKhU9hJSS/xM
2phjjFxXTWji5JDeyjNODSNEgGGZDF6C8Qm8FLToC67hyNJp/k3OWhPEvTyvqNDWSdWeMS00fIIt
seZkdCbzFca9LM1RK4nopCwzL5S8mAvdJSC2wwCOmgIpK35d3GCI0YTWubME7/f9DBHxMxk30FmT
So04/CnoyGA8mgE9MM9xLwmIUB/jbaQ6Vy8ghqYExSUTW6ButzgpbesI8AR5rcmt1rWkOZ3teMim
H/gENQ6jVbkOf/462p8yTMS4tFkpyPRNY2O+3hl9JhB2vRisdyjQoDNEvMacRqE228qU+cfoqUlE
dAIKlHkmBmTFrrLIqeGTwa6qykOfSp59Lz+pLVuoZ+qUNtcZaDtki7aAU8GgNU5rNEKeUW9f2wqc
8VXhJ+kCY0K6uVkoOFXnuAP25YKjT9UEPHmiRlbiwURbJDwbpbVROybCmTFi/jyLzto8bVGi+PcD
VyiNnZ0v51Owe3DJsrbAOPLUq8KLlXEFY/QqrpVwRgjLbz7kwgfS7Am6twFVKbvGOj7AkIWFQtk8
9GrzfvmMj0R/APP1YTSMy8M9FuH6y36AIouQQ5EcTxUmnA6Y7C/PdOR2tSIvNPwbgFcbj69STSxS
PNccnAJZOilPRtijHT5EkJ/uL/rSCk2bibcZuCsBw4zH8/GiNp3lsFtrbdWpfosWTSe0qfUIYp7S
+XUNvIDNshZyrqX5/O5U4XMYeQoq6rx9zxZknw2027vqIe7d6f8rMgGep91Y8MDan7SBtM/xTq71
tPYcyRXcpshrikT7TSvXVmzJJocMHLIZSwUyv2hSV9LdFimgiRSLCR0h83FwjYHjGe2Pq3IoAlpp
iWiZuCr4IF/krdV+HCycy+nbdvrvtiNR8909oBWgg4RF0LXhVCAo7995A+bA2+HdImnvMtwgER83
kwv8UiZQcb+wG+292Pkl5vV3ig+hs+szjT0kfYpIhPFVBA/askOQ0ElfFlJB4Zxb6lwpqzf60C2Z
lu5EQazxjZVi8YYTqXqhUkKh7qQZS0lH64O8RV4ZJKuKXikKWm0DB0NOG8lJT5GTuW59WtYJUqbh
g8wncdVqY6a8KO0u6UhOprCCex0N5/xhrjAd8xf0PSJW+8yLbgQ0KCDO928lnuNhIQaOxOz3+aFC
HYNI6gdnyQA2UHh6axFcuPtgBu1aEOS/ctaIEcE+XSULLbPgPPMiYZg2t5MVHQnqOk53M7RCcVNL
Zto5N9eBJqN7E19L500T0OynV430OPky7VcRZMeEpl8bC+XObUmcNWitAQ8AiWhZRv+CbrQvjYMM
nmrclSsCTUlrue82BprSvEIVOgtzFUgO6IhjLuMrdGCKwplWsacOJGkaOQg7uunUSFlUDXOw8X4K
eIL8ou60PnpFkzdDNIpWIxeRyxwgex59n1bqLdfFGxLByYbyr+mg8V+vQZnL5ae2NKZCjwcEdTpI
rkysLTlXQxpaMYp4Qe2Gro85AzeCd4Mra8Ikzl0RKGotqMe7QNiaNV0As1C6XxFa1DG3ybd2PkWL
Mzsb3Ln0dIRa0YoE8MC4rYXG1s9YOi3I1ur7DsOMIglHWfJyliyYp8+gByGak4vywkJaa7Gt7AcX
FQG/ZkMmI0iORTHctRIH3651ZWHv2zpUmu6sbhUWodlV8susAyIa2a/E/0CqlZ07nIfhJI4vgxIL
GmdqwEArThzCNNeHEDb8ghaUUyazUhIItXPgfu2/uoY10npP9KsYPLmS3hj0xGvNa2U5R9aROt6f
7SoXB5MYXFSIB2bQ1OI1zU8Tu9hfpGPs4SXZ9H8l8efnAP06IuET3gG0FfjA7mbg14vT/mdCjKIs
gHjKWi9dhSpI0HCRDpxfLebO0yFcHHCLT6JNbbfZM8Vd5Yz42rQtp4qEqamQTiTcIqGhvckK2GAw
Xw3tXO1d+lp0MdMQ505gERp/0QRnN6qrwylwlue+/oMN6Gny98LN8E4erdi3Kj91Khh/99laci0b
+STpwnrACxCxYvfupkZ2cOt0bnkbmBEbIi9ZXdqlWu1EYDH466YIWybCthar1PRmOHTXAECGb/E4
JfGMMhLBFO5FiE/lwvQatJzbDNmowJ0yZE2GrScwOdvaxXmsIOBWOyXrW25jCa40jZVW3rJ/AO2o
cEmc7lbiwd52h312oQHsmfWodpp9NLwDxSsO7BRXmmrGSYGb3gimbGlI0z28K7uK1STnkSuu6zAE
4vVXL/fnQvja7amixez78TeTWMNLZyeyzB1EtqeTwz5S59D8Phjgy6QSVDmWf/Q/P0vslBqtJC5N
yZl6iKIYhUeXJOvg8XNSbpEF21FBvUFLAJ/549Ek2LSUXSD+xlvr1wDFemakEv3LbECXK5qq2OER
C7+HO8GDLdZMSs49j0ob/96zlEg4iE1VPoOgRYJ5ZFlhlvyi7LjoNG2J7wXACnViAXMEAL6ffybM
ozaXRalRjqdFos7pH/MxPR3EzIXA/HHBkJEYDInY0UvChSOP7HfuHXQQ2ysr++5Tiq3buPvQ833c
DkTBd7DLA6PLRGGQZfvpoRluPzKvBoqeO1+OZYOsok+ygIg4MMVfKf5FEC8VKW2vooTyPL8cX181
oUYH10zmfDN0t8KASMOOtW+0Cl0xVb1lU+ersl65bYLhXaxAhdcxYmjLTLWztA+DhTt15N4Wibl5
ekv4N7LNDn3zljgiluEidhmcJAay6/aOc5D2LFqOxN+DOFVg+qeCbE8BazEAPhs9LTZPvd3kWr0O
NAqEu3xu9u0hFmXrJ/s5H452+6WqlKSNf9oIDG+n6rSTUt0ja2/dnJpJH/B5/zTjYYwMACYBUpiE
XdCXgxHEULqEbSX+uRoxG0AnnOvJzkJ7EPN9fjv/RKQbMvd2Ac80yg+q0OmMYUxAoRL5izsfOm0J
StIftjKQbAJ8wH0Sw02zzSIYUSWBOS88dQT+m0Z+RXiX0N3Q0vrkyMDCRi7+3i+OXyrAj7mEdMqy
dz7BK4J54rvn7DtEIdlkRNX3weeLUTm8ksP12W9/LjB2tRBlxYjWzJehVaYRy9rPHRWRH/x1OfH3
zO4Tfg5xIi90h7ZHOjKAPviQpJWDREpkNI79McmGonUYssf+LZuGmJc5ClUNr2/tprFgSyU7fvD0
VNALx0T3o0QAb4sc18N1y2l2xJM38FYu3V4HxEUf7Vahy+AeO8jgxA+ycTx466CUVZA3HtbnfddJ
bj7eNHwWBghKKUCPaDXVDDAvV93c57DZM0ehRs4TEXoXcGn8byhIOZY5EaWq5SN25rcHEP1i417N
9HGURG2RzZPeLp44uXH4duyavZZFaMHkqOe5VKJ61oRgs2UsLRzo90tbHlRY/LIhWgpvwQo2khPh
vfGRriZCDVoImwtmZ7yCkAE2hDft7o287El5aFCF6XBhMps7Tr4j16dPDJmaXkvSS0CDcpHAnzMr
0Ygw2E/tpjh1xasK0XO7p0kk1jhwZCPkEEJ4w15GR/C8+j7no7pEsjeT8j3OmUAHe8D6jiaW22bB
//77anlQl/9cOKGlFtlX+xv99RBwjHwlhEct6KEG25K3s1MlDPDWidaKHFsNx+X2lv+RNhEKBGat
VIwNJ4v7FQldD4H7MjUqqAVQ1aZlbhjG5nQjbEBog5JZ7IGtLs6uXA5/BkX7bDxbBQQ6muiKg1cy
KJZGvU88Van2g374+kKFVnvvnP7D+TMf6RswzPURjd1zxZEJWq+JOTHBpS8Av9YezglEZrbdd9D1
ztL1m3BWBaYr7zfm5Lz+kUv/jSSv15D5rcZM4zgXv9jXIjWrOwz4Re5FsjO426mcnwaDS8/Gxixg
Fgvx5ZsNs1pdWjt9ey+gJ+hZjfQi0fGfIA43Ce8kRSs1+Reuk5WhhomvnEIzKweVm248Vpsz2op0
Ee6RDEUKdSLy8JsFIlXqL/xF5EvM+MHaCw8rJgxMXDNgn3x4Dik595e60JmpFhEj2c9U9Pm/fI1b
9InMZmSy0tcBRrUiD3fsoMn+MZZsa00+ri14F7PI65ovE1eOQKNJKg4hFIoZf1q75U1FjzuFo+CI
7S92IoJmoZ6wsgAWXLozcDO1/byA3g84avGCIfGk2F40qko/hrV65FKMLTCDuT9+QshgROsjf8dK
oThqPd11AcN9ykhaA3hp01WERLb1IRJVRaIh122w4akl50F/6F3BJ2LqprXPuRET7kGZbvCgEuka
9NdRETfffEdupR+ZZOIzK1L0/Tx6eDLrxIuwfq84eOVMfigMo92Lk1TPdDtLtzwE64ju0pyOS/kK
hw6eIvvl9+1W/JA5pr0HUMtA3gMwXqjYH5mFywBGqQh6yok4WYhr6OrBR10OuSFw3+BiuxQLMZxY
q2kR2KBjYx8Z3gOu6sfRvHXchyeYMVGWOV6dXoXm8d8UzAyrq1MghgwLs5X77jNJbw95M4sZSN5Z
SxtavhFeSlkv4ZhSXuaxN5PUWgO3HOVw260LwH40ZxB+atI8bVyoF4MwmtaSLuGQrWEEAbGh56o7
qnr0TbrPz+ibOzXTXxgD3I6/M1C3y9x+3ilbqKPNZIW/h8ZOrlJc2wjkMwkwhcu/nbvG+OdSqlsx
idHrTBVKx7LqsmHadY8o9zC15aNK32+1dki2UG8RZXOuosqApViMFSwBaDR/2Rk6OCj6cu8prBNz
a6j3DNAfs5Qpa6xg1kXmJLS5tRex8L/RWab1M6WFv4JAFF9+0E8eO92hm3dn10xHxyn2pSfZBDTM
xMHLVBBbzTtrsH9M6NuRMFwWFDeASAZ08H2LVkmo3qw/PcoDqOBvsQyIdbCJr2faOSo2E/F4q7er
Vas7vKnXAAbbGYmngjYoPG5+NJ0bcuetpylel27GExQCjPYSJVgrsRDnCKdNOAWZTFUzuh6nM2QY
zN1RFKM/iz93QKWaNvUD3/aA90pverVtUqwgqW2/sFkL10YeJDUn2ZhmLqELhjusVZIRBYYnzFR5
EzhXSXGhsqrcFRhiFFWEWipGMVReG/55Rl6PmLfF4hWEWp8ef9xZj9D5aFEiiMLabpVsbS9A//3a
EvDoA16f0VVy1ZPGFMBBoa0DaqsAUrtfp0TyxAs6eGuxxfOk64QewlTaQYsBd67+BALOsZVx2FDT
9bUVm/9C0O8fmH7vSCSL6YKYxHHB2OMskIlqdCqgKEiyAGGSFqKKS6emkUMFouNvsVAdRKONo6aZ
741ksMOe8I8OZpgrlhASjo1nM6YgTOAdGYMdTnZTMYMBqd+jb6EUZfkyMYDPSoU9nzjaq4KFf83v
U4Nfk+d7AuSXduZK0YRrLePip1JnDXR9kxnN4xSrLzjmoZL/cToNkpmsuZGw+n4gfkNr1roO7JPr
WhV2vLifmpm3wk0BzNVCMI6bWXDZEeS650Bjvli+tvTGcZGsawFd7VYoYS8HbLmtMoHT0b7sOZ6p
KCzYewN+/hWrnL5wj+qB/OQPpoZ5qcz/wobP30rH12C2ckpU3qAUt+NrBWjIvE6IObTs8oINvgkQ
dz3IXSWQLe4pCkPjZqQiO4K/ZTMm3zRqzJo/DiTbtTmDqETcKUDoTxXYQIyGUwCboMJNry1y8RgN
v0qKq5TZc+7rp1Anl1hTYmMe3PdvuwTNPQOjTKrFo55cmD0J6mrH4emq5PtpAnjEZK9iWpZT4O7D
hKD1SSUQy3OoJAZLgqGJ/eELA07L03QQ0sqqhHx/hPn8M+kk6iG+ENwcBB9Hh4aXhbcWLGrjiEbM
saA39EeZ9yxd6ywyp/jMIf6gpkU/c5Q5JfgSxqkwU7ihKIdkBMYRcv+GqHHU2YNuAXZy52Z+VuGW
m08CGTzpRQwgw6L++YAPMt1k/AxQ/39wuuY03BA2SZfG/2Tu85Ct/H5l5fEB/tcJO+xHOL/ULrE1
2Xb5Y3X+Sv/AjIGt5TBLr0fENxj5dgLGnpEE+8B/A9/M8lqaqjdPugk2eczkR+vAQwOUsXrI21tJ
xcRHHH1QhBpyfH6/gcPJCbUwDDLIv9rsuRPtZK7W0uRViAYZ5ZDNBtr7xoqDI4mRXCjPceWuuT/v
EFqeM4D347VKFyC8Lgu0WaeC+0fvWvCsUgKqJ15sJcNFXur0rqBSs12uIO0maaVuSbqzoNw+wMR+
62osbMO83YbEPCoGsCutIVFpCMYcX1Sxet3zvuJX4W+XdhnDNKdi0CDgsCrwLJXPCw9cy1gGqsZF
Q1tNeQBI45Yiu/XMzmYUo2Cw1bOCxgDIl3SskO+gHlsoxiUhMN3mAnIWvX8jAirqkfyif/V/sfx8
b7jgGeMT/Rco6c0My7xaZck3kjDEhMo9nfOPdvfQ3olI77wdCKoTULV+YpxWZH6dGfN1/nihj5rv
l7JplLaB2c+qTMxfHmJB5xeedGGkxp8lFK1hHYD5mEXS/mTPS5E3VL1mQLxMc26LFhkf5d4FXmsR
OivCnkVJW85GxnjtnmJmEi0n3EUzth18HpMKECMwYLxrdmgRTWSL6pkVqfBFSCFnVrQpCH9dPdLe
0PxJFxy11qFgKkiNBi1j/WHqRqqupDonLLBofhI+GGJwriTdqPoaAIgZSEKFsPj1aCgnzimVek86
6OjQgYBcLdnRumtuTF34cTlBGaveZYdGLpHLi9XwzVZjjXuuCP+NI4qj4LyzF6+fcf1W98FyCu0M
eZI9ynQbSPb7Y1XGBg9ZFI1Ubo+I1LlSdxHfmxDwUPvqVamqQK2d8rSgQqo4JrmcpMfq3nnimkQB
OXJpfqlFzUdyE9TrA4rDCvuSUvxheFVaD37LLygsy16X7+yufQTuIJAofUL6KzrD/bfVoHYotvJd
04v6S/9/D8ARW5pZb2A7lrN4HO7QK02dZlhm9ylldoCfc081njJiYYhXTSJvbnly+QTA0tNc4Xcv
zV6oZwb95Dloe79fjnC0kXsYamNbbJsk+rMg2kY8S23xrC/rLQjWWchoNu76qVqM9RnhS+J37nUm
RwQ/K6X0VSOJR5Ee8mbVMwU/fvKWpMZtcqu79OJ9h4kfG8p82GyO5Iue7Q4mhHI1pud4KSFTtdTc
rNnottGstx6SRg3Vw9gPhRAuMn6VR/HrWGTynxOcIzNSr81+y04px17jgRG5TpPDv1pYNGxZnXlC
nQTEK8FnqKJ5DYiFU+ulVXsHQhl4OYymCWzMO5Rate+iQslNlc14e1Sh0jIcAZ2ANL3JlxBkAk/O
KE57akXtCLIQqtBUuoDPDC5w7xgaM+5snfQBAMq7REWg7/A3XtUuhcCH9PLL8ehwaJSiPjEP3k8d
H0BHlaueGiqbicYxeDITWHXMWDLKOsZ5+PWsniQq0Ulm6LOjksi/U2Y0Ut15dQUZjJYqWo6G9nK+
frBwfXIINK5Aco409vfSkzSUSCNOCWXHbWAQ9YYc1FosXFa9VIjpl1/yRxVhiSP0IUTHg7SOBs9d
+5tLs/ydQ4d2G51RlUlroucJgIYZka4jEU+x8lHoJuSbX9ghrJ/jCB/VCGAoUD8jhLHT2dSX/fu/
2BQnPSp8vSTqTWcDZlrgfWymoaCQtNsZEn5Hnxa/dEdv0vdm6fKRG0bLThrRSoXNtGV5pZVrZSy6
ffeQahUNEhmWH/SiIhtz6TF6dSksEddIJPjipVgzB776gbVzZXDw/if3FPuBKsZkCCZhuCS3tgm3
A2D7xig39fUK6HEr7G7AAL20rRx2+ntzK3M70ZI+QKvuPZ3UWkiERZ51ZgQwN+iFCwKRUx7EjCbH
rFcSP3c38QjvqGgELB+GOmKRYaWFIwNEYbxGgy6N8Rw3vP2NPYE+D6+1ZrZcNCV3O7Tlt90RXx2b
g/bYbMgawusV5cj94GXb1OB5hORa6Zb1MQVsAWSxR+VpXyvtAPIlOs8jmgdHaCHl5d/XDB59FUBX
/psuAlJUd0PyP3y6oJoJkBAra333N7wkMJp7ia3CRbs5ndtfVmbqrYVbkzLh5vaz1DG+m4C3wS1m
jlx6NCs3eUrBtecwWHm5DlIODrhgYGclCAWhKGvu9hKyt5IOF+kv6Y2IzexIDLQpt1o02rg1r5UM
wQDZBrBvpQcw2TDZ7Y2wrOPjnSwQaX08Ngsl1Giq9to4W0R7EzoNtgc397ftWJoWfBvONIm4xKY9
9+4kZDLRt7+nOBkV8z+lHhzS6bcDZmL36aC75OBRYymi4C/bjOj+xCwqbDC704KXrOh6e30rFc2G
QIQZxml8nPPZIzVVZ9VsH5jnH0QI9/cNLKnnLRgZLN0Gf7QGxzvnunJqbJ8Y5RXYAHX5b5mbvHWP
br3oBOIFqA8k3RnERvMot1v6XXJ31ONngVsoOd7Yg39vV7qvMT2/oD6txC/A+//z2ngUuP6ZBncF
ZHxAME+BDMwylO43rulN74oCm2fpti4JlXw6ySgroLdmCTMZRWiHT3zv8opezG3wx7biz6AWgRkY
UoM365p3Ysh2/gc/NbeX+XvcwNXlhYZT2W7wrxmM14t2SJErf4uh5RrZh4xUw7eeTb+R9CDtF0/6
ly8ZFq2kDvMDIihoQ7/Mp7gBxHgZ/NWdOVJQqRGmAmU2WdtLqZ91WXozShHPSdVi7JkEVv6fm6nd
zrfsncXCiQ4rXrQhCKIjZ6UAlNboe8vjvVudkag0PE4rgSHpDJF/3rydRR3uGVSv+C4zYJmPPKnu
w4Ev5WWk9B2onOruBtPpEZabDGV4lPadkLq5/ykxlMiCKPIssRFxBrPhP7K6s0oT2NUlXEncuD5d
41/YZdBU2i6iR3unZGTiYa7YhqZCkX73gvWd+InC43wX3IOgsGoHTFLm8FCGMzA8iw7EZuLep3ol
0a9YtxGkPwTp8rnsI3JngMT5ykgxhLi6Vk5tXOiM8KKP+/RiJ4/1zqvrEam79ekKYtK4JnINP9gz
xrBbam3sPEnL//6iqJd2eyoQ8aZ3N9CIZ2PXXxpwUCgfXxBl9U1fV3clQEJQVxjRFNFzrCUBnGmL
agzUwuHIz1YWQedjy4DO1CurhlAFoyAKPEAV00yJ7xACQaWVkcH6rH9AswHlUIa+F9fqw0Uxe21l
xeKcWjooMUpHw25aPZcxn5cfHuRdGLgHxjOJNGhkXJOeP/9wl4oTQrVJ6957a+Sk3/cAqd1v14ei
qg++ud8SUy3lZMkz+oLglGHR6k2RK7ewu+ARxFkLvAxu0Gyf6L1TPFNS0/buhiofEJbVEkeDf2bK
u2I4JkAUuT6VcLV6k/7+4eA5ZKQguKoxKd8HUCjEp70n6s8fGV8zqR40azx7vCDY0Pkt5I39VhVs
SjLYng3nbiLMQ1TRg9rAkFnZGxhUNB1hAZY8NtBvnstw1kYSodPbREaXhvvJ2pRRLx7pOuPuF8Os
ghO4opQkWfiUiAGzmpToTP3XdADMRKrPYfwcz/Ehg+d70Cx4UGzzgywd51rIhBoAMyiw14yuiNAW
yz1hTOxZDyY0mFTgMDgHS8z8vBt+ZmuiYavDN1Dkpzwea9AY7lF/bWM0+OHbYrpPYeSqZrO3JXUC
mQB1Q5q6q/6DL3y1AbSlKGMqHrvtjH58yRHdTwy2LDej9+CVg+4StOZKAgwSRA9/tEEadtQg9CYG
f4+g4LpnFrHmizLxS9+fl8b1Als1tU2uVUOJlsehvR5jXpeszdLxMwJ2DmCTIxxpdLt660kFMkUb
N2KM/3Y+R542gI35SRc6PVNTKgKy3yscYl7hAfKbcl0ZhCR7HU4WeIR1YGVC6L3or4rhSTsyea7q
kyB2gGkW63cXgKdAFwf9EjzaxG9FQya59nCuzVII6GPoggW+P6PtBu0HSi698/7lR1+7bRJP7kHQ
uQBTeQsd19cy+6zgi0DiF0b51bqGul3+aoeQHeD9VfhxA/sujce/WmAuTJs9JiKfCNSnJ0mtlqce
fjioLSWFt547irNB+9FsJhdK3ca87qRC6n9XZm/LvgOrGApiQe8w6rQi6TRcfb9tDSdTMlDcOaEZ
5spUNGnc6nZFN5SdFtqvZV9vttguX5EtfME24MAtmWBU0wekgC1NN5bS5hGxrd4Bok2yKtMeJrwC
R4iGnFfyDknbmEdGsMGrm/3V3a/Jqh69jLsd851yT4Aelf4PS6hB4v3L823qgB+CXj230rNBTyw5
NfpEroLb8rnrHSd8F4t+45/1/j0XVvLKntLXC3njGn+U6dKboFBZRbBFdupKgMDa5kBHeHTBn+yB
YesD9D+Yohe+jm+1EsLRyvGQw5mDvJFkrJCwEdOGyNv/cfXR+JZ9UwbQ/XSqeIzujWJ0Bu/6qvww
fn0vIggtyqxresCWkMK770Z9ALjziRoqI5CltZqq1aZb+GISikHwPQcVRTBxVdDOVnw61v1Lp1JK
rIHlEzrkcoUezPCtmEipXg11ssdd0/AOwocs75Rc/xWNjNI0mrWeTUxxxslIir0HL1KYf84n0Jpf
D6p0jCjPGo9OrVei4fi2NhYo7T4urnlLZeYkoVbAmNeyq7TiH6wSmq3POcSs15PYRBBwJ0HFyhu7
0+t6JrlZeaFeVV0tsV6J/snZ+/UFXWxP6OgjPVxWTJfmfnboYHpYrUWpHod4JoOfcosCN/G3/RoF
ssWDVdPVZgVr6kH9kBmUXtLV3flrak772qGgtDjqErEKdYewXH5F3UKP2L+hWDK1kPxkU0NOCCmR
AVQCCMc1lW+Edg8JWzUQ93XRig/ZTmlRsaPON+nkAeet+OYw/pUxk92Nd2Bi5JQf4WbV2xdrX+hy
cucoY4lFKkFbzt9HySJXIY4n/e/om0pNg/rZ3TLTlG3AOls+VgxvDtB18xnQI7tzVor562jedunY
sWTjWd3WRb6P4GVa2Z5GkxJTLVqzwqOebAs9fagWo/xXaablRumHLaITDevQ3P+ocFl8s2GNyd56
1LAzaYTHwCgsu4AFHXXr9s0VXUllmcayu70ry9WSdMItX/lRcfh+LuDM8zOMtLd9tnIWekfzWcQp
bQqNRKlU/otunV8BQng9XcfmDQAepY9SXpYu8/EWdGIAK+AX78Wraa3bVkcS8dsOMhvVHNicZl5B
c2YeJeV14OhiFkxOBTXAyZ9nW3wwlMUEcimrGpT7hzzPjgLkOENAOawZIpap+W1ovV+rkEhSEhEF
mlcyqyezNMzJSzWm1VsPQxrkwNCC+ozw3j2q1ThPGUxuDYVM3wgXRKIHQFuF8D3ibNj9/lZfcN8g
gy6cIgHusAR1U6H7J0Qc347sbNhgDd9etLb6Zw49MvwhVmba7NJhPmcsBLUWl7bfbzQIT35XLy8E
C7fo9gyUpFL8jfr2l8mg/fpJK6u3CCkuC958MMKyYKdD0fyqtNRaN20e7gPWgg2RlZF+GBwoX6Yx
oi54t+eX5G8nrXKZULSJwP/Amoym/6VZXWDN/Z3dYNDkuql8zLyJkx2ecSoUMlOuNVNCrsHhrSNB
vCmFae08x4J3G8QLIcCDsO3i0cPY8ZpGNISy5So1jvP/UXflnLIq2KKd80ou9c8k8Zr3oVVOq03K
JDiyZ352mQ6IEdrGSu2+2Sw77jS3o63AD6WmCd9vBOHDgqkjt/JErG87Oq7zS0+ZzIKD6qydF35W
qQu3WryxbTOnYfzfqABrhsXEfOY3/fBOI+um14oEr3dbTQroIhnU/MNny9kaRyiwq8Ci2XNDPK+Q
7dhnJFCsEFyX311Cft2BSJxpLrSygPmQma0jcqZ1t6BM/0KeCpEzK3OFdQfW4Dx7xd2Lpg7k4OTb
ddI4qzRmrYgMHDePb+kPLTAOmSst4ImD7Kr+ne4NPukc0Rsvza5SS7+CiFjQRmCs0nOE84RA+mF2
qaBot1U1h8jECc95JOUMf5VRkYlzaNSBqkf2CVmWfNRUm4/WT76NXuovH+CoJMOZ/VDO0SfQVRXA
sM5Vthlmj+dqc7bUTnb1IXvtq8WA2C2lmbwDkRjrhDDi1XjQVDNndibCkzf8YwBBMJA6hG6UV5Co
7jub1G/0OJDT4Hy8cHlIoizor5J1Ol7b19WlRBw/boY9ibJydNhZ5Fy0s9GAC4sfeObb0Z5d1O8B
0R7Jot16+PTqn9xxB1fkM8rahjHj5Ba2QjxzL4JYZzyzdt8L2Lxq80sTYOU0lveIvk3dbNvIHtCs
NXjA4LTLVO9mTOiEMbOivyxoCIqxfJIQnHTkRl9jPyYpgQYQWffGhtVkGVT3/8G7cPjp41gmsgG1
A05xOQHuJdrF9RysorDG6a5QmU/gF6mcfYNN7ASKIrA2lEnGfVedMxReCbN5XpCfS+/ZvnT7F69Y
7QR+PX0xGPcWJGz85oMlEuvQc/xrFsH1zodff1HsDfne7ZWUsVJym5Ff8kij1dSeWu2dpAYtkzqP
BUdGFi6xxcCHMIA4e7C5ASrLotEh5f4A4uRCfkKFFVwzkxmtM4RTMhdkArXsj1lZU2s1P0aUoB+q
AaXY/cmUYXH45FU/t4ML81/ZlY7UkBnpOF27mG9ovJpttz5JjGG+duOQfdouKXt4XmbQh/3F2Ccc
cMcDx95wfgXCKxKMkCLKDLTZAyS57AfAXS4dxtrj7hsWKJ0oVp7SHkPhm9FK3QZx3srVSmH6PVz4
BlR8IXwLUh3vykpPiTCFWIwI1LTrkklk2t94T7RSUMsPBrrUmSW79at8SoIElqVgat4Scmk6HP/i
4agdUvO22RjDBuXBuvBbmh0di/KOC1qce+LOLJLJJuWZWrW0BYyaXm1gFLiW5jrwlJ7UF5ZXYCgO
oH7sXRlsv5Ohus7tDT9xmHq8d0VsMnjf1z+JjjA6dA3zFxO2+yQkVzggr+o/ICheZgF/4+e9hsxZ
aPvMonB7s+21JwZPwxW6yQVjNNSWUduAWqfQRoDpNDW3MegWGp5kRpEHBXv6QG5m205SPMoYZOvk
MUCkwXYJwKvyi8e8m870aJHJIE/5jS1cBX3kDZNL28NlUklEKFUiQbNdXHftGyd/LM65Kw9y+dec
2Ok4qqGbTN2yUvfnm8IzXR1I4b1rzsyzvOf5E8WOtJxM5/qBh0fdU8O6NUx5osPf37OZeC4wlOdo
G8fsRAU+OWCi9jT+xoi28+25U4MZQWR1ghqAZfxYnpfgO7eBACzlsy6R+aRwF9IQ5JzfEOLQJmVF
nuqg051GmaOBu8qoZmFc37hNmFZ6bWC7JQdo4b1iXZCl1F1g1zFHN7COOiavb7huY9dr9hAG1WxM
hJF87oYuunIJOvclaj91+3Gq96O9YW5+deXfBmZTNUChmsV/pr32giwDPca/FdwOKSxsFaWk/aWh
BxstKDaG7VWBDp0YNc11VXAA0wrIG9FXy9pRMSnNk5Fvq5j0PrQXoikj+R2KKIsViDh+nsgvY34y
wb+BEzk+fqrFKzWqg/K14A83PZgTWswBqZyudRTLQVN7Uqom9bO0xZykEqlCSm89fhfkTzsEEnOS
Df5sJ2PSKPTV9oe0cJGKmfhUEzK8U7H4drTsIIuZgcPoFgsaUSxwYsZmKy6gfR8mCqvpvFyYFyKG
nUBbLqEwoS4oGDMY/cpwd6aWbaW6rLiIr4Kqa+R+Cyo4PZioaU6lTYf93HGLz6PT/svoFwkgBrW0
GhPff+ZCklmGa9MlnznRxcjKSi2SI6lyvhyht5o6ICaLSfHAHU4Jf1VG4qDs+Y9+ahGZ2YU+O4Hr
dol+GmuGVyoVmZ5fe7+tYCrC4wVWtFafpZSb5C5bvZ49sq59OIM0/Zq8VnDPsrIjO+sdxzUaJJ3o
QTUK1wiZk3DVxtvO39hSngNOxey8Hz15UEazZvYKduDWKJb4gFl0iurOAdlaDX3C65iFMHyFPCvW
n6M7lCE0DihZTVyAyCWaHBnWROk2L9Xs8DTwenwRY2CygLmbFFGoaXIyI7sh2+HDbwAzXHXU1IOw
0qpUF8Tnr4cWvHuoYIiju1PkXdyc5iLKvxw1WrgjiW97fRmqxJ0a8FJ6t242SLif4iZs/+rbZ+K1
9oUjkK4DaabqmN+bYFGvEUhzjuYwmWhvfaxaw/38BxVQD0L57eC9QIOaKCRDj3oC//4UJzY3sDHc
m/Kyztkv4geDE+jB1rrIHDgJRSf2VnG+jCmnUKkZbJEcx3647JEjYdZNqAdIphoiOMg91KutHWrd
1rtb3bR+y25bdPg0o7TVgEaxO7DxgepYxRNTI5KUb6auEwkB2ma33CVi1sdVEVNN+6+UatrCEFGs
MO1QFCs6Md6lVvv8xSzEyAiBNEzlmtQFtCmUwi0jA1QQmP2gPc1bAHG8yOpHu3mwwYUiqfjCdk0P
i2AC/BcfJbahUy3lPjlM3Z3YmAn55Vi0m82+0YoxJciyqVCn8QWvL3NSMD31kgvnTaRkftPM791R
wrx4wDLuLp6mDDXF3khA9DNQR+Pnh4MpIqTDjP/BnBVv/ke02AAkYKnQPcJAuov7wn2lh855j9Tg
JJLZS1LWrZiantYyCRMW+1/BJtK7vhaIMnZ16bw1EW4om60CDUfA+PSatnuI+77x0Os4e/yxpjSw
1wxqZ+rMqRMCpHXkTGsVn5ax2XsnSRhPQ7W9eaFAcvd+pG4mbCXd8d77vjM/QdDQQMAIs3GU6Hgq
1PswrYA6JtMhi4WAhv5eieHE4qWrM+GPrss0HxTo+0rotQe8aecybmP2+TAsKpj114RXnthxpQJw
Cwyc1L0dhAuh65TLc6U+I3X9ehINyDsevkKpDkIOwoAZLfVRIU8p7bp4UrI+KCT4ak8ETk/8mZdp
vZFm8aGc0weTvwVWYFyrpabePcZczmTAf1uIPbxAkE4WDVddPeYGu3wpOjNOojnMEIvWSgeqKImR
rqNVj7ivPinxXo+ntkCzY8+a08XKAF4Y8j7CVOddxJSS9THfXbPHmY3WrWiOV/mRShiyzjkpUu0F
y41a8QjD/WO0MEc+/DhFnshBTNG+BvmrDhVCE6ZmIhR7Sw90lw/epIoaXnb8f+iSsZ46rvdJCJZo
eDmNFlkU8loES1nO++YrNSCcGpv1CVY+MiXPatn63W/qwU6ZhNoGVJ3X31nyFcWskXSjRSb4PYGk
4kZfBd5p5yzXmkyHj96PB/gZKOewfv5Bp9XVhY9Cg2J1pgE98fIRlANw5R+X522QQe9WEhSQG6L2
JGMBwLyxVVYfoNWYEKu3N6NBdfzV1VChkynf9eUqwzmF30URQzUgc9RFSHBKOlOiDVLuJurpAkQr
j4+wJT7nyCiFSLPcTvttttKNryZB7pGMfv6qDe6FU8U1490HlisodXBloeGpZefGGRwNalSSW+os
LEGsH6TLcjuTzV598kf2zeXLkKeUsWkp3EFW/IZSl6bFMyN/rDe2+2vbAqhwZedXoWDEagMvGGky
VXRH0jeK2NxGc7glL53wtkhytAWrQpvZl6AdY9TBlJTd702pqFEOcMmWq6iXvZ5EBIZaBB5qKKZu
rP31/QCqi02SFo1MsNCbvcngpW705CoPN1eo+9Jqmhr25gr5OQU4A4ekMgnOEmwhNDCIZTlf04fx
S0DRYq/QjZ16mIFg2UZz1eMpOCg1Jrad0HeXFj4GvWzUWzR1HG3JPCKk7LPX5osHDkQXcCBB10AR
gCWF8BDY35hxTiYAPYA6XGXbNUyvda9YRISxcWmFGfOd7MuB2DHO4LiGmZ3uBfjeRJRNVPoTGfm/
p5UATxDCFl1SHVD1fFkdJdJqd9QsAHwF2kO8fXp+qQ68GbiXpS5WVC05Tn5F6z4ayGmXJcN3i/zb
HEKonJCTNfUnYpmF6LQyQvWhQpw9RQTmYMI1UVOn6hFTO62SNJpzML6wXXPjcG7MGr5cutg+Qc4u
pwGqbIf2cbHrk32SFNh0FtdubPmu257hx4bpE3OWifxfwTnbi9JBeOh0OvWktDmnezOiqcdQtb+4
HXFPTPea5Xxdz7tayVmusm2kIMKnzDvBnEfMpViS5rbBRkvK33I48Em97daUy9M5GtvM1r4kyrAh
hiRV1ZvQolTP7SZ+Xk7XJ9pWRfLV1UKlCP3di3IPZ9IM8MbxdapKWy30jdNo/4zz1Xed1xDshvQg
uH95ns+fYzxjNYWqyeNR+AULVbTFmvgXDPB0ul8O8+V30CmUnDerjlmg1qNi9plkFmE+G9UhYMz1
Vdz/FguhDhAEe+G4BxrDXmsz+H9j7KBYnduLId2UuhsDRRi4EhCH7jWivSGqrCFV/NbX5GABjHRT
BG2meoaX9i8W+LzTVLozSFii/MqZtyjq9uPHQz/x5XmKHXEhyEO7H5uwVVgUN3PcsDM6P+5+lj4J
AE2eldXcOcged8j5wlRDu0m08EvjjL3an5OICgUxPTF7DiywIFS6xGSLP5wk7LvvMC9h0AKVjtuB
Wn5a6F9gC2BmggvsxBjvunX7W8/r4Fx4VYRnIfTwrQmOVINr4cba2nYK3sD/KFcu9KLbPNY05fJg
3EE4xvemFfECIBtTCsY2YHWTzCEcuwLkLfveMjgJsUfLuZ5K3cGPlX4TRwhQVbw6poLgRfuyqPt3
TgMK2oOjdoDcdpTiJlxK2Wla9kW+U+1es/t2gB3x7zxdRnynLXqdOuEA+WTkpXaNo6ZstDRfGn1c
ViaDzDgDDouTrMqD7xp7lQgnxif0AW/63CSt8/uGXQLNujX0d7q5BtmByKWWsJRaxmP+ElSd9YSb
b2mgz/IFIxHXbJQplRHtbI3XvYbnohLEj6J928D4vzVrYFdWtfDWnoT23V49XI/Kb3lOegA9tNdu
svT22ON4ue0CqkVo1fILx33pc+/s3CLw8jwb8nUR7pOClFNMgkPAmg+jltU6ZW2MgjGV/heLuC10
oOiDbYx9xQSU5Ug7PXR7EAdgRJK6yJnnjqSV917nhIUpOtS+kkaZmtoMwyLyS6pI+a25QsP8RNJ4
Rid8Kg+DiYc1hkzkABvC1WnRvLjJ01H8rNsuIYJR6TT2/xe5fZHolemSTcrViHDY2llFk9q+krgl
2g49qSFRo4+X1yARBuHexw3XYTySDvMkQ6lqI79Q0Pu2jt5NBEcfU92wr9/SZTARfcbZTVDMC3y3
yhSKEJdeyPxctwOfRv5+y8Hc9urRGjix83hdv22CZsPlXx/35pI1k47cYwLI9Ie0lO8TeUd7jOc3
+1S8+A+CjTuNqCz9WEsTmsFh0zzWsY3H8JsPf+xpGi9iK2MYX8Id5ceC53PddE0XVCPAkGBGipcc
176O1oOAKUN18YEf5lDm0fTr9ZBaGEGk8nnuY0kK1ZHG3A/N43ti0FuGiG5ww/U81ErvTxxNVkfM
yJjgw7+H3eHXuy8Gw+818RRI/rIGjD2F0kqANRKH3Ep6RacF6n0iDmQT1oonk/0UkrxAI/FjFt/V
+vd4JDfPxAp9kbuxyMklXJiklwwLknXR7PIzfL2ZDUPQ5DxU+Pnhg3/R33l/jtAffT+DsR5sgW+r
ZJ+FOcR24k0UQfS68Zl510tICRSZhpRrpFhi9nhcrHSghqvCuPTMF/RBRfkgP62sOilvGr6yQmDP
Djh3Rt6MCdwaT47HlvnDtTff8vpTyDlJrB+VglkrbrBdEFvP4nqID05iUPg/TYgCv0hEHr8CNA1G
I4VQKLcAQWRZeORc+3dRejPRcwSM9q2c04AzdkcDDDaFUVg5JADcaYxnOUXgmLMpXIV5DjSzvV2A
uRgjbr1QjyAyPm+gsDjiSrge7yNqMvRQOjFl7doBOasXL+tV1mmtlPRdQXJE4grmjji5XemZYxYt
aR0jbwcaf2bg9RRd1i2oB9GmgaZjMYeIvz8CXjcMC+wmd1hw1GZWvZOxnVQApukOIyxkyJhaAJQi
0oopTalfLIBwSygaQJ/Senw2EUzVdU4kKeNKtBv+/1eq/szWbDn8Adh0/6wsKhzV82N8WzqTPRQz
crQwvGwd4Kqlsr1CEsfRQqvmS+EOIjgLtF/47edaw/GNIccAnqEbESCt7HV/IIR3lxryUHV0R+Qc
JwsgYRE+q67p1xnjAnGVX5Id6mXBs/+02KpOEAWszYuv1CQtZWAzIna85nha+vCTP5GNi58YxQW8
znYU2BMVKYdAGYmdV08MzIm9Mn6QNDo2ZTndkWD/1KIguCWN/3eLQ7jcshKjVKAv9tTc6E6bZXlv
vE93DMVoBS6raPiUay4kL/77JFqY4R17XyffttiFEyeur4DhBe6ytYDIS2ZtfLoOdR683hSNWNZH
Avt53EBhUkbBYY3sovzQsETka9mUMGk46eHqDBE9sbN5cbLV/gQeHizTBRkaDk6gQ/+TFXDt6Fmr
3UBdzOLeya05I6Ne3uxfPET7XdSZ+qUSBTFfxwM6oBOas3cTH8Vcg7NIyg2cug7jDw7sG7RVEBoo
QC1egwg/6ZK05REaBAtacV/p+bYYCfGdTHpgHCqN5a70Q1U91YyCo89Uca/5SpUdOyVBeWus2ngY
KNPBsLyQcAM3TsdW6CUnyltO2KXBhTo938koG+gyAbM9FMgJ7dj25/nR3txLO9ATYZ/RIkiJsWvN
YOPGoHy7Osf/OHSb94J1T10EE55J3f8PxyOUoWzZQElUBdDHzzgzc2zLLTrwgt7JW3w4wqilkWBj
onRuu4U7RjqpUnFWFwfaQbQ7hk3EgyF78Q/X0IhdMMn6lWE6Tqa7GLYoBEElunDLxzhfCdLgVb/W
XvgL7iLo0FK15NzQgN0eBno3b9CSiB3yBQlDEnr7mvxnBDmd1aYBUqyAdhhMvE07Aec7QIYSviOQ
4FqlFeivRzBXvupu9aTNR1BqnezbHswSxnEyVsTyhfA/SNM8WDc2Etp/z5YP0P9UxxTSiTRXOkUP
rY3cNGW6BtsSDb2urjKW4KVqATzxDcgJ4WJ13qhFQ30mxBMWPCiMBPvWx4g4lSWyyQ4Uh2cFzsg+
hHVOZSdSBsZxa6EegctLOjR0SyCcm6Xyh3lVdsaKyvfgLl1yDpSqXw0TIGLyULkJABGiOuJFGNka
1oZAhx9nWGVbz35dmT0MD8cp+3ii7Mk5tL1mG9N7g3MKMPpQEhpwHcsqFPu1gHXLNoQ/7R0cdStW
vVLOf5KfnP0VWTeHsmI9KRYTxwmVz6Kqj+1Nb754wbGaxZVUiKDHOURMe5fvt3sQ2PwrJIsgeU+P
MqKK3iI04r1y61x/N86DYGWaYnBj5yBGt22QsxJ/+n4gRLMWqnqoYTtV6tXCp1MQE9Xaih8LE8qC
Oayn7dzTNMOevp7opCGePM3QA/FWKZg2GIHMZsFSDFBnjYsBH5xLc++j7RbAzgBQgmtSnV+09QB0
5kWgQnO/9MzBP4RzAtOtkWoOaiWJqW20lcq4B6wfv/Qo6jvcaRyDQYQOQ1zRC3xeiX1rxmHgSgO0
de90Qh9+ByYOmEZL92t+DgdUGkFU5O2YvBdD1cFg6Cj6pxXt83QOcB7bkWf4XkxcMFEsucelV1BS
IbIZJPz+AOIbAlb344F2xyyUnAg/JJJEOhRgKD8QWMKqgOTXNB6/UztBGhScAQzNqgj2+sNDrLet
LTsUjb4d/cof13RyasCFoNuE9UwxOhPa+Z0QN/MsBOGe2aPgmbUkNVQFNPkBOChsOktR90T5yZ0L
AQ5+zkUgIiiULoTWs6yFTlYbKAnzaWTZgp44H3dTZJM9dHe6qes3Cbp8j7NUkivzzsU5hhxHNCay
bBTf+87e3mNbx/J7LsItm4Xmvq3dcbjKBuOnAk6iV6fXUbfIt0jV4S9g/gmGr8ls81Xd6IqE9N/q
MARuscs7hkYX3oFvN22SFIjGsBrPk1TZ2dlGySxI8KhwKkQGWc7WkbpQ6S3X7vTI368RPZYOB/Qc
w30nEKE4kaGtZAPQVF5AAXlf9rLyY00TEZuKJKKtgrTYAny0M4iJrDtF8u2QcQpTS5pYEtdDYTya
CgWP8nrUpVQB3LRzhowG8GZgPvUa2NbDBFCLx2C+1fIrw3OG5w2ZroM0A2W+xmPL72LDJGt8CCAg
xIamMEO/CvKU0AI9xH5SfSQV2/19WpjsSTzPmQU4UAdWACgWLqWex5ZOS27Dlin0z47kYhOAN78K
9C/FEJcXNeQwVhTKRP80OfdpNjcefisxkyFs1E5Z2wE55LSuDuWipadN/rD2KKF0qLhNBII0BcYv
fQwkqbQi/19ZEeFW3UDP3pDGSG1LSWWOYKysNYjL8dulfSScmvWh6RrJ4kc5FCCFcdUHnrLhRtTR
Cst8IyiWau9+pJCFNZptv/dXYdZw8sFeHVNTzm5i1MNyIzuhElVOQnB6jj5IZZh6zILqlZBmtqBS
X/FhKzmKzr8bmJQctdbAMlToH87ORyhRPrj0mvmSkbrHVX37YgHu4U8OvBf0XS15P5ba8W8bxMqI
pbeRhY0G8EWKaQhmV/d4ZIesZR5YpCAOJ666LvZ7GsM5GWD58DNaQSc+u3FmFm0AFfWbaBUyoV8c
XqC9v7rpBc+ibyJ0u6iHhxhKivw3iJ576J/9kQsxF/CQNKz4KEz5qEgy5HfxXrczhfustL0c5gxm
WLB8d+od5YoeOZZTPzXtSV9YVugnY4sOwkiiMxxYVOHhz6bzgyJKL4oL83ublgp0ZoPdr19PML11
EVyAg+xBjZPb6CSqDP8UCwtft5G7MnR/Uo29XjBHT8ZufW3Ew4XufumPfyhgytlH21UBVlvNfch3
QC1fC3DLZMjRv+khLI3LzSVFud1txC6VY5td8nZtC9E5Ypp850hwPQl52USRWyU4N+JjwZOuod3/
mD/WLNsTd6GUQCwQnTO12YmRsdjCPFdawnGwLCi428jRWkHYzL7JleCKwct9V1vXPnSY/3RAVvrG
kd7uyWJmTqEJDZ32muWHxlV45UOlDWNLC4eyPOpfTvssKF0KW0RAdC+g7aq1ltgQlH6IlXXJ4wA1
q07D9TfN3jGXmJFjX+hX199WfRCPZDxymaOOKst3WzX7VwmsozgDqxSH72l6ASc6r09/V6LW/p52
8lrbe6P2kWsiewC0ndDEx3gIJ0ONPzmnhYAdtNRdEUACSJQV0cw8KYlRKYmWrPisiHs0vOe7GRzR
RMKoOqI2BZElJ8YTHjX+FzZDelUWy8lzgjWP10LvP2lQD8DMSEUNgCimecNU3fakmHsPeRhimxx8
LdKmN7Kk1cZcmlnTRhPP3HNiFcM+mUIBoEHF2KEa14ju3hqPrJmroOjj6PeXMCN69mQQhY4I4+yC
1eQqN146NvmAO41NHnvis7L6rIT5LQwtbgkaDxpAlGiANck1J66PwyauLbd5XdNwUyVJb1Cd1VVo
B5ESKF2ch38NHe9kjZ6gqExPh2VQ/oja1H6hmlHgReCiJuUJaMIJZYrTrtEGJT3vsHpJ9Jv7RFNu
PVaoK4thJx9BtbKIrhU6oztlVR/98gm9yiP1kJC/p70l6w5T+0ZxnaCspmtcM0EOMzZc60BsGrlX
mf/qW4mtLhZTUM/iDe7+ZTnyc/mbziL8sXHY3ynps2YTVeSRo0XpXMlWbxvmZw5Xwbs/PQDKdnM5
TFhtdhXl6TKPz8NVfuubWwtEW9exWVLhpJ0SzP89LRk/PkyHA5yBA0+0sEuSsD5hogW16odvmw79
xAPF6c++kjaDKS+s3tatCj9tzY5kOlAZsRJzpjhSRNIQ/EfNQWLI9PX2GF6rWkvbXojV5RLAO+HU
eZTwB/z+A1eNmfu34Qj7IbFT/IR0xgWTVfI6uHivhAE55YMnLdLfAoM4rWCe7naIUmcegC6EiaIG
s4Hqhaw7CeSpGmWNzLxwKgzuc17zr7PNqZ0g6Lx/I91vXR3iJ2Wp9t5h/QcBnFNbOed3ichbtX2T
4WQ6lq9kqUpIcIfEmotoTbUDUoQ7sclOR2w1FUPZui/LFR1GBLpSmuGlctUKtvX7SJ2tiX72sstK
eYf7kliF38uxa2MsecrX0X3eLx2tZ/F7MHqFrS1TbXD3WxqMC32GIxnb6up9RdJJJBaXF1H4XTBB
gst55WyYCDE4swxrRds/cwe2I/jeX/AfSAwBZirAkeU1TIok3DLgz7tfU6it/SBpvK0OES0JOMw1
0/tMYanWNrBCfgd+L4r6hnEhTWfzKMJPmymuTNIqrPO1jwic54FaAQcIbE6rKEZNjtYGr4TWGT2w
ro5LjmQ/+P/ntuGm0W92dfSYO5Q+NuZka6Kfpe4GwzSZtBJBuA+Ncr9GxFpVMfOtZDv1FWoaFCGn
+tipvL0WCEMHuYLNlwyf9uQVrpoQ9s1Dj1iiRe26CvTVYHausr23PRhgGU/VW51q8CHfzt9lMBlG
lv1Qs+XM6ZWAvXIqK8yf0cYnflfQXNTnfLjmKL6HeECU5I3qL92nkWUbDMVyuypK8AA98IpliD5c
KP6mGblhplpQ9ixE2WrczxYbFAdCgw1Ru1UBs3zuahHdv0Y7s9wEm8XnEy7Z6I370Aepts5ItoK1
7FLTvQ1m9rID+4MzerhILu0R1DT2mZaUSgJByFQFrb86kdnqWicuoFdEjrnyYZI0Y/FCwVDjgS4R
wpjvMQaTI3vt2MCHNaIQBE9ElmLY0OjUbzQIVtU3+YolCpK1RSbmDLyc5SQYLytpz8WRYsE/ywJd
nq6fre+3GrO+fOsaTYhgLrv41Le6CTtiI//GRbaQWJ1P56yUfEyokLv4IVW4XicVS+gy2I7ueIiE
1iOqXxtPxuhVL/+pn7nNtFTDtjbavrw4FZIf1B539bwdi3IiVnxpkveooc/36hSbPRHKRffbGcKX
pYnlK5qC9+OQT/hy5s6KjV/MxmrnwY//d6kTIOM1zegj+jHw+F29ROIoveHfgpLem1VptsWmg3aw
zMWjZYzmuFFNy3HiFkDbIc04Y+XhWXL9fEaDnIRcFL7apSd2cQwd5/NgPbM+u6GD1p9yEjDjr1lt
2i7Porpvg6E4YJaySnAMUhOw3geQJuuYaXRuCCeyQcwvXF65mF2frAAR6nxTRcbIYtjmjmiMk2IF
B3hOluPxP+eUXtHYg3md8ZInbVoIg7PnhgXdFKez0ePBdafo6oa6TTwC+6944ZWvju2i0UEThIad
52m65MUrenIlUOi81wCVZgNBaEa1pcKygcaKm914v3km9sfmnSrqlXvwRS05j2mGC3mg/Lwudk8s
7qA5XABt3ffm4whXSjpl7/H7p5UKoDKqgS2V+JlReR4FvCP4VvsoEIJ/AtVSLaEFxCGsbbYh/MSD
ZDWvcnFErl7ywlcFi0pX4RAMD9xdYsMmkQ7JM9QQPWiuSEfZHgDoxQN8VOQH9TLyFLXfZQnarUUS
6UvGpLGObGyH4aZZWbYW11geYgwf/I/7Q9lm/3BWSNbCO4JJjEpaa9AHadV/3cyj2LIdiW7XMtTY
V6qARAi1/jL5VtyJxWyKKk9DZASr/zpM0IiZ+OnKQUTZ2mlB0mw1iZruA50snPDWXIH++Sh+dzwR
i+j757IeIKfY/r5+0mumTgq69asokaRfVRYi22WmJWavtwfm8mQUyvjdKFVfbMHn7xZI88hg9hzc
MX1h3tWsFEtY7CiWdqY3wTYGKROygrRxmDLVHKMsBjiGOANK3dWD+Ai3fdc8/2ojUQOo3FrQDAnq
HsjTtfYIdTgE1AOQYbNFUsL8p+WW7RX963K6jnamMDwHAoP6n1FGkMEcEg3oFD+PhWiBqX+60FP8
bbxA3FIP6gmPw3weGrXxtzMfBNEhmitWU7hD9RPBcVWTeK94e3E+6XPT5M8ye8CEr+HYH+jkqrUA
wUxfPZzQPH57QwtV/cEGUhhqmc2Hj7yl6PDlhgCE6WH6IgOKZ4Fr/ylUN4ecTRX+DPrYfRNhwTYC
5wVBNEzMzNgHR1r8pkPSvtpH+ZSa2USKxDZl3xgLTF3AoRuqz+oybAp2YfVi4KI7Y1pynKuRrUvQ
si/MdYZi+cZJ/gNwQB9q61FnGBIj55PQik1+11K1lxvO0Kz0psCXTWhVJUDm6o3idVCHhLQGPKEy
fZR05cdrJPGKcYgtNRhnEPOud9V+TJ6/3WWOGK8fd4rj8BMAwSvLnSRftxJI7mkCS5fN+sIgQ3/7
wOmLV1IcUGtCJSb2uiiuir9dJy+NNlPi8gRg6ci6UgG4XxRmc4rJiNX31MymGOa1JawmCpndxi6w
ArA815LjmoHhoOeubNevAzK3Mxq3c5gk7etvGBJbwVMFLpDIvcPp8bl7CeCXsuR8h/+qdykenK6f
jrZuJuqUDxVALb1Y63YadRrE9yKsP43EdKBVhfF314yKZX3eu02gzcTWe5Fc26osYeRCQx8HNwq5
YfUjQ1DHjLnu3VWBhSxvmjVAR9oMsN0c1DUu3lWcfzBNgrmjwn8T1pxhqfyON7TiB0h0whVd+pSN
2o65WW7b1ejSlKfQTwa8cAubWdpFLFTTSLwVe7WSoSOyhQ55Rd4rgIclgNUsmY95hu5e95g2A7bq
eQfE7uEqlnYHCCKMqEzCVRholfRAoCp/pBDGu7jvM9UmFc1RZsug07LgPv2VFWGDby44Vl1RmIXL
+i7zItKzaePjYgQN6Yl+aslQUCHPz+97gQlI45quRDV16mCcOFnoCwOybT4p//EP7afbkRJUxf4Q
V/yoxPHB8oNRikPqWEdwWt9KpW01ZYYCbRCSIhVjyVD4sXMtDzQS22uM6VBQjMbU4ioWDK1Oqr3t
e2ZsY32aORxV0AWKWEkWSacDcMGpKVpJXPV5rnMCDT13eH8u2tryrF+BUaOfqOiNBCgFkJhHe6+o
IPlMUDxXvaKpV930rMezFRy0Fag8AJkCBzBXdeve2enaW9a0P1oPy29vd58NHVKB8S53txI1FTe9
how9c5A9RaIPSL1j4iVnUUXPLz7qk+82wxg2ANOoXVRET5Aq72kGY3RPz3IUhehARqZG7bWk9iko
V9TzJBvICNw6Hx+v4IYKffZaT3RlbDhRXE8KR2O31uqfypc/G2Bi9KVmPwvBKMjV7P1ruLJgo+Nc
2Y9OVXa88LjjUz8jkMUHVLSP2KBSuYXmTSpKyYEaOMEHZhVpuCeFWbG2AH73vLSbh4mJPD4dJLvo
JowqrFdVZmFkw+2DzLZqGa9mi86UzZvcVt8yWNddSwMcem0tdIy791xJIW6a3nyQPpWZc+CI5YkV
+OD3yvpF/AQVuTNS9IRKJSYeiZB2FymieTrrbqWFYLyZus61Qy8N1Sw4C/7PcCwtFQFFDa29j08M
TXNz69NHvB5aF1uKC4TMvD5e4rK1wJBZJbelB4n9FItU41aH8OMaWl9oqYJb55cLR/yjx7wPQh34
qt3gAAKGuBpTKoxE84gsthB+tsEEUyduZ/T14XqYXqvJMM8lh5omtLbK+NzMPHmRqDjGjUrL895f
pcraTDfH2uOaUNIWwQzmzBtgHA++Fl3qBqGIEeeDMEbR8u14nNU/4mYAVUlXx8LI/if5CcVd9iha
oD61pZAB1Mob1ehkFm5LYXGKeHifO4TVBMPiz3n02dr72rrKYC1l0PwjtrsVwtq1oI7/uaDt+4an
uB7fus/Q5hbV3tHTA6geEBrc/WOiW2tjnzU7b7+2KuDowuY6/t1wPj4kyEZr9VDWoOlPg1WzVxXM
I93QXbN6AOWXhZS3Bk/PimbeAho8dRWTdX9orAiZErDCq5DGtMRTWKPuNaU0LXq/4Iaw+Y2arcBV
XHezyO4KZ2CrPcehDBLs6LXu3WhpzPAncvYzqSkwOkeeCJrv3ytOKe+VMKrHfWdJ4MNtAV3lStxD
r5ERtrqn//nFaGAwrPf4OtVoyFs4IKb9vajwz/I0PQxSrFEHzlCtT+emmP1RXF54Chb1qrWd5Zn4
Ap7cqBmFycjpFrBKOraBmpYLmTqGhCufD5l9CQgRM/ZCRN61CZ8RjMeo0b5BQ/A9bWPFtefqDgqv
lB2akA3a0d7CEZ4lVuMV8zwflm+TdCRSqTcgxBFXkZvxdBdeN1CVxdul+rX8X5gmHZpToAZbPFHG
lU+QUA34S9ZJOUvlepjx5q/dC1Di+/LMSby6UX2QfESONZQOyUCqocdsf8nLY+IzZB/9Ph1QNM2w
XIDAcAfFZxWurOroA7tBwkYTUUoTP9rE2E1jt4Pq+MQYhcSsLpWI48FTUg3a3Jt0ZO1NlTr0Vnfc
uHlgIajus6HtbaWaDdJkyzbpiTIZ0bYysrtA9LUzA9Yy+iE19hSAgx6jUlparOn8DG4JevkRvzw+
r+hSVJxHrd0OQ0meqedLJIcBnmQoelTOYh36v2HSFjKoUntjlFGjPvVQq+WlJGPbvaCImQ4CTvYT
1+6ncG5leGH0OHD0rW9avt5CM6jNdWS10oy4Sj0a71xa2wfZxGYDd55HlR3+WntCbFaDINUUGCHK
oBGv+DhAiIHz+WSgXLtQ7OPgGcG8BE+4EMXQpPxIS0mIQ3FA92qIlTsiT1McraPfQIVCqNRWbxWv
MvhycBoXG4JwgijaHj7xu9LE6IpXV3bm4kpV+GOHT8X+w21A2YyUrqaQ+NijHHTjOGUYHneuoPQY
+K8vSMvDc/D9TsHZoWWPMoXMIqC400CfXLqJWZbfhxBl4OM92oKpSar0v18xxnYA7eMhHnD8MFgI
W45peneWaUBgZeh9KRKNZq3s0jElQTbHadpzJySBM3iB20DwXATOsPf2SZMV9LxqzmW4vBFca7xy
XxbH14ZlpaamG1vW9+M4U8sp2hzGzCBB6M+8xA8vT+dAggo4d3I0k2nFYOOcvoOvNZFkBQjr+F0U
ic5BoDuJ80dSQgaPVO+6h6QzbrePTSqHYy5FkCbVfE/nCe3eULgY1rRWhGlJRMX+JmLxqji1VBEW
0gn9pxH08pDZMlvf7V0IjxXHKNBhOvvhsb298eprDPN7FJsDmrVh0OzqG6R3mkL9pBmeXu/G/2jE
rmiAmQ/Inja1J9HPFWa8SHeKUNP7OznLPRddpSh6isRYnZjUgBDeb0Q3yWTawxOOof/yeSrju8+n
2yAQyxIqYQLSdYvi3eOBJYzPtrDWTTLPb7sVeRxRRMjPjcJVwoKKM+JsHSVhvMbdyGthYvedMzpb
GoV1p0MEtE5ivgo++MeAeTSwbwMxAFUVjRLb7SyC9uK3bi2wxzGVy2zKKMO9A21/GlX1qWnr78B6
kD6b9bJ0tkDYPAtvOgoxQu8+w51hy5lse4r2+1ReUe0V8ejnnjoggEC+P5B6PNfH4k2yY8z61bvR
N1U+wDwkgYyWFiNa8KoBTqlPcxZjvTLYV/Llr8e1efO2JD0qTZ5stxla9/Sc+6msm0xB/alkFDB4
fvcus1jqX1yzG7hVlFDHBb94EvJt8iDg2ocu+KRhQidJEPbzqPt4SqKZiIud4izFrEiVFJaY4l6d
SKP19e9JdjTdQyFEl/H2o/jXxN1+CVT8z3x7MWK87AqWVkPiP6g3gBmCGCPZ6Nxu/ENzqCQxnic4
IgeddDn7vwJ1K71CfbiwNAu26g6D87B0g8qdUy0gOh7i9sz7JtpjEVlL7pqsrSMssFieugTXSeG0
kZRFFfZvt8YIC4sFkYtOe+fJDFr/ZWM9e6NqAvuxECzHev36hYW+tCLmL2roRfPFdy0X01ff8DQl
bFUfHl9nbcN3Z6jmuz4WL4StQOtqIOotyxPD1lujYCnLzyeKWqcj6CoancigbHswt3G+W0BG5zA1
vLYoLw0bu12wtkb/NYAORJNR9neErac4ZEZf54NvJmBTvnXgwcpqcOrj9jkGo5a5rEbQzWv3srou
wBKbIbn7gzgl4WXGhjLimIYCyiR5SZjz/S8N88ThylZlxjRpE87IouUKOD8j87Qr5ylolGMAl+7F
EqJjL0oM1Hf5V7TG5JTWEaAPlk2LKmToJs5Lac4C+Z5SXnDT+tPNrdWIrinzW/7j63C2tExBgih7
sa/kIXRdUPPVj/vBDXZTqygKNQryqqlysWywqtaw3pSOaOSd7GQ3nyzo63EgCtcP0y8ODslb1MZd
UbGKUm43VbYTp17LnZTKMhPmdeoWRPWrpRqnSFUVl98FQslGS4jPWBOtC21sCg39R53cRpWgMtlx
nB+YyYExztyVbnlHpL6giUzX2cM1qTz0HuB7kxz2ynbEaiXY5SZBnzS0iNWmiuQg6HqKoZ0TmEfc
xqdwpR8ltZplpcAfqVNbcUFH4KRt01851Ix6RfR5VgjRmPfT9JGEAj5dvc86b67lnXdNwWrB/VRV
3goNS135qMxUaTQV+t4avA9zNscybsYgyazwk7q2DJ0mPtNF3eZ7TuQS+aFZIzSpx+vpOOeTrsvx
INRuS+3MQfD1n7LdhLBEecvv5OXOehKeoc5Kp4tzWMoj2xEuY7awZ5d4OvZNCzsUJvUMdANMRBgz
6EN+0ccms2eO0MzUSANXZIiQTFckwgUTMx9BLqXvNp6byifxnSZT/CEil3G1pnXQwl8OnOxb29hy
2JInP8mwd5ZGuHw1kmspexNiAaVEYhrpeSBmHKqk7Zv0Fb18Yxq+0byJb/kAIQoQmJ7POjhC9b10
1+DYjDjS1CAwSNAW7mbfE3c9PN6bsup6eJ7+p2M7SUNtyj6qCUrTmVdkiv9VB9neFADnUTnk0BU3
lGxTZ4NCjW0YVoO2LnQAjq5Ad6WLUXsYmpZHZcQlZ5SRiIZxaZ57Gl8iyvbrGBjCE4GFoM7GSx+2
yCuElYNMATgjyUP7uq1avxXExuaQDjG3RS6PmI3o6T80l9iELj3MqrwnT21PjlG71HbGp5ZiIf2S
bbWAsjYCv9ow+3fCl9e0vbxVboqGgc+kd0VZ7dPEyLBKxXUfRRUdMzWLHA+jilgBTxc5SdZZ0S6u
8veofpz82mr9I1FasxSAdSqb5Mbg3d13yHHdCppseM6NGDoWL7jaayD4nkigFkwtPTs28p+EFHKe
aaxWhBaFhT5QkuknNOV2dRUlQ+SZn5/gaWyeXhRF59SyxWoHUtajga0OCG9R4DF/pWDQMJAAqH0c
NVMoIa1HZNP1avSi0NrAvXmY4XIwxp+Co0svspL1zs8y+BnI9wcej1aIBbjNi2/v93BJDLFqCgBk
xHXD8ehEmp2n/T7qKLOicIkMrkH5geLdHf9rCHpbuiKvwnA2I4f4oQ4TXKgBdL4ZlchKw+/p4fNX
W9L9fGlaBnjE++bUankNDXYSTFYLlhGNNdH5xM3GzH4iKIjT8PCiEmMniEVQ4Ecku1bAOU66cwR6
SROcAxmdAc7owr/X38qNoyle5jcznOFnqlC4mPNExle5ZX85SpNTe+KuY92sYEFp4vWj6FsGrksZ
iJyO4eAmlKjH6sA1W4OQP7849AVxRslRcVAsSxpk8X9Vr0P168OA4gjvPG6/cYYc/MPeviXdG4GY
vqCNeh8SKQ5KSHYLteXEaY0Zu2tJJwJt+m3i/4WgJBb2unWz2FyPC3++xtzzPMBviThQHO/oUiXv
m7We1fys5T9DFcBOqOI4QXAAsePu4XcoRm1fTUoN59RsLh/7VnNWvRaLlNDy1/DgLp088m0tO7KF
QSGuIzoDDQ8rOBXSoDixtkpLg0Vb/GDxDH6OX3SDnOynLIXLVytEVleYQqN229N68qLLnSwOyDS8
NKW7gHOSbA8Kcz2zmOqJCrY9ddmYEH655JV59THCqSuLjLC62cBPNBENpSGvf1tNhUBvFTAgXTQi
eIYQornQYV8FwKz5H4fG49sXdH5uYJkxXBTLNHVBJDKSgKaN8U/jHFKMizscX9Y7A1YUsNpGXTzY
uWrPgCji64+WFrgFQ97w5WJE+ZQxSHfRpwG3mxQpuAVUDMWxJhiP9saS7kdP/BAQmm/rNq/Xa0CU
XLOU/TwGaa1BEeZVNfMVx0kdevIm7aHXsMRRoBvLHK/lrjjyDXfsJeXXPu+m0dkQmjScEzHG5N+p
M/dJbRgAScabZIPC4dHQduVl9M/iH8xbZ44Y7u0qwKJ+g7PYg+IkGDHKmO/76IFt86KILcubwTaM
CcH2BTinQuYUnKMukuxZxhMWbydaGHDSk1xxy2MGwF6j52ssLJMcFZZ6fvHvFc3grxRe3Hkqzek6
IB8MLE1ZlYg4VNeWEiKzcw5TUqlnjJfIzZ5+Q/2ksfMABxKqjDjgT2rvpELi8JI9UiuVnifIYki6
mf7wCVEhRkm4SG5nQKntsKX8I6L1T9w8sd64c3xaxLlfMNopZ9YFVV3S7mhN7kkcI/EtNMaw/ilZ
4x72piaxZsjI0gZf14T4+9tXi3ECO6op4DoknkpTB9R6kxpsTZPUMNcgevs+0CtF3oitEXHGPHbQ
2xO7M4b+BhLlVfxkpJ1wKMhB92v4GSF+m6oSj34i9R72b3rSOgnUb0mHblih70+bBzsf3abGYJGG
Nw6aR+grW+Gdct7vMGKksed6/LnaCYq69pkkka84qNJmY0OEPRpXXuiGrVEHkcvlMucDbqDvzUV1
tDhk0IDkPf7LRxuxcoBA7kGOA0uXoSwXR08RfgxuuEb4WWwmKOpzi/cx7PvYePy8mCQmyVkv+eVI
MURR/2FvxxCTgA2Ta4avQeI/yw410cPXMm387IlBHqPlTRdJkpMBf7w+NLgu4gBm1JpFZ+wbTOBD
UAZJxRJ9f6gxjy2VERLL76ZkLumXCPmzger2sIwnToj67HzdvDp8CWTBXYh/AC1UD/t2pT1D2/s3
IUwSmA9OE84GEGBpt0dYqpJqectqoxIHM/K7aFgjak9logLyMnJtiaRUvlN3t9oeLVGLABLJWq/w
1GgsKfnq0vy2jbvmvmQzpGVcnkvq4DwyGU2OAnbMG1OvtVi32PmHNoeTwDtCjL4wGZW47v8teS8t
YnQ8qmZQTrbD2rTjAGHz+bqHZ9ZFORiJ0hKSJKBbSxh/bvFpJZDcC/11UTSmoOeEH0Fmk8MY8bOP
eg1v2mGqaOCLh+51GtgZLD2lFeG7oOO1y4xccBxZbBdpN2FCT2albkNRGpyrxCM5w7FvukX7B+zy
2n18ggiJCppvIZpes6t0c78sJWJN/2gYuc2hfo2turMLa3BMWbyP7MuVS45t159p8AePb1RyCxcK
nQJdCqSk4oyqfC0rdrCEYrv65Xtm+Q9Hx7WKIHhAqD8eguLrTainFjJl0PWPDrzdEenbvpneq6qc
ybDyV8XS8D+8B93GlbdLkNwrvXXGhjqVcPioWXuqRgfTokU+v46tBeVw4ox/BjmS9lgW78cFYZ44
gU1RCNwZ/doshhtDgCEDc3VX48t1wBFZ/3T4Cg9oKrOhSgbAwcoC9jaohP94Cxxo0o7yRMHUzjoL
NmOV6IJ9VBZCSnBri7MNdubQfagVxb7tOemlbL5BFqoG0jcEmcTEZwrLrQtzp3oNvF6nG68iv3Re
cvol3FlbnsFE7JO7OVrI+RMgJ5p/78wL9lrgMmfHiaF8GJzCAU4Kp6HGPveE6Zdr9NY9S+KAiZJG
9wSQcYVZFXLZrgbZL+H7rqg4Onfd8jLlwxARiuqrZG7xxvquyYuUJcX+9cdH0CaXGk04W+Gp7pmM
LHoINEqNsBgAHBftRrXrp1fVRVAxJr6RGncXA2l13iEmuV5Hy4wjUR7q4FWBz4rOgLDEXsssdeTc
O2ywy346gGWr/O5gRmH+NSmIsLTsKYlh998CeIsE8DulHbZCLpFWDawzRsaPiilFxvYBgRcasKx8
XyDWphedaXdaqpUAJLlzpkuY8Q9qgCwo26CnzpgB/SofddjKpsMUKeiMTA2XyXKbZXgG1xzmpBQh
0OgjC97cluNxyNKDeMKY11evrHYJ4dGl86pxIU0unPbREklHCpyP7FIWXtZq/F0Z30SC57WniiDo
qytkI6XjWxiqqx0ltaT5a5Tc0u2pAkjseeP24SklsDQNKiLCHfd5NP8CSvWsfapEIuNub60s+6aB
sbHlumwfmgpyuF1hDLIfTWuYQYU6R/K7qiHMr+WEzwAIbsq7XOS31QDMluuJKtDYOFLZ4PwxgT4T
BDh8jbXV24uCgF4/R1sL95GZR+RiJndq0424plZTDQuqjEu8JAHGeXRvC04OCRzdtDGdQO1UV9UV
T3lERiJHDntd05iNwqVVnTOqy9PMEhKvmWk55t+pHYSgbygKZVKjC5OeH5l6HVBu//eWBWhSSf2j
ez51OceZ8mQhfFNltUc3cLzmJqUjZyvbGVtNB6HAgY9zQjwt1gdk5iwLG/aDoz+va4iRdb3SiYVE
fIUbZ0aYxsxxPIg++ioRh6OWKlQb5gXzLdZdolUCBVzBi6kNAAlYX9WZ2rl+e8FeQxig7KrilDyN
m0Y6zebjfYPTLDhWzZ9obOoWCwDSQemI201/88glshKxVPL/h4qHxToo+bAHz8yqWwGwN9X1iHXg
HRj5yf9Zi4ittcGwj69VVFTi0y+Cq6H4lHRiDPNHRm911FdYfxBB8qHXvdmrVzeXq2LFvGtUklLL
OItdeyucCi+MmsBGkN5h3DfQk98+TtfUJAUXmvsHcwkepVUycMzFTNydy5ugqWjbdtX9b7JJeJXZ
lcF8kHr8fQXXckYaNp3oF/t5sJznXgVZ/4cHTaN5xG2dd5Atb5DuhlY+14aMzS4U1xBtP81LNWhk
iXt1LRIsA88Ti5U5d9kRfG3WO0larFH8YEObcivgqBBfkIj1se/d/v0myCFzdVIcbvGqz5EFIUl1
TJQ4EGUnZc8SyD8/kPARSQHmebugasFvDgFhO4zg8n76RCoS+6p4jeLueR6F36Wk/B0fSiLb5DwI
oL1jwBxQGjXDpeYefoGzFpK+NV14it+zX1itA2eJqINfxBGLHX5Bso5qDiW/n91QMKH1bSkANQxD
jLrxdWPgZjS2gqLG+OCIXYVM+Voln8Ppl764gLorNgKEl6VhkusUiUPB6QWrnOtohQpkH0ETXkDo
rb6LCC564g25Vydli6LmyRcvWxuaHNfL/EKkJwpBKPccdIrLtvCHuj7rGxW1I2J3h81cYk1rWPHP
1+lDKkHcKlbmE4q+E/uUBazQTS/Cf36xk5w+SdM6OsVWX4aFhimyUg3NamJmcaDVM5p7m9TaU6SB
86vK07/kIPy8mtl6BZO0wYJU17CpQ7L+wWgAKF7/apU8Tp1548JEV64HWJrwNesSbmcjAvndh9no
i7Xp+gbtREdBbFXKuDn+F4IJWKcLR4i52T8XqvhAMF7fI1ZoZd+1HCK4El67Q46FD3NBZ9dsA/7P
C11MplHC9SHqe938lEwO7zh7EBxbP/MNRY1WQ3vGuBEYjvWSqKrU57cE3sCeT/rOo9idKzK5Yzrm
kiVA4nDULUvJ4vaMB6qmCoNk2ZOpBKpooSKjFrsmJFcHKZaDQg+x4k8j7KUSYcRkK1NPyQnzkQnk
0zCipsX1aiijizvawvlNAV2691EjN/A9TM5gxHYj+lpgh2HBitUkbkHaCNYTGzaIzDxNagKk7zVk
LLONcdB2QaHsUG6ZedukeIhkpycW/qlBitG8LGHHrvtl+sfzDp18tJtrodIzsyd93H/wR8ZoK9UE
4Cj8Hj75n6mE1FaFvma2D78MYzhxTSlEZWbkCCUtYvYcBY5QcKPNLnIS97KnTp9ZQ4HneXekGk/U
igpRqRNOlPy0QCPY0hN6XFtXlAqsWA8zN0SVAYJsIgzoBaUjDV9qjVd+/ptz8j0iIRYXkFIXMBF9
Cv+q31EatZRIW4/VPSESTVy6LHHiQIX0wyLIBSg7BLBHY1uF6aNMJMpKQkby42izS1WccdsoLb/q
OeqzAtDCMDavXLWK9V87Wl887bddqz0NJRVTxHAxNU7u1PXXJJZjBAC4E5Pz8LYdQ4R+U8a0bm8I
HbwIo46xuzt74wuuPlmLooDseMabmlX+ysxCh7+yiQMYNazUKZ7EoHtoiPp5bVV7VItL0nHHE8IE
OE2ZDmKRW6TGZWaeND8BoywyFErhEP8H6oXFb4XmmhXtdxTJkhceXZE3cc3lqbpqeavvGP+vscmG
Jr2qH/idF/qMAGo/eBXp8JIIzlnNJ15FqT+QAxIihdSO+QhUDN19azkg9/+fz7EmwXGdz24yLxOW
khG5zV62/mDuPIdIo0jA2uQCo0u8iWza/x5tVATvWGO2ADcZnTlGVS51OuzrU++PY2m43hNYZ3R1
6uqCi8DYSEy+3Zu0HcRBR5ALyF7v4Ht2jmGZIm/wC1r7A1eF7hUTmBzokcI2gO1Pk2idkOma3S0d
arN5LOmdSxIB/FhdaoakAIoQQSPY5TENkG0JcIWB1HswuwhdlOL2A3nET/+rbkX5TQgtlEqxT7cz
YUCOYWBKbfQ10DhdHPK952s9lWdoex5Z6vnRzEmH1lS8X68PEBZsmpLOZCRlaFV3rahaSh/EZVaB
OFQ0Ga+caH+wjnTSgjSfdkofvgkmwMiYXbp8Kh3dwiksv7eQKD91FsO7j6as11oI/+9GyV3jNmaB
AP6B56i+AqzQKmPrvlGkoDdtMkBie5ga3lcC8Do7SONlZIlppI5y2Dl3lKoKEOy9zn+Qs8BGvelE
qxbc89SnLT1AkO+TTAoIA8e4lyMGtlZsp2lRcL2Nx20V8etTILICOXn+659tWR4zIdjWKqRD3q0h
5O09tyV00BkQfij7bAHdyhtloXa1t7gS6QkR5ixsSEZVESMOswvzCiU9zIskOx8Vj2fwKRYFRama
Gle5BI3ZAmi/VdkVAFDGRdCnDltx5pwSUVYf31sX9VX5RH2uVQbY9vMU+mUI3VK7W8eJa4CGbXEH
inxk6WVhgUVqmi4zrNSpMBqyCIqrsy63e3CCe9v7AosGHZsBOgd31Bt35C2Zvp5QMEwCEY9F2Lt1
SvvWN/PlC/vJHuwmOS3+wE+U23rhNgoh/yBlg5qVHaDCUuLTbWD4o5q+PnDRQCuLFCDR6MUNlJst
9HH5QXL09CWHLjYsCbM2i5Ww71hjn4FNlPYJBNSN5I21J0R9AOcXgmfR54CA+ofbUrofo+rqUAoA
rN46FBDLI/RqcLrP60NUE4z0wfWQEC3GXmJWhVuYUvXnBMcVi9UW69OhR1bX1wueuo8l6YzBPig6
+3bgRpl7UJzOMMxlhjkSQYl3d1guxQolQZiQN3rgo49SawDmSWs6VRrbS5VaXNToAr/XUEumXQH8
KIhN8zEZqZqTIRXzk8/FYmwLdXrAgm9X75+/XzrRBJWcwRVwXbY5+EP2AUxZP+37R2ZGGmND2jfj
jmkyNIPMNuu2gjAbIjq78B3eimY8e3ez+6jFMu4BkMIWB6O+jlTzDF2ukIgKKHG13E4CWGuaiJUq
EORD+C8U+g1duvjSBuqatIb9KSpnIEIUAZuba+VJY/hfXDO2OLtuDv5D9IyHTrLv9a9jNEYNgPfm
Ml4ayrvRGnNa59Zr2baPUxvQgUcQCPzobe3OXiPJcna4bjt739zhj1UE6nYXIAKLFjvwWddt9V+j
4mHwoE3wfsMOJ2FpnJqDyK777n85WqycsLgEaFtIyL2HCF3hPeQoJ9ig3IS2iXtVXYgf3bK4hrzQ
2rwT2MQ0uRXqbRlLtMACucdJ35OcaJClUEh5zxdXR6pJ9lYt8CiTyG9HntsXXcqJqjbFchqWgC0f
6pghnsB8TArOF4pUkPXt4GKRc/VKNt9OjQQEg6om7Yy7w4PFM4PsL5ZP4cCPyBUgqMXD5MRZHlfK
ThQyOLIYF+IIgvINk+CNc5HG/ipJLjTje7b7nJccHXvOK8DJZUF0cDmdxwMBsaAX5F/gE/i+Oj3+
extwvuYqWu2jgHhAtYDP+ULFnfHsnIDgqqyYe8PIpxAY7sa7aVUNXl6OEA9YE2k1NiGvl3p3ni9t
3IYW2Ft5qgPCs8Pe83DUD9BdFmPRYlZRUCy+YfSX2OEus8MkOLjuLzdw7jHWAAOsHaHeQzSwB/YV
OBY7/+QOutf7WS3cMUCabq157vzr8YqZfkDOTTMsPnnmp7SoMcTx7hgcv0ruDVTi8Tc3zPmGarpY
o7GmWkUcZyjDKAj94Po7m5mE8TM3W+qsYV2LxexrRrf7NaEr94hmKemkMrgu78axUvgIjoBL1W/r
L0WGpQu0/wUewHsy5nue4AYMMRqM+pkzF/s8grJ27wMZyz+YOuWdxbZkf+EXlnR4uQJPmiDV9Yh7
O59F8FSL1rBH/0IRBa7ucoYjayMRh4PtOdqK0UlTEC1YgZ866+gmLUjNEZBGA0XzSVpopEOHarvo
2w+f2fvQPOES5wkVOX25lEW6qKz/XkZp7mSC3n6Mf0CVsx6zraYtXQND9Dk/wET3MXliNkU2b12a
FFz01tGilZVUgM3nJwBtwW7d12DKJlFbFomBCCfvoPd/unu9DU5i+aQzkIfazWfC820ydx5YyOFa
n4kErHAHTUq2/xAJYUKzfqREvwyP/WvRO7d2TIFIcKPkajYywX/eE9n1wz95KLKxhGN8V+odKkVP
jX1jPng2dn7JLsU0x4y7CGdJlUqM2w/3dzRLFSzUTFerg+xq6ZwfrULJ1pIvoIt691IHBUTpF0Or
weQ6mnfTzwtBDe9W3XixwYxw9eNoKZNoXnnsFuLJBw1K+UsDAuQpWTFCCjd5DTfAh5vz8IwH7niK
rB1q3gRr6mFHlBuRTMESnikmYpdsuWK04N+7KzCDxNgAY5zsspCe+X0066q+K+VvAaC/DKPMCaJ8
Kwr57fGIiNw62ycroBK867RhRxc5eAL8ztq7RNcbJWMqIlFxBrX/fWXmxnUPRR4xF3BBaBXxHYjG
s1yx6cjCYOpq2Ki5iMvmHZcFXjW9KaMhnAr01Kz+tO1TRwr5k3T4KYYtn3MY0QG1GyD+qmZFg18r
G46uiFO2i2OCo0Ff9k2Hh1oyLjWg/cOSRvj70WqS5r1uraaFmY0SBHT7k8WA+wkKvkr/6y3cI3oG
X1V9tTd2r6O3V2iAc/BUU6QDKvxkMSwyupzOq6IFHwkH0uOllclG1G+iyonMH3KxQAEmYMukPTkO
H+J1D7NdJZnriCKedK+qGvNUYe8pw6z+iJBKw3e0GRWY/FAYWsZSUPhVpayn770Q/uPKfJJOa3FP
WgmmW5vxqGXBeAS0XH//vj+6ycND0mOVAYBEI4sSuhxt4Ll50IyO66U36aqR4uNxpCLtJ+vRc+wl
Unxz7rPV9jNjwd74v14/KH1Z6iwC/BKX14S9jXls7Fs5KDTRKtsoHJdGQ1t/BxDrWQiEaVc/TZbm
KtSix/gQqa1Eu1p7NJJpOcspl9asfDUYhgTdm+cEb38MYweyewbKoHZ95BZ8YX1hKC+gxOUnj4Lm
cwKeaqT4zg6B5mz5AQNoS+3sJvTKpxP4Xb+5Txemhhy1J7LTBKSPsNXrE15rDSWrrEAEiP328YF4
XSxEVwyaW4fUJUyca4bWCQi3yYaFz2NTfIP3b8MSf0/bj3EjcegcQMEf+EMRQ42uh0133FoCAbyW
au6Stz/VcPPEbZ6gOnU50vGf/yu8soXGIO0sLfniUQJXXXFhQyObvXBkCik1+DP1NBVUSVg4Acnw
RiFcUpkW0srpaAILFthz1jkkZdVh0BAvOZt/U+iuYEWISlCn2dKV5KlbiAiIEudMma4QWUaFrcAR
RRpcldbCeFmyyBvi1fh7Y8oQn9c6gpZ+Glf4fw25tEAc077IigWKDqpmBjEqr/EM1YEXad2EsAD+
d0XZIYQeYaIWERQXcj48sPDinrcQ6rycctrlpbkuFplFHYYLdQI5Zp/LWNu8hC+LmfaM/z/5NMGV
AWJFZxkPIpIXjOEhbiI4qJP376S1Nck1RsU70gTOMFq5fUtjqUmCJdKwO6bYoS01EGt7GXWNvne4
qLgbOZq5j+a9izOyvgmlB9TRZfc5UHhhCXFQBSKCOaM6Gd2LmWt6w0/zyQ0Ar2LCSrxRHrXUHGpz
OOM43aybJuYsO9xBBlX6a/Jwj+ijMsYeOnP4OToE9ZfATGotQT1WA3Pcjv8Zzzdjgo0D4FfE58Lm
OB7lUjh2r5iVjbGBU4ANfUqS44E1wiZLWJXztc4RU6WIbQHUGt3bl1bW13eMhB5oA6YDiogwRGfg
a44R3E5HVj22592ngGOCr3ZD+XYYvqIGoF8WWULpznpdHF6UKpPnIT02gAQkmfEcqe3O5oP7lqnv
yQSEgZPGmMKQAgTCA7YD7EYZpp8RKpthYSOMYdSaAoAnOTx4u8V7zyPPwkBbmzOPMlJgQJA9dYqi
CNA3PsShkWRsSVnMyY745L07Ge8r41FL4IrXu2KSHEPi/KJKblD2wmSH1kXjhR4gV0y1POpgohLV
PU38bHyzwH2Lbk8RykY0nEr9LOuq+JkAlsHWwjY4j8vWpYRRlqav7D+ZofWkOg8b3dqWoAJE6aUT
YJwWyqoXzZ98Ej1Y7YJzuZLl+0DUWIS9BOO5IwLEglGKo5tVIUnZNkvFfr01kHWxbF0D+kzdiYF0
mhRbJxrOmFINNDI6CA8n6rwvIBE+wqs3l9+0mbqd/IPlVaEKkEt7CosCh85V0mO6bRAgXCPcq83Z
UZdNNwkWUwBkfm9Ou0XUpFNQPBj85SChYSFck3pH4AMvdPwgWq5oWrq386U9VKMfOQDxJgJUe7yN
YnP+Mk1gi+SseEPR+JBXJJ+AgQ69q7RMDDRCZZmWV7OyIqXWwgf5YoGbxIwFj/Pzs6/SFc92RN7c
7m/rcUBFGm5Boyml8f7Sken9hLhmClz24jMBtSbs6bsQd5GoicSsqHk9WWyjucM7lfCUrr7bSO5T
jTJAhINB+O0Q8CtyS2n2nHS41GMdLtFBiCIr0KYRlCKTmHTKzaNNTVaXZYxEtxKbBGQqRfUP7OMe
Ye831E+SheoabVtGj3/piRmWT0FxRThFn9113Z8WFh97gF6keNYqiXhLRtOwWk9s4zGMxfx2hDrK
OaotdaGTjXjKiU8uIAEAIIzmznR+CjVIamOnWP+KL7WlgV1zeqeaLWgMpOJlC0lw1vbu0ve3UTsZ
5g47Fc3Kl5G/N5jmpueuP7mcSqgZdH3RdMiPicFSgLeyynqmwXj3hiZCzQvksd0BgQf7owFAzYW2
EcDAeHZ0/oRv0ZlEdScTRYJAArUUYOR8TcImTaCLjx7oDkeP0uiJ1vi9AYkdu8omE8goTY9J1jmd
WdpyXnUAs37szum7j6n4nADJ4aEnpEh7Oi1fpNZV5DpZDQS5n9rSRDiu54gthRCR/a3j1ytRQdd5
T1xuZx9itECnpdlP5FkbELbBKwlsIAXd8/NUcFBMzx2nkL6jAqRNXG+aD+Az8n5Fw4a7a8MyVKwk
E9JUMHPp1vR0GZjHCrMpmW2L31ZsNNNK5Fbl0SfVRjoXf4Act4hX4RGAK03LKjkaygHZXG+K5jqX
mhgRL0bEPF/0AKFX8RtgumqAXVkGLudL6l5lMgDyNRSXAaObeYc7jfaCm+wgleGPDqAsJOuojScw
HV7h6wwjizBHYrQeKrari3u+M7el3hKWTetHFcQNsegEuweHvqvokkaE+PlYicvvx3dwptTgLmL7
0bvC05ak/NzVcqREeHVGJw4HBGMyM5co+iRcNG1b1z0RLvdepW93eYIHFyNWEvHkkM49VJB5Jr1K
DFa0y2Fwn96sXbZ6WjSGSAZ7Fffmjd84eKAJFVc4F4L8moi0K/kUJFdPvB3rlb27T1vUD9R6jfLT
Uqx0IC7alm6rMflWtpB+3SFWe7CH0HcOdhQcxXWieJQTJ/7z/mvxohADgZrlN8IgUyKpFns47K92
aQg+MRGWRRGoB4BzC97WIOHeFS1BACJlKjNYYWy4iXn1+ZRRG0v4UmKd+xMAuHFtkGYZmn5OH/CI
AVFtivE4BW83ch2N3msIR3schdlmh9eYChySoM7MORrD/Sr1aWIp1ZVCXFBDg5omiI3emBkOHD8X
B2fybnZPxHy3JWZ+NVaenSlaxXBBz3XqjjNZHE3blLxz++PZcxnsq5xPZT+70lI02zOl+VQtcJ1E
nz+GAXDPnWsL7JtSRidD76nO5uiS39JsyERoW5dEOTdhj2ozvOMZuhvNJfFBwGAdPR9CK3Y689Vu
05W+mrNdVClb/zo3qe+DDx1mu+k/LpKHIFrX6ixjXZnXc21V97DlFT/fidP5xctw6st1WgozV6Vc
/z7lTXnW4U9nHlp6Wm1LdujSdBnBBcWDIXzBEKXHVcV8wNDyEVTP1u8WGUtfviE6j4J1DD6IBgIO
PrCGlAwXU6JVH3NxKWgrLeF8PN+LXrCxZE1MoNk2iFnhMybst3rJsRo0fK0Nd7fIsQwJ1bUpbN3Z
7AzTp4A+D2nzWnxF40KJMxf/VkipY/CASdUc1kCqgTaW6JAJETSWJmEwAFoHxKic1rviGUZKZ6sb
v5gWqIgSYQRQd0K/IlZyJXEdA2rmUx1ypsma5I3EFdb0qNW8E5yvnQzpRBqiFGV4WfmjFhWH/Enu
8XC8idg0kKv5EMkwZtDx5LmfeHPxujceptoB10EsFyu3VS5xmultKVoK7mudWrtyaRO6fZUUoUOu
/XeF73RXAxiJgztWYgMIWaBxboNP8aQJqNbsJbft2j8RXzJDgGk8Wak+pYoVGA+Y2kgi+Ip8em+C
3KpRKgtH5DLwJStacE/7yj8GoSRkhvoXBJ0XH+y+OmwkBg1LwFGDJXQkPnMMJyydJRINxA9Q1aZD
Ordp+9YYQb6C8PBX7ZhmyeSXnnPLxIkzKGXTnkvXHn3cxFoyR089z1296n36Mb/hy8OM5Q47B/he
ZF2lGpfn6AVps4zTmd7tQVPXq3Bycs0iDBtF8ap3NSX38Zg1HsKwUXq3LnTL0TNgQ+F3GgHk/czv
jSmk2VY33CfahtPSStQSdiFa4nPqyMITkyLTVBwrxsLDc+aUG1GrcbpikrAURCb0cSmWGi+JPM+w
WLCW9FBeY0hrLE7UVqSIEAkrPCiaVZSvToHg/R/4CJWg/j176aTItkGSTzfX5z/UjhUggxRqdl6Y
eZN7SVmbJF1Z6Vs3D1m4QJhgkH6HxJNauJc5AyeP4EcurwnDgiIqqTuTKEFCq3uVv8s3bJeEpox1
5biSQCFC8/z00tivFTHXSjkcnKhVbFwzGve0zTkRUDRUf1gFe2HV5yq6UIRN+UsgfQCJEXFhAxiX
j6puMGuCKPCal+IREHE4dEcV1OgM/eXYMAiKUq+k6lAn+Skp2IA6/RGrvVCmq0ExK7TmjFYjDIpq
TT8ezLq6JP8qtamk2Iuxry1Tm4z3OGbDKc6Hm7NzAx4UHHiQsF6U9LBCs4aK+SFKGdyRFZOFk8j1
HXl0rkpS+OZf1eEPkjbYfLUTc9z1fQ4kA4tf9zLUeLMQXjD8FkPF5kuI2TQQNueaxQYRahYkXoFy
D3wwgkwcLu0YpJmCQPB5YXBC5Hb/T9ANIrm/cL+zpNuiQ/JC7ZwWHvT9yYCZlAv2+iGwVuNtVwNd
wWysE8Gok3s97UzsTl7ucX+ou9zi/vtSOntJOGiUhqIifFS2ggArT9tOtpE9KpokQhRLJqKxyvws
G+ENgIQaeKo4shzqKgE4FIAsGiDFjY/3B42eHCqom2YTugsOPfQrGcO1YSAnq2zfummHeGUl6uMO
m1/zvMkmuZ7yieWv9qGZKcXzUmNfBumhzciMQT91PpfKVWVAsLziS5fSp1/A++862eIVpwd/BnSw
uiEX0mZTGsgiXiDQgOVkOMj2gdl6s01tPC13BnFPMxMwInm4jClNRm7eq8Hy0J41a0xo0RSWe004
iwTssy+yGfJAJ1VnvhXc+lrswpfcIa83Z/orP+nU1LbJNepyGwqjAhQKXkWtgRdOTsPGPfyhLEAT
gepLqQZPnIO/vLxkd7Uc1xvOQw10OrMCfD///nQeWDG2tWKi9dOZ79IjEIBwki21Gy3A+/9V9OLP
w3vCvC4no24dhmmlhCKLmHq4m3P+opd0v/nDOW38FxB+VcF5OSHSHSymg3F24Ab6Rcu+aSkwaN4w
hRCiFqT/KC4i0u/JTjC5vCjNqMDb5XuaUhzDcEKR0PAlV/8D9Lpn2LPUbGbyGTyeXot95QItIFAN
YIywULMdAH1wEX1AviZyzAp+NJNZNv475pBSEVxipFlekXyduMX8vf3QX6owXbXr3GRycv2ddDjd
WwwrCbTPJ1WNIM8wawk1ehZbAtwqP8y2YjqIYV6b89JvAwAIH17/qT+8btulgRaCPlq7vxnYgqVh
mjcpIcUzCUP8b0qDWQsDM16fuDI3hcpcMiVZiDkMX8h31PB4eoUo8s9tEQWe7D1dVGja7FgC6EUd
PmOQ/tTsS0ImSM/egL104/hdV+wwC2G1R4uX8fyC1fXcrgQ+CqObG7HADSjqnrcmdWz0YNnhj8Nf
/q224b73jbwlndlRx65Plr63EuSg1qeseWgXIUsQEBxUBeBMLWRFjG44fO9ILu+qrJKrC89SzHPH
48bqaI9mBvdwmHk7hsjmjaF6KNk/ZZW8WbMRoEYNMnVIAhb3TdMqHmDr4QWKXnVksRQrRIwyvHt+
fisASrnUMw+4O3YID6S9q2xJaqDkHJD46FprQn8OAAuMWngn4QA6dZpZgRgdza5CEVExpR6Gsex5
eMCKt+2AOOeYeXzjbVr+QP5iRXWWIGsY5q7WIEPKa68L5MDwYXOslnaE58JV7Y6DyYNmSH7UdCVD
a8KvxvPs9gqHIBOScz1bBEkAMXYcvKytOrDO3TzVsqzcnZVqWEekpCXJ4epbBe9HMwQ2fBQaG4pR
fP39S87G82CWLZMtZvl+X87DMKVykGHx5yN9gTCIsoNVhqSbD71ESRP1cKlt4EtnvExq/EeD/mog
hb5E/3RoUYNwFbF9px9bPegLBEfxSD11nFoc48lRwmqpP7YBNEHhO0OmPHO87iTNvOXKFHb+3Wwc
049RU33Se9EByXNyETkTm1f3vo6LszgxyOHpkocAPEu17W2+asN6rz0SVBaFpWtk7BZz/QdfypV9
saUB3QAzmWype5utzShIVHpnSxOEa4gAEKHLcXc0mHRdLi12mg63dJoPOYDAZVY/K51Yz5ehWN21
EaQQwLD8H7Ss5f+GYvPXqkuQKhiuohvzLRlln717G6FsSkpEm33Wj7SZlpAkWH5zXEI++R19+R9l
ebTFnlNFXOQ39qlZI5MuJzYHWhFZUKNVwC2PiD+CDGSMvudOY7B87aqmKi5WC/+lEuN73lifKP2c
n/M7R0PxVANAOjTOylyx1L1b/68bcOw6CL0GHuSQ0PZjk5I+kTl1GIxkDjdjx+cPDUZjjxvXiW0g
D0B/R8i45FYsmuZI8Z6003KBg8/NWsV4kgw2AbFdx7oY4/TzH4Pkray1AvxGvfRFCqcHGSfsYNYx
E/LOjG2baC/spNrn1Gdo/Aa+igr4e02gFEGg6ZeYza2fb4KmlOY9S3XAbUupTPz9obf8kjPvuUPr
7WH3Y7VEEql1unF51n1zFixBel5SAkbqUx9SYycM+SQLDt0hderK26zw+3tKdosmVLcru//3pjXj
H339K3sE9SQhoz8xOLxQrIb9lftBZZDJEDykD/vbdi0GrhaT/23ta0QYZaPjjjvixeL6hF4O+Ror
JT9croUqN/R3VWP76cESsCbg1dVPXrfZyBrKWmmi8fIotF14PLGiuos4ZObuOZTQqecifetnamAe
IxOUcFzDtNw32MXlYeFj6EkJXT1Bo9mD0n8y6lg2s6+nLI/NzYl0dwawEeI6aJDR6UYY14C91UB7
8z+VDhMJAGCIjfxvwvBk/xXMBWv9vVMoked8MspvE6jp3UEEJD5Zk+82r+Qyj953CWkmyzWgoNrL
1+VceXEA3M435rM7xbAsnRXZuD1WTFcoiGmi7PWyKAtnws/DrlMOLsOlr7SH1wyTQwMAPf1C9h0M
Q/o5ujKXxxryFmWFLE3qRrNRHAc4PWsuyObE4zX0StfUcyS/vWfED/zCJG1nE02mXEmAED1poqt4
ZHJp5tANbd8bILNujtbjzt3sTjw6HxRZ0jdRzTEA2nNq7JCQqegXiUMRrbIpIqEAgw4D0edcUSSw
/B0fDhA20GJmKAttSPhLQm3LIYdgkvZn+yZ+Vv0gK4auUalKkvqLYYuMUGnOfNf4prLYIcPx3qhH
owqwW422iylvv0SjXczoqLNwwsJhhD/rGDRXdeIHT4a8C/bT1wS7TzbjGzt1zvIUs0rN0evIvRBx
C37nD2HlRxLATMuxnI+MPK+dcwfOvOn5tAhUl4lLHmuW/ntvkiKvOizjty2PloaBZVm3fXqjBu1V
fEaepjC5WxyeCYoluGIJB0rSfBIPkmySSfMqvKc9LzudM2/m9O2K9kKtl4uNpSIuX3UGFVrDrq4I
k8IhRfzEQxLhxvSj9gc9DGOJ9VAamfjBfa4Scz+WkpQ/7v2ZlM+ZJrwfgLNveh42KSKFdEUXmCTN
l6B08FkWU2XT7Hf/hHUfz5DEvaWp/bM/PMyKybjfUjT1c16wGu6oQEi1h7ckTC+Jsw+7PXB/ghIv
RhLTuWte6XHzt8iQcsacxG1kEgqWv+2M88IswH4SikpKSX78We+5bB0pjEfqk41dR20NS8Za1THw
Fhg86aeCQK+8adlc4m7KH4aryOokyrSfhozLS5xV2EmI2jWGgjpP77ISz3WHO0P9z+0XhSKLntb3
AzwZR4/qixDCw/EFzm4k+0+w8fU3b0bDLF87Rf3Veb6M62b67SJoKGd1kpHaWdPxu5h3/jzYkoTu
X1++4c1ZB8ToMu7BahqG8vV+8DKI9ccnga3FsOUUYsnPtdBDM4BdkqDOfDm0nwDr9BK9oK5YAajw
r32niQnnLmPNNb+GiDZBDfmegmGwZRuTdBl8WZyzE2dbsa682jJSn/PaQzlQNgaoxGA95lP5ijhe
ibw+0fOdljru3ExDwTI6HUoEDM+/OMmW4lvvjyVB9cjGoP2pnHVidmQZuizS2FIFnRcdpoaYZdLT
4B2kmqUmOlOqCgVld0g92/qPONA+sktSczHNG2xoGeKUd7REQXoI+1+0qQ5p3KliS/V7baf0sjCg
6BcFHPyi5coFnDEErgw81uj4F3MnH9xECHidMqsQLgV/DFoW5JTgVuk6JQkC/MUlYQhfBst3JxSa
NUXHYSUrJM2vCNr6KUKLIeHoXwDCX0zL0N+hJp+j8AdcDZYQjKGjFsmGFBmnYLR07ueKq910PoWv
pDSYx/+tvLfzLt/4itcw4P3AmbGWfAj7yWZW2GEDvo6CTEy52zpyBg7CTkjJHG3OqyzxD72ReKFb
fh/9NoECTzM++sOZDNl8Vv3hcUsrWHiZ8z+6NRmV2O8EP3D7IeISHY3IbBOQtC3VyJh7wd2YvReR
skrats1hgaYSYed6tfHkmqxq6NKWWWhKw1hekVzuqJOMcwlHg26MpH897DXaLS5gYX2cwsIEYagp
5IPlFrJ88VgSEkMfMqgkaptJh2KfzsZUWLdoY1reA2H0yLWEAeoQbMyP9uLpXewHS5YcwkGxxJwe
Hw+3DpKG7OaQx2/I825ASvhwj2hh0pOYon4zN9OTEQxn6Tk9JL9C0fU4Q5pxL9C1lDn/Ir3QiXSI
R9n7XJhjmwXzTVFBXoRMC9LWhUl94MgyDyWsCIKmU3QR/8jODAtBy69wGaD/c6pGnUBdmRkFa4yn
s3js3a7mr0/3ocT0aXYvmeD/OoWfx6qRPy95bz20D8bDwdTVJH9sp7ycmf7KjZ21WsGwP4Jz10RX
o7QeVt8eCpsp+DrQ/5TD1IWJQ79HMPi/jziDWxDvFUKbbtloh6Z9jfK2/gRRo3XMuWDIxmlvIHET
0NG1yFMirGv8UP2bYpIPuNej+gu05zFWs/2u3s09uhCF12yLHDqRyOjkr6Cy9cp35kWcCgcwCpfT
nEmcjQD+3kmmQvY3ImJdwYrc0HhyMh+1OrSyMVJTELz7C954vCulL97YMIyIy1qmKg92OXmEAxdn
1J3cJtpnBjt2nmAheOiSxCfGO05iZ1FBiaOENrRwBXbo+9QL4sUAd1e36Sm/TXSc1qQtPucOh8QY
WvIz/1JvmydGaNLf7Wo4Lhb+UVlm0qbjrCK6tDfOSTq7FC3HK98HwKe5tARFCCwfOtLF4opdV6X3
FesxnnR1D3SaP9+Wk+N4mJLmcPVwxvAziO2+QgxaxabE58ihCiqCCvhw5hUT0QlDs0WIyJPBWXUm
hBF4IBcxmSYMPnq+3kSaT1KdJS2rIHnwi9aKHU9gLV3QOOdiqcWlfeEo/GGzoxML21qD+EkjpSAY
A+nu3/ruJ28kE+8AJztgxLL2owbdx9DkyvX27KBMcOOqgUqpUw+H1La3O51tz9CnBUi2XTWUAdNo
iqJcgBw52rktSa2v1naZgRlvk8bLcWtYZcr9WE5q6xC3u6/sTOsTy6HH9mgo+XQQGxsXqfT/yKWq
AHcBn9WdhRiAreGWnGf2I0ANckLPoslKfZ9GTCtC9UoZ2FaL3kPIAdkNeOt2I8lknJIgXiCEjnsk
L4CEK8XKKdUrStF0abuQeFO4VCIImTBXHgD/GtfkdJqNm4yhGhlWdrRkzi9KApq+1bBaIuocn6Z2
QEwjbOhFQTY6svJuAgAYFWorJxRsC68Xb42RPZQWkrqus/PnshKyhgU6sxWfMtBt6b59m4Va2cfb
VJSunP2c2QE56k7geB4oQeFrt7lyS7h+fg8uErpI36xsDZScZDzDAYbju8yzWYYp8gMyWYMW8Aa1
dkU73aNop3r5yIc140c6nSeCQuOMMCt9LT5iB2YVPna4TdVp/W0bydmvsxuCnltETbVoXTCkxfVB
JreQbZ/o9rr31/SD51dPBs79TQd8I3mFGnRK5EpAWYABphER0M8T0GisvoAenl8e5NvzQmPHTrlL
5f8Rqyqb+DbttXUpRKGvEjzyfuI2UUtpWpX5HWndKkIT5km2YwJmYGyWoqG4z7z3NncgX+LPPXp9
vd5uuNgfoubTgM0fnJKELrgA8GNYJjc4MXMJUZkrgTrfI37e76zOOKL9CJmqdaZMj2ZXWXiRaTNQ
Lp81OzHL38P0geqGo7X9oC6MSgGLXVmeaV7GeVUzjT+hWpcC+1E6NXomar+uK6FrVjP8+7aWGY3g
h/jOtBWRW95wadEe7RyJf0En08CBMYMWZtTVy07WKrzd0T7UzJoUUfLmDaCw/BxCeZ+8tAsanJ/h
J/YRkKpAXqu1K1Hp76rOYUzj0FjY5nXM+MURg4+Xh+CdZT4bJOlUV0PMgSE34cHegNUh4Lslqkl1
UlkFoCaTPcCX6EQhHU0TL0ozRFuUSUgYPczZCi/Py00+V54dNh+jF4NqRN4HY3kJkG08ONv+uIeb
kXxcgKUqH417ZofOGNE+0f+B/1DDbSvJAcT9wrg0YuDqyx7bBU67wVDdjDSkAW4xvLnALy0gQYw/
Hma1NBEbsJNMRhZoChWmBcNtYpuAN/9b/Wl1PffrVsZQT85BARrkz3eCrQVFUJwfEiWV/wVyMtT1
r+PK2iGrV2JppZfA3pkj7VkVnBm/bu2ND3Tjo5nUuOe/j4rCcmTEe9/bleEtkzbymCLEUNERkTiw
tBvN93KNxlZ0z2gE92M3R3JytH+76wWhh0aR3PqxR5jTOBkqTeDk0nQCgDCX7faUUWm6pLzM2mGS
cGNt2RTFwPirlHZKZY9n8b4lLg8yGB+dowdzeX4le6XuREtMV+klBTNxySv802lz1MKaDQiKIqYW
2IPDUT1IOlt9hRQ/Ws5+I2CTsDqMLNiWdX114ASSaEu6pq/jKdrqakf6c+7kWKVjoAaMRy7ZRvyY
v1Vumwp5Pac9ZBADCBDc2S1CTQulKtZp1wo9R9LBHCmg/lu6iK3e9iLpyFPMT+ValQJd5Qo1/3AO
6e/GX79S4NNvvzmxiApcuEtZ1xOn/DIWhPtQPjeigATKd8NqL3Xz8dW1NTQoG6ElbqUVHsgDdmNz
k1ICFUUoZM7O1mDvv9kjy1/Mn7gqHERW1wbqxY22iL7FvM2Kzjv38uXWjYVpLysM2mfrCkZGARmD
9kv3mQMyHSIaE6TaWNHru3A6nxFyE9TLvNTOll74U3AncpnaD9IVa/H2wNrEHGH+UimTgek1xNwP
A7cpIvwOyI51D5ENSvzSfIs2rjo4+EYMec9cmWeM+yDcAgC9qVCVi5mSlRnC3QvdQTyrWMoP5cDf
/jrWqg8IlZRh642SzmBCU++MJXh7f31qExt/YcfvRFM0ErEgzMfJnvYqGIFbZGG2MMNouMzAB9Xx
JSnWm+D1mPtOt1XnTmCgU5J6TdkMmVXzO5JH2CDF+UNEnoqQPF97e1qT7x37KtEwC+uwEwvMW6tJ
OPPbB+ZNUMC3C/BIYAUvnuNpE23kzpDl7v8nxVMBixVvm+V/RQeqPug0aHPrtNe+1wToafjAHhYG
TtOs4+cYkPipbYCQsoflwj6LhCngnCCWf597U/EYI8eic6iP5Qe/RhV7gYpY9/U+cYjyWnca0Qxg
jV9dT1yTGKKwReNF0RbKJ27geoaW/25gvVo3Vw8HC350j2qumHpjRieHlNdIHkh59NGNSUuQtCZB
oFaWsMt+MKgkooMlLEvzeHPvpUm1BnQkeulDSSMnAomrCLpz5XYXRz7yoFDcePLnY0m+NprmwA1X
aFEKH/6EU1tmPXNN2a2IcmhM1zb4e+vUlXShZPBGCF/U6KlfkZ2rDULLzbfu/PhnsqyovcpkEN2s
ZcWMMl+9yr+MCO2Tyivw3KbZ8y/OmsnuT7x218ibVYiGcsjYVgAqna4Fx0oDc9OqRzPUqfH65zsQ
vHmwdKn6x2pq4Ej/UZyWVTJ2t97HtBqo/CHw7N+8ahUJ6xnpxp2YRHEUu7uydu3BcqAL1J+jW6+U
RMiQ6fmU7VBL2/I14YZDK8CgVygwiMDqBtT2JQ4YFArRF8EQMKmKCgAoCSD8Z0vi0VmIE9Hj7blu
bzby/KpbVMfvBSoDMsTn5h5ge5TpUyj5gjvpANgKouB7uRZfzHldXr9+DIH3appcTCIneDPiGX2/
VwG4RdR0R31aHFbzEXX8FBE1Y+7hGLkScxSejpDHA9sDcxNYwRnjlDUBAI7x3SKsB+W2wJp1VZnl
ksHldD7UKpv96oKT5BlPdAlGsTAUqwj7r7z8AnuD9sfgiPRNjI+c8XMoPAVEEm1H8kY5VowXf9eR
udSsqQrlj3x5+9fGJBTMEtUTLue38EHKm7APktPzUMt0HqLjJZMa3CV46x2GcEKMa1YWqbyUWX0F
K2W/jMD4s5OL1Siq2ZWvxOyTLsSCSruNu3MqtQkEter6Ts/HtUsR1VRVaGxrRJiOfdfPUWAYglS4
z7scsHdkGkrdeg1Oo80b1bWz6bbELc4yiOX9K2Ata6IFcKdt8ZcQDcRTIuH9MZ8H7yp1ibJXxate
c/YQSjmfh8AW387/Y75MRQIJXLA5IbxP37Fecp4ataQiXpdEIl8UcIRezqnSXLeAx5bRq77AYffs
KiUEgmJnFtRJ44j7ucRJpQ4s2lgszdQEZohJiDJhhAEoekTsl074plJpzt57Udpg8pEiHJn9fr9K
tnnH5BU3o8Al0OlFBOQjUYw47+6IXsIXKzLArGdnKXXY3IerNXfGGKtjzqzcE1PUWGrIdbE+dIir
3ocJaHJx7tuO4+bYfqbcxAd6Wa5E73CUJnIUBceHDFXIYV6WfXIpAlse08Mdrg7Zdq9novUb/8IH
I2dw1PyfJVcWgIkmlJ+fWofGFXiN7RYzFhMFY0/9O9e0/et7jbNeP6ZP6ntuCK1vSkdlqt8H8tB/
u3yyKqiZa1eWX6yiuobzcc2xmIJ+AjAwqlD+CajHwpXIshYEBcgxZXI/K79O8+3JN07lXzEpy2mH
MlxycARIrerxZpf9lAhEsbzxqhXsvAjUdD1ef4rsbpLMoyChTBGZZblJvDyTjpB6w66Zn+jShfPl
z5aTbjsJK2xOV2TO6IVUZAaW0lU0HumqQPv23wwqvww2SM7kdTwSaQk9iU9DMNDQWDY0t+PR4sqD
fEMdKPY/wLAXT5mWic7gQf3EQz9LVycYj4nK3exLeyF/GEsWUVVaFrQMZJpY/LcJlu2QfhrrImCm
k+gLgy9GZSKn37Bpp+5B4wg5Fqk/mzYshcjQEdZ5ZLN/dL2iQuxOxb0FYPVmDrGZ9mFnpLqQ8v0H
AlshjFp7M6OBWggF1Flhk7vMTGkR+us/yp43pAfPLsAIWLy4X1mFlr/LMLiWYKbyyyrHIJtOWySi
/BbApjUvrZEou0jpQ0CRYLjDAdQRaip6DFs3rjV67jdiO/KDgX0nwNtlP5if/Jphjlm02dEHzFEd
VRxpq5XZzJ9yEbbsZrEUhhU77e58jy0nW+fm7KNLrIRJp0Zxa1EW5iEpws22M2M9hgz5rShr3lLN
geVyXgHgPFZKHphzmv0eKHv5OOmHAx08J3gF5Aw+1Lr25MnQEUhH1PKzAd+SO2K4VWjX1DG63vWG
Pn+bKG2sy9P3IkArMsSzljOCHS3a8mETYTUtUkxrM9o9/3wlPhi+WdwrMlU5rMWJpt0BZLqOHWMw
TgbqXTgXpw5M9ZvSr0NN4RW78EcRJTq2YXY3JxXP4lZTwJK8lFwn/mGsVJ5q2drt8SaQgn1Og18u
h7dqI+p4ACg/2qxHcWD+BYNA+vKHjZO1ZKygURGeN8t/XFGfsRbejFsHkQ9RjxRwISN9fJovFvIr
9jXin/dNt1PBuF4Xm3aEgK7nh5SVlXNxsc+mvU8tKMYlz0upOQVA/DEccgMtyW5kaTzakruxz9y5
JD97//kgx2k4HGEb6FuJHSO27+jEfr5Q4uZbJgtoZvkqaE0oikCADjQyYSOk2q8PNnnefoos1fow
C5bvQsQ9Qw0OGsjGo06YmvtyyEZgGEJVNLaoQGtjp/AWnrsKM91JRykltffdSgaKimq0bxX94sgX
Zc9xhyLcdEbtsYXQEtBCzI6qxNtlUZtFPSEktDnZacqrZyr8GqK2eNmDN/DWuxmNA4B9zJ578BSP
gaVoVf9uB+D3FpdOJN+sBsaa4U3MpI0OYjpuh99Ezy4m77kSWB1pi342qPv5hVTMmvMd5YN+K9NM
6EYMDpaO8kjKdjM47PFHwtimA/PlGL7bAm+PgfosFBy2UMR6Eq8YU7lc0i3W7bguXCpLiFkJgi90
We11lCf2FsUuMcxoOa9hr5lsFzi4sh/k8g6JTh/nPTMr8VbflElqNbaRt6Ca+SXpUCi6Y0Uw5Mug
tXV5ddQuuKuHxVq+OUtL8UW0GmvqkzprU9GyU9jXEPgKCSJyxIhMcPvSvqhFXBDhlbBgxs2Ay1Fa
C2C/X7Cv/ax9/Oy0KQ5/sYePyElY+HG4jdPtJtHnt/Jshhsio7Vwuy2M4uCpArsFWgk+e+mJzvjr
igAAm96f3PPYXXKYrdc9Z81rKnE0eTyeCWBFJeLdjIZQglq19VWzLqXrJnBxhjuBx0lfZDuoveqj
07gOkvQFj/rYImUhM6/WNrdMGUARu87Kf4fNuv4ZVHP86ljZV/VnG5b6A6dd/N98FAQScjTPYvjS
lwwft5QVLiXTBmCc/6u2cYcYwk8JhG+eRPHhSfr19L+KCXA+KIf2R2NVYEi8hwewu4aIwk9msAeg
o8l/1qDPsHMs1ZcD9HNtbkJVgq3PJtnA4Yk+k5K4vtSfULV3SVsKBitDkKwsgrZ7UXxasYNo+8fK
ozSzwNwe93wh8pP1CcUYrVMX/mrygBJvLLGFG9f6ZX0HSpe/EVXYAeNJ6bR+/A+5Xr1VQUI8rD+H
0O6ZHIXAuWevQxGPMk5l6LU95VtOuf16f1HyHs3XK6Kl5ke0tIPHFO6kkdf5IHAiKFnOohclhY0x
2pgtORIbJZtPq1R8OE4oMv7oNszLr3RlmtWI+pVQ4A8zeQoFgvJqUcsNorfirirocJOlSrArWSFZ
TUBJ4hCYAcPykzwI5FG3x4fq2hqVyH7Z425zK3pJwMlaH096T5GGyOAKppv+n6yDDqbjZDm0ufwB
SseIVw86a9HMcLTSIhxIZgXt0HARg3E5xHi0iteYPHuq6V0N/w8bb4eFRG/GIdgFjEl6hT+Zc0TM
FZ94XUi4AeHGL8edJp4DOaTgyBZloI4mcjUZINWi0m6PxjJOywQVfT2EChi7S1bc5gdREp8ls4qL
DSd2Ar15hbFSrtcDWWN7rkfGeDZgYc3xsY1cMV5hyvLqfqk7/CxVyHHkylaT5CYAUr4WRsyf/hlT
+BsLRGR7RGWpnrrNg2/TBA35He9xwPvv4IMUoiM0OklHbwiLhybByNj89e72qW0mhZMRx2xHJGNI
7qvpPna7Ymx2y6ZlSNsXZd/Pbrni7vKJUaSU77UOje1du0QIC3fOQY072sr7RwRT60GBqu0OfKOY
lRs22WadPbCa68zzPutqRnhnvXSVaYLr+wKDCvRXW6CtE8+UWQpINmMhJl/bXlGrbqJT5vtPqobT
ozF2QgWDs315W29JNF+13PchQqKnp9tUP+CBYLrnjQ5msT76P2corzFMgN6sNoep3pPFMC0dsPEL
1in0iqlaGM6pMALh5Wzzs/j/HmhI61duQFgRP8k1ovZmsseLUchvS8KCNN1FVAtIAIQnfQJ+eZ2/
sjJFBHBWILzfbrZGJolu4eDeIE6QJrGwwfRPE7s5p7dPwZrIaGXz3ZKek37NnOedQtF9rFnuO5Ju
IIgvqs6f7DVa/A+GoHa5idEGQxwaWrUGK8xSGjTpd3unh1PD6e7f4oowEnZdwbnf8LmDmrODXWPL
MdyPsnetYlR0Wb/qvJmIfxro8Fd0+FY1M6U79zjhJ24nNgjpzKWF61uEIsPir3PSIQKE3nmvQYB3
HBeuVHAAWathduCZFmX2+dQUy0WNIRWB2Y6wXNy6au1Tr/n8p+R7eSoBneUh9Ho4srhV3Ptcbbjs
hMS7KqJscR5bl0VnUarYyNTBWqkK5FwlY3Ou394vUKHlJqUNfKW8uiym99UJ+i1oYaMGEs+12uy2
NrS0CtW/N5kE7D2ARcw4TRGeOwXTZBYYq3+ekUvVJBHD0lXOlRBXRA9vqj+cpkH5XQxvPPUB2H7t
f12Bg+iM2hWYlR3GRelo6cbdNlRpqubb4j47swYt9teuxEK+bVFpOcxOxr5CAGJbbB3YrcF+UNku
13NIfm2CLxbx2Q1W2osdDUyn+fyMczm2O84trPjBrr4e03VoCBMilDsM8cmQCcMcvev69T0c6QPI
UH1W1YKdl9C3IEU65r5t2aMXgFXVarqmKoDpMSk6vfPKcDWOoq2kVg9QKmwkfi13dgwGTGB7bnmZ
fKbUA6mioHWGwoTx9VyLPkamOzUocGLnFkxraLxxiC45D/f0JXvScloIB2LF/aXMWcOQ1vtTbLSa
uf9nCCg5JipOR6/mFxU6DQ7x/TsgCwGHFStg+79ZKDxApTDEcWMo/wm6dd1eXOtSt1gQ7cm46Tgk
ZgnxU+IymrwbtOxtoKYNElHSNDw4tfztND5lppYQ95PlioyGxjEANL5rNj3AOvn1wfQ6zJpkAWRv
RFizqVkB2/XmUCdTg9OBDF8HL9L7y8IvVuSLa5hEcZzsGLb5mN5FU/NF6azJOiIHbOJ/3q5uqqSz
FeUpApgAN3o9IBfcIwY5fe5e1bkYk0/SPYsdBnanl5oSe/rD1ljswwRgGvvu/KyWU4aRzwmTLiIO
cqMsMpzWVxNqeT+nwBrn5hGNJvkoHRye/JgbwMZn6zIODVf705eSa8UMqd+vxIAmpb5cn6teNxf0
UXLqMkU29adQ9+rzLHCi8WzJxKcXRT/fEfGpxesBiVdp8u8gvN0ZnhSpIams4413sTLpc2Cp7TcJ
hezMUmAFJkixd/LkBzBI81pXnrt+pCe+iFImX8b45KtlbUL+daYRM4E+9Z0P5EgAnQ/yMvLUPuT+
VcDp2dnBtUd4dVVWmRhE3t7TUU0vy667OH9U57uskL4uenBf0pt5rQThZlmLZYwrqWAE0M+bMcv/
+9lMB0e4zTOdt0YuvJUVnDAk4SChlnNuDryprzJthK/J5TWf7KGsjfjHluJCTzFumPyhLhryL0JA
OEWCjm/XWw7Ft6XKPrwjE4rxUxKwro+NJoKY6IIWZbL8+KaFgMsqfvwXl8un+8UGM3MWEI7/1RRA
oweorOTvyW/0ZP0/A7SK5mDWV6+19CQuK2v00g3rusQlDqZCZPWOTbCA+/LXBva4kW7V6OAdrtwQ
Ej6L1TcYzbU+DuRMK1lfq23FL41cAKSn6szn9rsVC4NCl0EKlIRfiwG3gdLFk1v+4oAl473JCEk2
/jfwpz8YSLcYTOyWOfkrHpug2uJ+NrWvu0segif3IpfVzlzdUL6vVPGh0yYtH5wbzKWrIHqvpEcx
nBz+aHVxMGKFLWjQNvmw3m/eovOJ0jeeFczdOvH7h4JZEJ8ODmMZ0ydNteHzAg85jS6k9HwQ+o78
HOKhpYU5Vv0gkoFNSs3Kh+71DKeOiH+T+ck+UUYaJRfKEFbsnSw1yAN9L4cSt+jbyr/GrRR8T6LK
xL8W97DRIS5cf9sRfU8ktFQEfSeTmEgO9muqS/Ww+nl+qZ8TsAjv1p/d0+8Xyl+VhwFkGIRZD9L0
cYv35XcVC7kWrGKLAHcoHBi/nBaFCESnI/FXBFwgZ3BHBcBqkLD3u/j4iIV/oKCyNrTgMNlJGI/2
6JJTTGn59jZS2+7oORYn5q59AMq+JE/PgbOvt4Qawe6cfHWqJEkKrLtNaepiVIIvXmacf3r7vr0o
AABFdkCMbHh5qVZ2exnDWPljfqIaPWk7Q16C5ImYeg9i8DL2y3R7mMu3G9yeY/fAq7TqSipFHJbo
nXLN5+QwxnJEmQpw7IeduTwi5fLK+M/OIOqUajMrSngpV4QWAEGU1WmiBneoEXWF4mqT4Ah9hZP9
F9ffFyCZ1CaUhPdN7tBgg6sBf/dJGyhypqCXtA6RA+BN529ISLtxzbIrakw4J/htqLRlN/r7nFKT
tukfd7fDMOIWJZsWy8+CTh/taFNp3iKS7iQotLLpXfzjlgDbQYPpriK3sQFfVdoYT0Jl4AFhKoHF
QpULqqpi4vsvbOzvnXx6Ha3kClLN/SJ1/bpSrlM646ZIsxRqpf+KafWU/5P6bkFtMsFjCGTxJxh3
nphXLgY2uJvtxrryog+awjYyvwu/sBsuUfPE1L5prFOPEwlTZkn9Wt/+ju5xpUWdws9QTVTGtuJO
vbfW21NRGT8xmcfQ4R7AI4Kku5YxUmGts1kGhGMOQg3zfcDJuOZ3A1FrUTSMc/QePQ/pnT2Gac/D
/j5dlSLQg88i+7AFqjhSPR3XfZa5U/G61/O+vI6w79mvsBgHfFWn2AFjXafcC1AA7jmUyKzc4e5O
O1+UFZL1T+Sm8y6hi1nbVhq8TuPEVuAk4WxEXQJQ53iQMCUETCD2g/TBNJ2AzJerTIBegYhFJ4st
g5QYzO/N9vn2liBE9uXNs4fsHjvYANBs8lKKer8QAZnxX9y1vPGU4OOrxvMXBwNqAzVn5uHoqP04
lWvLUsgnq65Y3PKwhW0ywq4daPnwxNb9Jn+YpAZ+f27GnDT+z0MUbpjtt6PkvHUo0iXeLwqk6hwB
GaogH/8Tj66MfzwA8VPG9YZzPSpk00uTHF/obEmtkGOnrPPs8QJ3iY9k7J51o04PbRxOiP4MLc8x
anPuIWy+iuG+LJZNoovkguQj5Rv/8UKNCT4qD0P4vkrio1yZyXmJ04l5O+mF7+E+Mt4g2QFbQVY1
+MhSLswe2QvMMSK9qk/uoep8yTYDZyUu5BMpbgpbpOZ9zcZhZFvVtUThyqJSZb3RhE6dtDjxTee2
K+CNjbPvaW42pEmrceazYqV+yz5p8VpA7MvN559ARf1K6HMnuIzpAT6h6hzzQTyrfEaK3miUxklg
z5yKehycJOT3G4YyFxpOhG7EfBQlZsKnWRugOpF49PTgOAWNTSou19gKFbb561cLk2ZsjfJxxHAL
b9vC3BNQd6GQ9TZ6w++v6IJ4MZOvPjqvToYLLOUdmhRkHT97a2wuULn54FateLkMHBpUN7vOMgag
PVzZQJCBdtJCx4b+C/MZfx/yNWDpe9ee1xncx/fUR7T/PgBrwXOl1er2TCCl3gZ4k9knw/6ts/8F
CnkSNHvKsKNLWUfVgCpPMqHnby9Zhhme2rNKX+Nm3t3/dzwOXdrSrs57TaZn36bnNESBQ/ELig9W
ysjC0oJ9iK8Zn5GnEkfTsYA8w3Ma8HCLKZAYed+NdT+ZEVJ1509GJrDCeMq6hZOl9zG9GNffgQel
BwK56/KUsv03wNN4Lkbp6IVvklFwleIpfTUZLjXqqyPEzeIhfBHM2BJaBFLDATEbHnzjuOBbDUzB
hv3G4ngGWBciBKNInHzCdDYqeStXn9drJ/iuKSTW/GTs40ng7TzOdyPslG0MiipGevsYC5n61j36
C0ogvzv8FSHNWRTQ38M/3nO58FWFG9MzJ1+DNOURmr9c55XJbtas0PkrTCQEeRiQD1ZHdfSRMYRX
J2YlfU3S8WGOUhGYhrTvgXqQ+WJPTX5HL0UAsauxn3DNdBizgi23/2kcPgSzD7MsNSlt0Uv0T7PD
e/P4wab3ZQrMZU6ldq8IGnWLj2yXkOkvVaQwpfDCFK3cOTtt+rrknfvgU5yNYtkPUFl7djDNIQlb
hyiT1tKojcQNGVbhz+moYkipCgKrsIbC1b0sRGpfWwuy9gNWJB+TpGdi5rCe3DXea6Yc+ysQO9j9
QHR0JdaxKxMA6OrOcUm1JSSqXGKwzOpGx1aqwsy2lcgP1B9RZwnN8v3Wsww0reSJjnAJjuqIuhSn
AmcpiOoTGOWWStcVVPoQIjQL6dLnPJPp5dgAlrx+1WO6ZQ30rfORdphukEUZ0Z3phG2oGbkp0Brw
sVtjUfDpyWOx9enmJO1B9A3pzB/7PYHS6cfFAavVb8VCJxy/VHXgPD97Hv37WRXBocXUfp1LZBYT
UIbZWItQeHQ+sj1nFYpNBUkdF7nZfQ93Z6UH/P//6EKbOJPYaWgZea86TjsCbheqYSwZVwSSmSdE
U2hAqoUnMA4FkLCqN71KHky0zOpQaDHcyD5VwXnkgEyMNuoBTHsLktp6UOtVLr98UgDw6ntqeJbQ
1NckGUwuj8tqEPb5U82vDuckv3szZb+MLu7igUIkRl84wtApAG3kjZHNYckMm5yyyFFXbQj/X8z2
hQbP4J13LpGCPaOIf5riIGBUSlKFT8a2JqOEGHF+LI+z1fkixyMVHWQ4aHRm0XOQi9/2DE9o2sVt
FSG6BjPkiDzYNsXdF+R0YAkwTUN7o5mC3QOlxi5WC1TsgVR/80rkKEr+m0AeihlCQSO2h+iO/ipG
ydllbO0L88M9GE4U/xnJT4jXPIOIwijFScxqppkYfmUcYp3iNJBxU3exZQ4HEoy2RwOTyPcD7pA+
DTihMo9arSBA+pkYPXAnCxrkwRBisL63kzJuVc+0RvFtWWvMTk1xX6Z/OCFdm8rpfwO88wjMJQ2p
h0nxNuAoh8TKs1Mqp+qRZYslpy4cQ15WAnttiQavsgguqPksEV+BZCr2DVcTWs6SZF+XMlk9ml8e
p9BR67fUugY60TKLwxGtU+GJWcXDoJj1xGjS9VA4nBQQ1O9XHq9t8mv+zACBhsVWVdP4xsASUUJA
X0qVlii93OsW81CcO8c73DNWDW9FwlDSDqi9tzZ3dvd96Hw2kT0WSL18/Y2nRkrfirFBrrhfDbvN
mTTQpP/EgY+MHDocSeACuG3TlidgDrjP9S+YbMBeC42wOsWoVxtV87h7ERnjiZxYwZeybEuhaBK/
GshzZ6wxRCLUUUynbKlTHPNYv0ZsUnkhqiHI7aq3T3Heu8CE9z7XL9bgFMKBW0btMcf82Qo7zqzR
qrBsPTCHuRrjxXHKF9xqflQIrYVul8yBBxL0mp11svgpiiMEUkVEHdbeRALLkMBFOcrlZN4DzhNV
CsKCVxmHs9S/tcCBeGTRx0HKl0/Db8d8/K2Wqb66mIRct0OxxrPqw9LFCfy90lu0TIZ38NUyG4p2
vs4nv/c0xunWZIemOu+NgGSGQJwF6Gh9XRUeaM+qanHMHMMi//GM1gSicxRr7enHXI3RIo1wMbjZ
n+k+sEg0ADbORlMhl6SiXmnN9Aqpiific+TbPF7D276eIYx4CsodKXVlC87DaJA47/9t2yJJM3Dc
T4eRhpSPkGq2noBtJNXoeKatcqoOLt2irNNXLyIRtmKpWYze/pyOcl2F5EsdveajU8gHxspBgqgB
bILwaIHdvIvC7u3N79T8k+8aUhdmIt1cowDXz2iJ1Hpu98UkkwkZV1a/2+sm+jV4gXe6MUXOxlpa
bEfrmUfuwT04NoPaMPjJoAQmL8uIGk6ZAFpN/D6M1dpku+zJwdZ9z0oHJN/tQXaCAlzZxK/fIFtG
biT5YJHVJ8VR5bdLaqpY40/4saLYoPF8xIZwU6XF9FrTVn/7V5u9LXP/eZzWWAsepC17pRaiN2T0
yAcxx4N4SIBSehHoilyf8eQ/VWFxkkvZp8X8PvoJjkxOqRHjv/K+9Eyeh/k4CXt0OKG0bj53VX4F
ckLsspm/2/O5Zmfnq3BN13qsweXk9RUPP4CYjV7iJ+8xxWmXjvur/K046vmy/N/FTZP5Fx7W0lPY
j+PJ7FQjDmg7Te+nhG/986csnPhG9yAES1DHuNGRLe3RHS3+FcQ9gXX0yK8CcqF+QcQsDG/4gNLY
AD1khaNYVeizcDHhiMyxzT3Tpdm6c1OQxP8p1gfImIq3AyP2DAhF+HTAOzvIDO4qRfLcbygdXZxr
NVxVnHkn7LSXdzcYoUb+QyfabEY5p/hSDTMRcQVxxeYhIRsyxQFQglfj1tZPK9FbgbhfivGM52Uz
VpHSyyTCzeCPhsrXXqCYkcYfOdTJTJyTSLGjCvXCW4ndaPd36M2Pw6B5I9MYTZqYXk3eS25QEZBv
wy2n1RXB7xucY+7U9lMTzc+tjsCHogJE99NDoW8wNvXyrhnHr+yfjhAmg2CrwchZRhf6hLYouX85
UwcEL73tQnSbaIzkNWpcDosuv9LvANwSAhu9p5J/T6DSqqBZM8OZf5E+VUqaysYpW6q100Egl8me
YMKCv70eObJfQHnOyYI8yk9EughBzpxsQqf266+aQTrEgi28PQac14kw9KC2jCSnNxfNIDGf160D
bH2npKI5inZic/fGS0l7TDzKQNcNK/LzmaNMuassl9TI83NsRSzNGvn9FIAbsIcQkc8sFlj0Rj7H
xr0XzhZWb85uEiLPxtotzZtHv/mUk+VSefn9KgQ6uA1lI4g4T3QGO7YEk/kxwIOIMbQtOYODLYxP
DN4ZSPU68B+Qgjl7+xEHg6X1Dy6+QE2ICh2iYfcNXDTgsG0WpSVsTDt/FYUgOybEvmMzcxJkLFG5
VIuzo4Dn9xVBzJbj2ooDoIeR4qEW4DQY8UTdcuaQ1czWHa64xShE9owOiLqIQPctzutXX+3STjbM
oqBdkj5O64Yyw8h+1rHgKuFUisEElW1y0cfIYLtLGWAYjVlJBTrm0fB8/eNo/rHzdjUfQxLlkA3J
5kAYspYGDQXxoLiUAjL7zxXqCriApHc00Mmzksctt8bvzLYXHih3coqkWFcfpY6/61AoZ0+fAbod
Hwl/Kx6l24oiVjKjyy4/poDooune/SlrwIXQGXITlBL/C1vGhhcDf3NRe9Cmgg9WmCgTcgqiIRuQ
8s3cGz0GKCcP6Iy8MwHICyTPKBviXtTC6lVzQCKmpLs7EkSs0kh89DASjYyxX6QO/fpeIay6HC2v
PECljFWX4qz3vBzKn2s2wVoLGILxPT7SJF1GJmuLY9Q5q5FIKM3VgE7qurPl7LywNtmNTx3eb0yb
QBaTji5kS2MskkI7eRCnSNrkK0KYfVchtbbstpe0OntvIPThl1gEaoNhaS1nwroCXGjsSps1pKDa
uZSz9HP2B3/ric4f/dHDbPdCypaNb3dols4HZVl7xNCVqvKukCPjlvw89Zg1TpiVSargUDq09gjM
DqFBV1LYjSWRFfd4XAUR/wTTT+WSbGJX0jWRjCnhU7H4bB9I7XEraw+ZopVnXCOj+fdrUGEZIs6O
lTMSnKumMlpzklyDcA28BQ19tKU0TfkS1980QusvQms0G5de5Sm/oKP7EfhWimms1nGwUoF6uO1z
7NX6w+tgtrbZ03oWUxsDkEjILaenXDLj7HbjbuBw+jnlEAr/Z12r04QiWFQW3zTgOTReHzUzdbi/
n528dUfD+ZVjoiW5ldm+dHDz+upTmavtecltCTSGgEi5O7jT9bBDWpyem9rBRGZgGQP/+KZ6CrLS
6+lZRfd5OeeXmf05WngeDaDniCh+ol5gV/xT/MmXjdVsjencF3VX/ow2HwIS1rVGogIaTuhhcGAL
asIxgsCdggsa8DRBOgzmqlIJRLwN/D0BFimg2+ktg3XeER/65nvc/J4frjmKS5mzMN1hLRxslmdu
XRR5lWLlgNUaTY8OE5flLRkYuk43FgswWR6BTEGmcxw5nSq1nI/o2UQ4K9RBQ9ZWZNhFS/szkhLn
8cQARB7D/SqKDN9IRFZydrxeGkjdhAHqR8mqHw0iD/2H8UG9vgpyz+I9yangR1Oi5u/rJzHhFih6
Fr1jgoUZmXTgztct3uYltu7we8bh6wzsg47NAo+N0SHt/7AtCPnHdZV2EemAm4NAqgkbALCt7ay8
pEpt5hgXJCDtqvwoVBf9xqQix2rIWY5bE2Ou1H+YM4m+LwFDF2gglsxP5t3vG9liMcOV7GW+ExlX
8/GkYse7HtNG+iBcDQoqXLrIHY95gfJhhdeS8iQU1vTe7ZO8xc80yualj/P5ZcNgorxn1Mzxtv8Z
OFVFUpgoDEq8JNSXlX/F4fQksX4b0xBWGsVwjZ4z1YSWEoT0ZoZlD2yjTM9aNH/g3uciTdz2nAr5
SkzbQArbixhWeZretTqEu2qbcy8xwQLNumJXV3UdffohhZOvS4TpuWUHO1+BCunowx7I60KhA2aG
3aVFpSN4Xd80oSZlDvJJkiG+ziXhCzb9BsyxiPCjvd9HKnzolcIJaf42PJ8Eeehn3eUNafhXQRpV
u6woC5w80glZI+QwR2v928Rl4coSKxfUJsqLI4jk2W6KFrE8UymT0937/zNlW1i2kMYNFzYk6hBp
k4VP5VI/PxMycwLJi4VsqZvje59tTEb0dPut4GXM7q3lucoygOQ9QYUFkUAWrSDGhizbDOgOBphY
zbz9eDQf6ktC2rtRESxxNgCIQlUC5+1XCAxCU+TR8UlY1QHpHfIzTtuDqhksrxQZK1leqU8MZpnn
66XRiRh9+DgF/mkzsTk6dqxZVXleV9LDXNkJekrHoKlcnBmM52HqNy4R4mcsbUn/pC8bnJs2VEEj
AktOruPTfunN0K/IkVtwN/4raJLUzlVAJk9sObzwUmY0ofWSQdyKtQ7Jam6eaqnlrCJLxn35UXQg
Tfr+kPJ1Mx2BRmdtnRUEjuhTVBRVRxrHgDKfuJqHhcvy7T/c5ErwhaIFFoYYL/vSTba6Zipn8SoG
ZcGSjBj9fC8OitwXDelROpXI4qSk+KHeZx85vs/uiIfPab/6m1XPhaeyWwRjco0LK40g9qrFWqru
sb6R1h2stA2P5ImX2iSqPfv01EGlNYqtxIoxXovBgZT9vZ8G9R2nw1FXDex87FjgeCHgWcKQuEbN
7lh5F4qCdZOHDh18pM44CrObl+pj6D7ZmnWpkdi7laxKMf9DrL8Ucc5fJFLHifYTMY8GmgOWq5CX
k8QJGfEQhz8Q+Rx14//dzUXfjNDTeXk0uCPXZ6Xp43Wiu6b28zYvhyN545HOhxa8hVdVMoN3WWNU
1oaW40rnUG07dXrkSTwTsB6VB4fkUL919PH6b9pdBgu6cjxpWZaokjOqGxVY8wbuOtQ5hHjG1edQ
e27g+/HiBOibh1FsrWY49170vlLgu1RVSUeo37t5soN8IX5qtj01t/KBe/aaoEASmLPnRhdpstiz
hKY3PtwTntiANvbdyWi68N9nXff4lEBc3tF9qEwnxdKvVKD/AQYBs+Erk2rhK4zkkNIEd9z685xd
dWHyBwLSs9oTlAP6BlBwWIxKm5VJVGoPBO6UfvF2wJamkVQ3wD1k3s1veD2hFAuWaqcGW/0ybiIw
fZWH9GVzc7cZdJ86Vc0lLG6M5E54MVPTXgWPvFTPCEdnb2O7Hft5jN/KEqo62uxMQpNyLAZqVpja
IVE2Y2e2v59B2vxmrmyGT+U+eylTDhayWPAZEVjnt6zNTmVsk6mIIDzaKCnS8ZPWneYvcxSnkEDV
+v6yndsiFMLknoip9ACi8XCJQb+SgYj3F/gJFxBjKeHREBda+cPBQngTP6HKQQ9Z5Is2D7rkbhmx
0egAWnSGWzBdKx2PrMlBsDVahAShO/Id4O2nfNnuVlZ5bX+9M4bKmvfWrehojNdrnSu3JDSwJvid
mBXgG7zYUh225/Ls9QXTaqijZgEzn7+rU6XLiu+X9gOw6oB2TOYSKadhWlkS9KT8cIw+RjFDFYlh
0hvKtB58eUpjVyqW4kfP163UJogWULd2klydtkvReJYwucRc6MFgu/MLm4In5fth6SzOlJbAjyxr
r5W+ZOphtCtjex2TyK9s8NlIx/TkmWmKZiwUqtpItijVZTzUYPV+hlrhPFJGlWQlk6FnqFajEpWd
PxVFomFzqP3u6aoJb4boX8mKujO57sDyPI4Udn5NS44S3f2LpvxTWPNbmwdcNqJlAGbtXR5w1mLN
hUuBFfkjMGb8bgtSJts4FdP2PJ/vvV5kcbv/X3zI2KOzxR1SPLcMRM1NYj2IoCxQNMmw2Z/BeixI
pQCDd7F+ZpQ4T7x+on932Y702o5epDFz56/PL/TvCFIywUZMVlUGe7waB9kns/dXWl5gYapqx8dr
YvN9igEA8UAW49xMqYO+VSvgGre9zX4hIQUA9VqVl2vBClx80UefN81RG+sSwkqXaIqxaSocyw5e
djlJN14AfNMefTa1sjfFey6okQkJoTawSGnGthTHQffLm6xLIrDpQEv4B0lpb5E4HDaWpc1YOVcj
/0iRTMA9CsRo70mmnRx3yH11Lx3Ovwa3eS0joFhBFDcXhMAeBD5Kx8yLDSUXI+k/M8yOluiHeZCE
FPvf/DCf/fzaosiQJod8n/4NdPpEzQ/e5h2uKaDS46zoOtmdLD2eq8vDug3sA5N+JyiQFVNBYXBM
JcEAwRrivPmYjN8lmOYhfijHe7eZY1d3TbmwZqK3nKX2y8uhcmYwBFxHQgPTCK5LtaiaTb9sOMrD
MJsX4hGZrMljGqwBYA2cIbfJY5HcRtypwOyxfGhwpW4RLRfN3RZLZHc2FzO4hpr9WnqpLR/zdTNo
WfxuCdEuEQ1fqpOu0WXPjqv6aGh+blLeqiLN93+rCyOZQBjR8uaHcSOu/vgeJ/TNIAv/sqeEmybB
bR+RXjlugoCeQXDFh7QYYuolUwFBh2v6tKt6sQh6/hs1Nv0xM7hQhLDJSctRCaVaLQC04zWwL5Np
3IIcEZbL4p0s1ym8X4NbdfsVydmLLudyb7sAY09AWtsX079R0/RJvaOlhiypbbnC7ica1e4sC30G
RZLy7Q5Sk7hU7rnN8L3ctRi5z7pa2yQ6z9ogUqnuZ0n/cFzqdUC/ibCyIR4TewJipAwaccW/tw9h
nL0LO9qfaVwPTS9ePydVPeRGudQnHS6+UHNdWd2+MhIDBiSMoLgEy5HH2mZdX0juD4BkNTb9AYXI
qnTAPhmL92wtRVKjXw36HD10C5s8Rjl7msJsGX1aiTpObgoaaNg30x6HqE9XR339Qthpvdw0tACI
QCbJP/q17OBwdboFN+Grqc4ROW8UVtaYvHlwxbZVq/Qc6kfGHv7xi4iefH7Y5GfmdTg/uQxnKanM
8/0jiL1OvriR2M0FODbqPBB1BTvhcqzLKIrNdq4eEhWfVE5sFtBWrY9uSGN4Y9oUS+42HdQc+owM
S2mHk3+tefCTM/MN2DDr7sShYVudfjkYCjmjaCQQqCHz8Coet9TowtjU/edey6zhk5KE4+NDhmmG
rQ4LvJDUvYmUFK7mHxWgb5GEo3COQr2cwun/sCWPJiq9n0FQJ/j+9FDOyfulBgLSa2lrAm/xRnbc
Z6GsyHOyxqIojRd2N+HuC93uh263baEfY0wic9f4O0+TBfWkjWjZpwcyyeQd6g9a7//zREMYOYtf
+I1uqdt2zDtJvKr+qL/bbbN/z5J95e+BuBD5dnK7THww7masV0aU3cK+8KnFU3ZLXJVkdHx2VEdU
A71t/qog/vL/R1GacVcb/ssZA2RpAKhpeCEfLzBfuQjWEbILa4mPKe7GyOWPURZP3jRsDu5llZKK
NUKcubbNXcA3tyVvkwMEYGl78PHNVtugooLQLuXdf6xMWthiHsYsNvRmp9FWXtUh3I2/t0G2UrWF
xBQpLrinIJYVnsaZWp01n8cDuRHbkkK/tycMetGesv+zpjJqs+u5lvbqpLjXbeUqwNPh13KmDia4
esbkFAjDSOhsmCDoQ4/SSH8HNfRWj8oSoX/Ggn0+Hcdf4H0tMcYKzUQN4/Fi5Mt2rSil11p3c3Dw
C2zz0nHnTT0rdJTyBtuwGWVYRmBpF0G9Jnm9IISr1B1iX6bi52UEq7twTH7wnJ0aeblj6VcH/dd5
eCs24PgF8Re7uTtXQjD8go5nGcpDg6lG9CnuquT3dyX4pp3//78SGgSQJX6X+LdjlKUE8HFulfU2
XKDxXsbz3s/7TItd1pgLW9MgFA6MSS2bFeqpBKCOAnFfNtX53cuisnbG/YuWxL+5oP9exy1PgL92
YXi6FJTwqBZtx7v2ci2PGrWH8Gd9VrhAay7DCE9DcUvpHtQt2u8m/WquUgNUOezAsOHERkYUs/0X
/+HH94SAIcs3y5/rnbQngLGB/qjYEAbZ1XmiWNE6hOaTCcnXrCY/mqlGqCnMvGnsrJpkgqV8wtOo
DGNorPmr6zY9Bkdu5rSg/eH5IVt5ZtEyo4k5X8Jy9YlYeP3hmVoMmJkjH5jAq2WgeuL3yu0VePng
Zr9GLJYLsSeZMVl082Nx+c8BXA9YfCr8xvtwheGFw2j0RECDtb5L+kH8ZgSnPixHdV7NK9woU5xl
fgR7UHZFafl5D92Qamtip7cPSVj6BC9wVzHMe49msP8XGvw2XrfnLNulEQN8VwvVCf3hDSOrl6zo
DeIrqBeZyCbPQmTTQhcMKIjXBNb5JppLUVDYYKExQN7Du4sOjfazmGtPdmajIN4WHUqvEI//RGAf
iNU3HRWCbbGBc0yQ8RLhdo2un4sH6H///M+YwqeUq0ha/3KOvrIxWT9pFRbjApAeg2eTmNf+YmBs
D2w7gbKunw8W/fLl4IRtJerJH21I55EVw7pEnwB+3AJ1sa3+DyNabf2ib/A+2mJBVNAgNa7N9zEF
NDyXEXp7i06cAUQOXuM70qMqt+QlHh3crc226TAXsxYElpW5/jqno28GaWdquhKhQTqq1630Pvo7
1wAkd4xVAsZhtG2eeXhENxAiqb6jDyqmPrV6JAcxV9Rt2qcnm88O0l0qOr7efkLV80OeY9Og8KiE
/g7GwWpsov+tmwCA7Q3cIUKVytkyjMiY7WC9wlB6A6QnLGHi7yKhWdaLm1uDahuOgDE1yMeamdCL
oEB5QJA044Zq5ae6tZgAb0lSCVkFLF7evJ1wB208RsSandOzK2jWJKYlFkmvlGtDuvihf7W3Y0eQ
o0+R1ld8GWLmbX3yES4JjPV59+N7nv17Z09/e3920igLEL6xORbTxilZ1324DWqY9wNogF8IIzS9
kODg7MTiKs0XkSd2ptT0UDxpGZqWgkv2iaZMdRlvSPPt17eFvR0zZxlt52AXKZ3hlGVL/V2poBYT
QYSViT1xrGeMpCs8Vl0EYZRZnMqPXYsrwSQj8Q5vOZhC5OO0A7mGQrE5bMdjbO434DCcY2XtR3u9
TFXTJqX9a8pkTfqV0WkO0739oqEYXOT1/6fczMQmu7oq+wkQ1M6+YIO5jbIA5ATCIAUuqem/hXbd
m1eWPpMksF7tUt8CO+UYmvfGheTiSBVMWmDQx6zRALEqG+8kf0/1eiVhljsPAfqCfOIjALV+Fy3h
Z8kLGLgUvDsufKUoocHM0sFGnR9DoCB7rXva3hfNsXXh2FwV83p3XKFHZhroF1N+EubKohB2NI0+
YcgmaRqO5RpSbr5siZe59s4zPyd2nVIukwJOfYNgD9kIMFtJXTIP7gwl3lBubX5VfxJywGInPuO/
yDuDbaFkiIgvbkK8BZp1BizYLMKgTL/quHrMh4Oxy0zr/y8+zITkvM2jvRCatf8t1X/WB3+ZLm4d
8STYSvnC8DrwTBkTcwwWbHAe6r+h3upIRYuMGcjdy1nH38G6gXJjl3tqUvgB81alAWgu3wGQR1pn
oXz7S8gS0c+bUPcAGwNIVR8r1kbcL7jmpmJX+2sjh1klppSSuWss1dCw5JmlcSolVwHwYkYHMN9n
hPn7vQon++kvFM48Mb8WvN2hS1t4wPwPYVWiKrVctJvlAWKNl+3RittYyEYGx3gnlHlC2ucezo09
B9f79CecZYCen8aK6hwmxKEFz51maKkXXBVqy9VsAqI0c8Jybvclyf242uIHedtrAQVDEN4qKrrk
AbWHt1DUEOSTcbBYa+EC+DhWFwQjke2gHyKORSoY2nntDV1fS3dkX6RCKVWebM4RDk+guRSNQT90
SNtDph18mTPuhxx5L9wz9VxwUZnwwukCW7E17Y3OwbqnHjdKi3IWFXNo8OXbT+p1L5iDVmzQyS2N
hoacjBIbEBqRReo6uhHaAIPWGqPVN7q64yZNrzq2NWxs9B4YvA5UAk4h963sit7DdrWG9q0rHlyP
FRUMpBC1oYhWcnhTw97g8KKAiWknewpUPt5sFUkla/AUKDUs66wR1pxJ1odO2logg2olOuOKnCBK
jqb7ATqKmmJMBtzKfHyzEtspL2uN8RGHFAp8uyqKai4kqCJ7L1HfB94ku860CuZ8tVjNuluHz0T1
UxOAkzvHCxmdjHf43INX5gz1rZs4ezu4Xm17kil6j4YkrSMlIFIwAlxyaEq67IE3cQFWJrfYGY2o
hpijLTxR10UY5e2Pni6T63RuCZ2XGL9UWlZrJiTDZBUvvFIGNG2F6e452ps5QkRiWsucllryyosg
AQGkCo2xUFjb9PcgcBkpqEwl9foy9vjOMsnOaoE/2pU+1Jg8eK4kVUW1udtesWKI5wG64Av8PQX7
q/SXesO1M46awH3xbHkCzL3F8/t29YLh0o+eo+WdG8GIHVFFPQlwDlB3DgOisx7obhHvAa8/ddiF
V2Ehqhbpm827iuH7911ubhKhageaJMN0MRNDSp+LR3MNc9I5iBXTSiEewtXOoLpeCNDT1WFE9Hcq
srATpFmBefNprCaUKLe2d6QIJ84jd+dAH2Vk3mkctQTBVPyqsNQ1/ww2cIW3Rooe2ObnKC9Fe5ZI
TjH82fCK66YCiGqLANVZcYSUqBdvRJ9RRF59Os+7X1TxVS3Ii5eFgIxPnziO28cHSOsnkFdYuCBh
8PIYHkIjW+drvdKrt9tjMM0QI1iKPSF6Cqdko0OfjJlC3FJqKkSoxVUhxsLf6XKnxpJH+hFlW0Ee
imLMDfkYDAb0UrMTnAtBURPoVAtdsZrxCAeOdtc/Lz6EdxQd/ioxboTO8v0Hw470Jvy3Pp7LkP0p
Np65S1IlAntzUVTV7uDAQ7ZKequ3gV1wKG+z3Q8/x8/ALBXRpEaY49Jh7ijLlDpWf3h2cLJfUJcl
G1RMnZLnXeS9mR0OTHPhWKscQlif0xVF4DPehfmGpPn26qN13GPMYEQJmiUKgmrFIwp7rJ9GqAuV
ybTN9/8oAUiGKqGmi7R85icCsoVo5EVJ1aQIVYhIbLdA43P0RoGx+6aiagupceaJhJ9O4tPm7WsV
G+4Qs5lhH6wppd3RhQYYV+q9tGnSeDxhr3wVsrdogW1/Ky2U9gf/jN+jhVc9nzz7lcJpG+bPDRag
7uF6L4lh+FEmVDv5u4WHR3G/WdBrX79BRZOHPAIlX8IoDMMgvTvkeFplzaL5TRob6gy8dvuH9QrN
In6Jt2LEiGWp6kEYMUkc6j5gzZ9/Xq0gmsc1clp5wsHigv7cDvfuXEspml+WgKVO4tXZSlX2Z+i7
3ETem/U2joYDQCc38hZDEc8PJos3xp2W0/NJ4bg9cXy6uE+V2MhKpPNCm9uOe4qVp9nhtqYA+2QJ
djyGmHwoAvGvc7fxn5RELV6kR/uYHAJSb/NsFH87ebedcRPagBaakUYJfNB7MNkhcM4PACelvQbV
qcT8Ci/cCDNXC1TMhfpxI/bOF8Lp3G7WFDpbSdBDQfdkzNtAA7oBXHyXyv0ToQs4j/HhTrfMspnN
k6msSRDsm3Mn1GN3KkrGdZnyaHdWl7X4Z5X1H1qnpPC6UBQCUO8lfGtlz8LdV8UKAqyWLAN9ZMKZ
3WjOgbszgKYfRoDI9jS+kBc/9/hSko0FtVFQhnAyHZgQdXiVT/HnvJskorpsfy/NQzTkGfxK5cqG
e5l6fpU1o3v8T5zXCAv30aMveRttwgLzVdCY3ktuw0vvg2fQPMWvCNDlCdhzwWvJ+Nu1zmWjZY09
6OnyYAxc1rChMm3FLKRgqU9/AC2l7PKOEvPlPvPlls6pfUTHg65BxbmKqI4QDm8R3T66RDox7zkR
FdslPtFBn6he6DZkvUmX2L2YPPJAo7Tyacn6ha/KulLRSEe0JKe+U0tdJtTLIfPSSh6LlbiJlVHD
+4PhgvIEk+lmHHUIUYoO51BHuK/oVI3lsQ8Spfyc2r2ctXYOP9N32BbchT2nwUdYcXY4Lt4+WxIY
2Qz9x0NWGvnRI56pOD0JYcjpAS1BI2EzKd1s3q/LQZ51So8My+KfZgaqgOwZtfSUZfMxlJno6q1B
CH4LV8X1y05EM1uSto1aa2Z6dYXU4ZlYlZoo+IBPHcuHvd7+pTAVcnvttGKEWiFaY7XUq7VOkb/8
BQ8wHu9Eyl/qXAWKuTzN4khpZFPr4sdMn2Oj50jwBiN8vWONklcEMUGDvuaANFaEe/O09Nm9ls2w
ipWS1y87CIqeYbu7r8YwRDPLmjNdiTbrixXrIOY+86LD6ZfRBPtNHdPgYoHy+N0vCjQs1sipRCHo
kwsrCLDS2bVwsftE/3Wwp8UPTFIscGWwStVbA5PDEXuX7YsZ3tMR1K6aBgYn/6ydojGizLw6oXVv
qn4bNYT/m+7s9IOBROdFTPeMLY0Jw3ACBaj9/LZvknh2kxZ+K65tN80iVOQbhPRkvgnzziNsudv6
11qRkMsI4mdWHzgGMV7a6ybsLnGM4J4McWpnhCzQJDzgOHtRf+DiI2d9AfUoi8I++gz7+T/Ix38c
nErCL19yVzYjC+uF6w2qfaDuT2ozzbOWJpMlOfYQWLvguZZmbTCiQlZeid/zV52IDTtBmzwtsQQE
mGWpdRlUpj7JVfxdHPgLnAzzZtCMUIKjEgtxmPaynXQ6dEIIOf/GCKsYtRBr/24KYDTR6kmF8mav
zeirmuz95mjAnSj3sZAbYrGV/JU7XwrTq2dgE5hrSFLUQ3WaPl3t53Vf7shA9okt0KThkI0cQiBI
sUHHWKy6CZabOKjCK8lmqxT8+ci4h7sTaqR9OQemnzdxDehaI92bDsB6ssEWFPeCPYb8XiZTf4z8
2vKKQKK3POuqKmSLDCAN/TtwMiBRjP7AcFsHrKDJzuu9oxtFqGAK1sMZ3P0cAGIXCHmsWrDZUMXQ
PbHQi8Vb1L0G78yMSSxYRhVf3XcB+q6QAvtS8kS4nGSvq2sjEEmuQDGmv0K5iuGBuRXSR4zC0yY/
M+8QPlmGIw9bmKBox3bm4zvLxf2z3cVXwyBKwRfPIAsvfAAKJajAEu+FkorbSPCkSq0Y2Ov4NcQ3
MK1WGc9aKPQNFXkZ6KhnJONzifMQby8DatNtBfKyk44kjHeLvpFGMTS78FMcXh3MDU4IWUlWYFFx
Pu1yLAwDBS2Def98Lq/JbEkuw9Lk3tFMnxl9xg736SuHSTmsDbEtfgJMIvJeNiuk6sIylLGcn4Ae
iS+sDL1wr3MrBA1MryoEGo7lxa5QhbK+Uhlv1yzGgS7f753yaFTp+2JfD4FCZalZCSiOl4wg5AoQ
Yq4jPQz8TfVS777tbGAMZkqYvzHkXgXIszeEM/tnvSGAg6PB2Gk6QQskXrzy//ZzyzwJnvsGnko3
+IMrRMrxhudPS2nmfXERzrMOKujRwSR4ajrgwjqaZPQpTCSyz2Rw+DWOKhmv55BrtI07hLUaFhqz
YlnbXa91zhWTZLdGdROaASBpiS6vX+awIffoXXkkJr8RUiSkfNQM2oHbU13zi0xyeN2mWgu+QbkN
O71jmHUcl5D17iDl2Y2ZgK9ezp8/D3vmkAVMWj/11GbEFVjswW8xS2u14KcdZNzAWFuuqlvnCvRt
EgvLiTJaJM+4D9BFXHQUYJReexuRSwBs3icDEPFXB57CHHqnNz1J3vlckvWCEyQz23xuj9SsXV/T
dFirydGp+Jz+rp+nuBt5DbF1uBNWHQGore3fEqSTjgGKGns9Rrv2/gh3Wut+IXQa0BUyiDeuuTVr
9E3fz4dMmqsIomnpbFE41N1dUqmPEqiWFMEw6EkcaquFzuSgPxYKU0mPqNv2pr+4y+F4+tVV+y88
HLS1frKtRxJZwad19PYFnVrgid72wr1XUKfU0NNnKVdgPjZh8c61RNZQEkijhSal0VMVLjwWZ8QD
am/rZuEWCqvsrvsbjlb7H8bPVYGwIna83ZNrsbon3V4IJeMVPDS2MromSImqLs7bwcpuxUp9hY7B
kSW68Vxwq2QoAQqnITXDEzNXZDzxRAnHIGqxFwogQvQ+lhslplHi9Mf2B/CcKS5K4nfIcn3rvJVz
PPTfhNUCkDenw7CWXKDAOA/4zTUrjxj1fzsO2tGbu/Gb07cTQ6WeSo35tHOkxFjtCQQ/J2IDpfOB
s5fb95fsRmzke4LCtKAfkHAzdx2ys2kRsssprmt8s1eLjEueiEX7WKJWDeT1Mw8XCGzUHJqosMtq
e7W955lmArm/i7Wu/swmDME2hQNZ3b8ItRobZ6V9AdLfisn1JVhbsJ4pP4wH2yOOqkY/qVAQ9iRI
XGS+NCeBBmqUWjykfta81OvTcz+1QAEA7CBkWprA5UlkXm0TmIJOItvP1vPHA/bR4TkvG2YOXFCo
jsz+MPBp4A9a+s+Bwwikdm4AtbxvBaTwCyrl48KQTFm6o7SV5SuQP3+XWuM2WAu0xuKcJ9joyyso
hn4chzH1w4IObqKMQciljemocSQCWVetCM8Guhj45cqvf81qX5oJUryHAsHa+U5OU67bum71zFAw
bxHpbGNj1WEKIDRxK4A/JaJZLj4LslsWnfmTQbgxUzL/gtElnlCQc0ayVYqkj1Lvv8ZRNdbZRdje
FZxgnup/juJXFbhWAozb6C6wmeY5oQV033am+xtpsOcjhLt3X9/xRSRF1dvDVWluDc07uzMxMbVk
tI34N/E/j1s2iurnHgxmVJEI9IAaZCrZHinYblD9Gecu1Q+6XwF4ShPn/R6cv0Q4T+SccGZd4Sfx
irw/KGjCg4lPC2y6/eY4orXqrYBpMTcwK8b5mDantd2HD9MtE+utjosZ2+Su5jh19+UtNUVni0h5
GTkIwPq795ZiwK3sW6xXaSqlBfIGUXWiVOV8M2+QUkvPG0e+VhjpakWmt7bVvyqm5nS2KUkzhj87
RMuqtCe9NtHAR9cT/KRiD2UxA19knN2tAYdvWEBU+znOejerbaOp0QHw3i69FUqw71slNisNw9io
T1eCaSthzlDSjfrZaQ1LvKGKQmKEuEm6WXFyOuj/PHkQQ0WjT7t1aRP9y4CgkN+2wk7Uw6MuNmo7
ubfeELNHLMzNHkOUNr3NrtPOy3zP/FOPjW+Niqs3wQ8k6CABwJ6s9I2MLcAwVfnwCi5S9FA0m/P7
kOQhDItFxIgVan2CTK7e+TF1N8bf9gxc9Lo/FmDzsTM3h6vxL5NkbArfJTnpXWksewF+HfMeGvwE
1LWqcuqEAFwVDhUBAJjTFCX7GPE/ADyvHHx+M/lSe//1peRmw8W54ysbTg6PoLt0cycRaW76Zb+/
Mhkl89Dn/w9oUFDx1YXjqs1NFufSoKI8BRR2ia/yR8vjMbnnf9dTK+GfLu9ypgC/27A7Uf6ZTdjo
ORSUWK0m30VLA274fPm5ZvvDAMrwOhIsGM2oYGfcFSY4oNNNuyFhEsrOqiW1/sroxhoaczGgtTPX
jqdWXGQMRiXCvKU4hvNYvHRbK6xeAIrzDe/8VhgW8zu06E3KVd9yaoH659o08lD7heHgEi3YMm1f
jjAjDkbevXNvgamzAX2DlQYd/FzthW1MAlQVZCvnhgO/s3dJx+wSa2WpuoxVno/JaV1j25u/0t+q
XRni0IC+61zlVOxr2h3wBz6zsg4SqnrSH4zFnpm28143lbnWkNax1aVPyceXbCb29rrjouReZrdY
TFhfKnZjLPs7xrnzN34zdFuYTKZvIf1H0KeoEx8B3wAPa5zrpM/SYPKQzGuHRKcGclXYk8CsmVUY
g3dBQSsFkMJxS0Zc4G7geUYG4w6ReI8+rdbH4eX956RCFTy9ikG2b/jn/ql95jh1MW1uLAzMMQop
VB5pVIpeDdUCTnLIVWDMy9NJ/VG32sZtWn6iMhorJXYD+8c73a6JN9NRJ4iWxWfHi2s1qiCMD7K3
zDiP1CtKccd4UATw2W57kQGKiPeBPUalCdXB9yN9nAqQMVK7d46IHMJGFg/pXCqd6FaZWPwHNFhC
6Fyt/F4T0ahIeeoVFhBh1jqXgaG9+q2jQcLx9n/eMsGaavUZ7P+HF6xhV8e4SUke/OQBd7k99bLf
Ivs4fy8mGA5IT5Ge6nE0/ka5UfDBr85gJWzUKXr+PaP3Oi9txo8dn6Mj3y+EvqzOOVRl9lJWmbDt
akBIJzsLn3oESq/PZ9WNQJuSLgWNMtS1NP0VWiEDrQycbX+p9VrN38DPQ93v9DQAPqM6s3Hn48JZ
aooE2H59jWEnCJKm5ymvDe1keKZg8YNuq7FTN0E9Qc3L1F00WKWi8ARcJ3LWZ2tkFFdEWxMmoiX2
Timqk9HqG60Jd9LacODFhsYUMLJFnC8GTsNksO3hndd6ieyBwfMVVhQhoE5arg/wFEtSsNFF4VPd
RE/rXOCCeccwUZOfnHCFJVhLVz3jvpRErfqzzisj4T/B1xBAoB6KPIx/2fnrjd3S5MmsW9W5+krg
KI99w1/AHkpaLLYv3dydUuBAZ0l+JdZ6txyhbWJ9OTW+YXNJ/XdPO3vZRBp29kmJBNGInwRj21qQ
cLSWYG3E9AZVXePPrd4TJI3l1XC37YcYG8efIlUQefahmeIqjyb0KDJsJJxVHNrhj0ry2X2ookqP
166AT+yd1Sfvj+J6r/PPOEtXsbdCi5QoVLsAZwVT4B/P2Go9MgjPZ5c1NCAlkcxVGFdrDTHaGuoT
cS75LLq8KTCJwNHMmfoMbSkMFyRLF4ItOXQYKjGWUU3T0mrpsf8nWLVhVLFSbjHa5kgswo7y9raN
l1iZvm1ojv8UlvQFkh011vEo+gqatN+jNIgOZb51jUC/1xnbkYaR+YJQ9psRv4KH/iQ4v09kqccf
XQzJtZabJon7sH+RG7OzymPPSHhSqFb7YTuCUQHtFeBzrwm2Rb8tOGlN1wOkT6voeocQ/ZR/4YVp
hmbmqr17NZr4r7+fmT+FpDHmKVKX5S9ZOf+UcGN1iJGesp4w8zpWQG7hwGlxwz6gRJ43pb81ZZ0w
X/Dk7vV/mATZrM6GPRNjGOooo4qxW82Q7DyBeBZhannpxyRwfzM62csIfNhlutJQmLWIASjqKx2W
0ToZOWol3+vkfHpY7SIMY4fRRxXkc3uCUiBsL90ffTHXVwam7UWtNNO5PmU9mOHlfrwQ3FCmJl+h
MZ8arjg9X0eW7DaR0rA9qrx9XWR3aWUgqHmSBK0L7ZPD0eCTEOVJ0A07pWKjpuxaTEUE3s2urQqC
Szsn9PIho1SJUmc/JAEhmANgbC1d+EiQyr/9gnfTnT7OkZNtT0/ogqgN4go4OKR4tLu9gsybdPf9
YijPR5nq9zq6g8LdJuDpAXVSVagxvKweOyaZ5Fte+PHkhWC4ANdsP715GbIS0JHekBUYjGPb7pqw
Pn8tPm+ZrN55h/YntN+wYI46s+jVeMcK1vsCrn79u/s4j0Czs16G9I9VdZVi8Olh9D6blq7kkDYu
u7XmxePPpYBlmoXvcfMbuiJin62iJKYMvKvekS3zkK0soPNctJN2bjkn8flNHVF+uRJH+rEwO/mD
s74DcYnw0UCWZhYlLEblaYHUg9bpYlBA4Pe7qg/TuHfprWwwaV1UmjlARHvXcXFzG9uDtwHMWkFM
+fQGpUuAkEpWY4IO7cVYp04vYFGRqTNQhKsUoMPeQE+tdChWvv4/Z42rJsBxc7hcOlPUvzdpz80e
YU37/zcW8fuG3k1jTVaz73D2jvrTLAoBl3lwl/qJOkT56V60tUHSi2JtFgRhEtveTF7yemMkOCrq
6Mn0sf+jBw55QuljfzRpb6PI7mPPXfOAoSxzXCakQQt3fBjC/JSVzKkRw1Z2vCs/DnviL3Qz3e6r
W1hzK9Sv+oH/WSFJdkAcRrduroCo9DrWbyqs1UE/+bn5X6C5zzdpz3CoI58g9MtACZrwNmAW9C6Y
4wy52sCw8Jnnf98CM64+rBLnhZcV03eJQNi5PXLfmEde81+LE593Ve8qIa/O8GC+yUZ7Pq23LIPV
YTUMinr0I0qQGMBbhvdDX7vN3zvgoWbUCndRwfSmhiVSFN0NDzo0GinNEphl6cTCOCLIVSxRe6Og
mtZEzT0nQxf7gWvFlsiOB8CqniTeynNDKNf3FutuYBmgZjK0EmoXoi8PXI/9ZbJ2aHF/MirLawm1
/x5VfSrpkw+ma5V1rVXlDV6t0afcgWXOa5OuYbfTnVtHbQlseOD9gBco3qetaoVFYD1fZhSoqojd
7E+pr4jsg9oNQFwsxBAlwu3AzPyvqFS3B7GrdGt0KJYsTkwGCAWEZmFBt+7BJVOqKAckrzYch49f
lV4e6mEWB7a6v2gFTgDXbXYqKPv+L3RoS0CS1x/hIz25eLQROJ5aaE4jhpdojuF/sBZeTSK4H7Wp
SKlZDmjNTBX1UhoMwQjPt7fhD8LtdGX/LAAGP/HkFrzN0ws9eaBVMQFWqX+rsoJV0aXLU378YYTU
Yrr0I0Fy0eeR3cvSfnYPX/bv3C4JHXCjixI8BDDIpI2BCU6yqjZ6rGe2S5Y9Xz3M34IH43aQV509
DRAHC1bgCiqEHcrlFHG48jvyTRW1lQl+AtFXh/148p6zFkuKNGmIaHq5Z4NX5REaNe3tIFBW9rRZ
nkjbqmGINn20FAs+6GVQOJojz1XkF1W/fnKrjH5a9ZFZs+YmjLsJDK/wmPJRSWkyjAgcQ41wjxDs
Tt+tye5DPc43mcMFysTSLPgQnfc8U4OE8RVvdo5LtzXhdN450Js+BvOQIqgpEfxWH9bnqp7ejDmf
HTDRknLKCtQxUdgfVrTFp4tOamXOESO8kWSyiR0rkvhRQRAzAY/V5sLYYEkDhO961UqHS7Qnbh6Y
BHwvsT10X3qw+VXvqMR4HJTitQI4R3QtMyPtT6HbsFyKuo8c7+bVR6tAbQFKEH2DfwTvER05fasG
unxQtfR58P8PjoVZmck/T/rwmr31nHRpsPZUA8AqsHMO5YrIHRdp5egLwqaIb8KQ7XgfnxL7RbmQ
Tv/9+EbrVje9qO+qnoQKu3fDjJI0HbKNkfR7kPW5+LIhNoZaXXijGW4TGbAzwpP8CXYg67b2x8Z5
z4nxy0yL3mHSVw0eYiAohV276xN0UV0xjz65zmaabkUpjHRYfehmfktdPJ2OWt6RlrzKPuwuCLUB
n3IDfl+TY8cg+/u8e8vIHUbqbI1ZHUybrbVtssYMgPdETwQZBWWOvwYquIibJPDTWcb++bgAxkT+
eCe4lcE0DjDQ9F0PhyyS9zKa8MmCQRaQGc88DIeVM+NHT2GMo81eg0pQZGCMYL/jNYx1RPD+l9mM
X/gWtu2gcvYp/1DjEDIr2pYT84O0I4DszFIAaMgxMrgo0WpxjoTFrbDiTCa9UjPT5Nf+wb8xYTeV
KPub5sJVrmGl9+hujT+QKS5ideOxejM19XgwQ9LL5Y+uKxytxdtHauP5Rn1cavYRQYcleCkyhVNm
JoZMDsBZxaQJhGsZJbPHCY0NK+/KMqGr2n5NyooDN51BFkjNuL91Z6aZ/8WR0QCUxg5fgtrA0Rpt
k1n4yjDfIOrs86ic7EE4ftqAnDHJmJuJTw0ahJPsR5v3YZARJXQ95VJ7NkKbMxwwCK+bxS1kpcM1
lCSlcauc5v/8SPW3uzg81ikDXce9evpMTsCsHyg1aFUR9yEIFU1KIDBZ9eAyl5Q6W3KyO2OhlpdI
fFGX+QUN7Jx/jurPWO0VOQen6TTz4VIgVWHcFU/yJf3sk2MkI1RB6UfnuBSWG9xdiDLtOVJolTob
Kk78qyhzfFJ9zRDOU6vQHG4D/mCrXwrtMWjfB0n9LHGeQqCExmfUa71JlZyzqt386WX7yK+0me4k
n3SuD3bOsUTec0kyPYpCnTHEz1RPp1mDCV7KXuuYigmgK0Jhx3ggrbie5/jvloBA1SPCyAo3I48q
tSAZ1Cp96Pcal57vhJAHXfQ9S1bXdNN08ZsbZ8CTswHHsOupG3Hku1BGGW5RQ+G3dtw2aajMtCPw
YRjh3SwOHAokw0EXyE5JEDn0Q8yVsfvg1j9RU9Rq/JOTvSi+rwK8WZ2trwTbD1yR5qO3GTVvhuXB
/GuHH1Y3+umEgy/0LzpHjM6GwosyzCVpp1Ehbu38Tm7gNqB7Z0DtgCFjGct9PIGekilEXh7Jp+kH
ghewbzhgMr0jT8wM67y0W++lW1FRpx7WZXlTCjRMQ20/o4/2n+0Nyw/1wyiOr0B17nWE2jPILFmV
wJJ3+ZwQqCiQBcH6rZuJhInT0/KDY3ITpYVx/ZrrVQcfuiyWdzfTNdqSQipyJFPs2XSb2vsfgsWi
G498sYhd4QaMz3pIHqJMIf02UXpa4uEQiAM4zq6MTmw9O3rYWqKGGq1Uq4uE+k14A/74xgAIQnQZ
BqwSY4B/yG294vmF6dJF3yyi25IuUhfDj+zG7Te04MG46DZfdUqAtkgKNPk6y8e+LMSj+gDMg2bm
vLN3lCf+3nimSG8jE+t96t2+LF2IEwWpK8saLMFchNDg8SG8kiiVHxnviYixpnoTDdLQnpsef+7u
i/LCuljwct5EQTcVgkXjaWZOOd0LwqVqO8LazDS1WWKVR5nL+Vx/BY/czcM4eavBSbnZg+HmbiK9
9ls2r5naKe1HfiMz4hHSEvyHcDM5S+hiyNphwIxvcq3odxCRkN5z8XqBDsNUEU835ETni0vq5pCd
ygFRg1xVoAG5Pbc6W/6/6bSu8xAfZw2JPB1VVkphOGG9Yd4abwC2FJvrYb6SmC7hSD4tgO68W7uZ
+5xTnD0Z7jSglShq+wn2hMgVsoP6rG5Wjn+smBSWZ8qI5G0TexvJN9CJGfYjo4qw7fNPUAnfnU0j
R54fbyh4TiCA/RN+ScRsVGzXtgIihuZKZW054oxhxLgSJG7UYoa3oRDKAMTTaZ0hKY+bqLsN7z1s
tpAaEq/UxteEeNs1MPb0T43iZcQQ02aYGtcbvo/1EL5+f/pZMLW0XJhBTROdpYLRt8Q+MNjePn4f
RvDxU4Rzp6IvEA02qzfyX+yCsyhrPcLD7GxBlFk3NviZbMnhKWs+PnlxRoZfMio9jSr28AOVF2h+
TLj0inFKXqNM0FnujtOZl1q3pnW7HE35Ojdte9/NdnDOlFIMOeJ7YXOK/mYA3heKsgIg+sU1AhDb
bl9uQ7XEKby2D+BFmazOvGBj5a2nNFpFdw6fOb1/sO1vHeCU1nJnY2QefkimRNJMba1iyYXLY6fm
KGEV6d1Pn6DZ7wA+8aMTVLsn87gaDUVvRvTdU4XBWOgJV6Y3jy+AoEteqtLzofqiZ61lmlF2g/uP
zwPKPCqgPOxXrlArJuT3m2/y3ygGsPQXz7VENrsaF0q+JBzA51yk0CfUIIHdeaeihc/sdLyTxc7w
J6sJK0TRO12RTxSj8RrcP1lOQl/8YruNCkaV76gqLvlepcLCoEg54B/XP9xHet9qefKMU9OYVJyh
G9eh2hxiNgGmNKN2WiS/QBQWFgV2QIBWDRcHcPGPUgv0frLS6Wm+63xBKONMLOShB6j+RZ55wZzb
dTD/N4zn8La1NgFU06J3vIydhB89BEe3KNRW4eDp0kpgaTSnjxjSPx2RVSyB2D8YjsyQuAPwWJde
ns4Qyc+dh5X4OWlXuPJMB8SSk12nYxFMwKNq5EvU/feu+L+nFrBi9y5+NBdAEcDHkBy7B3zgJnD5
ItkSWrwxWRzZ42niJx0rrcMmPnfgfKGV5wToGpCAIyNxjXvV+ZXVRbSyUeSH+reFzH5NETU842eA
asAA0F0rhCZsR917USQ4p732Si/r6eID7xAGKr2eqEhhlL9hsYfUlDqtQrTIYA6urmkn9NmkXcwf
E8hMGI55JkD7dz1trFvgNkvi9HVA0p5upwvlPafxGKBkZCYFQfFBAv5kVZ1r7zquuOt6CRiJDb4W
rPBDA80BqhE2TdDNYib6HBnAVtCQ1Ts6XCcbx8mTihKBgtu5ITTYEjqA6NQGvHijHF03ZMzn/HXU
3ZLHtm5Md6z+BEoCEpmrJY494MNgI3wrhOw201p0vjTtcgh3qHKiTgudg45uvwSye6laQQTYvOMj
pmq2CWkq/lm2teZsy0KSGzBT/ublUchXVb9Y8ft1+A+AtiQJeI24QNxDWCQo+eNWbRskgXw+vVJy
qjX072f/GiVzp4Is7vpicneWYJetSJnST69iYqHORr0921vPgduYhsVLwzSl2CHymUO6kiLn9kks
pxJnAIMEs02CfW0Vw8HuvMC/mpHTP7xPclj1EjQ+HcKlA7ARHy8qcr009dW9MlSmw7ro2t8y4LF5
1VK2fZlCT6Pt4rDuS8cT41n9ezspHfgccNkd2BWdtOVi5Fnv+Q2S4iWa6GLEdysvemTraRz5XxUT
7pCSPT3uHHGViRlE34sHAsh9r3JtR3siuAmQLTsxdoLmZCaxEL74pSmbFIzSzONgp3BNhRDiZW/C
lg3twT4K+W9zFzby0lezBdd/JZB1xWV304OersxMfUFzIgijaEKj7OzBSvBt5yeShMxFdaOyeB05
AzkfrqfA06NcDdYNuSkDHgqg6d8PbLhbuDsros/gnY8KYV1bO9x14tCAChQTO+d7xIQNWViP0H2s
Vj9xrRNfLb+V99TfNN9iX7L+mvIzB9uMXSN/HAuaxgZvplytv4FlzvEvwK1CXtGOf9jYfz+1csfb
+9Vvywz+YYH+0t1GuusUyehq7rIl4T7jO+YciTxeBOYVFOECWSy7N8UdCp3Rol8fHdDLYtfRbtXF
WN6+APXmsC/9xoEZpXWsbefhvlMoAaDQmjmzPRnthkIm++wrRvmT90ClZi3NhHvsrpBziGq3sGxP
1bizm52QYsKiyUqCGfSkM37SsEVx9GaSp8gGk84mUt+R1MiFCRKg+xOyAFqOLuwHHwj5e7jqC+rA
MRYKk7QgKSdHyAa3BtTc0s6/m+sPMGSYz35rLkGff786feNEXNr808gPDLHo5TKRnqBFTgM998I5
lhmaEoXBRyLwHAKZt4waJk5bHrZ+VAEYyM9PzE6qkRynkEsuw2RimajHkhdvC7cv2oy0CNS2j75n
IG1ltGbV1NmMqzxwtxUw45EurLvhJ/E0bxGQ++sutoRREA5aGB6bKhNRRNStLH5s0+Yfq4Q96Kd0
Q17ubcjU0M1la3DdUnVm5Wm+SQtMMtZ25WqqCFxXSDO3Sy+EbdE7t2U8gWdZoq208iSyd8FWdTq8
alGOed+z3JNqqbSBgsyjHX8dKxPsVm2vSxyTYV5k3ISGGhXnmJNFl6mFqMSslIzhp+UrcXuuirJq
Tc4GWh6RfrbCP2vwtWu4LxftobDVucbeEtWB7Z6ZRtRK1q21f5TSb2yCXRICUYrjC2vcx42zmLXS
ebIuOB4eyVlMYt/K8wMQn+SdBHKB+aQ/rOZD2nNsRw2TqEpSVl3FCHW6Ws7RqY3vifVwWOEZmzld
M++xE9MK50gZW8vJok65aWpyu5XczTtMCTXVv+oiFNz6R+TLOlhAiVDhhhU0G4N5auYK35Nj9WSs
GHBsW7Bia3t+nDRuwVniXUXjoPJBSANVtSjzNA+53EaEbWMudyL6qZPPHOVsK7Thqra9ZXTSNP/E
I89bNm9KarvUZ6UD7DitPJ8xXY9CyaNGEYbuuOQ8cfxV3wkk8H4Dk2zhXUUC/g7zgvj3oeDLaUQP
b7mcOvPFIZ2U9/WtKomr4YTvPYvH0FtsIoWLEx3Jc8QRRFFtnq16fUFSoCb7g6TML6ks9fQaTGcc
ycyaEjaBFlHX59x+jRGmPqir1pG26mhccVlUmX3zF4+m/MntcbW5esQkrJUeCurvHOBLOE67eO3X
5DYPR1Yx9i9KeAAR9O/9JZt/JiirKqUsaWNtybFncDXeR6mTd6mLwajdrBr6Tl4EAH0cAeANNfKb
ugs5NBa0IsXtP6SYKOylVntHMXBY4kj4MLb4kNJucFN5+DVxv0Ml+h+M0qYFvbl87saeVEs/AJu6
zkCeXaIUmJnMW3fRybqEAHFCXpmvUdyo6i2PLeOr/3YTdrx+4hkqp9pW5ICzFA8OTPvgaWe0EFdk
nqboYC0MXk9DsA/LQq9xG7SEasBkXVTsx5uVSZvPpisIVdWpoQLtnmHecIHFW+kYEipV6l4Jq98t
3veCXN5PsZavK7ObiETbUV5Y58NOEoM7N1VbjBVdMZe6eSn7g70bgHzbJfvFErpN3uVTnA4t7BV0
Sbgqm7Oc1/w0+n0VbrmwtenFkoCzL0e4a9Y0g4Idqjx46h7zESB6/Z8vwtZjyyz9L5KJS9LmyEyx
d0Gb1bmQ2Af8UIAcLfQaRroRYMDZ/C++yXTm1Vk/JxKZFeE6Q7ijbL2Ip0Olf4AdxbhNHDR/wi+U
oTFzxqJEVCV8XReDxJYosYFYmllJkiMzkTgq7vpHjRB3UP54yBm71AQZvng4NVXtjjGTZGsnOORQ
tz2wNLYX5aEvlDtJa9H1dswn8aLGR5t4AbjWY8n2krpSApqsJFRbY5aniFTlBluaX4monWsfkFWF
qNuJD2ff3zC8UL0xOy7a66xPYJSm0TM/4tjPiRiDZZpHh+6T88uIt6UT8ErXlj7U5wQbBLJppjE6
KvLWCS55bbIr00pR4nBPURPC9NsuQv8jAjp1PePsvAM/C0I1eY786g4V4z3k+jk0B4b91wt9HNNW
dObuZYZeeER+q1RZjjxEhaMCe1bFrd/DLoLa7xJ9mjlbbm7rZKHB8VI8Y6PKga2pT2bij/CoGxJB
iJY4MykklarYFTlmaGvdTzN7A2Emh7OQ6mB/3pNRYV6MbKlHB+/wZahzqD0KlgaptZz83DcVMvPm
WRucch2OUz8xiKckVoD6N/dhjOSdlSDo8PSqDZbkLGWP1lrH9IzWb8x+BgfVWVkjnuFAZihBFQB5
X255ofxaDOPSJfTuNvBQtEnyIRPiYXSppOoqaU+ZhK+fBNmeENPyQB8Ow+42xAIhue5qrCLBnjy5
q7voKFE2nLRTa/nra3KFZKJzH+5z9Zr6r7tnsnItBRWE84hJi1lRPOktntdN8YtS92IogSxladsP
zBqZ62qulWRC7rBLmCWjjMFM6DhctkqNRToTnbFhIM9vVDKSAxbNMC6FrDm0eTXsSbKEHqMxEgfW
Blrs0ttQ1ZqSlxSJX5TPo60zyLEcGco9FPyLkujBLWwfOGr+Pw4tyJxhLKm6z8H0llQVck19Yzwk
LjVqL03quY8tVv8YxSRUM4gPeZ7OI2f4wmFa0WI8ZkJJZ3Eu/kZ4+mq2cJ8WA0lCtrgIjI8rb83Z
0KXaTdpsW+QFzUJkCfSPiZhaWG6ZzUfoNqNtPQm09hM7/cQBqE4F96MuLvoZ4fjEE1JlcVa+RuPF
KjUhhAVw7cUmXmUA7KBa9C6rX+Jq3GEIHj2MyIvpf93JhSr4VdEbjZ8HTCNoKd8bQmf1CBCl+Snv
o9+aqFDnmSyqHq0LTIVHxIZHmD5Ln0iLl14zCEkZLuW4wA7pvqtyw4KnIjL/vfVLUOAHEnilNYtd
gjXd/Tz5+xTcZIF0hMabwndnFVk9XZXLlTQMVyd/9co8YUMOr14q57GI8VOMsEfWct1UVrQZ0YML
wwkR54MmjK68qO86oC+1LQXZ4R73BZXAU/UBRU8c9dBYzuBr6XG7wwuNsprpUE8lJFc+kN+PvuJ+
CMoHlsftRKBKNbUt+9Nx0CaekaRmqrRGjZGQYit5sSdhHEg6HzET/Kss8Om68WBz1ndbJeprWU6k
QjhR3Ot7BdnPEOvgDmGFtcqbgYioaaZE8RZTSFF2Dpyq11gdtb/ApbYHzi72PNiLKIHh367uZqSt
QhYaDzpn5Rw+H4ZNhPwgPk4Qkp0lxO3RbOf18k7fjIU7UAvsGa4wWpqM91sHLFvWJP48ZJi/M3ts
VOxhmTTSTXzJ9wuumtI91yv/An7HFrMP3W3aH1MImekWeJg7WHM9tLuTaUVuqL6gVMl8ijG5++0l
LGKwkBmHf976QHr+jSOMAgVAsKvP56JkbV6A9nRiyfe7SRYqTdSU3KDj7VZK+JmELhWrLAzE4485
PFoZiI97RPPowSYU3SMfcRwGwyF3/G3oniYYtqn8MFDk0Ti7OdV02/ODPf15o2kKoqRjl4ySiuCr
dM37cWAwiOS3QeIhfSO6RUsB7yCuzFXSLD9sVuZV603LFOIiSDaAqKey+x0B7MllI83JMXphU5Sr
TxOLxgr9ovhmGKbpmStWf4UHqQsBtOe4W/s7oSFtQzdr6gkZs0vqJGdFvwSUN8bLZbdkZMoxrlsi
eKEkQWB5tSmZpxYAwUfee5+AoBRFZB03Fidz4mVt1rGGofjD6/AGCdDxdg+c2ZY16r2rcqKW5swW
+VCWs8Go4bGWvlegrx3vEhDsNMvwVDSRvgG6Ehjs5ya6zRHdLAs3wDWN2CAVFK37zYjF3pJqzYUV
oEdKHHZXIP6VWUHqyLSnIzNGv7DVz2BVXee56XNRk2ksXCDNOvPMTvAWucWq+dsjtDGPLaDtspCs
EKVSHSntUASCG8Qy/a96MQdlc1J73GZdAtPmaZmuTpsTwgDxeFdJT02b6R+grgD3pOQPg7YTvtRO
XMq1mwD+KVWvStVmtEE7yz9b2igFFPy7/YgjY38aV6/cW5KRgo38dUkskj2r+UEgVrq4IQ7hgtY2
HDnYvear9gPfgAD9bGyBgVjABI3gVDJsWWgy8VrHWJ769bZ69YjCJ2oy0KMOHKBUAIoZ048D2K0Y
nGworJ2hzpBFGtrvAVUGYlIbH4fC7DbyV57vOUr92Y0E1cuxGaum8GaUHpfF3E2jkwR9u87m4dCO
6OR0NPgMWivFc+R54p/Z9Ej8L+9cvAxxYQ+AFGo+fdXo7LS6siPWxz7i31gwMSlRBE1ruxKikA6Y
CJ1ERR2u2ZTdf8hPUzyMj94dYImalfpnRztqf4gF0x2CAxi44UI9orHP6Srfty2Nb0cz8Vevk3iI
GW6ZrtAa+j44iMc82jixGGk35Q+2pICuP9j69vasFdoywI5uybg6aHstT9dRLN+rxMk8Lnt77SfY
VS9HQW/leuBJNG6pV06xnxAsxcCTKCbX67Q8GJ+3+1+iScYWEI7d+0ou49luAuFpoLwAOaQ3bJUG
byD65D29J+wuBdAPMU06RO4X2eeI4sv6O0LB2GM3Ccti/k/tkC1km1j2v/7MpT3cyNWLV4laQmv8
vFgpKLXFQycERx8b5do5jAk+XM/ofksU7S/NmW3V6RNvQxRXUV+71/juzrMGNQwhvD+vJPKSECJM
5kmAFFJ/1YJDZfbuTgrCY9KA8sozmkRDRXrLJ0Q97sWjPifdC4BXK4XTyA2rKJUO1pjabEkDcgNE
AbilCIiP9I42EQ1nu/eGVd8tAqiXgairqn8pKFdMzUttHWjj5TdKJu6H+cKRVbtqw2E513XApP/g
fy2RTfZFcrHoRoR1lwL+RIDSA/4C/vkZGOJ3bxjJfBqG4AqNHFcYf96/cyJ4hkITpExi/lwKDd2d
URUWecLyG7JmN19X25IVb15vy2NYrE/rEuvywXzTtlf402p0CFI94NRmWV+qHy+Ilx/cn76r4K7A
RbhKcmkvO5skdFPJhe8i+MBPhfakdXPo2MnPw527u6NIwwifvgPfk4Y/1ETX0D4cEarCJzQZ4HJH
hfB051+/M4/CGPoXTpwn+/Xamea+Jin5h4EOv9zeMELIMgIG0FrACzcNQzb84N12L7LCdSyl/zgA
1nN1nilDni70yWktMCjc38gJNwl8+KX70xKFF5nRoo2Nf8HcemK4aTEz7zF1XMV/wYgfrNLz67j5
GCyeNMet2cbC395835KKehUz3ZbYXMbhxQwW7TH9T7qBgNYOoQieppCeGKTITed0RRybKKO0TC+k
wXuZQWbyrpNzuYupIRRMw9veM3UEbLoh3bKNkdctMhquSiLI+PTRyI+w7OTVF056wAQWAXhtCN27
Cx4APWM9Jck07HDVcV7upPHHgqeLQvNk/1UOrH+/a0r+Nsn7TgR9NpQ9gnje7jiEAabBe0VE7hSK
G11LSwYD21G/2L8Fi3Wey2D+otP9bEIkpUPZB3iRGDy12cjExDW+VOzjgyfPsRZuU13y3kXzXh/P
mXydMGxhG5exoOj3p9uFjA3t+C0UEV6pItRAxN1qTLxfAOp9DJnMbl+zcUPQbvkSCZ3mHgV4cBTk
uMwsc96FKB/Sh9xi4phIoRnwmpmttjJxzwON8SFgvj3ghxODLPVlrLz/RqFgAquhPQEcXnothfLT
9CkIkKBub8HcHCOjyMfD7GZCc4U3SsJbbb5y765+iyKyDHkwVZGq5nJi3mRhk+E44sLjY8S+iBN4
H8pEhIcca1bsPoCbC5a8lITIXsS2YqdrpeZW3dzMJGmE+0fKRGuMrsAPDOHWJPOT5BAcdBNQTUKu
xCawP+vn8kzDK1ESMX2bx3Kslr4Nn53KVTVHW92ymMSsE8Ahb4+8vXsC5X/N5z/RrcUJ47PqsUyR
0GWygK2PPIQ4dLzhRdwu6K/KDRe9uO4mH4bVCIC6L+ThnoL9yJ5IYaxnxvYLRHrSWzAXHzeAxbV6
iH06u8XyTHPvLVKngFWr3yLY12+oikSxp7XzHfHD4S6eq1i8MXdjiwVtc66lUgd2cg9X6/4i9gPW
dB3exS0ps9wDDFRdrBmd49jOF+0rl1PVy7mXjtIzo3NZzA2TAddaUnw+aFZaHdL9ye4OJ7J2OT0X
Wcr7Q2fww6uWt7wEli1sZCRjOsj++VjJ3JZ6DWA0vMmMcCxDYsIJGrdo11aCvDKjFtDLQ6Sb14TG
W8vd8nvnvkmTZoTNBJ7uBPzVaHwWIH+8AFXGJZIW0PbhSwaVg+qAALH2Dm83J0x1MAhDz+dZg+vi
PI3KaNzHl7mKne8fLaOPaxVY1K4vc0H/XpLaYqAsNsbNyltxJXx9tv34wkea14HcVkI65nYAf+ey
AOBse1tBC19QleAoYxhm8w8b99WKTw85coQAkxPQZpODZdX7g3PLFRSVTpPvi+7WJ7/OmAY7cbbb
KqEHegsEq8cLO+30BijXe0PCvVNR4Poln74F3HVWOKUowwLrxKLGKb+3pO40DSm1aWN2mmk/kfNA
Nt54r548aL0KcKq3KHhAROctShD9ty1rzAQ/UVQPF+vV3lpO7Lmvs0OwgJAPxnPnoCsAKHyeCUZ+
zxyHe2doKY7wHoWqe+EyLLLO/xdKEluFYkv/BsctgVej4GpMu4qKImWV2dq8pnlS4EessH4pCHMn
TK5l3YOPObMSQFBvMSI0bkwmpN8pmsFrbDkfc9F3ylkO3JF4alErKjQzawisDh8oytG0BevjeLNC
VKMFE7K0L9OS6q8r/Sx23yvdYZnvvOBXZh5VuRP3pQ3VylN0c48nBSUaBUymcZoJd6/CJXikj3Be
npwFuDJOByMrlLLQtumwS5cWxeo/PzeGOSWv2yoJg35ik1TVagDHuqTL8H+T31UBeTPLnhxdBzpV
tk8VhDc1FKT3tmNcEIYWQMQQoAQc/TmfJe3vi+3QUy23AB4kSl34+y9bH4icJeFqEFiSxRTOeY6+
Wo7nay/bKa1euMKJRkt3tzY6yEFRrAnY+TtIRth5t1G/RTAxV6mthP5rXU4eGE+6cPrPYkeB4MEM
gsovMqcv0CvTakVdqNIh7zYJmRhCNkitKnPI5OBNKs2CE/CyoeEib38cuASh6/GOrjanMm+/DhFy
ttzr5pd3fAqmvOKqjursJTodPssl/zUn/UCSqObCWad+A5f47VIrD9WGu5dye5Wq4TK++6UAfcnM
n1ueJC9MppBCvSjo5cT5n4Hd/D5BQka5xMaZmpe0/YY29zk889EuvYhQTyrFRohZnD32vjeZLnoZ
v4/lkRmEe6BgB9WvbOtgCGcyLwxWh5tM469ldThrGI8PB/QCTvcem7TJtgV/hWd9iXvgJvQHRxob
TmiItXaNzccvSKSyisHwYNdh+gBXhlfCoaOaYJheClkQJ/R0s5Djqg3oI++cl6YGsGIwKPHBQFEZ
apKe0SbCIRiOwY5l2Fuu0YRMcteSo8tJxgIVSXFftswqkbOG82x95Z/ypjdLzR01Tf41klR4O00M
JudzMrZetFIwfCR2EBhqg2//3RNrxwtyF6qLL543Wli+7PBsi7z+dIk1HvQh8wDPs+eCbljCTGlj
QvE5phTXHxkd8A3CqG3Qs5sk5nYQ+N5oDbj9TQ4JBtB4pYbvSmztVMLwo3Z4j25rj0G3In4kJyWS
G4Xg+xe1IUHVuDsJGa/hZLnj+0BUXO1j1vYWFD/l1U3R0NzthV7fMC7pZzPbGOV4b7Us9IOMhCW6
e1adK4GZ/XZy5tsN6ixWJmx2LA7MqVwaDGMwDks3W1ETxi7kfavph0PUBh5XpL5TllrgAPYLnNIp
maGJ5gHcBT58TzYTxqmIDjTGB/t2HnigGYBFI6D6a4oSuJNtXB8CVkboZ6emLrMG0kIpAuwANIln
+lQIMcP9IbCWtBgPPL3dwVImYQ31P21fk+EUROemgv6mhbHIVFdFygl4zwCQhijQ0JwqjWakZgi2
Mg8kaXAkitPXOdW2JZ4RVxhL8cG3/9Q0k250Ja4LGOAu07ZWazTkjukyNtWTvePjpxUuh0Onr/Z+
SWd3nnonr9LoblRb0prEP2n1wejJJFcMxnk4KPk8JhCm9uWDGU9rax3WifEI59RMF9Wj4LCl2CPX
WE47hpwg/+vPC6Lg8Cxx97qWVqJqTomvAVwrmRC5kIOuVnquVXl5x83xhsIwkWZa8OIErst43+L4
G8J9aPTwKimqPW7idSz/ueb0HTH3UnJfNmY6ArLFHl1p01FvlXiEr1oPE880DkfG/0J992eFl3nC
fCCkXojfrFKxI2cuYsp604Vx06h5Qjx1GirGzjsDZq3Tt3Xh82VZWKlNkHZkw+fHSmmXrL1r0obQ
pjfPXihJJj+KBKd9QT9GhkPBaItszN5YTzg2K1G9RUCCweZLRGSx6F0QWjRUStct7fD6EVz2w2h0
ny7QlQyE+R79b7c+hpA3ib7+Ld5iUF9VvZ8y0WEDFsLvxJwuXKWVA9SiIY5GuI/WMz5vqcnfIpcY
lhibiMy5FbrAYtbwb+h2u/NijkK7U86839mLlO/Yy1yW1VlEIFwhs27/CsCSpnyI4JX/ZXzZoees
Z1QnScKD1K8P1/XRTlYb5QOMsa/TUa5klsynUTqY9wkH4d3+OmGvVDIgLtegMZcWdvRYHC7yTWiq
ZTAifFnIbQWtc4yMsDJKeFlHpYqdp9MChuI1kiUklc7tNJfxecHOfVD6dVzMm7fI68hO+QvCIl4C
wypXhpy5FvnUp+gKg+1PMLhicl1F+tB+9iKIlkGQ0lyLFtvLYvRCsahPpYi5wiUYBV1Fd4ELyRfr
TFaYWpHX73bvw3Rlp/MX48xrpWLrui8nf+iQ7+z8V/4kienCaf8TqlKgX52b2kWs99damzv78P5X
PWc1zi0jAWfOdFu2EeOmDhxonmBwQ9llOLZIJHPf0g3xUNbggDjjMfwPYqpiwmkHKunYA+vYEl6T
flGsyNptWx3I5AeTfqq2ir68G24h2FFqVfHTIdiARVuHFDR6CB25jSbT9QjRS+LzWTq3rhNc/Rwt
YtupF9dna9ca+MbM69lccr92SVzkMz8Cst2buyjcN2+K++I3+i7XHKK09QBgLrgLcF+nA+1WQx+r
RPSmohODLh0RuWfSWx8ohwI/NnrPhVwKVhrXdoEWGyrqQgpQQEE/5f5WRtq58wJp2ujegNUu8/Vs
6A26dn98hMSnpG7RneGyJYfTEwExmiPsZbu4JhOg1+w0wX5F7VLG6cglmh9BR4lfopF4C3FrjeMX
6Qb67rG34fqHpE7LYazTRrDNa5xB4PTh74cfexGS5IhPvXYRa4xyDiEkvz9JYAYvd70dhFh467Ii
HVaAGnlkNnIOgOzSKEmJzgwGqKpprU3qT6mvyiWxL9CNkAQiDI2FveARPPrdoURu4CcmaPYhlGK3
U0vhDAy94B4EbxtQMfr59T+FZWyHcZlqNBfyR9diCOESX/fd/8/KX2mbeIjUq47293+xIR6Fajtz
ymBBYvtbnRm78OYyWUSGGqtoh0kIPMoNd7Wb3prog1rKvTfovzr4teDVH3KG4q07Q2uXkp5hV8pE
qRE9jym0H3YKSVJ0E7diZOcyMwWaWokLouk7spLvY8Sb+mYlu2WAMUH+Zxo5wU24djwUeQeIgwyi
ykJx/q6JNhYS/m2O8ixvGOwqcns6VDtdqzRpAHfovxcTUNJQkz5eX1RoiXb68bNUXU7H73BKEeA/
F4M6PMIH00YNN4RCjqpvW3lZ/ONU5uolsa2MMeW1P0dIYD+S1lJUSJ1kKeXCVcFeGE8O+hyAElgK
FkIjqma0ZA3fRBPPmzW9i6z528gaZPGspRi/w7ZuoJBAiO05yUN+P0XOe8FyFzrTa/J0skch9ylz
BYPsy+TdZ/pbfZQ/qg3y6cHVtflF9SbFL728J0FkedwnYc6e7uRlyiQe0dfPkgU/ZZLdWvSC2sUa
bsEdcnX/BV/2+5Isf9y4Xe8X+lgM8e3ijai7j8o5H4drJ5iLeTgEIvCn+dcDekFJrKc2B4nA4FxA
Ld8inE8BbjRKJBadZ6TYCSWRwVUJiLwlMB5UCmoszujiv4QSDuaYH+Pd0yVsMSocNTPxQqJLkKfU
aVyPjJHD202SDBbYQ6d9gVYaqPqvIAXB/YzAyIexwPeBspueeEHVtn75Om8fGOCfHaa9+pfIteP9
NsT4E7T8hrPXMiefflq1CfgIEGuOTH9nyzVpOsQQKO4pSJLXZ2+NAsDfsVZMn0AgvSOew/n570fS
FpaB7eKAq0R8T1NXrSXDOSsMWpCWkJAd6lbcZbFd0ItGlBA+tv/sOciNKT7Coqd+FaGlO1WdbMFy
xiKaeiwpwb7WR7mRleFIRNg3kwb5Wc1vZENGTJbzaLD0zmXDYcQ1JvBB8HqD0J5pM5LmIoLVamW6
aThf+fV+WEwxTOVZqnoZkN6MHAkVBmtFKjwV7HH9rv3tmjjJUz8NFEIGN3cSEkOkypS60cdmwzYL
OVzn2NWPtXIeZN+kSEyyF6vanyMxPgKw0Nfj7C6U5oW3ZjQJPjjfrU3TyrW/2XoaZQw8XmUDVYtm
5IMij5CuHU9WrG7gn529CxIQYVr0+QLn2j8XPee5H+Piz8rjX8KDXMDnuCh7jHLACDiTIyzjW/6v
G+WltdOX8U6nvx75VhrJg7VBQRigCaobodmkURG5VMfiUFZ5FsLhnXoez8zFrxApmz08aQh/m4xe
tS/45qcujHnhwfscpB1/ZW7C7D2iknmjzoQWe8EaGpjz1+S4gdi8a6wId4FScmYGsgGf6Nj83HFu
A/ssUTJ3q5krAIzYr+ZOZkEgZoedhecpfqXjp5HyVjftQBhoT+ayVYeN8i+S9WRH4lItIk4seCtU
+LgAfHjFu+VakqqCvCRRKcQyFUFmSkhTPB/25/UbVoR2hjsPAHF4fnmxkFPGTyeTOejj2RVkjlG9
6vOiy9WpFrxn7LkPhToFmdRXhUnoqyiFJKobwM/ozZCrOv/x7rBR3wlIdZem7gx6g9e+M6Oq/+DI
DaNhZFY40vNq2QSjqRa5VuDEoFt65Qv2/rJymYbw+WSxu8JFJSssgU7OZIzeFZ0/1BJHPjNPJQ07
pZO7ebno54J8cy5pc06f8d2/FoZjmQgZv8XrQsNHCm7SkE1vabh7bd+eWpC1MjYj31bxQQcrWBke
Ooc33vh7mlD7ADUtRdLUxqN5UDNiqsl0BH6mJEWNRAndpvTqkg+9wR0LlRF+/EYUbEcVQD7Ux3Lm
vYgCcu3oIhgqHnPKCe1uoxbfyr5tuCM8ar5zSw/BgJQJGOygHqrwJYKohBdR4gmmiblD3qc3SSWQ
qUpmzx6n0s9O9CloFWvX8mG9/h5zPaDYsDAPOei66jphimbdCpsa6TvSquNwLMWNLqY0QC8vKM0k
CVMGkuq9vHO2uxxRMxrfHQILIthZyoCqF/veLzv2NTIAD+s1Yj47aN/0RjTnVOW93uqG8VuvsCEv
3ayqU4fZGzlv4rZMR5MM67Zcx+6l7/3APLV489jP2R+V3/i3ZxZZNn8gGVpHt947TYVPQCsGv/gy
iWImEEcKSruUxJ5CbrfK0UOmO0JafI1Zaoi2OtfJRYF81dr+4Maxlx+OgSGnyxfJ4A2J6GkbX4Sz
JSNwf2+QCK/J14VzsqOcz9Yvzy3jtgqyTxOBecDhYFpc+jfGYNBykWfkIh9IpbXfaB9fjV4GesYw
8GCZGCqhpIpNZnPFOwj1fo9g98p8ci+nI86W31/PtosJ8wf6ADwun1cGqbUrvaXqEMSNrvKA0MrR
LIW88vDBVSJl37EHqUuOmGDGCcIDmALwCToj3ogTPNjm9vDIUaC+na7WbprD+KXP+grt+onX9dnF
qZxvAJ0vAucio438IJnHAEOkfXnsIkKbwE4St7MDf/upEQo+u8A3WcGYFN0e9bOl6kVyhkco3lkr
awS3M4lJoVdoSfzu6ZP15SuBpbPC96EfI1gj7qKDmqVMO+7AkmFa1ao6PQRYM+8CeYIgiaOzZdNv
8vT9epgDctyff77SnqBIuB2Esz9rqdFD2Sg9CQy/zXMwZAyB3my/rEccLbS6Sx0WrSjmOamhgzhx
eeuaOvg6AHvj4UKNHKEsSLb3uyvbefbz7uHhyfKvi2NM/VNep4ukrem9NDnqfBZaHHw4nP63+yCz
xmJbGF1OCLuHAkDvEGk/uYNtb7ZHByYjw3ipenrABwM/lhNoR3kJ1I98TeSOMqNceIuZB3vpFyWJ
sWnVLfvLJmKXb0ezf3X/Ehqt8CYiy1spqBik4wgxcofEFkNBlD5vurbjlxDL7QNjWkoUHlbhEuda
FWmIFezw3La8Bzt822OBxjgb2+A0RLe9Mbu0sbtR2R6ra120orkFBxEFbFTfQb+StHZhpT+0+zdf
uUHNplFTnJZpdpXHygire1CRp40C4uc9fBDwb8nYlM1dBX52gwG0eQnYgD93+WjB2ZYB/6bKBowu
gaKZfZMcNwLMazfbnCriT8nzKP66XNBwLhEq+wLaW/QNuXgSXktQcm8cZKM4m99w+GtJZ1pXrT82
k+nTowRa6Y6DNKr/D9FMVQL3geZowqd8aa1HN5mN8H3LDeIIRKxKYLsiGqrqcw/1fQJ2sJxhpvZo
hnf1A2XlTHx9FZS8cJ2+tQKnb4MCLp3jpocUMY8wPfqS0AKVhwQPVv9SWTOKeksSg/8Dn77cMrwq
hGTMYoIk+GqQZko2swQKD5GI7OCTPLSC56tqdhkNv+npyeDw/sw2HfhZRarusatGiZNm6LhfrI6H
NNcYUbNcKBJZE/QJjgPsWSPRN7w9OYa8xTjZveyhPBHxKCTzIrtrOzf5JQXVO4pGdR4zaiQSSAVy
15VDqgyNgPBfYEORA0HrkQcgUT4lNNFpVWehw1tX8viHknWvoWC2zcmJ/Qs0JF5613NV8HQKqMIi
y3c+1wsHDKsPPBpee3oI/A8HFAWhrufx0KIlHi394j1yXzBym/VlcmZKUWxqyTsExZXhiNq44y+4
JFOR72+gyA87Qx+R9g4i06XekxgLCo736xal2wihhdz5PlX52lwd2qkz2IqEblElL+d2P/F3M11x
3iPHvNOSM8FPjqktg4UxqWdOWSr5XjJ30LtCz0KUylnZERUR71/VV6PJ5gTxDaa+ZmGHVAf0W8wx
ArzxvMGw8V1DGoRVqOyrh6U6jSLxZ7N9rkKu9QxsTnBeatu+NoC/TEdE/pfKqzikxDtTgmdHw0Tg
tfKcZnj1KcKf3+7sFTwqovn3+gH2TSFLrmdMLNvaA2iSR2nhN6KiQgv7acRaFM23u7hg+u56APDr
ZGOW8ZvHhpEs9xU05dh74d5qHE0tH9uNw5J+P+h3Y2h5H4P5Owy/8oGF68RrjFavvQQy0lIPeb/G
c+pHjB5uF0Id1bLvQkMUGIUAHl7FAZgooHcimJ3FJTZEx7+8oZQ7eOKceCh0c5FKUhFxSFtc4m9x
16IJnceJPwSKHzR/8EktpfKE/C+kvFaRPRIZC3iNMJlqGQIUjWWeJow8jXVMIk00EFL+x/E8t+R7
K+Mrm5bm/qgtaqlHm5YMOTOLuRYqwVg0pEgqCbivwE0OZMmOPxAy8wEcNPWmmhDKi3ggG74rj4LB
puFEKJnGriRlcCshmMztN0FK4+sYOLddgYGI18WfQjPWMvLlEIG5J+g082mbu+Sn/XTaM3Djb2qc
fZ3FWLMDDLzP2m0LwUHak064+PXRDekT16ARtvoR8UjHz5UJhc1XMOt+d1kKwqGuvNpQA9gmKnSD
3EK2TGNJUztsZk7TGVYC4cHW4h4LHn7tF+LA8U406NZ5wSzCk9rndn+OYr2/zr/I39tB/DLh9NYx
cQdfPMd2VslAufTbeSgvzCIWOSZiLt9mU7jrHCqOebArJFHawcA9FS5Yci5htxZSoBfjpHwD3RK0
jP5XfmLqpN9QmZIDbHr6bbiKapiyvKKuixGxHJ3tnSF6nCMpEunvKeSitF9ttaAss+mVTvjbbJC9
FAHF69/6tcxQN24nPwq4+mW7jbKHfgGdZSYUSERKXk5XrT36/P6CSGVC2zPgFJin0TJ4whIOv6a1
NOUFmrkTUlnthaLNJrsfWvuWtaWqqttssjjs358seQ/VTGGJLdqu8zPs4PvBPydaPe9BDtoQ9wdc
vrkCBMgk9gI7hCsQ8oKybE7K7JOEEdmEf57hliM4X2sbOsC2EBtPxAhELKRUx/OffwA/iw62t/ti
ZtooRuSVVt8vf3WeUVJTnA4F6svt1CN/42k0NJetYTVQNoxwdxHWi8YjrgcQIuDqR58U0RU/IJJB
1Plb8dU9fG3FvhbgiE84bW7rEsZXrxTsyRXNVumUkqkHd4PDU/SoHte8jwmnT5XKV4HVJXQcefIX
nU/JaVN2+BWuKAisFCnm8TUlx5pIXVV8M7kRgNIGFn9b+Eosd+kDO4xRWlbc/7Eltv3+/f7NzbTH
zbRA+Cb1tRzqOgq5t+VMb3VbySnMrj9WuOzwl6HDl4UDG76RnRjx7NmZiSOQGmX1+1ouIhsTLkvn
54V7Spi/YBUbsjsVFHEofS8/dPux2cRbyt3CPEjqrFlZIBCQmEjnea+lWgOC+QE5hXEALm1gLFfB
kfdvI66J8tilfSIiWDEILiUyNZ20YeVLx71beshy4/qK+t0rFtxtsjL8ikrX2Qv30F8Rip13zjO8
3Ik93asJFFM3IjjR3xW9PAfLJ1pm6D8GMWyLTzoMlPQxxVaKMkvE9SzhIylu/Ujs0m7sEzUvAgJR
+/fHZShQKclRvPylGN8DuY4J00My/ocMuNcFHABlE7T5i3nLN3hxRAMdGtQ9K5PYfMuuyEuK0ugP
yGbhiGsigxhJqw3sLaPzdZDDN0lMwLV0eGFAJZBKxaAl8v1vTst5RIQKvrr6hbi3yNyYjLGaywJC
V1N9wkiQI8p+NH17ymFKht2iq1uoIrWwPPNgbspVnpk+gVKYXHhV31AzwUpHeMyV457Lnru/+iAu
qnccTr+LbKEGB0vF94BwCLj68SSKvTYKe2UXUwoMhPV0ytl5U8+ztcd2au/yZNR/NDnjJxdnf6Vw
EXogjM2SITPw1690oE14K7Vcpgc81CW1hqEbg+ZZqgdK0bY1QOiK94tHbOyf0VnzN011FcKdx7Vh
BKUT7vrTGNG0CT23ETViHCtAdSMa4Pp3zmJOA4pEqDkYlSMgak2i8H9xsCwTlu5fnRxPDVYx0dBN
OH0uGSGzKh+M5q/EsuoW6saIy5y6gaQFmQD7IEiNS8EO9LTVz8Fi6Mpc5mqmZMFYvoHUGmGmeAfv
PaHthnFt869s0aHZq6nTD5OKpC1+na0vL6bfCD/jYJe174UT+fZAbdwwTuzb9s8SvPC2dzhMUlsm
rx7DudgjpOHTZ+LnmxwaYCAzKr9Si5HFLATpG5bOFJypyxMv9y25NZom7nD7ftylwlbbxaJ6L8pi
awd7/OgiioqRFqQS2wM1mbAZpe9rT6CHiq3J0RAMHDx/AesmB6JgLuq36sWZE8Txwkr9+BpSQmU1
5nGotdixj9Uz6Q+zdXPEQ4X+lWm1cz+n+MM0WejPAYfrjyAxVXTVP+ZS26Wu38KEdKW9kB7TuSZn
m/RQfSlcjtiTArCdEEpcOM/AIA3B95kjVpxp9Fy++dJf3m0QRDcUST42QV2/1GYUixdd+/lauOzH
uLuzMm5bjAnInhreAbT2vGioqsip+Ed3zthl74A/1FWPyJEeltjI+OC7zongwSPWjNGYNACWR026
zscmd6uO6DMPK2wn0auBYu30lCARJRW0jFeTRlCI7G4fl2zGP388lihryaTQj+gThwTuDYoPf3wT
wu+K+ILG5YiCbCi45afpiWelURkXHlsUii7okoWR16nsqH6ZGCe1p1fVsJm3URM7ZWs6F4vdO0Iw
pfnCo7ozwUUAjJoLj8ncORnNV4aISrucBJwUJPDHi9cFoDWjzU4bXNOG7Xe0O8aettwubhwHzi/b
YxIjGJMfZd2LVBbvaf99uMuxk2Y8dbPvb1BXS/ub2+oZS1wkUttaWgGe3MmkurhxGa/6nIRMKZta
lgWeN/c1OrDKQhjBrPZNZEQ+15JwJa+VkbNtdu2eofg+npoUPNWMUmWRfM9SXU9lw+z3Hh1EtTpc
KNJyPcZ5XFt9PTIUFqnQ8XE6oV6x4pSZRA9LmQ9PoCPbzX65Oe/pTddJQT5Og1uXPqhg2P1/4tDO
qj+xuUGkOOLd2KAWO6CdRfhYxgG0ghA3nqkLAtP3Yy7gLjyUq77RBildyitF+VJJ/uFuzI/hwWjK
9exQQH4KzLMgklu6TYkY1dGIXNK426ZB56rliVJ7Kf5DuN2n10q/CoSh1FIHbHGsJC8spm16sDSe
Cw/GU49aV+S5bgSWT89AnwGJpnJd419HL5t2CskUPoknmDGMEEKal7/hEAxETVTtdbhVKIIsKitG
bKxYmnZwMzRGOoRWRO0JlIsjZD7DM7s+74TUbLeGX1ZaTJybjuizfI00FifDpPDHJdO0iH6jfeFM
IZO7PzAf1EP9xGBgqUAlMZS8wte1pqt4H7bYb5l9Qyy380asZ6+D1I9EkVawFiQQ6zHBLqU75/pu
cqpy7151MgDr/7GpE4oYG6DU8MTsTw+ezUKVxRZxDbFwhqkdpt/47R04AXP7NM3M7aee/TJimTZO
siq9mRTgOWRH92+OJGcZs/dQZai9ISHUwwXdWvOHNP6mHKzedxtZHaqU7/yq5J072/8cf80oxVWn
+fBoloPeurPwtO4uSbq+6nffUMHkRKj7Hc0Dd6+tVMxA/4DVYGq6gQj1sSWLFHOEBZ+aPVT2/ZBT
t9v7MFoy7rfHdthqukJubiX4XAxT8ZEz94q7j9JxzEluD+YYxinLOhW7QIeZj7RlgW5y5wiQMR+O
di0YX7bbRlOnyYZx1PeCekNzo0bt7uBGQ9OqytclSxOGUYcC0fnn9gPPaQzateZdp/M6uAjoAaqF
BOImnkJipdBXo6ECikcrT/o/naablN2cV6HHqZH545BGf4x3zXkS5zpcgMiJOfrgGrFahLov6xiV
WaB/jfOLZ7Cp+fvBCRXZ3tSC4Iq3Ambv86QkBxqCuKX/B00xOIGIHVSpErnGNRpOxCGWIpg1qvf8
Bal8Bqyi4Owfsu2XrOHyTkiEtMsqKZ6/IHBSznSIyLJBIAyzuRQ9J95nkQ/bkTe8P3wjB8Ymq0Iu
EWYrYBNuTyHwFzl0zVGy88cv5NT5MF0qBAgquKLdtqHZFhCB6K8FS7xy3glWOSF31kzvO4KZ+njk
ZMoAa3b0LLjVPdeioia1BIqe+4Ex770/7pki770TkqaTqZFF9cBXdosYiiSKZfii8b+aw33nnclx
SRIB3aL0KaUu1Rfcm/8cBOgR0CIZR2vjSJVxQzE1VLr4q7B7Y7+PEg8hG26agj5p1zNvV8nK/7rs
HM2obzQW6SF5QRHFVeAg3q3ZM+A26TRzgOIgzppaG3R/AKHZRvueDWJOMVDA04D7O1z1cL1w/lwc
kmcDqmq9jZO/smtyu98MYoTZTzeQ4njtIpjIZM8p2mS7KCB3kROSPNqGdug1TiLHmuqR+99RLWhu
qrhpExsgkTPIdj96D+Y3USvEW03Y4adPFY3mWiHBo46MqQ4chk43OEYuIeLVO3OyeRR8JAniIoob
oVBNMtOxsACjRusF+bf1xOBcuzQC8mAd/S/+q20T3+E2+DB2ZzBq7I/ZoHNeu6f+m2emUTIG0GcE
mZTjY4kivKuX7VyoZSVFfbRJ9i9lXuh4DFVcT85BjiwdScCA76+z41h1FEz+R3yBGHVIMamgeghp
YzpmWuS1xUYbMyc4rzAOU9YfaTJA0DAOPEJ9r3jTuA0oeco1nycx5aI8xxLSW/+f/80tfbO4j2lh
zTUJZTdY5u2BMv/LhdREUmClOnKqM0RdtPq3zYHoIBP1N36QU9HPIEe7dku3WMGErpyj4u6ZivEl
mRNvWqBv3f9wC6OIEaC7nydIS2L6BCdp6uV5aghDoZ+LymUysqtc0ww0octPYxe3k1+fDZo/osMN
tkGTy+jxlQyk2Ty/CeZalqEXaexEVDhBdaZvIS+skN3n0WA0i9ZLI1rdFGpVx4QyQPUanJ57sjNb
eoIEBW0sPdzQ1kmyHqIsHLXPj9/EZypgcXjqkul41OLcVnCj/NTQRXgWYoSopBFE7w7BZT/5C57e
Se0Caqfm7hhUuYAhptVM5kDNWjK6ynHo3pgBhA69EcB1drUfAsvJKlkJw48ekjz3+g6FJThtRluR
ehEtilmHuOVg8co4XnDiLX+cbFWnic8wgf6xRCICbiT6vHbjJbJmnz6ue1juYXBdy7lBBq+Bpy6v
0Kv2uoQvMIim5bnGkSengbN0rY8lswfc2WEj/6SiTkivWnO46+Z5Rt/5VkNxnaAyxtAAXmdPlgn2
h9xJsAMe+TR/GoKnzYE9zkrAsatWq4IR+IEq5gcDfWAVmrRktnT+PQSHwrFUthaK56QBxs9PldgN
KifanYK7N8bW+5wQ9c8KP3JFqi4Z6ApBzQNv2kWNSv4ZFqerderC/MOLmV+Noba83vG7UfSnkyPy
2sLIjp8+MpUjF4XODf5zRxjkm2TW05yt5koNKL9Lcl8p9bF70HNOlk+y321pGVkPGoM/98r0WZzs
wlDYeTAMPvG89rTjo6v98Xhy69obg3fm3X7tLF2jtJBFWAKmBroxtKsABXWwZalfjlk2bcLC0gQ+
bE5kVgMDsqdvrqDkE+UFJkbLt5phq2n8t+qrlbzZHQP8ih4dVPn2r196kkWIpqHPcN8eouvqn7bQ
OLecYyOIGnHr2suav+wM0P07Bs8cH0qt68joWf9t1reUzP0ThxKKVTtslXz1ct9qDKD8lcrzunJ9
g3+tw2vc/3Uq6b+of4Zh+iLRtpOxV0pSPxvmMvGQBxOgSP68PDiCvhQ01qHeHsMLbpH74ZYj0G8T
lLzxxzUdDIokU4K09ZBtLbvUzlwP6XR+eNHBv+gFY/bAM5r/Ls44Xn11degSWwMWeKDJmNN6d//v
Iy2nTohujUXdPry4yxJJGfp4Jq/QnX41BtZcrh73kFYwevtvvK3LetSySzsWkilR6Lw4FP3pJkhM
bt8ET3fmdvCsc6yqMtx5C2QFAj6W5L8QOtvtuHcdpsfFL+kzsDATgZUk0czekTLFUIx0vAYqiJJ0
pugQhqUENmGFl6jczpegp2Pu/8fXP6gJjazwLUKdy0ng6LY40X9AJFOSGv3jtmhVeFSqEjsFg6cf
ZWXJ7pqSqOnfsp/WIwyl7IXd5IFHPOWJ4T095JvNa0RcG2WJ9LlEb64lGoswx3GRETElyJiTiXnB
sgCiECbIz4QOI2hMNLyBcaXcLwY/AK3JzVRHdHGngsPkKi+uS0nE7vRgExQiNDHMg8k5aJxV98mm
MyxaSK9OOBqYDPlFR06AwVvctc4PDKtYAe8H9L/WRT67F0wQPObLTf5DtRr4Qag+OR09c8yezSUI
1Cpq4Nelmq7Kqo+DuFJXrEWwKfHeNRps/uc5hcZkMDhZTAZ3oSxAfOsRrnVKS7IayFsf2YUuawNa
Mz1qtwFv3G+w5hvOaQ6k6iKqtZvgr51qyeXwc590KeKn7cG6YEAHWzQvOVKWazH4ft7W6BrU9pUZ
5Ptga/NgkIY2aET793JqBP/1CscLzl1iynh+2B+2yB3SiCdcwz+VlebBoOZPoimZ505K073r1UCq
KKkTRyL8YkY6jQKqMu+CI3z55DWhb5WnukL2ax0axm1Y6t6mP0Nl8uRH4G79ojtqe0m5684pRB97
QJgh05/J5C045RiYNhoUtiC3a7MMGitDn8eR5HXkaYEkT4LlxIIbgfUo7SXBsKnU1Z4vC645gk8J
dwA1NryMf4YtiTelOfdxvMsBNNoOgQ0wXuC6z+0L9k7/wCu6T5lufofPJZ3cLKsnb69QkR57WjY8
Bp1mbm4H9YmlL+9cpJ+hcnH7CyzZbOq5JJWumkVTiJ1Dx+yuTG/QqOt/PxiDzKNcDT16PqjSHChX
0aKp/DOqgmVODJJb/aoE4P/9j8pnUc3McOHq4KqTGf+k7yKz1Qs3aBO+1CB5oEFz3bDu2o5q3ST2
G4gDAldbji7QiL3hP229ybdoi3nss3t4f5IEKtOBLJiNywwkFMJuUG8FYguIvT6VWbRFoLqsWxpP
eRDxkF5dZeN6WPwUJK/FF80GZX1enP5UstljYsjQWOdyhTMcbKuDEeooiKmqbF7KOtIoKguNxQh3
kGVlIKj8z6XPh9H5nYgeRx1bhGPVYxNDfxkCWuo592AmITodXYTx2Iiqmps6TQsZJRST6ztsCsEr
EjJJBmqt8VcNuMv557nvvdg9QCS+A+5KJKG1oHy/lMcxW/QtZl0Hvq85iaPvjvf8ECAW+vUYM70a
6rWNFmtfH9E7gmJ2lLcL7mbmFaW1FYdHjNKKvoDFzCCUdoThKVyUN55ahISNPpMHEhDmKJh+CYOt
r8gpPPKuUxI0WtrszhMyvdPls/kjfQ59546eXrZSBFqh5/da3cnNsr/iHXbh/S+RLmbCKNpygcJ8
nyHh7Pwy0CbdMGDpUOQ/YzvGXuxBhDBL9EnFZQreXB+uP5E4Pw9pczD9ITr4W+KBIw23DR0wptO6
w4ZC4n+6S58Cn4ZPvVLABHYy5S+RMfYxdQI/PwwyIwBk9ujQtF+LfpFh3x6OQG8V0nKd/jwlu1dc
p/c5qv7rWVQ3ZKbw1M9MGSs1P4S/LIu10ElJEj/qgUMLZivATCJ6NNe/cxWM7ge72jJOZ2FvZIE9
pKZ0WscE6Gox79h15fAa/mct/JRBQmTyx+ZvIKc11FuC11yPHCySOnZsPpkW3A4UTKilOIisYeiU
sbz2m5A2lF/yTXskmX7BnH4nTbfLpOsIarRZgUevSSx/8cNHrwfhWiBSP4kXCUcEoCYE4q+CklUM
0KvQPn5sOQyb4ecal5NapPj6yqzvBncGKOckktTzYKaKudfNkQx1szAKdAKkGEvw+812BVqRmHnp
jshmm0HECkvcwAKoiZXPXzkDsDTiwHlnXRe6rUe3HGfbB+/17dfELa9ChyXW9o7JZ0IydTVmBX6x
MUCQKUsYo3fBGmR9OWV3sdHtH9YFNL94b74V/Z8VGnTTCvlUerGrHKOp7ySJYqlp9EyoaJYqoAJ6
zXE7fUdZulvoZSXEgwMIKMnlL6X+/x+BTwzI3xeHTOGGVXf2CF6etQ1CmmKNtR2ubIDWujP5eHY0
BT05C5bXFxdCxG0bNtSp2VbGK2HQWX2ecCvj1BpWmzb9HJTOuDNCZCAlCf+PgKJB4yNY4pITf1TZ
0/VLeoAzLdZqqcJS3KXuFVbsF2P5Xz0Mb3nw5HIGndIMPlhA/j2wHKzqodc7MnHquDVwpoBRpr72
YRqO5oQUJwVLpYqRiou0K4WnHro3+29HxG60JWwh/fDaaFQTe/OQVKE6QmE1czCEhFejLumpTgX4
ZuKEXb+c9V30XvcAtbMORjisNsuZVGl2QNnbqRMK39ga2lGRE48z6oa6QxTLG/YmUoZNwp3nr7y3
4Ru/mYdEo03ghLgJXUxvwSZ0W2cz/YSVuYA8EWe+Ka2SoWc1ZkOdReuo8nixNmQrCoL5KdE22BKX
Cp31aRjNjhG10X9pcgi2erZJnRRCIjveOHY1Zx6Y9eKoWlDOsFWUQ2lbr7zlM44rl4Y0YQ1Dkd8R
EP9FWm8A1/H/sybwXz97vhlM/4x7DSQFwkqCU41+3P/hmZFGg2ySoT7iMmyudpqtBQ2BJHnEHTG3
Udu8d+Ia+9AkanAdBTxq6LXNowsQpTMttYt2c5a40mHN2fp0/EWsdUlIitu7pRe0RoPie3hCXjmR
DKPbwYizR/aG/i7udq4wFuFeM33OtfH9g48GpOOKZfImVSIWuSIlRvekk/Z0gaBqLEFO0fvFVjaU
I3Oqp3poexDyTWimiXxXpKsRO10Zow4WXUIz142s7+HdILDk+hIvWIjbNwSDv+ceu0YDal3IZKYP
otPtWb6c4PVjTVQddGEXj0q1Nr9Fv/3t/srvs5MSea2g43iCQoJAF/X1K4HiFUGF6dl0qMu1DJX2
GeMY/bqe0yFwXk7G3RQjy267/w/E14AkKgTEulbYDZsQj/8MQJG9bWu6HRH9TmciTvH5E+FSTRCw
7DyFg0E17++7Fc7jkRPOHh/skxUnFf78Ct+rs6/+WEaOo860oAF+0JBa4NP7Z1ZZjkT9Q62/UIRG
g8lEg5j5FcWNsYijQLzIyreFclRzAB2PhQUuqY8/AAbLDckQDUFurDxhkPNGVu7Rd7onShyVRS8x
2q8w22PIw4FxM3OvZdeiE1nNviDv5KYDCSvOG9gtj6S8Z+Y+03rZxmzmBYVo5zGS5lPEKGQjSAAI
EAo23KxzU3Z+eocZFisUF5MHL1fcVoSSRmcBpCt9bkhZqxZc2Wm7IA3DA8Y+Zy4nHPx9MjenArmM
BqIBewT2L/mZWEQxm7gFSGgGwr4uzgJj1G3Tm5Tfbu1fXo13CXO/UVkAdmQJ7Fz1jnaQBQq4gC/O
dI1dI1p8vwPLoPjwKsc6uVsq3k3UV/PxZ0k+IOn0g0E4tD6bEj339okdtPoHTslreX5ILnGUhS7r
Qr7V6TX8bSQHdjjRxfeul8sPOOlG4HsVnLluP1aRJzUnZ84n44MXxRRiSeefuACt+y63RTg1zqLI
/spgzCpnwm8YBzXCO/K0SVU/EDHFltob2EKAEQYtp1+5PfwnzHmd7iyd/TfvW1bGlawZfnv7FWQ0
m5jPwbZ92bZciOm2b59T2HSopnigc4intor+qN8xNFruhQhmcf8XB+AMu0wGXDT/PXRDeovy7fuy
NYxNl5U+UCikGtZtGhxes677VXOjxrx5eiCYqPVHDkiaNhCkXpEPV/cTtlsE98lIWynlUrsA8WHu
BDWJCPY52rVxnHy69g2+DIUuTmgEw4ewachJYMae76kCFoK8Do98FfApOly/th+XldTfRipTQD0L
YVP5FIGKwvCtc40AlHwyXRLgc5cCzWZQt4AGaMShnS4Pl52IHTGplsLtqnOQIiKrFVYuKurbpaNU
H7Vcqwn4y0m/aKsY/P/HoTN8wrYNnnOoA2oTR1zkCpg/49AspgX44OaGMdE56Isk7Ce2QNtbUYxO
AAJvXeFWDNbJymGZpC1YABIIKmPOJEnduYIQrhEs60gvNWPdww01kmAvVOPAz7b2X9nGMNzLLs6z
UG3PcG/KJoBqh3lym3lgyetCgNgtjUTy8nhVdj/GZchlwD0b8a/S/Jsfj2dJT/DwjDTGxiSuF1dD
rtuY/ub2rba9hdaMjaubZMSwy0BVAEJKPtYtWfOJfuIFLaOncDOmHVr8mERFrHNK5mp7dm6AzmCV
GYua7pgXAboNUs8rsuMpiCx3c6hNDd+SyB8uAK1naInsdajUcDYEXPP3M5Wdt/NoZCoiMCBR7lr0
JhPPgQTep90ILN1svRy8+SEINGr+6n4AbftnGfgQYxcjfJzWFmZg1QjALeqZIJy/3NYJfE5P9YMy
G6iDh5IBKbkzjpo4w1zHUjNJfdWU5XNvKr/sTraCudPjRtESpOtS7zDh1wZlvKLuFFgGnvfRLfwh
p63snyetrWTt5r+gGC91zuDmw4+KAuXXQZieQ2kwT2G22bvsQgElVhYCRCnBbjm3gLV241O3Wk1V
a4HzyRNBYdnUny8xLvdLVqm41OfnMlSAtoRRBXuqaemgE2xXgmwNI/19WZfHeiwQBUT1MsoJVOVq
Q134+7ZI/S542fxg/Qv8opPa1zewhoiim7shw/Lj0+WoG48G1oZJZXn5V/7aGr+woc8nFBa8+Eyc
JpkofD03GrGiVFga78+bg52BFXi9Fx6Ugbg5hWh+laiH4eVphhjSJlz6iHLd2sp/5YTTjzeVUYVt
rOZoj2nAxcR9PzPFmYMAqnzBgxWXSlxvoCAG2OY5+LI96Cacw8qYe1FQ1vnOmcT5eG0G5IzfYyE2
G+5pnvZpTDzar2qhC+NV+n9QYywXTC290fyvDCVSoAci+j+N4LL7Dd3cGKlx90RIo/Kp5Z/jBXBE
9potAjUW4CzxnVlvG6BZx5SYxUTiCnxy6/1xzvrKoz8zBwkpCobm334r/QtcJMxwks3Pg8pH4uYn
gVtEzjb0Noi2wvJg27JQiZVr8dWc00fQrih5fQEKNdIP7IdoNScfJRW/KOO+Pk47i/B9BO9x2xUj
fE8Cr7xXqG/8tJPJB0ZR1+Y1+JcGSpaQGmDP6E1wa9mpNBZWYHZZaWNbyL3fe7yTX2rbYHVNfO1x
C6ucUM/Umqso4W9hRyRNgqhz7yTJZxRyrQqJmTe5lYidddg+zn8nGg9QXa1qR8bU0ZUKcBiZX756
gMGJPiA5jVM+c21octTOcB1DvRXRhRRtqrP4l88Cqpq90l/w8gho5eGyB/u8R8pit+jC/EyFuBrj
IHk/D1NLjFAAGKIapvHo6Df5QfX53gJGoR0ui+ro7jCSkAzeeQcaw3A1xmw+nxQcrx+NDYgTNtKh
HUQFmBpTMvOFOOyEEcCtxoZxka6XdjHk5EpC9XnHHMbSnC+eHtYvw8JDtCxyd01Xfnnfqd22V6NH
sLlf9hqcqY7HnObqHFOA+zDX9TpYpf0fMUwu4V1eV5qnCdCG57ogy/MxJPMz+WWUpk2gJeSr6Uat
tYNXZzux2ee7ZxXIcJmfDTZ0tt6Nj2/7jX+QnhMx2D6tIJsp2LQq/L34+tEzLMD5sDexHRSlpwL+
lSUkF6j+0LGzv2VZ5tnMDM9KhJoxS9L7HbmYBpo6K9uQJ+TjgaRTFtbEBsOymgSYswCAN5UB3xO2
0y9wPp4ZqCUVB1NQ30R0nlqkf2LPHL7FDIQrdOatPbG9qhne7eZs+CiaIVRJgWENRNg3oa+Biena
ADf96V3Sw1MByR0HLxVnVfb4Zp/V3f8EeMroiqfRFjiyHNe4Guxfobd60dkdMssXixa23jk9kZxx
TLXtUkS2DTZu4rV/RF5ChSzJNYRHwHaoDRQhTA6d3eRfYYMpdyR1Mu725JGFEeGPPyyzuHLCexjS
LPvXpQxCDXbBWYUJQKKvf5WTASLq2kMpCdxhVRNJsjlVHUQBnTpxf7AFOsSAJq1EwvbBWoJc0gfk
vpqr7emiXt4V0jieAFW53voSchqf7ZCl609nD7oaX3bhGKX7qjIDypN5yb4vX9lxQqXgzZ+sKb/5
cAm8nU+oDU0k2iVfLy90tgFn6cq8qbo80fYMmvF4KkQL0C3zxDF/4z+9aJdKgv/5VuUtJ5m0ABl7
6pK5PxNVkykHLPJFcOWibrdLDJ/BPzlCWRAEDT/vWv+9K0DbbQO50mCBOFpJh5iKHD0PwLGCx0vR
GMHiphWEDqJ/9+gbWup3TpyfgqJf1s9sx5O+WTk6oYb79H09fKERd25cZpCAwkIfqt7GPzijpGM6
kH1CGuIE8CGApAGctwXqaJsanqhZlOpAt6/SDMd4pqxHcDUFp0BmcuLm+OkLkPlzTqYbztEG9Txt
vN54uJRWpgYrVUVodR2xVy8gZlRadnPgIAKci1rpXq7yPf+P5MmCAUsBTyEZRKWql5gkmOB87jib
qHkPwOFKzvI3isFuAz6E0xkkySMOVXX5b1oKl9IUtd/NbpI9xd2Of1eOLStHEJWigQ+7zVFo61O0
/gIYnYISfiTBYUHx/CPWpowHVi58tGwVECdBuBUHIEaZNZgAczxKVO3e1+Vwrc76yQwQH/ICIJiX
UUf47P6bbWUTYQu3mhnRQZqfYaq9LgNl9kFQmEdp+Ivo1fp8Z0WHAfru1Hdzw6eo3xTHy0AU7u6p
qTd1H76seH3UWsiyZojAN8vh5HlSZ4v8TqFCXW7inl/QzrsADm/Os5RYYS2lQog/3y5+5bod0/oz
nHm+fzEndGT49gmn6O9U4okqe3lnp3LfT9Jz7oweGkOj7wgsOdnxz5RzHoFDjeXFWEtd1cxhmm2T
tKo4fMjpdK9atfVC8LULPOKmX5x0l0re6a7p2PfHsf1BTnE5acqTxpG0UejiZGTUSJ3vK/aW13eb
kyy0NyRSbrd5sWkxATOwyDzD0eI3S1IxuxsVym68/GYO/6WKWn4ddozLl/ASsTt5ZIpvVtD17rQc
fObPDcTnFmnLeaBWBphx9G+v40TbRKDLO6Vyp0eHAieJv+oc0rVeGUK4GV9Plr8vi9achd0w8k4Z
HOIN8swBgmx9uSmrleXDeYMQOprP8gaxZMdIcfRuQdfl74y00WEa+ru5N7h32C4B7jV5GGBEPwaM
3n0kdtvXRCyrppwmpuwF0AsWHKZeYug2EUOMHukDVDCA1og0vy1haj1W69USZzRWTKYy47Y0yaII
hNbrnXGU36FCj/gTy/xUP525ZoPlGq+QP2Ufrv7GabfOU3H4BP0o8gGj92QrQQsLIOy+ahGiOkeh
Gie3M4X8HREK1OtPFRZ1+Q4FUXreWO5BE+vxs7Q7DOAciVDGGoyBUvaOewEm9ngIEORRqrut8i/4
3+aVUUwMoxIuGX8WSN1O9MLE4Vjfv8VpLoXwRlRT60Zt8RhRCWL+es2GBsVlZSVoQcEgsGk5neAu
quLhjLsbd5A/qGSi0M0umBZVUy7RnyCwL4TixyWlsksyZwWhmPUnykwHM5lER7CE8S/wLC5NbSrG
J14ABWCdCnuuYTyKvtelmc8ycqyrJB3FXDcv9x8CE9xVsXu4mwF3Vjzz31xcY2cv+iPUx6UOpu0D
iqtesnpRunksDZkN8fKBAEP/D7f7Meimy6tsRfYmVfD1U7sRw2ThYF5ApNA7qeVp7RWc07UPy9yG
1lMqzHueT4qtReBBhv1VSc8NUjzqUCDIQQPwrpxJltPxDIyvlWJhJKZma5vjDyeKrvi/0GjCtaRm
gWw7+izF+r3Q8iKYEHVpS3VZXYezKB2RnH/SPzGc18UZjc/Z2N6blRRFHmxj5m1jodwmDJwOWF3m
hBW1CJpw0WKW6MJ0PLIDdnKrvz214S0bZx0R5ElJtyadMw0lZ1TsFQ6jugGcb/HBFu+Zqn2BqZnG
VTxukmiGe1Rz5JqUdE9zyoeGpW9ZlDZBW4LOssiaMlkRUg+C+xjWx8dcOI5YPefyXZ5xNmAqPv/f
hJOF0+7zYxms6BtlmUAptLZCqXnFW5iR7wbRSSQOS286JKk77kaHSlmf8iZ9yU4IlKdtZS5ILrzd
Iz2kGqCTj3PLOcZ65KWYj74NL2Ky/Beq69sX0Y6b6G2WckLl5OdIgdQGBxklxPlqs9pzbC4d+510
hDwbvdlndgdpWr0oAuSBzigLaqyZ7NOuaHspdnmN5Jo4ta7mcwkn7hRTy/ulxg8LdAEK6hYoMihX
LylMeJnTVnoIVN3pkgtP1VBsGISUEwoAvNos1V/55agGWw2lg+tqTWHNhKauJni9r2ve7UdVClOA
CzGrL/ONHjHSVj3mxItgmSAgQO0A2wHXSA/V2tUJsOmSrS5G4VAenYDXuy6nUxNxuHuZnjJ5T/8b
ltHE/xg6F+sopf4Mr2c7b9IUphyxZzhCOskWckrA5sxtxO8cqvA30p8C3qti+1K9p1Pk2W0CXT7X
ZExeFRo3k/vHOUcT5QOd3fbxj09OcMyWQRnUUy4MMCOYvvNk8sXmsp91YLnTn7+KD9s7PEG0MXO1
+ZieaDXi0U57clrEe6edRy+ZqK+5+rohJV80oD4Ga74wfuPIzB129QwwZ0t1r1ENr9TfLKwJP2vr
ObkZ/SqXkH7E7gAatplCs6ksXtEPezfyTu4176pmtrYKW2pM3jgphTGR/Qc+exAEg+i24FBAb/26
vAdFUc2XiQtgTxyFexh4/w6J8g0uisF0Kpl7l6iPuU+nr6ia6ozAW6DjOhCLTUZJGcKuv33UJC+1
Oq6HQQQOpI+O5bRptsfcAWf2nGiLlnS9/NzKrV1WpcP7I8Xs7pduPPu3TiDF+YkV3pn+ADktwQuy
iM2gvUzmt+z9BB3OBVUbHvubhXgfM+9FzBE1DFEWBFq6DzgQGmowHk7yoGmeC+PTbAMqcXT2nCWm
xJurNrnToa6EHqNcdFqAuapT+LWlmryFAiMu6ZrvoAEPIPB+/tkIWTTbR5PuU3tbapIGI8LEuBvS
GQXDHg7dqGBMcBc81eq2BanbH7R/8j2NC2Mph9If7TzK+aPNYnYAA3KOaHk3qHysQOeau2xkGGmw
JMFt9/2JfNM2pKDAEXU3MYkBm1S62BzKiJQmB8n13/MWm6ynvCkzfeBs04Be1DPV6G5LJ3zDn/fz
UrvS49KOW10wGAmJD6A54EB3TNwtapvfAp8U0/3t0zanFRj/RhKnThl0f3/hAlMpcBFvqJDdRF3g
AvNlQWAbU4tj0VjkWeMhEjT/SBeU4zTZHZbEKiUXhTlgXrU5l0nnq+UyrEFmZjh8QWkTtc1CZnCf
Z9S1niPsJEVgACB6taBaWjtl5odc3Sr+JgDycdu8mxyD86uzdfzRJyuoClizZ8N/8CNNpXdyuxBI
MSFk8lxPZagtQiILTibrje6sPWCSRZx6P0WiTUzRhaMKbu1OrtKjb6BrTsg9MfgZUhWeUkEms/gq
gnXSyQD3q6RbuPtAn9Jz4hX6INpINqqrzgjjZ0/TYjl0sFTkvKWTC3ErlHGWBLj+HzvnVoQ9CZ1s
vZa81hd5FET6p46a3A6KHLmZDtnytO+fSaH4hOW3RbcWQ4pu1OLUSADoGR5ebvHoT49NvpuHUJGQ
BwkYRb7ZlfUi74cNcmqRY+yVSNDQOnGAPpOpqGPgRcBZB/99dktH/Vq90orlHFCTSi5G/tfPivw7
VjxB4POntahjs2BSeLBiA+pMTYiDkGhQueCyKcSBNNCckCyTaO0Hyk+5IXupAWwcX9zo1wZSc3PP
WRNkeHrfMCeipi4XIHn7FyA5mgo7Fjvlz8hLtkG9nKd49OsP/GfWdRpoR8piB5jJMlD+6wK5VLYS
YbphKwiVZRrkbPv1i8dD5twQ6DEuV0ycFPthhfA1QmTK43eyNhTXb7xdGBnMcMb6nT/J+q6yb8xN
RZjpnxbhSjNi7GaAOQK+tpAANcof5I2zMyqb3wNVsyY/mJ/0nfuz3+RlvGf94heVsnMu1ov6Lxf9
ZSlGB3hwlGUURbXCBe+FhQAv0qR2wMcWwkggvG2W7X+3rRbnKE+TbpcJxWhwd+E+GUWlg1rjLS38
YWuInaUiSKz/UIpy6XmE63t+lmyp8lSKwknXZD+r32/xzaIoduViO9tJsC10f41m9vA7G+hxULst
ctVvD4qdM9py3hYYVmk53NrVTJm0tn5uZ6LF1PV+os4mXak30M0Uh1xWPIOxAB8fDChthVq5oJE9
gz4PTZWhlRro6iT35YthZqfEnp7qb+wQej/fdBb7MT7uNDqw2bbRZ+x8k5BPQoKAurDe8yGKbsI+
6e1Tlqfbi26m2mOjhb//vaTZZhBEyW9h2fOta9ObTIM/X7D3QXM0mUPhXnVRxv6aRyjAd3NMPC34
dPPn7vS5aWHNipTSXXXjmwHIC5vDOR0ixCtpHSARz9mlS8BgHKcbwNsm/ZLNujzLvZJV4/1NaAg6
EChqll5EJ8vbXL6r2SxoPibRbQUH+UBF20r8gHRx2BKpT/OgHnfAo4mkUEJkJProhLyLvarWpp6A
3XCut9SRkvBrXZ+20QbkODzyweBxi0DyUybmdAjFCejUnqLNSfxgaL3zJKFPK0qqoG9LBve8+/wk
IBa+5ARSg6XSoqfmqp/Tyls4lF4gig7bPPPcbH+XyUnVKke2N4LI01fhkfjoKIlJyuGSOIFNV4me
gAAO3S/3UGzAKGuCu+YpOcKciD/cqQ02Oiqw2DgwPi55U1TVGc+oZ6EXUsxpamwJKGIQdU+l5qIy
JMReJP5xr1Vgod9JpowWlMAdNsQlIptwbJgjvMbdl0rnoaK0Fk5rMvWnaBdAF8NMZO0JsYX7ItDk
cJUvTZIMMJaOF84yGxNbldd5Jrh9Rkv5lDRJVL/7RM2fYXyi5C+Ec85MnVCgSTL4IxMXnukMKA0h
6rOTGy/VltsDoY4XAoCDcdypLOpfGPdhNZhe7E1k+bLZqeQ7vWM0FE+4MKwHXH1VqH8fKyfqFA9J
JDksrWL5q8JctCTYHwC8wZ+mU8ats0Eqf8LHofPMB7PVynQ0z8ueIOrwuFYuGP2Acs5rTXyb9y57
Pb8CX8r3z07ae6e2R9j/1nuIkTUF70+TVxGoz2CoRPrXcTMseeep9HCTi/elx/EhPqlPytO449Dj
djO5r36CabKiaIKeSxbk5X7W8BoygMYqc0JTMZUqeiWzBvAaj9AQg/KGJLOIfbeurvsgmVDd4GZU
yYNytIWATujWGnYaJKwt2JCBetKg21twOLPi+Fo42kbYh1bNRSsYfyMNquanA5V2PakB+jFtxhWv
La8s9r8FXmQ0kkxJNsPrng29BKC89BoVPfBCgbnVvPFdDyLdg7wDRKJeIZTZU3mHgGo84cbqg4p8
SLHPlHQym9QTYydgEYQBJfVcn0zz3WIWpr+tDVAjDSfK30Xl38hT+Ld+CDmix+ablJfUN/KbrXb9
ojhehXjzCHGuNluAl/qK+oKaoToGy4SN5VABfL1WpgzfaXP1wtzowxuwDZ4PW6RXhpEF2VCJ/Jsz
gFJqmcYPGp7ZGYq7gH+VLvxpHSoGEQDHuDKalARrx9Nz4lb30JZrzwcA4tvvxCKoSnSy7kmugKqj
5RQWlvsR/A1jQfsz1BY3kBprHcCpiFGEA9JXFj3NeQ4RaNZulzSZM6scS4dB09fPzM/ZRizXggxw
ZwdeSIq0a5RhIlSmw18i0PnkifZYNkiza91M5/uVpDr2LN7D8Z2L8tvxhAcGMyidPDYjKfAYLl0T
IKhgu3kE+2vCoq9xfZN1piwnyXAeJVzNf67PKMh69oiYKClm74VArsv0InBz6XbYU5BeNkJLqkG+
zIjeu3prQgrexHhGaIBl3t5gPQjkC7tB5K5DJcZww0a0pXZdazQnK7JuUe510/P1UIM6MWwFSn+y
oVYaXwcUfiRxMOmwnqLzZNWJcpvchZas8anaUB7rZqm+hRiy+t4qlNkGlPD5MGThpvtxWS4JZ0up
waqd8w0AHglK3Wz/Fr8BeIatjkdbvPsjF2dkxnafbZSewUUuiFaCZcdZ+mTHpVDx/iR/9gIcLuyZ
Ij4p9z3bA42e17E72F2bGv1XIICW+PS+SacAciqip55lB/GToM9/NwTN1KKRpMKO9e1kOYJ1A5DX
PeMkO5l8FERel0URZqURnWP2SJzGDMcL5OiYCUnwJZg+Nl6ZMHqePYvR0akiM9vLkFSxbFshu8r3
NI8E+FhlkIkKWW2sCUm/mPp+ACEYd9o1RysDdvS848SzOrYT1fDjKJ14ASDHd46jXDDBcKYJ9zuG
qrNDDmuBmKvha5cMB53gLnCeBLBoXU4kr3/DfYp3GyoIWE2QD6XYOoatmAooT9zioUK21r+WMswt
FQEM7folJp1dLv3kWomJskghjn2/fH09z2qFgWWulBfbHQhlQl4veEOjCYA3Nx0OFve+S/R9y38x
ad6QA/5oJYLYPgtP4fxXP0OzvZgHhR4TJJqV8eFh0PlV9qGX9shdStHVaXR6ePS9kgmKerqj8txR
weFXFDmRnKQ62WZeQUQOBfWxLq4n7tAnJ79/MXb8xHrdExZ1Mqn9F0vyAC5Bpd5vYyvcrqUKEFrq
MqosSyiwO5W0E7rF+0QtibbsApHXm3l20CbOPQaO4vOLWkANDIrTyuvXW64+JmB05llVX6nFsU0t
2zWmdCbpnYGmuIZHEYWzJ+gzXE82ZoTpt/01MMIMOm8gwQNyvrXlNRt+5cYq7EXs9K/n7NUdj+Ic
99E564u13+0eWEkA9YwP2YWYOBqOQLCWBigzYVN+Hg5JozUxva8RlwGZLJ5SRfOLzv38AOioafq1
AfDNmt/Q5fX9u1gOfRWxOQtxWHZQlbj57+3Lrq2G1PedksA8ixNRZSyKPhZ4I/D/tCaeKv6IS9b9
fZEBPeiYIleXEc+o59lemdHGfHwEpVctxjVyuEgoo6fCIeiR8x5RXlsSAt6Zd1K6o+D3+ZceWFQ0
yhQiQdP2SjFBmYtd3q5tYuk9vJDafyiADdqoVPfkak3qa0zviMu3ZXLKfB0/H7QiUQtJhf18XJlH
Vh8No22xP1CUesg2RQplWwD7xQhW1As5mvA8FGCWSxrOqZyYjOvb83vyRnqUQTeKOF5aDg/FkhLs
kTjmqDVRUuYvT47Bb+Tql/kTIDDO4djERNpgYlnRW3I0EYjMKTIAmPCWv23gPNcgoH1gy4d+MMTM
vzAh2KTjlOGw4H8/9M/TTtqNBDcdh/r9TERUs1VApRziE6CFwqASjmB+Clca25ZAZFpnvl2vKh6/
TW6HjBImqu5yAx7VlXcDdeDD9cSk3UwEIIsCLmFo+djj3zfrmElLyNTTYUMZMvwQBWN5GkKWHkqS
2Tyqmx8XkX/AvGvJciUcTKJ+x7ZE3klm89CME0mbYad+CQOr+us6kizsVwrM9338D++uGTi8p0eH
pDKat340RL4N1K9bEWb7ZxYmHIkUNNsGczIQtuE49yc+AeetoRWL2qAQsBgu5bpZyC8CfnTGDbM4
xPJJOrd2/k3CD0h7cmwEbCkDam7Vx/vaN5VdWAVx/TSADqPnJrkCsp4EXrtlVGRQJkZFM9PTS0u/
MGgd5VoulSnGbhArUlp/0FUjF10zaDTMgUUnwmlmtqNqKWKK83kSnHciKjxOnp6KwCaC5B6xp5gn
82RRkdk7gxFCIh9BERgE39eHsJ5zLB1JUmY/PU1V1VYmydLIxZ+jI4GOrdcsTY+R/PPanszkM46K
SJQ++Y1sY9OWVopDfkMpqz44/5g9xBeh97Llw06iBGgOF7dNGLFwR3EUJmF5RqVuoohuf5v5zCco
JA2pPH+ZfqmAnZdfGP16ZMLXVulkv5ysXwiiaDdsIAdgfItLCNXwxIHtrZXFJxsWWLmQC8eUza5Z
PfcLQxL6Ksvo2L7nzDsBJXQRhiuz1PPMr8S5xxSAurEYs/nlClwNV/GZx852JWm3jZEOJldfIi3L
+7JMwInouGWYS3mMgcv50xlE92NH7fPo98h/t01AQg2kUx8tsKsY+Rt/sYPPREqC/LizjcyQO5CI
pTiX+sTfHvFOuL9f9X/OFCA/RfdaWaqa/JnPnzJ5/c8sYTnTgNlnw4qK5a3/V3K2xbk90KzSoESO
F4VScujqYLEPCWLVSXpYhZb6FGqHSn+AH6ZUxk9HqUnkftT0AK4v3AZg36AM4G53M7CwbjKYSjbw
S6q/5PFNunDQCZiqzwy9fkMZRtvXKKNR97qcYlGwlPu+raMCPtlhEWdGWWOkoCiCOiWwO2moRl/6
n/ugV6lvstz199qh0PqldlmwrIkvZXzgliTuUhsrFBeGzSObXv+mBXxAbdcti5Gy+MxTi3Q9ri8L
FFekliuDGHy27Bhp1A+kLvgJb/FMxCx+c1+lXAaJTKD4/4edB8e73FHpb3avgV0pMCeYbbjt4dSw
pKX8RvWXBVWtXBXwCO1nCBHn5EBpwLS1ZCECSnbFCrmrEpmttNyfbh6tc+GQhwLPrsszmGwsstlO
zofN/J1pulqkUzOSInUKtwegj8ePIQ3/pcmb/2SCuLbIWlz7NNafnzF4ABTrm6AjguX8CZ15biv8
DZPXYBwI8mSYnDHd9cyo+Gck0nHKEYgB5NWZPv0hbUE6lD0oNkWtPbZQn91cPphkIxZCJ/mrQy0Y
MYdEoiwtrTwGQrmiC/WQtGRsPdx2uQvOa5Y4Rq8tcBwHQPxjLKIGev2AyhWdg51roIDpByuRyrj4
9FG6rK5PSQHUEAn+gA6ZnOdP6lGdCZH/SeFAsyd0V1Bg10jpvo4wzTnikqW+BxEarP+8J5XeHluG
BYCpDQ6WjQGZO1TCuyAR/JxqQ7L2ovdDMJvDteAT9vpSVCDiZU7euz5grvXSoeBjuqGWkMnua9TB
hc3bpdAja1u4JjB6AOngkvKTBvct8DwBBnNtWKyhR6MM0X7YQ+Z1jS0S+qjodvYmB8qN8/7hAQ1O
r7KPPp62cz5i6qZK7UBsNql0terEPEaMFBwDUYdate3Wr/UJsO8dhldxH4h1sPUNGCmexVNmFad0
/m4V/Mmc+RdDhzYMS1BUUs3ZBtaKWv3Rb/kPT2uwfmvCiHEOePhZ/4/dFxqUnVHdov/XLfKkh+eI
CTtv4pkymAokkk4pX3eVyWumqMjWORgHerCElbGBhIsokIJyJ3GddcA9hwl/trDM7jObFGUhv/OG
mFMU15zpWyxCvJJ6pJeCBTiqv/3h6gM9XIa+Avqjr1jqsOMVlBxM05LOzMI/ZLak2NdMv+9/eLxL
yLJ1mkgVNYxIwYEQ/mrr3IzOyZKmShhmJZOwuwo8fRdwPowEt0jrdx65mWOzEQEN3gSK3f1hOXgn
RLE6LLLlxmwWziklnxQGJXgK+edYm3GZjVCp+oUa663O23K6PqT0jJSBcdXeNO7ENPyreUFR/ikn
g+WvCfyCufW3OTbHMXV19+4krXFLGnSZEiGc/kinftjmlApxdvoektG497QeKou9VD/ZiP7wHt2O
To9+/rc6DIsmJ3iIhRTLHnN9ujF0nMCLENORHI6RVUxwgjcTVNmaQv6ExIJv6X3qVxCK+mySo6+t
MYWxKqoYh49saxOY1a/1scR79K+oSFS+ND7m3wLDMd4PDd2xLQX6XFU3rClfAv98XoE6/xvhObUa
TOgc7WUkySHA9AqKHarreqhHv+skwpije/+mq8Y21HmvOWM6OgE+lmYPAquRKbbH+GHu4O5TSUlT
w8ACmYaj2NY5iI1SWWnzbQ==
`pragma protect end_protected
