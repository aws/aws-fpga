// Amazon FPGA Hardware Development Kit
//
// Copyright 2016 Amazon.com, Inc. or its affiliates. All Rights Reserved.
//
// Licensed under the Amazon Software License (the "License"). You may not use
// this file except in compliance with the License. A copy of the License is
// located at
//
//    http://aws.amazon.com/asl/
//
// or in the "license" file accompanying this file. This file is distributed on
// an "AS IS" BASIS, WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, express or
// implied. See the License for the specific language governing permissions and
// limitations under the License.

`ifdef ECC_DIRECT_EN
 `ifndef ECC_ADDR_HI
  `define ECC_ADDR_HI 5000
 `endif
 `ifndef ECC_ADDR_LO
  `define ECC_ADDR_LO 4000
 `endif
`endif

`ifdef RND_ECC_EN
 `ifndef RND_ECC_WEIGHT
   `define RND_ECC_WEIGHT 50
 `endif
`endif

module sh_ddr #( parameter DDR_A_PRESENT = 1,
                 parameter DDR_B_PRESENT = 1,
                 parameter DDR_D_PRESENT = 1,

                 //NOTE TO CL DEVELOPERS: 
                 // The below two parameters should not be changed.
                 // Changing these parameters will cause place errors for DDR_A and DDR_D pins.
                 // When set to 1, they will ensure that DDR_A/D IO buffers are correctly instanced
                 parameter DDR_A_IO = 1, 
                 parameter DDR_D_IO = 1

)
   (

   //---------------------------
   // Main clock/reset
   //---------------------------
   input clk,
   input rst_n,

   input stat_clk,                           //Stats interface clock
   input stat_rst_n,

   //--------------------------
   // DDR Physical Interface
   //--------------------------

// ------------------- DDR4 x72 RDIMM 2100 Interface A ----------------------------------
    input                CLK_300M_DIMM0_DP,
    input                CLK_300M_DIMM0_DN,
    output logic         M_A_ACT_N,
    output logic[16:0]   M_A_MA,
    output logic[1:0]    M_A_BA,
    output logic[1:0]    M_A_BG,
    output logic[0:0]    M_A_CKE,
    output logic[0:0]    M_A_ODT,
    output logic[0:0]    M_A_CS_N,
    output logic[0:0]    M_A_CLK_DN,
    output logic[0:0]    M_A_CLK_DP,
    output logic         M_A_PAR,
    inout  [63:0]        M_A_DQ,
    inout  [7:0]         M_A_ECC,
    inout  [17:0]        M_A_DQS_DP,
    inout  [17:0]        M_A_DQS_DN,
    output logic cl_RST_DIMM_A_N,

// ------------------- DDR4 x72 RDIMM 2100 Interface B ----------------------------------
    input                CLK_300M_DIMM1_DP,
    input                CLK_300M_DIMM1_DN,
    output logic         M_B_ACT_N,
    output logic[16:0]   M_B_MA,
    output logic[1:0]    M_B_BA,
    output logic[1:0]    M_B_BG,
    output logic[0:0]    M_B_CKE,
    output logic[0:0]    M_B_ODT,
    output logic[0:0]    M_B_CS_N,
    output logic[0:0]    M_B_CLK_DN,
    output logic[0:0]    M_B_CLK_DP,
    output logic         M_B_PAR,
    inout  [63:0]        M_B_DQ,
    inout  [7:0]         M_B_ECC,
    inout  [17:0]        M_B_DQS_DP,
    inout  [17:0]        M_B_DQS_DN,
    output logic cl_RST_DIMM_B_N,

// ------------------- DDR4 x72 RDIMM 2100 Interface D ----------------------------------
    input                CLK_300M_DIMM3_DP,
    input                CLK_300M_DIMM3_DN,
    output logic         M_D_ACT_N,
    output logic[16:0]   M_D_MA,
    output logic[1:0]    M_D_BA,
    output logic[1:0]    M_D_BG,
    output logic[0:0]    M_D_CKE,
    output logic[0:0]    M_D_ODT,
    output logic[0:0]    M_D_CS_N,
    output logic[0:0]    M_D_CLK_DN,
    output logic[0:0]    M_D_CLK_DP,
    output logic         M_D_PAR,
    inout  [63:0]        M_D_DQ,
    inout  [7:0]         M_D_ECC,
    inout  [17:0]        M_D_DQS_DP,
    inout  [17:0]        M_D_DQS_DN,
    output logic cl_RST_DIMM_D_N,


   //------------------------------------------------------
   // DDR-4 Interface from CL (AXI-4)
   //------------------------------------------------------
   input[15:0] cl_sh_ddr_awid[2:0],
   input[63:0] cl_sh_ddr_awaddr[2:0],
   input[7:0] cl_sh_ddr_awlen[2:0],
   input[2:0] cl_sh_ddr_awsize[2:0],
   input[1:0] cl_sh_ddr_awburst[2:0],        //Note only INCR/WRAP supported.  If un-supported mode on this signal, will default to INCR
   //input[10:0] cl_sh_ddr_awuser[2:0],
   input cl_sh_ddr_awvalid[2:0],
   output logic[2:0] sh_cl_ddr_awready,

   input[15:0] cl_sh_ddr_wid[2:0],
   input[511:0] cl_sh_ddr_wdata[2:0],
   input[63:0] cl_sh_ddr_wstrb[2:0],
   input[2:0] cl_sh_ddr_wlast,
   input[2:0] cl_sh_ddr_wvalid,
   output logic[2:0] sh_cl_ddr_wready,

   output logic[15:0] sh_cl_ddr_bid[2:0],
   output logic[1:0] sh_cl_ddr_bresp[2:0],
   output logic[2:0] sh_cl_ddr_bvalid,
   input[2:0] cl_sh_ddr_bready,

   input[15:0] cl_sh_ddr_arid[2:0],
   input[63:0] cl_sh_ddr_araddr[2:0],
   input[7:0] cl_sh_ddr_arlen[2:0],
   input[2:0] cl_sh_ddr_arsize[2:0],
   //input[10:0] cl_sh_ddr_aruser[2:0],
   input[1:0] cl_sh_ddr_arburst[2:0],     //Note only INCR/WRAP supported.  If un-supported mode on this signal, will default to INCR
   input[2:0] cl_sh_ddr_arvalid,
   output logic[2:0] sh_cl_ddr_arready,

   output logic[15:0] sh_cl_ddr_rid[2:0],
   output logic[511:0] sh_cl_ddr_rdata[2:0],
   output logic[1:0] sh_cl_ddr_rresp[2:0],
   output logic[2:0] sh_cl_ddr_rlast,
   output logic[2:0] sh_cl_ddr_rvalid,
   input[2:0] cl_sh_ddr_rready,

   output logic[2:0] sh_cl_ddr_is_ready,

   input[7:0] sh_ddr_stat_addr0,
   input sh_ddr_stat_wr0,
   input sh_ddr_stat_rd0,
   input[31:0] sh_ddr_stat_wdata0,

   output logic ddr_sh_stat_ack0,
   output logic[31:0] ddr_sh_stat_rdata0,
   output logic[7:0] ddr_sh_stat_int0,

   input[7:0] sh_ddr_stat_addr1,
   input sh_ddr_stat_wr1,
   input sh_ddr_stat_rd1,
   input[31:0] sh_ddr_stat_wdata1,

   output logic ddr_sh_stat_ack1,
   output logic[31:0] ddr_sh_stat_rdata1,
   output logic[7:0] ddr_sh_stat_int1,

   input[7:0] sh_ddr_stat_addr2,
   input sh_ddr_stat_wr2,
   input sh_ddr_stat_rd2,
   input[31:0] sh_ddr_stat_wdata2,

   output logic ddr_sh_stat_ack2,
   output logic[31:0] ddr_sh_stat_rdata2,
   output logic[7:0] ddr_sh_stat_int2



   );

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
RsTzdiOfx916A3LehW7jTlAVcvtHG19E6eRiu3AeEu+ehE6YAQX5Xi4AV56pFHcrYWRsBDzR3HG+
cexlyjtsuHWrY8K4XwbbhIS2A0X/AtSZZTszly/YpM10qoi6dEbrZH6LqLsiIEGXJqy3xhMaoyg3
qEBGoMbUZ6+7AlaU5OBFA748h09lqLoDdfv1iO4Ke88TwbYuCuRoMnAkS2HmfSTR6O0zMLNtj7AS
vw5Nhn0vXDmVP03oj2zstIl3h734CpCMy1MjLglX1t5T66AfBkCY14ZxW8gY1F0RrDUbXRwZZAK1
hpEfcJ5IuzhpnfSVkGy7a2g9aEIhHNdq6L5BhA==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
hENH+ad+VndDcX4eAhmDi0WkcfbtfpSjVszQ+JC/cAx6Kj/3dSycAm1wfoJ1cMaPcdZxX9Eh/E8z
v4ePsfSq3Qt6bceuftSvuTHXUNbVdQ4ZABy/TWUNpAxm/yD3DLnAf8uVA0P3aEHjsfSLH6cBoATi
dpSSC2gP30jYH+MfkYk=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
Sf+ag2BaqOJB7QJCnMkAkX2ZD7mS/R/9i4edtFskmr0JXLk3AAP8m0iDeRTiu/J4a9ZQicQ3E7Io
Wcsqt5QGRCZhLeOxxSd3XgkSD+LyiAdE3It7HGfGI1uH3KK9Fu09gBlV+Vh37xV0/yJmulg28j1H
C/hzsepOSIuNCHF1W/k=

`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
lutnuYufITFn9KI0i/9PbtD96SQlq76fJl/y1oD7M3C8AgIiSfG7BAb1csNPhRNREjghwXRo6z0H
ZOTEOPh1qQ==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 76112)
`pragma protect data_block
cURKrZD39TvtL2Nn9QptDjGWIPOe9WRoYfkARc41S3yEjLlEhkxkenMcOfcHUsj7ydO8xpYvmOL/
tNKoRynGQ8YTK2gHVzjh500lsOuLefI75yNY/Zmo7j4+IN7UpaZ6Gz5DvBTkUavhyt7eZ4euC27Z
1OQxXMzFVFgfqxpqXS21PipUFppeg18CxxzVZdab8EoyyaGFBLZqbBJ4xphMX8kx96fDFg0tJthw
M74m90rAr6+XDPr1eq0M6dzQTmOuHheZc176sTo2b8oMd3/hD7IbcPs8sxZ74Ivh8orFSyudOu4Y
aWgIFqoG+ieBm1e/9y90OriTz85YgVtUAHBxtym/cWzg4yO9XwIBqvJ7MjHTghS3+YEykz5GtGBo
8CUTzEI9KOpdzpiQadB5H/D+MfkyaPF/EAFLgBumgraLb04X7+Y+ELUEjop8aZQVnS8ymPDm+n07
000XZJ7qyIXGQnWrbKc7VGN4ji6HvfjRNKfBViYZDtt6V0nJMsQiMZz/6bjTq/CuyZuFjudaUa5M
Ma1pdBizpXXoEuj87Upuqtflj7KkSOGOehM1f8oh2IM54p3DGZSM4DwLLJgZrlv+TO9uueDwYkGz
VjYzPcnpQ/s2QZIQ3iZqSI5wrPyGCNo6cF63UfDS4t34c05zt2hp8ksVWUjpMYAIgf4UHiC2aUyl
fD4223ilhLiam7Sd6oG604FfAM/YQzGMrLFCln4c6FwxnLBuUcfSW2uqA2bNbJVv9qjONf79Wl0M
OnYdKlThIxWKlHu5MtPE4ejXCijrW7YppeKfCQA8iw9+cn35P/Ze9ckWZ9+YAj+Qn56+VuXAJvSC
6PC1auZzms9VRnjjsvcKB2jll0Rpy+29OMPuU5eOCG9hbNI6kPYQpiNGTw8FseaY+3DcOmzQo4Y8
radxzJPUSYwlYuFo4ITXPmbSsqW+pVWXZZ8PL5412cyvOGsvBR6wvLSCvea30UG/LPI39LSyds0j
UVI/XlARwI/P/oBDkYTD2awB100pDY0qGXFzHFSi+dzcq937AfkxgxVFuIAfq7mbJvwTKZpK0A9s
RRiKvu0lDP/iFAxhKAYGJMuOudGK05PLX3r4isJcI9LGoHKNGWXElAIUvivDuUKnbkMLRGuRyP5R
jeEuriG5TDcBSOk/V7At+P9w4TVEY+NJCtcJ0nwjFN1sROqp+EldRGwczOAWlMj0Iwl19Qzr+0gd
Im94q+fDuus+zjtqgeFW6i6A4crOcwmJsFk5Hx6TcplHJFg00TuC04w3Mr2s2hVxAyo0lKE2Uxhr
qsLcqtBiPaMDzhX+7aTyNqp/4F5qfMHQffKcsUFtek02BfDm79Okt2Bw23Tr7xk04YG8TQJ4W6y5
FsrGU+IzNDUAbTqTcbxd3nXWPfdFeUSODNEue8UUzQQ5iKkXm2byow6XY6zvyt76fDl4NpHTPgfe
0lEUpxvWJBR6fHbi4zOtHx7j8N7sKRxWyaT2juzk4WvTQiTlgWBSbiUBrfd7OnRz9UBuUH1H7+hA
FHY7NgZRvD5O7nZLM+4hyTlmCCfS5GVLiq50+3JVMV1uV3RVwxoEc0nO8x6v/ZsmhpAWSeRUE+G7
+OjdJGJJgKVjTG4TGsYtNgnqcmRdNj6SUzztPTnSnNl6333GgongD0UsxAo45vp/ouK0PoL2SV8A
iF7nuSIIuGTPFPBGP+1Qr9ZS+OiN6yE8YIHMFQXFm829OICpir5hxa6Z+JJVLOxGTZZ1KmdBilvV
b/EZsx7lPhZaeEuRicwXZLZH5cMxZHXuhs+00La8bc/DCxYLxmCIAJzLf1VbhtVUrXQ4ZBz0HACK
YmufskucUBf/fMAJTRC75J3xypxWntM7DGA9mSecAiUs8m0Q1kJH3dLlfBaD8Df8kqoshts6Pu9M
thz9te5XPQRT0bHlBpbMqjKgga+5Q/Z34/SKJbF87DEZ6OxbHR1nConwZHLqOqYzEoXsB1IFlQ8g
41mZSmEJKcgql6dIRJM7ycbxUJOFJQFQ3KfvykCyZhfmIiAUWuTmUCwnMOW7gQOnAC0QAkBd1sHi
cqQ0NqW6OSKTXM22Rcwu2pOMmHk0DYESWo2SUFw2uViNz4V4I0gko+GG5p357Upd0JS4dgjj8ohH
+8JSAafm66D1vL76NCVvZkPoG0NadVT6PpEK0T00VC0VydlT+CI9SnD4XeMzwtHmYBp//ezb1718
oSGUoOHYuriha407QByPtidi8+Xek5Q/OGxEd2ok2WMZaRPnCikYfBB4mcK+nGgqDz3DLVyIcaEO
8NxWBIyFwZ31KUCzNpxgS+Zbawi0EIo3nW3qLYyQdTGAbZa/SzY0ZgtkNYx8gJMQThSQ2JpJJ9E2
/YLNAf4c8D3UA8tigFOyNEfVUoMYigJdZ0d705sItfwe4+jvpdCzBgXYY13wxFiPlVk1Ok6N1WJn
UO4y5f/Ieni9C1NrQNsgzY8qxc7SYrxN8bqmVhqgLtKFln/oMQdNcEjopizl2ZnYCGCBd+Ni1n67
jL4zEIcRf905zaadqDznsTC0pAIAUOGdvtluSF6/qE+l9Y+Y2rgDkvZB1s1X5dE1eus/1vdZ/Fd/
e7n+AmP3VpGf6PXyJstQ7ha4suksLxNroPKMSrBUocAJZJR/3uXg2BQqroAwfexzncRRKD7kVvnP
/7T158CAGCK1ds96oJg+bxk2Xho804jo8U62ZyKdVywVR84h4c3uNHRFSkEhzyg5IpCt6TqFgBFe
Z8ejJ1o6135is5MurUP2bF/y2onImkXG6bhmM8fal6duhtpzTZO3CAbemj77Gm3bFHrmtQODu0L/
cEbt6l5VEfxHkEj+YCew0z56eJ2B01N9mJLVaMnVypteRLWGXIOUp/J83qE9Ci4+L0j0rRQMdxZ1
aLzCdNDBLq6bsbduO8EPNMCmwlbwKG3nxrA/v4c7ZThj/B9RziJehWI6MHHnDdvBieRvQXBAjaes
bg+/FTvhpuesEsDK9BfUEU3vxc9FeECaQh64mCKMcX/w/SWhsa1kt5OLdL33GhBgH/N5Kfe4Z8q7
UwLCqKvAu/ACmM+hHecku1eU3YsbtMJOkNhNYa+hXU5Vg41Ud73ipVZvea/v3AmjCg+oO4QoyCGE
bSEjvYCGmYmN8RApeVFgUt10ALs4lC6fAALvemt59wHuXUIasTFZkyo9L2DmehIiNcjR5S/6A7gs
12TO1BDdlVv7Joz58n8cHNsNVM72jWlHZIgUv3ddTfRMe8O4dDSzXGThiWd98GisZnYmGrHyPndW
eOLgCkMmoPzjvkOmSlS3ezUuf3xGt2EI7XONUoAnxbeXnOisJ+OFJ+zBI7NMBKHTQzqwRPMOW7fd
3GreYT/8xpXcou85bo3Yth99WtdswcV44VJ8Atw16jCSHzoE4ffL1ZcbOFtu/+ik3Q8E/HYbud0g
c+l3dS13JYUeWWcHb+9TWeXyaBjhXNcBVgt3E2ZQTGxmdK20w5h1sRILcy4i00JnfFkfd9z3AB3N
ostbRohdu+hybjzRkQNAiGJgldOYzE1WQzIXl/Pvle8GGoG0Vcl13lxFNkXZNL9MEdTli5/UmE+/
EBLd6dhWcU2c7yqfj1D2+/vLQS9YiTpRQ4OpTRXGXqCCO5HZ2GOl2voMqs0Gc+7KsJWrWUbptS5F
F5OZASvkuMjLXSiJe1KCreXuACHG7tSj/8rXFdNuRbtrOqwbWAQut/2WoujdMe8P9+GH6Av7dNjm
Der2CG62Dn1a9H+MV4TIfUwo+Ax05FbtVibOnAcgaadN8CPpW/jhceu3xoRDSsW18x8j1UPDYN6+
P9OO5GkJ5GUA/jIJRV2Wx7ek+Oa8KrCKteM3DY3eMbYWRkGUa1sxfHDxoWOI2bNrdUuF+l99n7K4
2xHjK9nFDDp96Nkdv+viA+dBmFsme68ATLZ8aFs5O3MOq3xazCy3yjsRyJkrlJYFD/EegViwrXRe
atHKn/JFTNDHi2h0olvwDxmX5F0JbTJWbdcjBEB9LIRp9tJZ5vDMXWN0pbK6eyi6ji91nY4ysYwE
jAMJE63JJ+NnRMBW/1C8EpujoQTKFNiFlfuj2mfjFHns9NaeWJVMxyBRGwW3tu/sKiy2NCRPd8rc
Yjgg/oMAR4n/p7dHtwfWeGdYHOE/JB5t3mXWQ2sM30C/MP27VjYEBPHbmuT1VFxyPjR/0D+bgpey
sjkaT72kpnxFp0Zo8J6kl0mpDUK6kPxQlu5GdPSLYbikG01HE4WjN8iFVzUoH86CxMSS2ZJ7jnAV
TLYFZShAalXtVzBcDoowTURL4QZY0oIccVivFkZNHKItlpQAcYWZz92M26kD9PdMbq2eSID2HUoi
jlIZ1osaDin4Nl3cSU/CsnmQjSUfV6eoG8p6/cWSzsACJZOjKjq8PTnlKm3krdJaHKEYu5t1weDB
f+YrAOspnig+OT27f67V87dqzppLka9Zc5c+fZTAivPScolV0P+MtPw47X+7h8C58pJa3wLvr7rV
vTfZsll68x//fm0TTDb+1rO+eGLH2R5G3zNWX2hD3e5Pv/Dfy/sngq2Gw+FSS/MdWTQVSniQEa+E
5vsSy70lNTOgG0HJqwsIl9/DobucfCsPIyFqKvTTc1OyaZ6O1V8pCmTRk+lx8OBpodHUvoOyGefx
omkmA22KENigwzn8XEjRFTP8YBecNsSv9v3mbuvo5IotkfqRVR7yd9Bxn7cqB7+5Qj2qJjy9qoFI
V/mzuOJXxFEmoekZqAtbaIXEruaojPR7kZXz9q4nj0TF9tFSXBls0cCwjPARv5ThXejiDmJOHhFq
F6DbBUcfXzDmXun53bSD3JewU72eVE6PN7T723U5WBuNiffjIGZYwgzGSYNzkv7yR1wTNfADx1fN
Fh77YLsZsN0p2XUbEwFuw+4Ge558UZqj/YZLVgv4naAs+9nSHAlrUix7zi3eYTZLnhl+RtvtMVLF
GY9l3wWPgvp+X+rLOcbq6gNMB07YSqmYIf2XP+LP22hE823BXBm0r5iDEfpEPLQY+XzJeLAScTXg
dDNPHZAAcGD91gKGfufCGbgq7TtIXQw+UMK/z+GTzkr+8sPO4kdyQojaJ9HxTLMKHmHz5BZ+uJXk
YLHMOGufECJbmrFzL1PsMhssG/Z0wN35+qRtP3j9pgbIdYawjcOlindXuuzLhdqOhG1G09jO7KB1
G9DTL6REJ434MUnmVZiCUQKIQQhChfv1RO/i+/lG8yYvD7BdF+DxeUK15l55dGssgPoQkpXiIQox
SBAapfJ6gCZImWBDLLfn/lPZPBCnKZNllqtNqp4HihoALOexxGycPwenG83Jkt+A/C/ULRzC1mQd
AqoRfCrtp5MAVNsYoqK/XJk0XZqNBBijd34htJh3AAK+QXw4EQmwMXFx8rV+SdkO50y1aPs9pFo7
P6mGZ/Q910HwxgT3Hs0z1NsOckgjf54ECrH2STufH4IUf98ZPUrb60+Giw1SKaY7V+0ZwWFKKIaH
a3ll9XYgdn/C63PdFuvbGV5T5SctaWToWi/Xj38Vv4mONaK7J+qBS4LyDq4Lp6ZwD9/ZqyZFonI7
jWa5igyTAA5w6Y3jjbqlfX1Qu3MK6ybFVDPytrRukr6eNNabP7xl/AfXpVSc3MidfPyBkMmtp56u
PBF9ggF7vAMp4R5AJQzdhn0NR6K1eXMkT1cUVtI/RYrbDwqy0JtliODkBm3j4cVflKRcVfxphNxA
u7TYL0W2g4NujqvYjH/oI0ewcA6xXhPDrO40AMn5YENxA+UWxgL69tPvUJYQb3IjAuxAlK5kiWHz
haU9r77STaUGaFsnoy4FMuG6Qtf3JqY1lihpLnuwVpAjylspBJiDzEoCjiulxt2RIx6cd8ilJ0yr
/jFTNPFTcR9G1nCzHLEPpCgkd7ukQlbCqBycKkfM5GXw3cDtSHlAqQFP2q/Z5bbzUrS4It4hXiHg
/wwbwloFSjvwNlPqzSPCOMkrTlaL07VDviCtyZBtKmxfCRSMCV2KP9bmIt/Aauv8WXQsPu3XY6C3
CFXkpP9sRvnH3BeI1QvvBj+WAKnCtI6GnI5tldFDsPbj3LxFGOxTd9vI/pER+J/l4U6uiJnp0Kvt
O967ol3vonmPK64pJi6SY0qRCsLtFc0R2PEhHiPr9UMSku7h7c6zMZsEaMxCIKsWFN45E5/UZ4kH
RivCbHXFDxVF0h1mgW2Gv4dx5lT4YQg1uEVXvu6P6Sp5wSfxJUxzkAomJOSzVqoFBqUpEE9lMx1w
IyZ7EA1Xp3WHAqR2Y99pmwIzLeKoL3iakzXKAueOWNKo6L7YKos6VofSPvEv3uNSdBxrUaAKy7AY
HAwmArWfEuconq6ul8rNFOACgWn75BpfcKTgntKrwC6Dp3j4PyYGSvi2UJ+IrJpqVZtLLFlfJwco
TT+ApL+LzU6nX7tk7Pna9Y/hxb/32K3i1ZeJOLPLoPqYpB2/z+FePjtB4XfPAOIiGivQpXj7gCYx
qyLEpvgnxcKA/ybvRm3enMpdY5MD0wUFgPJyBneGsJL8uGnKy2ZQXy27avbG3iSJG2nxa/4KvGD2
xNSxuhdFoPWuexlFE9JrcZzFI/SuZuOf6OX1X04Ia0OH9ZvuXwBDMr1lqH9vca96dmC6QeSHWc0a
aw3Fdi6NEeKyGGL+QPx6z5r+ZHBupNPYMhxdhYtzRBdPdXyKB3H7ja48HIOvovY7QgZcP4zNWeRy
2eFELrUXNDkoaGWoEKbuHYnsmYiFyQ3+H3Xjlpl3CSIOS0xVqVpSus8jhchyS40rga9g7bhlP7Aw
HHA+afPUnK19c0qOaunYqeOkIrU30yHl65xYkQp6qvv9RqlOa/0AY6AZls8DpezoHxcFsXRdlf3K
48dJhlJHXvds22MCh2Z8G8+IKPLgY8kUOVt3mFJ2Qp2RikgxIV94FPhxA2fQSvP+Ts3cnwrsC9Vh
uXPKk+wvVuPoQU+8AULDF8nnKa1SWagsbxf5li3wPCr8yV/gdRpHV8jaMMMxMr3Ez9uLOijGbKE6
zBwUgGl3+puVtbc7rjhpvQv+ImaSVjJTmCOhLPOHeiqW0p/Eax4Pq20j4xwPDpTKMz3grY8EcyXG
fOyfPJyynmUcFFAZLWAd0JPbdEQCEjBm67KbfN6jbk3CnqYlTBheMJB9tCPwghZnGjS0oN3gdJc2
yz5nVR/Rsa7bl4oAX21scQg4veRULHCJ33kEh7F1VEesOutLoNg7aQvx1JZElZb6CwGa9llu4xBn
Y9c/1Ay5oFMdwyWXRTzDPwHn66uk49gMeB7Son9tbMnzOc/d3TcVnE5v5XR/ve4NgzUTp/u5A1VB
cKhr1O8xd0QlKZVb6G7O1x7qzhYQTOoaN9icYRcrAKvuxR+1TSMf90A5EtYEar7uH8yUDxVhuIqs
lmdPg+KsKZ+QiBjuyY7iG8JcdP3rXbK9MqPigmOSVc/zJ/6DWeX1l7VIW8i9E1KHwXwlXbgfhUz0
i3BXZFA4qN9Kz47hLwWXdc7xhRfQ17+LdBccREFxVLL0Z6qnXyp7FfEYP50slrkJ5pJ9aDD96DPC
wQbzdbV8TNy8Krs4DM9EXrp2DLzas5o4bTo28rpQS+bprlUvKfyKOqymUn3mCfaTJ1FljR5wNvC9
WWmO0tTmNo1pSQWv8FTXVk3+0g0rHy5tBqZdF0q0AszIZeC+38uszkpsRYQR7aVdMSfEY510e5BZ
ecdS8XkSUDkS/RRVieeRshxle3gzXoe4Otsa/8sNwZ2rvUA4Z9Kz7bbRI4qpm74jrrFS4TPYtIal
c+s8gtKK053VQ0wUsYdemIIWqtTac/pj7J3MUG2vLxVyijHMJCEbUvcdSJSW9ffNjx+aqGkyVtsP
VYxr7Oy7dqf47bzQ1lJXo7gTeV0z3diRLfXKu2BCKAPHtshGihPH7DQb0qfcKqoZZXz9ae9fUgo2
8gS/ykWSZQQEYDSTte8+WF3YY9gi287oN9DgLRElwLt3lXZzEExmKcyJxQ3Rc9/C9eXWhi8rKHWe
P4IilhT/80NlXxzMQ8k84+iuDTg8BHoEmhEZ4YiOVArVKAo/ewKbE0dNcsgDCuvP/9miCJhsqir5
3uZv9YvmtRA4HLJEpcU9exYaLz4nDcIxbL9/JWjpAm1R1Rk1ERz6ky0YF2xPzyWMTpAe4WZdkUKq
CmvW0yrk7ZESKInGtAZYygKJxsgLiBTZ7I0aEGAISm7SSDlAUuoUbyaaizYZSGnB8LzxgvYb5mHH
iJgy1Rq5j7fnExHKVj46mcpaqPRFi//rv6jQOLEm04i5OFpOrKDxezciNvSOc2XHf+XxH+c5PPxz
9yqU/aZQP8HPIh9EFbaHWp4axIyqY4IlGO4wvUrlG5czpSYq/OrC0g7iMeqGxPQQroQanwfSacbL
yqkKHtc7ub5mRFJtOG+qMg4FdCYuVWU6VO5/KTin2hPbkqZqEyhyuOKN9zLMfozEgGR98VEAZeYp
ASME3rVGFLwxdVpkZbE9oEnlzugeWsDGI7693cHccdt2/otinV1VaNweYCH6LnRLy3I1ZRfLMYuK
Ofubj81yEVc5zxAID+LJTwywVtv8t11qSUI8r/+9ZN9t+vIs4Jy4LauZx9JHYLwAPhbcrJoS5qXk
vdlp15oYKeLk71BzLZKtdy2t448sSZKQ78GON3Xmi9j4+bQ1SlxTnhdAz68b/JFpG10FyTkTa096
60rockzJdxBMIDjNmGQQFv0RcQH4vU1rH5hZbw61EfSHvn8sRcFtm3ta7Z9Zh5Qf4HPen1nZ67PV
oVDcPfKZJ/XRHl75R5KKeIa+FcX8ZKOlbwuSjPfa7i+eh7i/XjiWbYJoPqAi0FPO8SxpaHIcdb7i
ulWZBhbhIW4jtWpGwmZCT4BUaJhcTj+vlw03+3GGoMG02QavBtOyRzpzWkcv3BJu8ixG1zq97o/m
VocatBCvHEy8Yj9pGbSUoKcL6LFd1hQjMcawtxW3FHLndlHuhnpKc2X6TYWD3RYWAwM2plyGmKEp
g07zV3Tfg+6HYI4PjMa9mY88W//Vpsct4hHD29sxG5kcnzdWVzuxqj9YLRQywHLPLRo7/y9PINgT
My+7PFcgR4ZZ8oekgSXyq6BGesVaNjzBRr2IPIq3ZzZSZLrp5z4NQyydDAVEjYX3e3MQAI26MUTo
UmJ5DxBsZyOxOTZj62oiOF7ns1ym/G5HQB4/WbtqRuS8jgKgPVe8T2NutyPQaSLvH+VlJWiZlQcX
r0eWVh2/0Az0skOgFeforGMtant31+O761ERfGmauE4lRmbtF/W+1nuiA62yzGjJPr+K7jdfIleB
rANW0TIrqilbayxuoNh3TSoGA2Fd0OGh0y9CVWwGhsfnuYRaupTWjvNBagTUXxw6siKA5I8Tg3du
RS7CXLcVWsM8pKAsYOGL5PWjrFM648Os3x6fl/9MbJGhq4F4wxiZ9zN0+q7DzrH48bJg+8XsD8e0
aaUry1Sw3D/T6+WkYUXYrpfjVEiUCB9Jtnp2Etw0UVRk1XwPxmylM/hDmbzjS0TeWqXr3LUkHBov
Iptwfh2K4+KRqKZpciagDev5Qo85uWflCF9Rsr243c+ehMSZX9gAKkB5JWDCtVhMlzR47maGThsC
TxUvyyE7emPFKGhQ8H7Q7Q4tYWy78kTcYCvF3EqyWT7q7tSfgIamWhC/CE67p02ZlH3Vozvzng7/
Y8zrrp3xdIAkYrgvE7JcHpqZfS3S+/q7Aosrj4UPWSFrOi6GCj2r2bJnXXmZYT3ju8Tseo1il0kf
hSu98awvaS19gPhhiN+3Y0ChR/cPM7H7KdnEZssfTahDMBCMVDaxup5IOvKsI+rwyuKCoSInE0jT
KiZKvNlwc824rtad2MOsm96+ofagfkAGv00t6oA65/dZWeYjzaasL25I5VBK81lzuoUWaEKnUcN/
+YH52RBCZ3k/TTHBfK1Rmj/eb1XctIIENnT7UA+a/SZoss4V2aVg8nbsVN9PJwEnbcY41V05qF0e
/p+vyEqEB7Wdc/ZUV0iQTfjxgOLc4UY0vmV/WRKQopuaGblR0NbPcCahE/vqWnVuV+0lnsj0GKKk
7rEY630Pt6kGRG7OLVU7H5322s9WKaTrFV0ujcWk1RPMN4FR7wiTY/fLfCz+jALJnoAfmm/S5oPK
RkSQB+EUMYufk97GrTz1PVy5TDesJnvMGw5sZn7tyVQZb3KmEKr6+MTQSTDzKLJTL7oCIxrnOde4
jsoEazW4/Jtu0KUop0eugSJVXZZq3cDmYv/jCMolGie9LDOE2G7q8HLt9JfFegNZmAClwkXn1RSu
1SE3OKSVtsxniFl+UBTbbAqjTpltknI3FNZXl4L4jhC4Ajqc8JTXGW71HwmLwq1J8ZH3JkynTXQt
u27bXt8Vxj7vKamheZvZlsylfWREIEhvoU+I+Wq+kr4KYKhaxjoGB3HzDMhJpEPapH3/Ky9MQLtW
n50b50H63yjyqpe0OKXYoJ53hmH7zyxxJcQuj4f6PKYOM9kXLBdxg9SQaiN58WbuIDYnM54A/kIl
HcDIiSF5xcUrmReXFtMr9y5xSZvqnC/pNlIqtGtTE05f5nalosP4xF4CZHKmOVM7gNC3nrg/LWVC
3LhAm/7C8FNKueHG5aSkDBgAtYGAY5ARWXu4SveoBu/gfuF6fdfYFlb7gjE5zd5BpMQbPxMEfq6w
EtCUIMCorLLkJUbb85bzOJPx2Qh2R9NAPHkN+pmFPExo7jbJw3YmqtQOAhafIq9CRmBUnbZmmnmj
QxzyP9RU3Q+2HnEjU7pkG/8/vfTUAiQyZbW/quM5Or554+J4A71vDi7p4mn3CRgq1OnGXPHeb+Gh
OzYnmsPTB0QvvfXfFGPN0FLY+x06gbGIF/LSUQtqSnhjXDVgcFxTEeyGJHDacC1Ugya2tr2l2aWj
K95XyXtKDgYnaz0Iun0QrSKQcuWKhomRFyFrPgAVaMxGXx9Q687mJ5hhWcV7KxmMFrNLvfXYBQc2
t2LPYMWrLK0lmmU0TiQn6o2afRzlylE+26EAdzcgbWLA92a2dNY2488OfVAdrMLy2/3GVmhOKNKT
g/3KKPippiIY7o0lKwp8NqSXFBA+ewkPmLEQSXKmIslr6TtKORK66NfV55pCGp2Cme9Vb+SbEKEh
ZPFcoKrJCEAmSY7p3yJFr1/8T3gA6RGGVvplsBff4UUozNrhOwJCMaj/aCINpwtSJ2ulgwQl/2fS
4A3qX00cS1wAeX5tkZsq+pdKJ/yzgrCMutEH2uDvwbGzrW2F1pm89MPvjZgDsxJbCkKjuf6Byngo
hm9Qyef6Tc3CQz8HUtAV0af7gFMlP8027e67tefYzyagqS/ZMhZFVtjMERSdx7xfrn8m8Aqm5XmI
Ek6t94IzQAnl9SiNxf3kSLx+/KxdmSg7v4e2VrMY26dPYDwgWZQEWZbilLJ3EWh5+bmIgOFeR4HF
7VkajKixD2DTjRIGRLisiYR7YSoONSGd9lCe3cb+5oQgunL42rGLQ3U66jLxIr4tOQWa+KJ/t5DG
6uhYltg3QMSwbo9QjxkE8gSDbBguPde3ocMr1KJJqGFGa6r9pDd6zvRzzBjltfZgjEWqtkFMFKmf
X47pKiCGcyRaxnNd+EkZilQ4QdEP8/3j3SXVDr8pwvTVqOHdOqRiZQwFRd6dSJrnHgVchrYumF2l
wnA0NNC/goijTz1PfdRbMg0EHhiClaXbvFhHcXfnKvX4PJDqvIjKFvV5fcSElc/rMV0ifrdyFZPs
RQPYnu3guIxIJLmUGxzhUySoOKAVoz5+MM+sEk2isaAUU4P3q/f+7aFLxcTTVJSahqAypkJvNCiv
LaGNuExJRd1oQ7AjxboHqZ47dhoqD25hTRL8mQ6KU8GmTJ/ySnpcbiGmj9LZpHKU6DP1p8bCB/xr
NOZ5qc5KV5WHJOd+1LRpDevGMKY2Ju5+1Un96Crke6OCVzaDvK+W8ZZPU05nNOUcTngXlqO9+vnt
YCiCZcbMs2aYPoVFdR4LUUN8VyYpZpRT6xpefGMms0rT8LSZv1lLuNvZUbPsD8b5aLmHkYxUikQS
0/6yAj3GnxOd3VtSiTTexVK6gQqUF8AlwMICum2/TwVzZLzX6VPX0Nrvzkd7UKw+Tt4uVqgKNkre
GYNAt8a3v5z+UzZyzUOEw0qwM+9SpihDCkbfKn4bXPxKEVFItYQa4PEI2MtpMF/a1LSVDWQPAi5x
ZC1Cz1tuEF3XUDleG9m7azAycNaNHuhZyCENcPF+wrXd8KamBLPs+nbQiByAq+TEdkKTidKJGb5N
St7SunJqhlCM0NEr3LP+B8z0sXqSxZ9laz6a+iU2dbw5QBBGRSClj0FAAx3z1gRs1xR+1TCbMllk
rFGvCB/8wWObcxzKPFyQCef0/qqyt+mQN4yJSZg8xT5LKcrDRVmi7UZRQZpROV+PaKwT+1E6PgEU
l20mgKOxBeeCmiuIYfw2ThWhGslfJmYS5rDg+SF+DUR69HnWd5XY5UPhl5imFVeTZjSLQ9Eq4vRy
odDcKAHzb7CAxy3hnITarJlP21Du6JFc41zDKKAT10SYRVav0C9RhK4GqVGuxs4zwZICIcZ1L3us
gZ1Px14sKSQ5wZOTIFF0MU1G+bajStXvUC/RLZcYwaSIwQTMXvRdZw/ka2+S8ocV0vdWjV6bs8pj
1ss8dVhS97H9eIf6gNUnnEZUXGDYwVRyD6VoqI8IxTYpQZ9bAoL8ISxaZwArlC5OSoHPAG7TE+4j
fbwnCt6GMsNETPepirvSDmeb23IN8hz/RwIsICPHYTyWoTUwvSX64pXSGzq4MSE2PkdTdpraRui1
NabIfzbLLtKvyWIbCUNlUjkV4HIH694HnGPazIw6xA0HIGmMNQaOifg8FJCS82qKHyXvUBxK71P2
VtgbqTGVorjxi+NUlwlCqHjX9tsBRsllXeTo4Xie2mv5mTaSSz2NsyqMEtXoWnxM66B5MzeSfEFL
SeZe5dZYDbYvs0UKssbmXRybC36XjAvNMoCS2tNJYy7q5UswSIVIgDwGbPwkZi72me9RMKYvboar
CebVZ15bOXeFeJ7h12dw0JlGC0psTk5Udcdc+W3mv1rZtHcEdWIQ/dEwzVRMzOft44Zr0fU7OJp3
a9vJQIjErfQ3o4omzao0l+6LkT90R7vDN8fQDkLNdNSc3g/ABDrHGg1n5JKixj7HbknbHkjPApp9
3eb05ixvoOtDSs79U8GGy/n/d8j7e213qa/Ty+vSj/jnKhKR9DRnyEatuE0Z9xNPC2RNdQhUC0kC
gflNKe8duvHXBIuGf5DnNmyJFzre1cdiSqkgKtiXMWLdSIiygG0tmz36IAMiyNushxbAt0QpQLt+
odr9HdRAZ8gnIaRaiwwddME8fNDcUYItwP3mrfT/1Mqr5vGNX1RfVaOS/7mgBIGB/3sf8QhJJ06Z
IZH//A3e7OiLGk6KIGWfvWmehYjkVeDN4E9I6+Rgbpw6GutCLluyUXE6RnRtE+d6CC8sL3PouIXi
th2H/IcHGx6pmVKsd+Lw3vfhCvwXNYYtcNrdn3XgDvs5v3jt5AxeXNJFT1+GZdNzBz3zJm9YuDGf
D9NS5Njzaiwm6UMy9hpTtobILNYTGsAAG+RnypzReLdOBHWaydlgFsbyJQX3q0yQ52+mzVX05S7F
i9xD1MVkkjQPO56MZ8z4/xur/JDbFakZqPfFWPdRjzjPTJLEOG8B4vsmTygdNNP739XxSR9B7daB
/WYpF01vn2t4T5W5TlzDISxkFnszth1QK1lEWU673BNatdJ8pWxeQsD559P2YPrv7xZxSvX5933n
GvpKmBE7zueagCTOKwy+W6oQIVxno22lUw0vZM2MTgW56WHGG5CmW2tyDSjOG57MzcIZbV9ac3tX
eC3CBpQoJ8X60gu9Tc+pEK8fOAMFfvLAv1aD4G2W0AmMF057XxTvqP/UEprA3JhWDTQ53zDTIO7V
U98c3Hx6dTCWqT8ElyaH/NPE0lfnooHDq1aUVrqBHuE1UoTJDGcgh4OmqSxcRxYnL66GpsFBPyea
2j9YCav1Ak7hVlj3WNisFPYgZYieSzeoly5eVceKoV/Os/FYYtnahELgXfi+vG6w9tdJ4HVNNHGb
BjLjIv9whoyionK4z7PWqQMiHIGepVBXbFYsDTEKEweHnldMWuSYhxLyYM1k1oc83MxgaE96DVcC
ywaJbIfRsz+aT02MxshwG5tHGVb4FOwcwAb5f5FiRXtRmm9Obxr7K+/GLhliS71TrZH6YH3d8chy
Udg3oCNSjhEYsk5iN0/MvnPqo8H6Pp5aFLGXEsxz3vcfXAGPuUiY90echUuM4qnDXVIQnO4MeyUJ
0iUA0d5pIoqb7/fDh0MdiuB3yVgpfjhROKMDX2GgkKIX1OuLWHLf4+dtepWJd1EaH9yqVsvlbj09
4Pat+tN67Cmb/moe9jJPJ5qkJz4MQMhywnsra7LedtvDGtrS5gQnCVUR5PqMG0ZWVCmRZqvHEIaS
l0Hqzw9iIlxVzE6KDOtKTKBLjakfWEUs240hqj392pVaD7nLyKL5v84X/njy+pTb8FxyR35ALh4I
CGAJiGNUKNeVoZLEfnBOM2WNNTjRmVPfkBe5Q2Zli7ixi1/hEC7ehk+w2GtD5OC+8hs6utFqAYHn
X4gy51LxoYWl7JVnTShtbuDj5W4Dw6R6D3AGjDADBbYGu4fu7KcBfcuuCMVcil7xh/2z9/IbO2S4
KTDMAbxlQ33wYCBEf8WmkhFfff+ervgPTiSOR13B/01BvVbZSyaPNpYNcWcHjtpA6SVkSvP7wdQL
rmRMysY7Jhnh4y48PC34axA5LCDgHlkFjIGyjVCu4zd5R4rn8kjDcavjmlEwaIthm3j4/f02Pu5X
M0T/oLyFluvISSpYTEJDPFGiJAWQ1wfw6v9fo8UsM042nao71PQJxp4VBUfFMWi9MWCCOhDzp+3J
X+LlIzqr1GwRdwfjDZtGraNbLMeMXrgPQd714JBKFc8DZtCQ7vpzndwweTLJIcn1ibdTXu02ACGu
Ta5vh3mE/v2fLd5tema12bJ60SOXddUCBv5kHdm2hBK9aM5DBav+d+MVLutLYEGmnm95MMTWM4JZ
xQOBvdqWKCT2Ghe+9FWJWyfgoaoB1lPwgWsIsF19CVf+piEb+UNqxRtsG7Ikdz1/WInvsSajlTYD
Q+N8ENotGYn4Vdut/r6+kPbAMHmJ0LeaKVCz9YPBcjdvA4P5NhIWGjEvoijL1NL5HC6QgFMvEwM4
dZ3dG7Zj44iffpD/AaNA6ZnYEOq+TIlG9gkNyUvODXcqmMkwa/4LbWRrdIgn1eeSDIj2mAR/Hy6K
a2B8Wz1ypfdDJXVrO97aQT2eS2nrNjxXCvnmfqT/KLwk6iPEO7YAjanlvISu5iwdA7Fe+UJ0y/Vv
GTygf7ew1+k+vXLKpzHpLp/Dvv+jhwcfB31qmi+SpP5ohbnjyXcHILQhRPM0s97FkEsZFiqic2Tt
EiW6MDfDjtFBsShWBvGi5v03tCfUGp1+U1DdumWzxphF1fOFk6I4aC4PxhA7vrhqIB/Ur35EJAy3
A2G70WhyYWRBtivtzIgnolPRf1aXVeVUl0N3xplNGgcoYOIABIHVYMhtQUp8ZGJXr6FzR89p2fs2
mOl/Jnw6a+TRxFEPR1APj0I+t4sDRlerqbMFFQ/uk4cyK1O8nFe1/nDkUnTHWwppHVtpOPdY2bL0
fuxIDyzohWH6v6gVLMrj4jXgy3Mg4B6EXXk7maTmK8uZQUQwVwCwThJ1eITRxi1Hj5zwtcZBMIUJ
5MWkx+gE4pOUYjaMTqb2HAWNpLg+t9VnijQV+FRcKmxGXlbOjY0M1XYRBw4z3swkgaXz6s4vCD9j
I3QS5gEI0jf3KaZ8nogi9mIHoCqQs35ZHXWgeTn4FoQ0LzKOXUN6lkD6bavFK/EmYU4R7MituRKm
bDHBUSy7b5SIDmWVWOz9Fnymf7uXyOmQRU2xmhp5TGQNfXF34imWF8Jy7twp7aTJHmHQNn85krQY
5TllA34Tu752tNzRbIL1gDse/YqvDewHDTIPH7dxIOHGTv65monDMaSvU440vxt0tmW87yvN0sYL
7YFJaZW9IblPcu5xZH3FSkqzpNMLdCWMsBWkc+LkRNJWvY/1mCL3MqRGGw0c14js7KuMvYVV6JUn
Zp99ZIeaygih1KzcvifkPO0+2USwVHO0ALEzdn3dESVhvg7NrBugloF9Sy1c/+Q47yS3Uae7utLn
EEbqdgPQtZ0Ixre2tGJctWbQkvStiL6yRQxjbymtg1y4cJdAfOuvKghTFOB0gvd0nTqrYQaDoSZA
argP9MdiPleUePf44DrAxb6WPS3O5XY5Z4BZEnyw+1Bq69Hvyv1+4KNoS1m05XfSQb0nUKNVutU6
dhN2t52AQ7HcdalZgjzLnHioHaoMzkLgH7QdPW5gxXU5xzRXjxJ5xUKH7NIyRVaR0xt/u3vJ4gz8
DOnU5RiLVsnxotVH86/w1i1mgoy9/5U8PyGMUBhSB95Do5d4boANrzsRCUhCYeA6lT5Sz8eS0Ex6
4jF9N5CEM8a+vvDnZvHdaa8GzHbt/ABs0Rjx+qshKeshUDLcYfy3Dp9GoVwHfD5x1xZrJ4url48z
AvC8IazJpYTItEe7hUPkpobRq5bhGDTvPAh7xKcYmrYVihLgOXXpBV/CRNYlwRMRSW3oAChhu11n
h6JfbEdB6nbj4JbwNp2t3GB/rSmJiKDJzQQKeCCsH/YXD3Ks+LNMSrAA7A3hjKkIM3iJ4dvrsOnn
zx0gkTFt8KuQ/No6cddLDR472uuiYaVTW69q02cUMw36Yucf6WxBbr5WHhyIWINOgqTTJCfrmKCA
yHo67eU7GM0+/oIbLBU+CHh0NtU1iHfYE5C9UxFoGh4874Xq09pdBDGvWNQq7Tc+BDt8laqbE6IX
42uJ4AR2TLej3Lo5ubF/OjCJ3JFT6c+NX7R8IZFYyq3v6ysdOvtgfoUIoedr58GTIIqJOpxsiX+z
6hNqGhpS9tNgZzuWv5Kv5WeLETASpqsEPNB6qm8b/u1GH9E3Z6vEMAR1AlHQHalC8VdW0AhG7pSF
83CSqBHdv4buJYsA9T/ntONGrSlROwgPTu7qSLjoxJWivJ0T31fIhXrPAyU1UKLgOTBn7DCJHzLc
RoLV31SMoZckts70Lzt0armbbbzBGAS7BWOWHXpFdjlngrfYd9sx9wJgnq7+5Q1+KpmXNfEmR6YM
+80WT8MM/OEJZC/7bYrZIBFBD6A9cNHJ5XZiLc/tB1RwliXg4GDrt7BkUHxtQTEI0utkIioHP0CO
TPPkQCz9V2QSJX056M2YYoHyFNGfR5loe/CZlIoRPglkbuGmfFPTj+GYz6uyhUmLBJewYEoIxYbm
4yHN5jqrUh8maZDX5KMU3VXX/BGazfLsB7nQWFZZMP3xvu/G1Lp5zwpTxObiqlGvKXlihYICaqo1
aGc/OLUbI39/8Wgj+U0f22lu8EFv0kzJi9TDiqm1gRt2UqCU0xPcFLyCBEFphTAg0QgcMwYqGu4B
YiG3KSJGSw4AMNGWaJPUfbh5ChZWsed/AaHd2J6LDcDt6UrICo4efJAeknnRNhk53tNp45PKOvCJ
xlZtJ+3Gy0IATPjo4z0lFG7b6avKVa0T9TP6lFvfKWc555TeGa7sYBCjt+OQjkZC4FeP65erPnt8
Q5z6WgDhtlaz+tmppCkNR5c1t3XwwR6jXY0NSi/V2xtP53X4g5Ds3+G+Sy8r1moeeSgFg0S6Sy5p
/WFAbJzVXDrzcFZ+5RqwaRGH5mNJEHIb7qHls8s9GmVHiuzcQSrf/l9i3bMapX37xV93z0SRcZtJ
JT9/d8dYcbkzvzyW2OzCjlur6x+U8PBABRsy1zYYSZQlX85bmIzDyj+RJOuVg3BbebnN5ZGV/urc
mGB9W/KQPHnnreVXtDm+utSKIIAZgt/Dn4x2VKl0Y1TZGdOWWA/0JeOqTZV5O1hOEsyou/vmLj/V
Sl8BKwMyjBvGxX0KsZBF9GkyxE0IfD9k0Dp/4m7wJrgxV0yt+JFwmgkNsIntNCjP84mEfUlTnkgq
dywjPxkAQbu//COVCyEKeIAWhuy+K+OJ1PMgBBGx8XGdECYrM/qbM5a1cghMUQi4/sOGeyGBUovR
mWwQEBhC5y5lsktwnfwjcoz73C9bhTkNFA0l1j7aa7Cl7+e37recRTV+ujLSM9nVGHQAIjmtspka
fA3ZGlTBCNuQJhctsT+cqxAdWWRg1a5i7uLcO9vSK/W+lg0RBzavf1kt79s8uXOx9VQ4CCJKekjn
Nia6G+r5YVQu9L6fanYEOOlwkj6tBcKVE5O0hQQKh11WKS3pnm190VJ/xx4L0vxL9PHwTuYSknRP
6CcFwMB3kUhZDbqU67gOguaepneHNCCDpgCNI2JPJ8GSuOqQZtDRG3J4x/CYxAKCkeCi1+UG1j7+
Y87Caemb+ID9OR07rxXat6S3xpBM6gSanLqTCmc6zP+vsRQibaPrYHiE6f14KPtRhyyPZQvCd4zg
3xHSVFVvWbHKfFXPWwLjQ8OjJSGN2tUXHGYCmGDl4h1R5kO1zamQTGg0sbDMAD5iFsL/hPf7CLKQ
dy8VLFgtGw0+nAsXv59chmOVcS/KCppRCOJOUhEz78eWCTfTGnwXWHJNd/5Sp3CxFUUkfb6Vkddx
yqwDM4X0xRRuunh/lk3VMAD2YiZlH31qzW79dWXDGx3YeNbTpVjCoGNrMpiH2O7+syt3dx2PxnOE
eTcJ0Uc98jLRG7ZtgywH/m4r8vFUQgFlJhhT6vIfwzXB6LVusW3oyyMPn6csjJqyBN47P4HzyK3W
nG4DEn5zWj8r2MuFBMAfZ40+krlY/5zKeRaKgybfZen1pFYJBHseoUc0nmgqotK7R5hwsGP9sFJ0
fdwuzfcgKObbsEhgUJNq+yRthZpdMeMhHXuXIcREp0BrPFpn78gXr13JWI3XG1PPgAVlJiMlfUqy
2p4RsQb2e7GHsTSDs4kA7ND67RXXGlNSiTV02zl0hyu2s5YxRVftxt6Ly+fy05n3MWTNjI2NW2h7
q09f+th/dLjDYcT1r2EtWEF5dPNOelFRnsW94f9/JthzPxqgnr8O7RcX9xs+QHZRBJXDT1ghagPx
z4fNtwRk4D76m4U3mtOu/Jwz2KJ9lUbN3P4uHYGzsNC+Qh0WBBRW5fIX6fHRsVDpmDHIH2dhSAkC
g6Rv3mRChlmm7NxggaN4MKXdvAmcdrlarHH/7OxYlspdAuH/CyZH0bmu2s+qLddVrEd/9xFy12Ex
din8V6zC5fr4LlgoAq647sa3URzIYFahotY8d3tDpmwTGEU14uRfOSqNkfPhAVg4jud02wWvdQ8y
RBkNhVlZnDWyJhTuwA3wX6rwJyoRhLCMO1Hk1NygMiwOesiwOCSXYwYy8pQDjgnnNTXmPJiCEHsn
Mm8Cem4gZfJKyla3Hicxa2BDI6vjAM/3BnDaARSAP81H8x106VCh6B9W0o+s9e1FFGjYrMHFo+HO
rH8aNANtPXGXuIO+ix778uPfC/MI50s2JKdMS1q3GmXLP61VDQjagOnC5nG3hgsiIoVYGTUHGP08
xbiNwHTHowVRCK/MV3UB0mBoRdkBnUhVNLgFg+l8vH5NJ8WnSz/OQ/4OQhRKMmjTZzC6hxpsCKqC
uNxEC2JOLlgoUPBS/QQeEl8AVFFNS6cBWUC3HYf9PJM+BH5/K1VyqaONHYuo5efVQfVEx1cr68XU
UK0lAF506EmwtVT0JCVUs2+cwZ/ASmylefsbox4fYSHv2u+J0GlVaBTJdd3NcQexS36BVc4J3zCL
QQ+F9dmpRmxCBJvrk9qlXZZCF+twRp4YcqJs6eQcmPNkMpsFTI7Sr3C0WhsLy32L1eQ6smFgR0OG
AwVrfO4Bx1Y3NmdJAVP6TuzmHD+IgrfWZb8yx958QL6Ac1cTGcqCSRWKZa5/nEtnt294+/4g8Ixw
qlm8KJ0TM0dt2d94vQX4LZm2LbR65oJr6ju7bTwyMsb/znP4dcEU6Qe6Vsw55rwxzK9qglo8HiOp
paWRNZkqOiJkcKUTRktF1dt0PuuXaRF4mY+xiDAsPGUtT8V38hl4WTtI5j1lHMRJXwX/3gavsQcd
C7avrIFWg3ykKtHeVe6vzYyOZQUDpzR/0sZnQmZwrO3GnsZg1dPTMiFmjgJpBo5f8qb94fjHogR0
IWuY8k/SLOcmNrtb9UCox/7eirccR85k+KA81Ekx15jiMGViU7N5sLH8tgqCoyyWSTI7ZcHUDb+9
/1suSTg1fQ46IJtOTgFIHHDQ8QN8JvGYeB3nE331Azb1LQ1N1fer8mzVs0fymdbMufYDscdMBILY
4cjHHae+HKFZ3t5uy8peyFOQ0YoaCGOrtrrnpoeyIl7tm6mkNxP9KufmT/KS/EQ7vNmdZDDXrzwp
TNQhcR0aGvxVgFWX49OBvez2JUX4UVfJ8mAKKX9osrejG/LcDcVBSTT2HJJG6x6oY7D8MgN5q0BX
HwphOJoi89jQlRsr8qJ7u5bfdtKCagN84E3PptB//r7cV4vaZ2pNd/cWq0W+tT9vmI94JNzwzxwp
GsJ+ed6qZ76eq0NSJNLjvO9WTJnTExFmpJw8gmOcO0Ihgem4akiHEX9H0pfW2aR7nQhvqpbsU+Jf
ytABbOU8doiX5CMIQNd1nIegRHFAFOW/TBtWf0QgPqy1tY+lwDvsWGjeD6/4+toyHWS8h8UbyYb/
8hTDUrjfXaunbYEPD2kC+4HLbrim0Ovw2SlVrf6s3kSLVkXMDYg5epYzwLMmdOBRNoGkl8sjck22
ZUzcFeQqEK/xEvvpBMQbXskwhN6vZNXcjkQ4PjJvAzCOza3uys2TxLr9l9TU3LyMvQIfYMWe9L8G
GMtilEozoG6ITI+D9Y1NYLZruMFb9aSFsRoo4wjBhgtt3DjuFWjdAFSi7V4cZ7+JtaKyYLaRJMuB
qQpkp17eMpGpFoDFYmjnGROaAhuEMAwmtPXWexa8TO2YtbOl83C1JHTPp/tWAVSMzoaSphO3W4I0
IGfGaDd/r+FOBjUjU4XPR9+DTNEEMJy6MOSC372G+4J+X0clxHbpeGJFJiFtSOjwEHcjPa6IndGm
aSpNbWgRn2MKdbVyhbMctorTs+37ZL1r4MZ/dh7ojmKZ3RO8tPMpxqeqKQgeqSv0/zMDh3mGTkLm
YrYMKImrOIb3loqK4vuurGarbjY8tZu46lg/QaYpvyjJFdOhh+WT0hOiMp+0rhCRlcI66wW1uZ46
qFMyxyJRaVdr8kYkekcyvJmHrBVtFiiWc271osJFBL7B/xOUcbIniUX49cVL5mPtWj0/BO119+oL
tu1QeqkiIZPY+r6B5ZKI8aHDv3f0qSfl4QGeX53dbRHyQ+nV4zcOho4rlh7wcXCbuDdXQEL92j/Z
3kJd4qWNwWW8qkvMEyosm39E/4cWJ1JQsnV/1w92LvXL7gwy8ARyF/ThqwR8AoU4cSuZn6a6riFj
Dew+ciqatconfyRcR7xil3uU8b7omsb2T3VoCaLZmfQdaIYbiMVRmFL1yilUbIZqQnRVC/EurKm6
GbkFkGXnp3PdBVK2liFnJCrv4p0L97L+BHaFfNbQda0X1CZwkh+JL7UKVrch16SAsbAdhEcTX3S6
sBv29WE9+i4Pq59iwTd4MdDetfRWCNgc48YlpM2fHjp7ujyTabuRkG8pzA8l1xEhyEVxnDSICW6B
jj7HGZAZGKExMiNplTwpVppF6MIHgdgNBX5ijiGzOmd2wzPUD3fh76q1mQ5Xqpb5MlPWSPawK9l3
SCa+cjevdBfQE1WeBEZ5h537fD2MxfsYloDmv79VW99HspvTU7Y7GOXi/QisjfmLyIVI6c4JQciT
YaY/7sv3FZASkVIi4Dj+Bm/gVnp88ptQu86QoAz4/Govcg2DF5odNjFBAPRYoU47KzIUD9X4Cz9D
T981/CxbaQfgdgc0JHUXejUhbsvcajI5/VvPUogWf/SLDZVDswWgcOtLtP9ycrnYUDeeugB/Xn/U
gKJSKyykKIqk8sgbC3kOGwIj4oUZstASajeJ9gchk4m2/FOA5V50o5UKhDoVxA1n1eeyLwdFXSjB
6oKyR9rB5MUKyxfcLRRT1vgnT5Ntxr0LlqfxTKiYtt7rf0tXHVIWgQlXJND0nvaR967LYIJmVPY3
OR16oz03ktU8uKZdqFzfGE7t3FPDbWqlYscN3WY/Mkri7lHqmkCxxwUU9WbsMGgHkGn5BHXK9s4K
5dyy5csgxoRPIYnkH+I0KIi5fr687QXyY93UHSfgfQC9wP2ZrvgLM8kFvjupKGDTYH4/HUQQpcJo
ZO6isqtpzkLp8Qjlz0jLdD8VekTfJz5U16kRbcHKpEkrIffkA8Y5luQbIftfP2yK0tcQ+97otf58
zVYVMCNxs1K6Uyko4TWNTUTr7nuUhiOkP1fZsx5YAIy50LNc/CC5tbq17A5kLxwHul4os/UwUsrU
55w7a8L87zoqlk3/gwUNWfMmujbZNTjj7cAxLK3S1xVf+/3ipW159z3PqimcPLZEsaM9gc5xQXVc
1jjKO/AA0Z3v9O84I10l+EkidamqtgzwiKNbq9MFlumCxhq1IC5lHnRx3D4yTIyI/hTs6L/PG8zH
PbpS6RFfbFHyiDGdWaBEzQzs+QPvYCQKmFTND5+tjmEOHJdpc0+qX//4Bw64L8K16g9QqXbt7HBL
hrsOJ3PQatBMjOyliGb5KOn+2kuA+nLX1wSpwxOxtyF+uPG7e7GRRIr+vKu4d1Nk7iI8kqCWHI+Q
+NjvOg5eaC+Q7s3yciVhMst9nPVIWMbWgG4ldoxO2R7y/vb8XxBU5IzfKzfelDnOL98Qea/oWrK2
Efwk/HRYm4fCWdED7hpwdRDlDxV55bV6B8SzojAiX+25ULmnBdGJ0/BGdtAcQDOozgJ0p5YjsSOi
oXhQbjkDSpB2We6wiTv7pqYPa7565Ec6aLmhAzkiG7P95j02ReSzXYMJh6eyAGNQFAPRpCAsX0h5
UjvQdjTdzW1A/3b76WCzicpn6nj9N1A2vgkjZLLd2UWCt4H+jXmhnbfAiXE2LnOStMKMY6EPJevs
SEtPwnfcphd/ZH0WxIdvaw8D2NalkXOpqvjBRQDue6zT64YxRDCgqE6UdwmqxHQ5wkxvCFx+1nOH
aWGKMASCOOxtwG39b037w3IoLEIqhD573qaCxAyoBQNTOJzvLSAzg4KGyFA5iZBRpHvj7aVrqPtg
CvAqeKFQ2qDfbY4gB8LkvoQ3byWZX/e6SsqnPp4YTmCa3EfrUt8tH2aSWTTa2zglfCUlYTPUIbhm
INBg0BHqduFPBRM5LoGAtNvog5M2vBtE/Fnl4Jc1P0ntUB3xSIJL/plaTM7GNSrcTh4iW8eD85Uk
9Oc1poXlSQChYgDJ73Y56g/vr8kxrIP5ZXgxaSFD1tAPUg62bq2lpqif9y5M5s3q8aW2+ys0QGYC
Gei69jKcVoIqsB/kUMfhErjUbLtegw4UIAzwzgZtLkrWtu5i/09LiZ0rKjHk3nbP7h60uPZw9BHD
ADZRcI1k0ekcw8japqlXxbD4NTacKRAn+sbAjhHt9ouooygV3LGZm/dId8rnoxXWw7p5Mp17pAtd
IYG9Rth0MGT40rVtX61Pq/sGP360OW9IkN55EZz9OwPdmXcvPcR8JHuay5VTjNbGDzzp4lgq5glz
NAL2LghbCus5BDAGRwmiqPgqHF1eQEsLfcMuMh/TQit6OtBNHpIU9e5x6UtvnwiihQUz2UvTkDVT
k+YgPzXgQCBAsmUup9/5t/v2ID7C/TaVl8iavto9kfkk/BuuOWzuTl5Wts3B137N+XIX8AfeT+ub
Z/c/x1WX3CDz4CIxzOfYL0Jmp1/gf2O9oizm1FO4itSoXSvEO6Lm411+RYWvvc2CwvJDtyNaSutv
/ENg1vqM/Jw0awPcldDfh37Zz7KAljwkD/Qdg5uivxoqjG4e9Sdkc/RVInSY2GlUuCXop+udV36G
DbHik46OriZZc8HYiP6pJkr5dzXE8i2gDBAQSqt5oNZUcprE2g3AbUEmQC70g1gSFbQxNvQLdDiO
hA3bzMebEWJmIi5nLzeA/wKpngf6IgnkvvcfVoQNedTu+RTSuD5HNyKH5KJR4AwXxLlylgneFmuj
3pzO/JiuuX9i7Tn7h1nZAecN/2GeddJDrgRLj5twu11SRMzH9FpvdjBXgYQNQSNBoAdGaVCjXA/D
ZglFVDbrV155ajmGeweov88Edl4h5LUoh/VPHzg1yvyP3KYS/wravPweOb8taop7pSPvIRFaK/CW
k8gMPh3HXrga97Y31tQLcb8+AFynsA5Kmz0R55xxtfBXmYNUToUi7WD4pk3kJLr4oGXQrjrPeHBw
WbHfx9dZW/w06ASybgxpZ4qSK2f6t3rT4LK+BR4MO3sdfifklmklg+KjxRgqQz/YCa00xLvK3HNr
msB0wRmPjC3U6JIww9uq7ONQb8JakabqRF68H02sL55Ydn7aFGxX4jSudhaRIv/bYEC9Y98LK6rm
NKxL5vSGcm5QDFmUSGGbqbZbuPwlWdF/B0/ub/T+DcKnIECSC1Kva8PysiaRtLrGOP3lZUQ0rE2l
tzJEwhJqOzbesAC7Ru/XY9odD1xvwlosF4uw+x6p1geO4Zy1nxtHTpangKfa+mYeRMULDlR7NSPS
8TgP5euOnoyhkCjXL+ybKlSbB53bLoI9wEPBau0PbxN9ugbZC+nDOIl/pV4bBlRXwS9GJj7fcG++
TK97fmFEf4d/pP0VmMMgNJ4TA89dqp1y2SnMDa/lKxTHwAE9QUxsxIrne2fiWQxXL+Rk+gwCdgRv
+1zvXzTLwBpyGY5IVoRu5iDJSsDW0qJh57HOXu0hWPIZakzxz/XgLbby0em+fzxMhqDW4ShUOna8
o373/jsUrc/lJOvj6nVVkTc5nZjMq22iP6souENliOfaQ1eHb1LeqefwPhzRJ41FIvOtuR9HyJyu
F4NT9JLv31mwFtNF90XmuKFLmc1B421WrH0EYXmjTx1mNRBaPLoedYURZwToJTekyIB9eKLe751L
LVAgLZW/nm6a5QfjJ2ATXeSg1aI7v2K1aBjulrULxJ7TIYRrVAR8dcji7oQlWDrCToMLKZWawSb6
awm2GMA2ZxLnMIVNpDJPp/vjk8sp53/CJlbt8vfcS861fPBRI0CmIfrkzHxnsd6HwaKQJuETachQ
t5hNeYqbzSjQcRpLa7AaR0vSDQVtBtcTLDv7HMOr1vtxSkfDGAoBck4VBN/ZQsh4qte+duFpFYIT
BsmqOCfZpvMy0QNBWYEWcqwvEF8rWNtC3c2ziWhI1ysIKHvuW22HIU+GPjyqmxXnk5SDSkWa27ea
aY9fxcBOjngkqNGzlCrw+M6oDdIMSpgRl+B5pdePK+FijMqYQoGK7yAGvLvrdd9Tg9AG8HMPYGyV
yXhLEP8wjzHp2uaoOD87MVrqH9d09i6vCInhYDTh7eWuDOqbKBKC5CqP0jIHIi8HzhHdYWIYoW2u
y4FLeu+1rJ/MitFog2Nt/g7uynJvW7huNVm1hXHMTnqtQFq9pBOO+6FZp9ggM+S4bHJ7GJfXfMdG
XourStHpTm7R0MYyVXhy/i2pK6a37VL3SVCqqJQOvdNqVQoYp+epMu/ewu8lPgcbndlIPU/vejDF
JiiVt2vYq4e6KyAWjABgKg2rOrWEUu2CQkEWxmBvRAXEU/mkNv2+gPeEVCO41F00xfFC632kl91j
69lqO2pJOv7AjkSdKOWHvQHiG6DETDOylGB3H22dPsMfFgcjniKhiZWpbKLOKWoKTLQgTHJ/L3xT
qqg4hR0aeHaokaNnmz3IR4NhL4TKMp+eH118OHcJgK3z/AHYJx/CRFPbOH/SiXeESMGR9fG4XTIZ
RneroIYWZToDelUdN4GW+g7FMJ/3/oUdQdU9+9aCB95n59qoTTslQ+en74FQXjnWm1//R+An49Fd
P99MzsJ+nr3yZRKLdcmSi5rN+41qQNps9Tu8FBUeoA5dAOCZ0nq2gxlRcMB7mvKROmrw0Vi95XDY
HuLgOBFLlSAg0VJYpXnZGjPZPtykszC1WxRL3wvFkwnp/6oOFZEkNooAkpJwfcGpBvzhgBK/Wt5L
nPkAPydt71WeuH3ymm8oxex0+wkaOb+GBKCdfXMkHN1dYVdOX82yoQO/pdJbqtMw+/2/a1nifpn4
MVYg51Z0Gv7xD2RbrHPQpO5a1qQWRBSYIbkHYKYX2e6Ewp09IqxeF5uMzzZUSorI3H30mh/nqA8Z
FBtqSzdHHh7enRU+BMav8Wv8SeF9udgsHlXcmSVDwjQxzbg0qrCYtIGAacguc8EgHUTrXwIYARlB
un1aNRLBQb9PtSeTqa/10HjpUlO6jencevD0nBM/eYrpMGFuPzxDgvC6ZdvAPbaJs99F+QpZpPFu
LB8dsjPhauT3N7qazPgeMgApWyiGYBJ4NOBt1yJ7NOI0H5yssExl7iBJxoHU7hXLzpFxxYWbN8Lh
wMIBNchw5UpTEqdl854WORE7QSxK1FSmjx75Cu8obQwkjA9+5yecAqdFllg+4aUAdTghv1FbDIwO
4M0OHDHta2v05Mx2wbbJ8eMxbdSHH4gmJnceaFNFTa+pSDZuCD8keInNLx48Sehx6s/HEpHR9kko
Wd36UG/T8NRh5jBL+FU1hUz9eJnHO5kU68uOV5+pluif2ySiYlTsjXhyoKO2pZKlIR0wNxIhir4H
y9EJCOwP2uraSHh8OQYr83fAjWOLg6OfgKdl029fivqt2YNLfoics838rXnJ020310JsBnryR+8q
m4L4/n15DTnBMNacesxtPxpIIdWAaZUOH37UMlGdv4wtnrKBKfHhk5ctQZIn2egSiQfnGtvkWYlr
3VvCvESp9eHnOVzUGKLvWZdAWRVhAX3v5ARiJwF+An/0unKMNil17NV550ZQVbn1Ok2tICNbgDGV
M5Hp+sf1Mhvc92VsYE+YT7fDtno1UyITGnvlbX9hMhjY4rz7ydw+ovmmQKLA4U8jqQO2EsxEnEh/
Odii291wJwwbrsB680cDvq0Wiy+JqqP+ZR+TyJ8jf3zCGp+me5V8r9YI+ywttrPQXQXBL+J2O9MQ
o/lo6ADDRYwn31oQaMW6g9mkyIRO9/1AObuhUK2q++gar06vHkcueT7d/rgac3vfK1KC1mZVFAJa
0tNjUpo4Feke8rnArovXt9cyMt0yv2WBTiPg4zyk5RZyLslpOXaH8yy7+//B4SSIFLe/tcTo3SVi
TtbtM5O6hrGR1HF4PjS9YI/kGqr3NO1ii+Btgc1V6EcES3jHiEgadMzSY96Uf4tJzoT1P/LEN+5p
HyumU5WdQTDos89aN+2Tn/kcTMBxGg28Be2ivYLhP50dEV3nG9w+r6PqmPIVI5W584zO0XMMJOOf
aU/8t0w6BDznl+rSLJCRl+wj2B/czdGgMlGsxMd/US48vqUAH9CNjAfwmrB6Rg9VI25p0Q5PMcfF
x+zfXonL+u4dALB6fYyi82re0d9F/ZS7NOPEODUkl80UnRFbOo039PNMGQjnIwgDTR0IESjP01OG
yfwmC6Y8+okonADUTN+ILqpGTqTzymjLdsNuoTS4pKNjZyCGOUxwQxb+vuJu5ltIwUCTV10X+2bs
+Wqbi05SeZRlxBes+QJN16XLE0/mQp/obgw0EKeFtdgJB4ogrLg/EaGGKDalCMVKWlMEvqSbZarx
gOLLZHO4bzZc4+GuzoViF/hWpB6KKHS2IJIpNC3dPMOHkZf69CbBn+Pybwu0l4fZIKfcgkpJ+c16
uGgwqdhCoqk7PrwzaZcseFkH09hpsp92E56PQcpvDVv9fN6BZtBZJXgbrV59aOFxzSxO12NGJWfi
pMguLuogNIlRL1RNEhY6xUqiZm0x4o2RbbA+Y8/9YXYlLKuQBAxd1mxi8NjcAil66MKwOKNRE4z9
0+zhg+vWHL2WwoZ/GPeYBjqI28SbLAcZk/6voDX6A/Np7P+r3On1Vyd05JCARkEyI1sAIMrSkhC3
cwvw8W5ctGCNcPU1dqtrzi8YtqPHthi1T6+do1kGD5LF2oSD9JdL+Tsm7dCxyG4LG0HKdc5NBOwa
fZfNvbL8ct5R+4jKnqYEWrXKzLHSdNOs8XSvPJF8X65wUxypfTe1wLkpLwkH3icvINLlNlAUyrMD
LlcBrBep7WDrQ2U+5NJe7dD6ZnsDnFe7jVLNJzooVPR+l3X66jDCJJ73cTq5E2BE2yokGhdMmfrS
gc6MAARi8F1HlJDfYP1XQZL7yaog8EtBuvCtjatmYK5MKOQ4MKStB9dkfwhUDO723t6RCczV2oEl
AtAEdj6SLBzttmD7mBoKjIx4Rb1i7yFZWofFi1UKMhGvuhVBkGvh9PFLlT0gua2Ra2C7GAZ3ZnPr
iRdywvtAkAyOyGFoJ50eCGcDybIpnTN0n/lPDxg+Nn6XRZsGEahkvPUq2GOzZ26zeXLEaJvsw547
S9nwZJthXX/znCd+pdBD+i7CSVGY8LmCl3ze+gBPow3xGqdTe9uia7oVoBaVEmKdTrtOPGkn5IFf
wh80qn0t9QB+HiwSd7aMPzV7Y1ngOR+IF5FRwRxfRcqMqTWwGqh/VE8SKBWLFHCTlo0FhqYb7hjq
2Cf8864vnRcjc2a9sDWvB2VTZ8iaGw1TWCN29QPnx01dYddF9tnGi6KS2L46ryy2u8UkPrnd/vDD
NM0XrysDqIjRe/5iSkiMAilKblv4xg6y9cW3J57N6Ta6HUU8PrL7nUmfKFIjIE+fOOzDYCk04g9d
CG/R5T90nnsa+TW7w1MTCH8l1siCXzzjCNCK2N9T1KFcZFNhs5iGRS/JaKJGEv0+fSHJIyUUPACv
2gG2fmc1unkcmCmL2a6xBNn3TneH5BhnK5oOWFERVBdbStlwCxFoJZvrQfjFVnIGiCWsgSdvATS8
fWsJO7qTct6Nj9rDeHlGYj7ZcLaYexG9EHpSHxQAbtAtJ/X4Qd2B0rYPi08w4X4c2MVCoSwn1j1d
5Om82lhLMgHK8i+CTs6Dw75X1Io1b/o8vYYfRLrv8nuWkXRDOndFZK/wtI4kPEhLYKBUE5NyiUBh
OiXuYhqV+klGoOwPNWVGYJotbOvsHZ7bLYfILTb2+YTnbrkNFwkdtjFMOnKKTiW+Ogp/L5zh3n14
QPFah3RzR/8p+a0xJBN+Rq+wfYNwwtmhjoAxBBj5yFiMHeVMfpMHt1myj35h8T17x494qjGUQgU0
pZELc1m3fx5igDeIE7KUVFNC3GxgaV6rsSvQ4ErtRKd57EkY+/2zIe6wR7A2LgNL/eUY2RqgiEc4
32s1D52wcWeASSi7LRFpjjo9xrXTBvIac2zGMXgkf68l9gt0MF01+o8Dw4B/hI8UoNyrdidBVS6E
xpWhj2UqIL7aQxbxrVbeZV6vAe2EyGHa6NYjSGgDHTJ2BxXCTlSCFDf8e8eCiE9/3uJ7gKfTrm1n
yLeFQWbJuga/4GwKypEQ2YECpDVIVBj8Sibzdr+faoOkoJlTxAZbSCTZcBOxxNeic2xUQJ+Tifrd
PwxoJmXINiKCyKAYScqAozJFczw/IeQ5hkEs5zQkw4sYQIBTKAxyoWPjDUjJ2Qaku4u5uCI2M0MF
w9eCAXNSoyO8anhf5nDPB4qxtBfSeJlkJvhwlUWcFmLp5ZKf8ARTcqOI/1Y8zDqEbT46dQkJ9fq/
64ittmGJoNzqtF2VAMa0rIjSQmBtgCQjQtfnZp18m0729ZLeulhbV0ZkUam55RUnRsm2NEccsVP/
JMyMGvkZAGDfd8FlUSHchMRPlVHizNFUdKjV0+7joUKfP8RlOP6wF5sJVkNi/T2NIMKX0h+ulMP2
HhtxMPiFev5d9Lbq1lRkZsjhfbFvFjGfCupDZvAJeMhgpQdFl3Tu94GGf8O1aIDm+dZ2jYK/1m0A
uRAZYsJAgi5+LVlRgDuppyfpLFrxX7yge9IXevrgWSpIXVUdriXKb3of1ibHL10Mj5nEoRIPNUb5
K0O7aw8y4iRNOBeKAouoQ8vJQ93t6P+e7Xpz08kmJodt63pYJsLdsz0aFd64C+fWmGleEzBdUTjZ
Sy4x08dV6O7FoxrHbS3L7MFjfTJcFmInNytT5z5dvMrQVQgxgXY580nAYFy2WIa694854q9esgNh
k0DhBkV6zrlpS0RC+5qsHj3BsHj2O0iONdBlrjpjAhBVw/fkAAB80rWkacAhUP37rcuaEYtWoNkD
2zGTGcKOYLq+u/pF2H04T1KliAPZXg2qwdxHHLl6TMxCi6Cysr8PbWZ/w69OA864NNzFzGgSughg
ugQhjQlUVYWBEbER3wsx6el1iTvXSS3Cn1rJmmIUlFSylgnVY6uur0FvgcFerQKmQLdkuuldEM/Q
aURn7uIXnzCHtEiOI8L2VE2NKmF9c29fHpNX16VH4Qp+zFIYRwhw2tTxzcyUd6VsK2AgqnnhvWf0
0mpOjyONrXJsL5SzPWC6mn1c3ut4Zy+93B8L4CMh1LimJoYqBwxd5E4eCiNODXx1NCTsfGHYmJCb
RiUVrZW/3q9CD1JYK+sobE0mw7Y2VRj3wQv3soVEPkhts5CL02TKc0d0HyOZ3waevDclQnEzFO2t
KFYq0pTlctBk2APSoe9W9eJT6OZ/1+glxwOScWdP/uqlw1f65Ju8OOpBI8IO+O4PtI/W5wOJ+aTp
paGtKw2u2e8da6JXH+e6oyRvVb5wQpE+oAtuYLktrbq3x/0RhFrdEmqa0cEULPdrhbRN/JCAsLWV
S1WEpNK1edvrodI3sPactkEV1/ENxleE4EmIfaZXbD+g1lY3Skv+KCtLROdFMMnJuHebU7KexMVI
MWVyaFJz2qvb+aDyQciL9Vb6irwPQkoYahYJucsA71l4NSNDIOYSNLFUfTdtU5qzS1UZaYThg9md
IvgFDkQn1vtyXKnEpg1KSM6q9yqNXZCjjf/aLKrOxYgB9vsDeb09CXeahKqSrWHUN6z2uSpGlyUC
EYdTD4zTGbpWa6gfy0k9tugfcuFCKal7MpXZ1pmKxG8CrCeTIRT7/JKhTl9IxaMTAkFEBmWrAOHc
rTxPUdKJujOYxmnr6pCxAFTQButw6xOE15J21utBNVogvkp59riWYF/iM/fezJhOS68o/JazKelD
qF0SffwjWHBS9SvKnCMt85CHOyYL1UxYIwg/uhV/IHpiv2kikRm0k+tRvwdyGvnIHtlWxPWFTTIa
CZhR+pvmDZfQRN7j3yrQVMC30BqKAZws4TXGwYceXdi7uuGTi7dhEVIzbBCKsN/EXtttylif5FwH
lXvMfinuQuE1dlYVl89S5grrgpWcNbfLYC+7sP70LXoUEURjWrZzM15B0c9omK20U+ttKQ02oG3j
IFvYbLx6Okwt5Za8zzkyra39INHXNFEVudizsogPzxfLT9OwJ4NA2AWreg4TC4yz3A5KkFq7mn2n
YzoN/AtjRaR1gDZmLSY/ZgFPmdNFv4CG5HFaQPUYDO8ov9gbO3fqb6wEaedYwQMarvEdp+wJ9hp6
q7csqwRqzaYG0Kk/n11VjbDGRUX0sTahS8frQVLb/xG36otuGPkHwGUZPBslNv4OHTAC3OQ7YvI8
pWi4MKfDB7elRMbVlh7SIA9QFetliEYiKfVSmGj6Htmt0g2Jtd+hiYkQd6uO1wei0kDChsbaJUvb
CEVH+RgS96BA50A2cTU8J28Q/M7orPe1rdlGEngQ2PB78faPz4VeLhAgcj/lI2kX6jcXyixQQqM4
wlP4qXnliuqn8Oj0zCwkLJqCuZqrYWlVHfojJOyN+UajnQ+kgwAk3dGliKoLJOt9nfRXtPbHeBuT
sfhV9q9OV7P0R4vAMjqx/oOi065N6F7+1x56K71PXbP3+fNZzgMV4kF/AJGTOowe3p2n40s3YFSu
AhA0Y5NB7KuQ4UheYkRJdGxOGav6Gz+VwC5yT0pAZUEnkjp1XvHVhKTv2tLTfuClFfLpr0lufHbg
8uqznF2YMuPClwEXAjDLQlqwoCeOwutL8SmdembiiqpkysOt5zLPYkjl3zmAzcLt7nNwIwxWAyHD
vElKiRNGFF+vu1tIwrwDDXcGI73eTAyl3PunmpBHudMZndY+NcoLTSRyGacf/uu3Yb7dIL6HAfbq
ZJY2UM3rDM71hswfmrGtJeM6mF3Gyl12AnoC20Ki8snv9bp7KMFdIuVHae/NcbRwb6J2U9f5HYYA
RnzA8ZLHONRBnusZaBGuf4tjvpQyESYheurdoKuCDHLa+7bABSds61lT4RjEKywYZGIBzzO2XtDf
pXoYOkGsNMtNtCOjbsc2yuUfrXPRhaN5YoEhg/kWqmj3T1pptGbRaxl9ZVn99p5Mb1w6USL+HG3T
PB2ll3hj2Y7aKLjGXtRmnYXetIdDOrbRSPmWFfDt6LlyoTfW1f9nRbftl5Ez5GFi93VmGSwcmsUo
85RgQQ/4TuPr5dSmg/OBaEYM68a5rVBIGBXJ9nCe1Kzx5FIcbH90ckboic+a8SZqBIq/yFiUYYGw
bY338Swx1bx6fHJdLeAp55+M8X580P6zOQYowhPs/KV9XZKmXi5kg13BobQrUEVsidyVWWfxyPes
AJ8ANDAlENynELtqwtaIRb+/HFVzZJFd7KDqrpIb589Ie0C4WMZjGid35yiE2ApXe9+HjlCfZu/S
/LM4/rhqcjtKMjeKGyEtPnEWM/Qme1EKnwODmVNPPkeFoZcApNhgDMABu+Ly8Wy0YMXxl9VNDAtN
SpUCAsc24nLXghbVW240imG6ozbwy86QMm2xSnMae60T+0FVAVN+VmwmPjRR0Gs2okaGgR6Jy46z
iJR7sSRO4AoBaNSyjKUH7RzzV70PB3+280Ql00/mKYogVVy5DtUeoZ0fIK51esgUyiBUhF1P/NV8
UnUl6FYmbSAjDGdVTrY5Rbisb/3SXEWo2XxDb1Smxg89GcdcSSN+gY0Nchq14tBFFWK7RpHOV4e6
/QHKYlbnPIbuZQtBkzqfIRDRN+fEjWpQdBHZvS1lCeEWtTnsabIuGTp7kk0yTU1pT0mmmjS4G/Za
F7hesO4Nx6FNO/W9C2o0eak81fanLXOBLVHHbcdrFaHetzZFwD0dhIzHaa5vsDyZjmo7CH2LGMMt
cpl6MNgGgTr41DEB1plaZjEUS7j6TA/mCuIv5397XgSTF4yqPjoYZw97z2EVk/td16AR22hrzyxe
Dw1pNZZIPSJweiCdQGS++H8afJQ9feqf4/4O5W500BGPpTTzcsdn5VMKl14xLArWSSIbi8lbpPpm
OINTtNu0xj61YDvO2P4vIe/dcNNAJpwgSwWz97jD46RE9olDL9ZJcYS5wW95M0UB3/vTUwOMD3G+
xc5e3OCBqTAReBVmpew2xAz076lybFdM0fBhCj05p9iSV2hG2eYYtocEHLHSIJ/7ussGTzgs7d1F
bki1C9rQzzeMpbtlB42ys+4FKjkTqRrqcJBEwg0NsfO/tk01LbQ0kXaoSM3Cg7M5CGuyNmXKtRx+
HXPFuNMfkGFne74u6a+78XEAjTir/E+3Jo659f0nIy5l4gk7q2An7cvFKKK2JdotY3/HJ2IyRP1o
Zl4GI4SwN9c3jEEE98qI0H4/PILqqd/owoJiFIBFHiAoItQjJppeEoAl4tpVqTdPM1yn3dKDzkGC
uTaoU9lR7QhtlGaN4IWDpDaNiJ3t5/adx52S5SkO5v+6C7F4EwHesf/MIv4i7TF58P0UpSEl2bL4
xGTwhUhQ4ob62/xgg/MWpsUtWoAfXa67TGzuCutmST1bdulCoKp0q+p6cqEjC1m1VDrnJlEbL0dC
/rF6x4GWEbTbBuQ5mzcSqm5WD+2UH/FX8ftFJ73Js1wPNKmiWTIYpodjKXcsgsiAhlG0L9lXlN6y
Gc+pF32rUi6O67kBzaULCzKoZMyvAABKb4g+G9qQWWwEFDZLOEeihT8mW5ok2wofSjiJxO1LpmRl
EcTrKh5wwrdsv1eMNVMNL+qlyc95jdArIuaozGiTb/FMpHVdxwqIpjnrxK5g5tFvvQg0GoVNscZu
nWcK6CsJQ4Q+j38ivUNNe0GEYQZ4he0EWZS+tWZVKc7hxio5SsyHg2KxfLymbQU5FLFuiUvS514k
QtAunlqLSPbRQM67G9lA5JGh2jLTc3sdKMGod/FWCfSon+Tf8zcduQrluqX/VlwyTD5sjMTXta03
8+0D8E6vVZZSaQoiw/z3YpXxqbNvgjeE4QVzH8oxzUi8a1UwnDEdnebckFjgAby3EM2HPcOUTdqb
ehQLR/ypdCCZL2nCZgfQN7zySFW/4vPPle9TRKHfveFcA9Fzlt6QjQyLZbRzWLcoV7PxXYaw6LvN
9qO4ZoBNL59LPr/ESGjPockKoizQr7rmAJB0xQT46or8D/9mE9vqOdP6dt9QjbVVDB5Izv0dcWAY
8+ONXuWNKcdQ904YFKK0Zb2sqsCD4d4H+e4sMgp2U69mDNgX2K7gjSC0jv01ft4ApWowHG9NHoNM
gB41+KdfXaqv/nu+ksvs7nwzKeaKz4a426qixaS/tdbR/422keanXEi9TGyeZJW/gRZdff9gs6/8
6JbklH/XvljFL5KKcZToyXqn9925X8Pv1K9znGw/C9yjcwuy8bSiH+y1ImvoXA1Q4jfzjUjTTLGg
7EWWoQV45y/fUfvCk028E6nx+HgkIar8/fZE52BVOtI2QKWxtU3Z+dfWU1p1bFXCgLDdd5hHyOd3
xOp8W/1aouOnxl+P9HthMstC8zTHrx6NDQ3bX5EUhNi51HACKT0w8MZY3pEFJ+Af3K8oT6wwaZLB
I0KoLGbFIhqgOGadmVXEDP2t0IadY2l0SZy8Itfd750JXqv9eSJsASILFL38f0bKIDmN/9P/HrgI
d0XaOLcHbDKJ7hxcowaJtU2Oz9MIf4+FsBUc54CjNQNCWpM92ed27DI2375hOwPgcWKIORN1Usq6
SKdv2zwOAOp3FxWIYf2gtrKD/+Xourq49JSFokuIezm2IigZaSRk1AAZdmXkLS6Qd2XbUeuUwOXN
fUTnvohbdJJVkwL3c6AAmALaNJhM3XMTIMT4nc+jAVWVXHG2PBp/+iiQ3hcHUmE90o8QNTFvwZbz
olq7x9v1PcbGZ0EneHRrWSQRn37Q7du2wiDM37VI0YmC+vciv5pwEmJFJeLHcgcGW2pDW9ZF47vJ
P/mSVqeG87xdB4gawZMBpvsvU3COROc5sPA2JOwflVubgQLMdPrNfQJdjkUStMInqQPgXazd0xD6
g+q5rx4X6pq5+SjG5ovT0vT7FLD4084BCfra+TQyHbaSg/jTM4NuJPhrnv30ALvmXDyj/EzeuPcs
DTVUEntv/xuNjDupVPDluETUkinI2JtNmUn2WNpmaJED4BgHUDxIqpIqm7lgpH/DsWrgDfuLORCO
f+1P03MxnYhUyXel6BvqPs2a4ZUdPGdFNfpUzWtUNl/FjnOtEQ9Y1uDkOoC7FGEQMUbjxMzdbaK4
4oqJdWBlj6N8sFqJLcV94zJUyFwxAnZNagt8aiw13d9pDSRVylXcFeXsdis5jAHAJXkbMswxAPTw
rmKjRViI5MDrddrh5nLqj6rSICwvU0vv+6fC2FhZPzie/0ho/8s4wvZ8A5S7/r89w3wt5SDkgmxo
7xn6HuGl7hnI8FfCS+BWrMAST/F3mFl9BGAKP4HBb8e6m49c5IGAN5f6dal/MR8w3ME8Za5lsIvQ
ikF6AEpihUAwC4AM547pDB25VpvT+SREwiuADaQcmJtElmV5BFUVhGoO3uvhWN09YeDacHjlkt0z
OG4E5FqpsoT13WVAjj7In89XEowvXplHmVqOXokjX2M7+0htJXFgdoX7eZo6BAkQwa8BOz9Z48fZ
2IgNkcvACVM28ZBiuC8Ymtz1cSiAmkS/QGMIprQgeF1nVHkoFt2AzIbNODTD1L9yUYy0RJhwqkgg
IrBGdWlLWXf8JZW7ICFpeHVMXP1KgpMr1LkbFA4v85lgE6s+/HsmRCAdC3n2GlM65LL6CeECMaBq
XpuFVxL7ZoXVW0hlRPp+aDtGOYZ1RrCx96S6lOp6c9eOwtr25Y9bSJ6911fppUJft3EmuK2Cqq7n
TGqd0kdqqKV1Dvwt0XTD49wrTm1jar2c5AmUnk9lbSQDgjzPF03jkxQfCu0HlGUdAmbC1Fw0LOJG
ENsl+lsWsvc6AGg29HXs4Virc79sPpO90NLG4Ru66YEwUORe8Kwh6X9JxbUiL8rlsK4i65xkxE8o
L3V9eJhEmH6xrZDbFeG2W+kTSHw9v8cqpPLQgQkdfz4JsPcf8N0lc3mDeqdX8tYXytw1S46heMTF
L1XuRpAIkMk7lxuqgExmZtyBc3pGeCFq8/qlLsy96OjywnTCv4VqV4VioNkFhaKPabMGG47Q98uy
jdoUG5yXzaKtzchuEV8uJ4E9PNeV5TPy/GBG2DVmh1tPkQH1P0Hpt9OwdAANxZM6bveVexE9AT0w
hhxx1dmmgT7ecFLijtH2qRcHbfvRxpHuDPngDg4w2UGBuWg9KWyvFZmZcn2l2pDX7ebZPJJfPVlg
svmhlbHxqNnx0tKMYCiTwoXPnHj0KkncSgX9uiYXpeUr0XrwH+j9ENErukp9iQ2qxfuyx/EGY/Cy
eWoWF98VWDmOzflwF+m7iVCL/7OzPkMVvQWITHN6nDmFqel4nLzkUNCnat+iPVz4pzsaWQBxMv7O
5nJLIPUPUPk3bBJM874VL1b9WSiaienpnBZcA+CgyEbpri5N2RiQtF2ItSATc2U4jMjpTztRF9YO
ORJ21aKegjYMKQX06MSNSSnLTy56BmAxuvav2eSXfXCyssq1sxgoBVVb44WYsvDhFfbc8+B8Fr4k
dJY7PPstDT94+jtZr/m5SlvfQ62s4rUsD1G663NresOML6MIHWseNzZPexlAxtDAFKck3iJS1HOV
62fHO1F1VT2M73OYbT3e9TVz0abbx2hiOR2t4oJ5mm0t9mjjNOyTQDoPK7DexGxHv+eR4WWysMCP
ZuHzKMXK/cHvXRtPJBJWg5w5HcbTemgXmrlF5a6AV7+YKUdaphqhvMt3bsgIZns1HYmsbnctwkvF
mN/Z24u3zkHUX5/QP+TbPcOBYJUJQcv1mjYfVDLbAf+FIWqsrW87Tor9LnXsdHZhHLO9V87j2t/D
wjK3rYcrzRdb7wEVEjKURcfzqVjwh+ZcEhlqVnwc2HbfjvTKeXJmcd980xpXyqWOn8aXilBPBh0x
x8I4/ASL3SKjfunuT+vSgW9ruNAVGaztvDlCD7bJp3J6BqXUiknBREdDG8nB302QsnN5JpuoqjMl
XAU55yoq50TqvSClgKYa54Tn8QiFbrOjUvzIgtAWqK3kxeHscyQf67LQPlYI5VcqaH4MQuHpRSXZ
O768RXc/jDCYULoU5y+v/SiP/GlKd8/k5I97mOiPwDbAComY5+xjZocv1XO6qHj5HA9M96SjRFt6
5cu+ZD53XxJ89UQ0RewtE82CBvv7DA1Uos1adyilrmqs28UnjVyFS26q5bv+UuLzrE87oCUF/G/J
Yi+FnG/XAu2YQbkMwkWO5DT7YJlLeqPk2YCgL90S2AZJbvi9WAUFDotnmZDtwttSCxO1VjoewrrA
TlvBmz4x02E1yW8IZp2ES5MnUDwnj8co/a5h2h93fqrnIN5krbBGjzBv4hNu8xegRwki4CAmFI0G
Q7Oz0HCyqzmMthQVSu8Ho1xFCE8gLIM0I29YKw3w4gn8lF0lee5tYFzLX0NgGM/fVuKPpcRLFviz
9Qqco56c7N+1wCKlsAoTawxAywLu30YdgUjT5mbZHBNG/QaPcsAJGfdcJQpz8h0JhA2SbGSBFafN
Tkd30B7QOk4NMcsp9kLrsidYraWtcG3Twdvw8cyabkDLq+mi4/+jFzk7lH/+98pB1DbCjs7ooWBD
Q/BNJgGIdqLvqdmkzyZIj5Qqal+NKJxH/55Kkepc53L8Ybqin4bHkoo/Y5BCUdJk7ACiyt8Ut/Lr
oLtVX8Vg+ttySetMo/AnO7T9B0TNhg+Va5N2eDrrXFKV+hNCs7Hags/U4+XrPx5N4125v156+dyY
4PuYf1XIINAAoO0oZUoJ9usY2pLqcG2T+9Cbc6dAtGNVY9RYVrN0BF9VR7erQYnD57QMPXuNiFOR
2uH05MaeHMyBrJrhFiwtSw1s0Wmr169JeeCyC6TdHHlwB6FvjKizHZaI4TM+pfpKh1XPThMYKYgs
4FhdUiLy6N70YBjJX4EgbP7O+gho+PL7wiuKWOO6adBiNjdlhP4OKALW+J1Cb2DNvVqx2bs8sPvG
BpQw0b5fh6CmVySWnQAqnmc3bYNp8Ilds6RUO3Nt8v0VxK/FkY/Xx8d7S45G76ZL61uv+O5nMIOP
9RM4covuq+G/K9bjDpgjeKS5tQwpGgvKA1XTcCD77/4ZDLgf13THuGMu7zszy9ADFhdDCuRB67ey
FyMJ1LfI6vQxrgLruKRnfScYA9ydvIYq6ogAeotnPl6GoOLIWLceaM62S4I+jkTbv30C//iHe4EO
1FGy9y5GIE/IEb205egCXGLDV3+eOLfrvoRjBoujztXLGA3taEo7/dt78t3I9FIli39vT0Sw/w1B
wKpufRm6T74vp0ZQceFhqQamnydy1piAtfHD/BK59NzYEsb2wQEtgxbotE4VkD8Oc6qJLIRW6jxd
aguNiIZjRjjlgQDdB0clKVAldkdrC9Y2pm2HHj0GY5HDcNR9T4LPdlW03/T8lRH6h13fXUNNkh/k
t24bH7b1kaRALLyD5OW69aLIbCNMdhLG7HRdaQrk6rkFUEd1xpKTCzMnpFJD0jYGVNQ5IHvHKQNZ
vgNURW2sZS3Mru4NoSufE7OUi7AasoLNXPr++qKZ0/imWPRzoO05y8GTO7KYn134RMA7jfB8EY7t
rY5ZFqFvda0xNqVQF9FnXObd11+o7G8NhSj0KJe/JvzcPBQMW7QQPI1PUsW/TCicQnwLYV60qLQZ
12n703bevCCPV1smmvD1Sq+HGnenD57kBIxn8j1pUPtyg1Xn7zEAlQFYKjLQgH58fKFhb5i28i2m
hhSIu1G1fUKMZcBWcR0OjMnrKZy5aXaYOzOAnxWBp36pPXQvBTN4T6oYNvnErUlstKjJDHKuOX+Z
9mhBB74R9HDzr+k+XFLA59HpRB2YALH3Bi6KWS80ptQF7ZJMNe0PrLZ7sLTcHHcM/NhVyEEobMhO
gPkFocgg/82EjUeKPK3YFht/F0S4m8CxXR++1vZ0onINuPrLUa4C4hslUzBGoAWMhEGPwjUPivrC
0Hab29LVxdtV660BG2eRWWKm4vw+dBJ0jaydOzRnu6xjkyaDBoLrLdEdRmaOIHhiyebLoXRuQnKi
t+yFXZuZBCt+0alubCD2X+rRbFWzUssTyOzynEHoJMPj4ZoCGjCPtHvVHvYpiDgNJpaQRHueAxdt
naiestSIkHXmteDb7oiNiHFnH9m5mG0U48xrUyLFfpI2ZeunlJZqNvb6gLOJm8tqp7DgGk27TLAq
qoaEDxokruC2HyM6x2Av8fXXY4W668AAESt2LdjV1FAkfB/wqpuIZs4nTGnbnWwnhTWwp43CR8zL
vEDQBUku4DAadvaleeQsoXJ9p/CcLP+u5fVDw9HxS5A05uuXyh4pyrYHBkOcit3YgF7W/ETcYJCW
3869zxPqc83mVOeoH/zXzRVvmJL5hIs9aFLqyjhhSlnL0dDrOtChJEtwr6/v6589/ZuJypn8muCg
okLdYZu9sXJCU0V58D2SXz+0soDMbywIqPqNUlE0k0ULJfnBb/Y7bil1wjcS4FWBo+HONY436XtK
3oT7SYDno24kvvDMVYP/vG6Ciofn1FuPAsOFg418o3tMig4yTigAQsrOQypQ/DsBMgsLkB1YnBdd
815Oz9Sdy1mrPAhQeLaPZo1Li8P5g1qbD4JvhPV5F2Uo3ZPlThCzDtBedt09vvmWNxvU00Dv3otE
fQf12dzI73g6AzB/odHvjlft1ffmPyzp0/yRaqEFpjZVNbdN/Q1hitvRHBpy7UYOr/WFO4hDApiu
7uVqnpOGB0nN6N6u/aCZCrRhOTl8fpso06ETjNe4Pf34IGBj8OZ/YlgSdDRP1GT0fh1flyv10UAZ
bUar7etQvPjv+9ggArE6CJlrDFjIlIWHbYS6F+DDQpBoZLBrfAAPMyu6l3TSR4yNhjoxWOmX1bfa
nwCttTl3Q+HMOUk80kqcJ3/izOUUFcj8vlFABzhD4e+Cwwj6pvmAdVnuuDDnyTHHdpgpvIS/P2qS
WhDLz6ftswj6zZcJCLbfi1HmCHbAsilr0H3v9oRXOSz2zhTaaN0V+lFMLU1qsEI8UAel9nPxGaSO
bfaJgKydoZ5JRjQYignZ5kI93bCo5vVLN6Co7LKstmPd0MnwQ6PMYxWPJvc8+nms75uTHy7GTIwy
mtYm7a+MabCY7OK2qqn1kA4n9+a/dnlbPYspf5+ntAMCjGUUmz8pWhjrUVGuYnhA8gJ6Q+93YVxS
W0yODBjLYt0H9evtb9Iu7XRvzP8/5JJCHhSeYxACAwmvmK7heKwocLV1GeYsZPkoXkcnqTp9z8Ov
7+5hLf5GJPQadh1z5orwxpCOw4W/DAxsmHV8b6GA0yLObTH8ms2XfCO/c+slR8Tn7pvmGobfMli5
eRrBt5N7maQsF0VRc4D+Hf3+rW9ppJNo0t3r8ciocxLe8HFlgMb8MvEZfYuoJuCRnIIequx27gKB
kyspT/YBjFXRtrxv8MFmDLXgYQkSLS4QbKK8qZ4+/l7uoPySPKCNGPdyOUaT6VRmaM3sWq6KJybH
3X4wn4SSOrQ/t2aOo0TVeaOodin7+ldIGe9PVy/3IjAgB6JpKiGM/10h2SMEvsWhinROzGFBunW6
st2L79VtTJ6qd+MOkchINAZNVLCAM59/PE9e+7u/ZdD0ezC03UPY4D3maZ6wolPuv29RCpbn6Npp
vhgnbinVeoHsVbexZrbc7RIivI9CK8eS/t5TRtPD+QFoiyKHmYtOXjmAW6l5sz/Y7lu53Du7mulX
62zqUAB+aufrFexMfvBiOIr7K6icBIedgvjZehgX8FMXeSSG2SMBKkC6VMBxUzVZvyTBqj5myNFX
rSbah62gEOEWImp8x7pkwkzPiVm7CqLexA9kdB3mndS8wfPvBP1m76RwiKqs7Q0CmWP8tBS5nCaO
ckMV4H2UApDTs7b8+iWlhL+V3Ddx9g1aQquv4r+0GAaFrkLAybe3mAMMyVgm4MpyN+m8/OcoGo70
JNt9urb5ZtiG4tksV3BEgMiykPm6BseIGZC2cVoKwBieINXcvPH1+QhM7JEQp9PGqzRgbPzWEyvh
Jy6nxxamR3dSihYjletU9KcHBZFxbsQWDg0qx0vkk1zj4iQDpkOEAJpzoO4P2RQzjiB+JWAIpeWy
FuLot1CLMIKSc33V1+VkqPq/pzDrdlS1sURzTN83ZIDuoni/VYSGZNCZ+yQ0XN69CKJIKfwvBye9
7dA12JSbSM1tSLBcnHg5q0NMxT5IFnIPofembBhKXa+Z+m8lZ3rqzkTktd8SMZDPKVb592FBvOdc
HvLNoKLzpx1L2Nc1H9hIE/oN1ecozFziGjrr5COKa/oLZJPS9PHPK5+3hgknVqoi9BDpvyI1rMq0
v6DudhTb0cauFPyZWP5x1gScyA5vwXSPDB3xNNQCsfs6YACoKw2dSzEMLoGtMeorDztwgkNtTblo
YWD1CVvmnXMSg8s4nND5an1V7ScXe/fVFLeQHebE77ThpvtLfJ6lgchmT3PIJJUaHFGoSNOPC9fn
dwdEA3xUmtGfJmuFGE5VbHh+QykoFOMpvY4zOTxCPSbUISEYoRp+R3n4tcxkwA0GvWtiVww0pJvy
togxJmDl/afaHmAlPzScJUb2coicUOadLj2KxbyxU0T3uAcbyx6jOUIMiuI++TFb0/8hDZ1IT7Kz
LX848CeW0tQ7m0bWMtPONilyvg93JcXHX6hNLHpXduZyaeTAZ4MDb4K4h2yey60jHPBYtbtYm99c
emd0uI6WnpWBj6rsiqG9brv3t9+Yz6fbFlvPieutgAIjwJiA7WwiSX/1n3T6+sNiBrEjfcjGBzdF
8kWNaKdV1B9tFAhdDiuzH4u7YBCZftOy71Cvkb+B08hPQvq11oCM2SMehvv7Ny/vdCcq/PoDJ/Sb
9enrjhL4s+uJLy++Pz2NcJI/60WB0nOru2chjmtspEvoNt3k8wBwotRhA5tPqLt+UqEfWa5eRO4e
FGFdn4IRsn08agunN3I0oAkorvQQYRJS0fjfVU0Xm5OP/J4gfPwpqMPk6JRNgVj6wDv4elmoiHB3
GFfYJ3P8jaWeHpJPfl96PrUY2pmnUMqa7WSauQVGCAEApxG4psmdJVwF6wSj094pjylaUK9d/YML
JwPQ75EA6esvXODOuU6Mv+81Og6jaH+Jey4voCurTomSO/fN3VoY3WrQvfcrlx+Odlg3xvrPR08W
hsP5e2FdAc+8UiCsav6aaDTgmuHMMQB3+3fQmgu/LSA42RtV20rHeBvHXB4bZeLe3WYn3HJl3gOd
QPp96s0qJyrY+1pMGMXsjVEUbNXGODMZB0EGbeu6XnBgx2f/4cUPgBlNtIZO3SxS1QcTejfJEUlS
YWe9bmTorD91OOOTvZ6q6rZIqF27sOO5XY6xuiiwSeb4Dy/JpjJrszEESU0BJar13NUByb9qXCx3
yOgQzIrhEQcDslASUZ6jYlayhVlNVfhRzT2Uomd5ZVegVJroH42qrQO6t2b07JvrFJm7zKYBhGkY
x25qg7AfthcS0xCB0dSq3/JF+3dK0yigZPMbCoEUgdPvrXU89tQqlwRShJoPY+t7Xeh+mTPvehN9
FX2Q0+xUwg3fF5bDe4t/tT3vzRgT8B+Sv84ATFLL9844w0P6UNHxFs4dznVwoSSyM3z92fUJZNi5
grUIbJ59UQH9EeF1YT0LAqZA1OWv86vXvnLoj8erJcTLhbGZnXvKKMR9+jFR3NdXMEHO3gQtsjv/
biHd0eO28b6iPaspUS3JOJfzLHcFlJUmn/ODcz4LGk6iCGpbFqm/qGpEF7A0HUG2y/+S9VuVbyUL
UIzSoYkso6OGErxc2zWoZdbueZJcCGA8Ku3z+UF17wk3kyaE8TxbjqS5CR+OE+D00dQo4fp7cJIk
1AMQuJtB8FUx3Ehr3/HxbL87/XfHdmmqYCbXg86Vk+OI+S0VQsJikyEK6cjRe4/meFjhFZzlTR9B
aH63mXpLo/B4i7zFct1bY4Cywqg5ZBC0JzNAMesKyLownqRaRi5S4OXBji6Hp93sKOWtdE0f+lTd
vYZJSSLfDfLJ6yAWXdT/ijAV34hc+eyPxcjVLuZ91FvGwh/L8+ESOUj6nLew4AC5wtb5cidERrWa
p/fKd6rzHJzLvVDiBDoHAkmySbr0HI2q1IxECZqxw4DTHvxw4ihYFX0ObBndpc3aIXCIQlqnUFPT
rYgABliTkeMtG2aLGmKuHRaOdB6QmzVnoEzbLdl7OYhQGtYUDjIxrxGGZsSySc4bFXJNVWUGqic+
fNVrLTG6R1sLfomXAChbYHuNwoNON23zecs7gszhs/TojmNDmGutldY3wIBDcoYOGMUeutZ6qT9H
F8seprsx1XU2CWGN2UmQyFrjgv2RDTlBUuK6VcSYAlpt7FDLCTGdoW5rLb5ehFrqqWGqiPNhzUK1
Pr1oyhmhWRdxdsWIMFrATbdnhpKbDTjjyCz9puWCR/5r54/axnmTmSuc94Y/Gbt497AheQQQnZa9
B6iVM+QCVxr15cpR20BFF3SQg33xELoQI/E5R4P6bYPvu5GlMjkOngcKLSRkJu33xBCtMR+28dPy
Wu9XnqgU1VjKS0tRXkyCq/LZ6sqqCGyqqW46qurCNLu9eSLF8J+2Vx/IQ0viUHN304FQQcqIzr+x
YsfCDm07J3eVVZHUrzsWVgZihdCU9o8ANZohR+xBDi57ovxMrQzhFegbdpTi8iHQwEbJJt4fMmOt
nLS44d8JsmsDqJrFwXmgky23yff2KKX8CBKnzPNDoxne5BoeWlkkpHWsMcaOn2+0rsquO6UIpRFt
2CSnfpwdG8yDQPqE7GoGsz8wE4Gg2297WZUwPq81mfHf4B+B2GCW3/4FNUhjhZ/ZkGMR9ar+EkI4
UxCRAH/5D+W8Wta5TFZ0BDAOS/ZSVVCPhO/XzLzaExCtv2+uxOzzaDURaAnDF/9tTTqAulLjONUo
XHZYaRTNxGauI4fzmQRMJq2xHeHLt2V+UqyoH4JT2IXGL3mXctGqCQYiqRKhKmg05hohwWEXVT9L
/36NSGkA0emMdjxjhikE6i9afMfljt5KvabwP15lrV2sAoVZ3MS1rU/Rx05TdtDk5jXSMyMTV/HR
V1gmcTeS7IH9KDun+YyCrQFlTVU0NL76BBr+wedYRvEwcKSGUMhDsJQXzS+a2WKnZqwKowhcSFk+
9Ho3nM+Ep/kT5CGT8nW4Uc+ITkfsxcjyxuwen3fV2KKT0fDTJDyeM5na65iCWSA8DoWtRQVlHjsr
vydFEgSuMT3E/Dp+F5jCzqXm5oxgPbZIzT0GVBw3fwCOFfxwVOPzHBDPMPr0AWbO4t0cV1UjqaCu
L2mfuH2Bj0GOjHcmwwQh4Ub8fgVBCZr0ed3BndCGHf6EbTKlSZuAheHuoorevurlfZ1DzPJT2jhI
EERjhPIDV033zxkYMU8fmiMHp1Ux67vmeG2dN0FlKS0ZgAVlc4d8W5gMm8uvy471MywRwONOEfql
BPu+Z/ywSOPff84vKtOmBfqbWDj5132U61E5mamLpIhaeCTj2yfy+c+8dDQ0mfYQo3MsNRjEuWyW
d0ukZUbtRWKSmn/c7n8wMnsaCzg7DaimTYTv0x2HaM2oeL3y8XTwDTxwHfrb21EikHxZTd84pjV8
VehxDgwMdCZSciHk8tR4uHly5Nqn8rUfxxSnUb/hyfMmwGbmxj26LMdkq0qCwnv1U9c77W9CmVdp
ucieumY11XCVRjZp1knVMdyH82+G1UmYqQtJXJg9qGKAJGgHHbATWIYeOafsLy4vlEbyArtJSp1N
Wt08gba5tgLTA+HIya1da7Gpp1KF5a7PKJylcTosx9LIKgVe3AReSk9kIs3O8Vk+lWYDqrWwTk47
Gv5sqWGmyItL9C9gcy+Du6vnBi7kVDZaL502btDC1ewjMXolAE+i2AfnW1jDSve2Tb3E6XTFOSfS
r+4CjR1oDEeQJ/xxfD/M+yd6T46dQzEzV+3yHj7XrChGHYUhDkISY/8ojT+bgXiEABZ+iJCNKF/G
kYkXjOOhh0G2hpR5prxKMn9Rb/lB5UO4Kpqgfop0JKIJ1aQZYpoW0XfeGO/7OkZhSFJuYkI36fzV
9EJLZPY0P3BK0bwDDVKm8HUikvtG/BFKTQmDSRlSTxowdYEbRN5MwNnwzF53qFXtYp2tRhea/VDx
0ZKR5/DYHvJTB2Xr+ltS7wIOJbPBgnnX6XxXQFI8HvOG1kvNhhZRpnbmbFO7FKlxazvtqqQ234CV
M3Kv9dRyBjc8JCav5V4sDRpx4BMRk1RukTMXiGBANaAwPOSNuAtz5S9X2xH62RfAHfiZHU8oUP9N
hy4CcS5nWK48JFJ6pRLqRf9w38fDOnef8zSZw3eH8uU9m4ToZf+WiCh0DlROA3PsMNraoakWNG5B
NYxmLYkVL/Gasx1SD6AkNO5gP3UimI4FrCuFR1uE9CJTyAJ6de3L/IQUCV9mEMMPCsZpJfkLZJb3
2MXwuOw3+nrKmYgk6YNN7ByXVxHWMwMCAKqtxe9XYaLkAFzqlULH8DGGz/+EyY98a4KbDhFr+fLf
1js2J5AhTKmKmVyMrrmK3Y4r3ZS/trS4woVIULoguRh1H/eJPw6HUt7xDwlCXVQCztoRWr0Btygn
k/JEIrkalL7ivz7nYDJaYCpMXhMIbWb7DmOuTLNSU+DiLEON1lIyYNblr5x0UAF9pPU9CNjQMAZ2
FnwSmJgmP9xPHcCfzBPRXt4ZhqwqqQGOgGp6eipn2RB3bFDAy7z/VX1EGUFPjigjUC6BNV3wiPvu
jBUuE1MkLX5Uv3r9fwwdaPojlBnmvmYHaY10H2Bz6xbLZPbKk16BP3UzrseN573+SOUy866hzUHV
xiAXuGWjfoBhpU1m+/AcsvFSjhMNEm+tXyDHn8lyLcypW/hwT1s9cCnOAYOXZEf2tQy4TtRKroN5
6xl41Zvh4YsrMhgWIAAhCk4QkT1OzvVRkWMYvpdteeLl2ZhiF0qgzBjL4Jhu4TkG/MVwnX6Pn7Ej
Tz7V6lKZNaR1uYodtkk5NHHz2igFrrjJ/GtrilflU9nnfc7TOoctGUQhB34j4wsTHBPiwieCMoz9
snoBsqu4QDL27XUlKR6UTRWgB0n6cKXMrcu8ed3UuyIwKqhISx3rLl587woCdtAjagyVD6AEsn4A
JIRq6NcrceCy1RSS5rw4OyRgbL//mZLbpNEzLcoLx1XKUoFKrTwKykdDOPt2GV2MrlloHg6tq9x7
nd/pDKpu/zNx7Ir3XMAYWyWDRayXNo4YZbz/jmlaf3KS/nKDtrxAbq+B0OS6HA0Oo0blpxyCHlBb
XdtXv5QlT0W6juMeh6BoTNsG1zEmBBEjgAx4MV+DcoL53eQwtKRrr+ttSNaOHhQ7iejHwPTsiiS1
Dr9FRyAIwZogxmZTU37ttJ+uOUZSOBJaP9lhY9Naa0xz9yEyYWmBTCsc0yk/YN2IALSfu06TZL27
tPznRHINzZQeAvdjXl6Fpxw4JGoPKPWXqVs/fL9t06Etn9jqBoQouqgQ+h5PCSbpfit7jFCp9qMC
dxGZsmykKAN25QOmdO6Nt67KyTtdg40zgTeEkwWSj4fGrvm6hb908nMvYAyiePcstFqF8pEqlriQ
ayf545a73MQVJLQgFG32zHTnpIf8xd1/MkWOj7OaRJcmIxcm9q/VTUjIP7whOn+FaTt4bvTsmYnQ
WBCnqOsRvogx+1tSbyGvcWyqBqIfx6nAvv2VOySazXRKyPhw4+P6ZNbpY7GwMPqsj/rCH7n7hlWD
4ufeH4Rv3faMAAxB4Il/fZGkYRGuZ6blvxn5LMk0I3M8CNmdVT5T/QG5wqE/2a62sCwqdMpOMoMy
jBhj2YvadaLOj5XSAZKgfJUG57sm8U40lQJUx2OicJ+MyqQLpI802r1Y2kPmaDp6vUIitkDDbxXC
jqreDrwBhe1AYDVA7vPUolO1q2lenNb3UT2SCSw/tyrCPwb13mM97Bcx2cZUIsPryKfsdyK2kT2G
R7KZUiIo1re74AkVyoaFDqEe9YjtD5u58+X2KbM8j3knRQO/QMuJPkJeQ7KBq4jKJzltg7spj5DW
RAJwTmo2hThj2ymTJx84TPSJebgdR8/K/KkTLMfJxTO282QzZQyi+1GHFJwdl25DgmFDkQW1sKaI
Lio53Bd8b/9dOTT4pgG0srbIsofp4K+JT4DPNnXjL6vRDndH3WI1d+oUqbENRF2xiqL7Tpuw3nFw
Kgzy3XjGT6yWplfPLntfy74ykCLQRW98i/CiPyPyd0PIuhqdo9s9W/4vc8bA7f86CWEhACDqLG1N
yVDCn20yudPT/9QezP0X16BFVbjxFnrSyPg9ZTRCN+aRPKKmKgLXgXj7hrkBur27EYPs+WocoiLZ
B45JEahSyupNll2QUzq+tleK67heUk2uhBt9PIIfIo5uXepnwSym9JBWN+94nSlR6ZKR8r3roLJ9
G2yY+5V5Bs0gyNxwhqUH9ZaFs+aIOy7GDSKrvGqFbGT9oBieA0qmYHPrv4fbb57Xn3hYXelPzkxx
bL0FHLXyS7gDlZl5XOkLLpDKyzxK26034/0QINsdllflQ0B0mdAAN4E0hEuW25BdYR2O0EmUUUNI
O2MJSQCOqb+tHnKo00yI5YyUxR92dVb5APSOsKr+5oJ2SJnPCqiBlIjdWM8Ak7GZuCLRIMM+CY34
ZDy9UJf+WNufO4pmDKAP9zfZvSpzCN9wK5tud3Q0jsJXCVRR6kN1WcjDpJjs8Z4UbR9fnLNXphux
hp5QezFiX21Ew0nVEvzag2hOokl9Ha0hf7NI2JKfbWDsdynJoIftRp1F9ZlIL0n/zCDwBVFFQVDB
K+mn4IR4eDCcCu6SHzau/LafxM3IR2HSXRAC9PPhHEBJsUv3fl1mFvZ/QHuDnhygWWWCx7K4249B
ZTk4aDBZ9ViIcs7ABCN+2Qvpc1jJwtzIPYHinjAopmHampxPVZX7kpu9W0/VVnImZIgvrMhDVv6z
+fsf5dEY+4t67cWmSuSe6MkMDo8rETG7CSxYr+J3G65KpJfV+FuyWP3NCasCLcErWaTrK0ShVLbv
c27Xneiv6rp5iQlK7TnkSQ1coJtfjt0KVkZ1l332WWC1yDHoSOQkzGm1ibhj9CsqjWxUExKkFo35
tLf7l80jy8KH77cGHHPAT0HCf+Mm4q4e/5jsZJRS11P0jUbGog8A/ufT4OQU4PrvKK4ammnNAHR/
IrWYn9MR5RgfO/xVFIr9fXV2lSrmzixRK+tgPzE3RHO7rrlfVsyty24G941K4DiLhE86AiNJeADx
LeGr4snImP0gKI1nJWmryu/mRQnqUU6o29uvJrddsD6scHX8H5M9lHDi8/1WMxUr3Q2Zw5EQdgZD
vQHArOK7QTBlWnT3YPIaccwYU9vtj9QgGFN9Yq11NCGv7dnv7rNg8c0JiUUtrhv+E+lCKV0bExc6
FnEo33yOeW7cy6Lm2MQCXGdNE6csPvRAuOw5r6elC9h3w2TZ3H7QDY9JzyF5Ca5Dd8soJ5We/qP2
XrEvKyvAnhi8rxzK2Pgdlef88upjc19p2OrwZ1+/jf+frTpfQY+zb6bbnFl2XZCVRk58ST6lrOm7
hWI2Peps1AkHevZ7W5if5bUpZramFNj2glERB9uWS+jbap2yRUOSXdB5dnYjQhrOqYNLPYi8KJUV
lsG3FvTt8h0Ie5revfClfy1eK7xB8/yDgRHWUEa2z+dkGrQdr1ake/F/z12FdVSzgIxqmBzi53ap
R+l/oc+xJkuEkFdrR4prb4CcoW85uLBijr+ejfW31J6jfxLOJU+usF0zF+Mvr0X+psaepPtvDM6a
6b3gu5zmKHyBiNQI2zcOktrltVogn7f+23VsaC86gtMSCrSQ0bmSh6ZsZFBTuSj5/Jwr7AaSLkPQ
DtbM7yGF5clZHLdlzpjr2KqNas6cQD43aRqA+Okq3+T+6lWl+LTomVeUYs0iq5aMMN9mLLnq2Cnw
7UUGqXfOXXRD2cJcm840+uSnR70NuU8WOzt5OiAl+4gQFD3YlzQwMsUBScCLNQNEqGMJLlRtajfS
HIEsR06O+jnpMTMwfdqiG6rD/oYcXu7acN+/leU5VmyE6KeLLMogGoW70SMzQ25ol0lGmbZyl6wA
/Tt058u6tp9OA9pHIvhbPfbVkCN1oWCIkf/6kZ3QMKjSdKb66Tsyy28NfNOYyEm6qI//Wn7cptBW
5gPB5QOWaVxPw3JKfx3bRagu2IloDXtYPXXfXv9+dWM8Ivd8vwT8hIKmqoFgMi72B1xb6UiQwMct
FuVqJ8TBjv8KCCh6o0iyEaZy1NprFZnsuv7t/+pFSutAnxBxyXAxweeqxTBkCAebBtcDAIwHM8df
ONrpYJVGRF4S6DGd/R96HbagE1Ay5ck5+BcFE0xusLtYJGRFRSz7rWlccIV+Ek8+3HqYFz3C8D6R
hM1KqaFdxA45+uzTe1Tu+aied0lwOmLVuCyqaKHiIc0o6yoPiiEXBYL5pWFx08DgOxM4F4UIdi32
mpyHWA+y6zYFq866T+g7iYfAtXQ9xY9mpgIxVQDvRUMx7IPiTEfcj082hEOkIaraQBt8E6S9RtOH
LgnNEcUtGfCA1MhKvARqLD5qJO/KMABeRPgR1xITA+oH0zenYJwQbs7QYXxIJjdgk7bYZp2wOoqJ
B1805QXJLPfRa1A2oEHrFWOpURO2dixtD2AHOVqwEEYXie9qg+c6TXNs2ZcNa0eU91BbJifrpzFg
8ZOR5GRoAP4qXpdlbiuHh7Q8Tiaj7x2oEx/AzsC68mjdpMcka4EGmUt0UT8NSARHKOxwFsCYNIc/
7qdWIdRrDEuAUJng+TB/R2mpoBhrE8rwu0GEfyLz/vnvb1XkaoNiHKArwMjU2v4I+nYGEfsxSGmC
GfI9ntfA0HPwCVvNWZw02m5Fag/I5MIl2KTisa83bDFm2Qp0b8qN3vrhIkssAjjr0jmZZNr3MdEC
+mHajLn1tZ6H2IbWTczZxEtweX7ynAdN0fIgEx/4o5gRz/zDFgEAPKBGNjqSMN5Pr0idZvAY583x
Y963oLL29EmPm8A6GbgD+dGe9+GQCwtjDDCp2CTzqN+f/YG/WMarwBmBFZBNugHwnvxKHavOlOYW
5BCCgwI/rZTiFeiliLO/BS8s77AMABKrff7Ky5rZk1WytClcobMqISD5rglpHtwXh67Xsu79sYSW
jVL2uTBsz7R/OWYEvwNQppqJ/n2eg3QfB1ce1h9B/lpkBuEL9WSRpAJuFQxOiO+xbyJPhSoL10mC
SSzZjyW6286h848Z4ywM5Z/2VmD+1vzFsnx80r+Qh0ULjWVcx+z8Kp2RAlLetVms34QfkBSkUWJ6
+Asbj/4VN2coklJMDwd9r5ZfhqcK9/9yKX0uyIRX8TBNMibeT7wlLZABcA9uraMi9o/0pDhs55R4
KQbBOomAdOxASkoBdzgWqI6I1kyaSmsJ5dLsoSbYA392qMMiLowYvFL3LwBwM/H+CEtcQI6SEzQS
Jk/NWsliB5PtVSfHvyp9E0AbJqRvVmIxn4cB9oZQURqGl21YouMQ89GV4JWSxmwc+a2a3+OJH5Se
c5F5MPSKczKv7p58k2UJlLBhiktOyscQ+PK6Y8Rf0jtneC3Zn+iQ6NFbrxhbAiFkK244RZ9EkJ4J
eC93ADz/Yy6Goary00XY6XRoeQb6slMptj8l8WS/RujqfR2KnFwRh7gIyuoXrGEjbBwB0YTL/+zG
H6GphhIdQ1CB/eMXvYAjNhHRjEm3rvD1VtU6uiEq8ZLe+IkCqGMqd9c6cfJtz9IS2C+1HXo+xWBQ
gr7uarqibFScizgZxFWTMw3+S9C1XHeJ9/MyntuUQzDpaAPrZfxnReTTSF9zfN/AIlG4NdUiAeIy
mA1QGHWj6zMvBeR0YZYroo23S0/TB6kIe1xdOSYeBTIrNsQCsv82oT+MYMHnx3meiD5HZRQRceJ3
9f8+naFyHuiAtzjY+mcoobiQ+BtX7gEWyzGOQtOLA2LpPU3otRGzRXa8yGcdO0tp9tKEYWMBtM4D
pOwho6iWM1HFhiwUypTcLw3myaD4aHPjSirHkHv/NSq/C94tXRAfoVWhG98ktaTahOsikK3TRIQK
SjiJ0+P0324Y0+4GpkX1FdaeR14N6BxDVevrifA5mpW9Ojuf9fJ9MrE+EUsWjdvTUWtgasNiclTT
YL02GvU+IXw9wFjvkdu/6WMwpIBreEDRhuwidt+SOqVJydHQhHKcSQXUPsQ+jP/MtfBdV0UcnoNU
3Xm+v3qghvVXkjnegK6QQiqoBdN4fek2f2QfaBlJMRkpA0mXOdKBePB0RF3l4bVxA00+3KYu6/EY
Msn+pTwZZWtGJ5ZKIs9PNTTMU5GgKnCnbU/IcGoiEI9KcJL7yy4Qke/Ru9Oev5EHlbnKr/y/KaMn
HR84ZHv9Wp03ATeuLv1Z6KZugW2XfOIMpZLmpDNEUO+xRCvXjSjNPJoyAxoZW/qemqJYMn+4apuW
/2kXqoEVF8zWXtYE9sqrmC9sn+11Aw5/NcK4sb5IWSs49baHdbbMuS/k1lVLqDnHgb+xhNWjyQUn
qKJ2ay5mWUm4Pfq7oom3DX55wCBvtf1Ru9YRCeB7E3yphIJGlI6gsz563cFFJthi5HXtpZAc52X5
dwp93WmQI47YUu1cxfaQGKxHZxadbHZNXNEyj61mUWxLD9MGDbC5LkbTDESE1dR3GVNuL84igP7s
AJmg8R3EMTHFSMA9BrQ4aohMglCvLpt7RbZNOuu0ImZs9APtOrgsLkUHSPIGvmoZX9SOnn2M9BoQ
xXFAhBGbPXNFBSDdRLWTdS4rGZmwtRhB1+hF7PZurezB+57fLRyWfyr/vkc7EHF/28fjo6m/CNt3
N1CaoyPEVrXcBVkuFg9cg+bo5h+5P2pEEGzY2SCKLxqLMtRnAC46wZiX7tZZTahRphEJKjF+j/ol
kS2J8yhvtu6VsMmmzTA6gA/gBMHt6SQVEvIgHLNHifZ5fgPKRtjik1ClWKr24KOFvzSt0x4M/iYO
UsCNXuPs4DSf/QGKVf5obqpiyfI/T1ZadNpPjMCnRzdByMcTAAokzsvH4Gns0YC1wQQU4l9ftxjf
hnurXRt7jkHQlwUggqPr8u/5+fVfj2o7ARALXs6kymSWpKjcGE86lMMQk2pOA7HIAq7Qj7Z+Pkn6
KhoNWZrqTtexBPLfIu0DIPtUEdJiVhUsFH5sI4FviefT6hG2WjQUZ0menzn9cR9KN2/7tcWQ0u8Z
fOENDfjKmTnttnQKeMFFmSn3j+g3dvni0db9YSNGlBTvd1s8PA94OomWNo6vqTSqdjGXu38E12dU
aKBqUvvTEnDjYoXoAyvv/9BpCzjOjfu2MxWDzMQLMpAak1bN0DpRD6MseFr2Iqeycstu9SKvLwmh
fxlpz+mJIQ+hmJWhdioBytmBItO6cjtLHVT7KaDVq+x5Ib9WyrLLK+TuP2HAIjB5alJoae2vX8xz
ltyuD8q7fQhfiHOl25hP1RnZctARLBzdi7QrmTPQvuJXCEA8MEUHJy7QC06hLO3tHAw/UvKjufwI
pKnm4p9huuOuKL63mZMuaC8LiJCehL4EU4GDOopJCSV2wGlphVXPsUGn23urBcaX7tHCYVcmdFg1
AlEGiCtnGs6QH+sQgouDWhbT/tNId8SJvvmkQku0DkUr5jzjtueHSkZDeQ7X3UWhu6fdZyBZaH98
1AaaQ8F6nPaki6HQemVC0tfzQVubkna0roRUPaUgZ8wZWI1tqsk16sLwKpKBgrZeyaDi9TRPQqr3
64tE1rb9sbMQKnM8UuDN6EQmofABp0I3Nz9guEmAQK5eFFRHMzyDhNHMjTM+GAw027zhDMJ+9SL9
mpkD+qtT4bG1jvvOneQ7iuj6i3HI0hWMwSgR6rSRwDjpu7rmPBvW9Gj8ci+5l7H9xtueZ9RMZr4Z
w7A4eYeZ+lG1Ucf23yccfreQDS6DIhMzb3P8uf/h/DQ0A6sCpALP+LwoaVhO8nVY6OMDiwsKsQem
6hqQto9do/sugH0wzK+wDh486jD9ui2zl9jTnE8xoA0H733t1nLGpUos7gAFrQnxj+XXCBkNvGml
lzinVtkpz1Z1YAqpSzPKxoJsHafrxfvLhNZxGGi8cNPAu2IigWeJfqykHOOqw4Ylc1g4ZsDOBFkh
1CpT5ftIdD4yXOwi9A1Z7PQ8ieo/NXkNgfYoeu3TEogbnk7VGp0Sybv+BBWW/jC0j2aYQtnaeuTP
xWbC4IK6qT6BFfR0M+8rB0+Uu4xzsuwdz6IJnucV6nJJLYwBxiYI+wtyZfFcxncfjxTIudFqOgMy
hLl1OmHZ6RYrG6VsgdBJYI9pvJ2UDB5pP5tFGPT514Z/8T5LBRYMy4gAMhOeMSubAVm5jCb3kpUp
2Mr2hwRR5ceHy9HxZr9Un5JVQ0U2deCPZzzffIQjVIoScFmiaTW2y1VKXl2f+EoHCfvA6qXbof4m
ZAPpP2qtEhgCdRxCzrC0S0/VowOxMY2NSt5OUVdwJ4uBDwBYM3rL+xpORXcUx0Q9vEF0rZo7kif4
WolwtpqHiDJSw/FSyyZtbJhnsGkAaETvBQc4gpdoAqhw7Wo6vRsVQg+bIEV4NK1rlgPHydOUiUnI
tMscBfbqoz36B5ErtzJjrmUR1PW/sx7M4TzAEswTrRdAGd2ZznVPi3H/I47qBGysjc5oWhATO6xL
adFBZ9n9JIDy++UfN8rD7oT/X3AQ+Rrj4wWwP3egUXWF0b6T4YNnRXOSbqZGDNpYNT/Rx3MQVzsV
Jyi24hQ4qUF1taKe1JF7IU/mEHw8j4uXU4vDTG5Xrr4489Atr3gSGcHHbdvpEew8Q8yCG6sBi+v1
FepGvQhMWX5oBZy+7ISy9FngUddvfY0e/4KXSwiRLJ5okQEqCDmeSPOkNiZWCl9ISJLQooczQcl1
IRFdudkljQ9XFrvHzTuVyXE2HdVg5RNadurtu0nRJWW45uXAD4UHQznWov8R3zyd96jDi7mZZUHV
tC5EVJi53RRoW0soQDPZGGXo71OLuAJcdJNUMUGCC/Jf1w12Xkb/y7g230Zd8MQQkqzVRTQspB3K
GCtMp1xtfFRb/vlHekYMY1zRdBdfRVnDJ8iu9UpzLiGBSporAKIaXK6rD2tKV+/KbA0MnGOHQhb0
ZuQVNqbmgdnWdCHXPq4TuhBe7vWZxQWSPp13aoiU4e/txlu0f6wzpMWCFplpSXM9rsobh0pTaGA2
wwIRm/WSbaNxkLaWAEbTZGhuN0AQ4uplhtmzM9nlC2TisEFCTZ8wR+o8nZkcQFBSfSfL97nWyWa0
lj7ivm2M0ZSejF8jBapEZOokHbr6t4l+Tugvpf+0GMdrUqWZSfSFNla13ZTFXmt6ta01yYenNKKj
GxfokbR7gnH1Aq1q0fCSNcJNI4lgVfNDrQzfWN1k53D4bHLEOaw7Kumh3xMsZJZZOCuhKuSi6JRn
jecrbBi/a61MfF3EEwOkyfXa1pCojWlyL86jspsMUb3kLGz5WGUbZLYwQcjPY/Rw1IHPORbKRw4Y
wGiQHmgjdenYKOqPXwPfLtjahVj4upe1JHEl49iPPa8t6s1NN07G6iFCJPbjIT9eJCSeBLgtoQ4j
hnnMBZ9Un5HFieRRg9KovGOcmKivIEPrPhP0xO3p2MceHGhmAu0flacbzXBp+ETmi/fWLO4/8vAm
5ezjTpRbuzYECdCRSJRfKHggpzefn32k8GBTDZeFt9ZnzuBiX11nlX7z56BpAJMTIp70jncKFMWY
YQppYCAsVSNE50sO+1eXh0pJGz7/cCbH9yNuehlgzYH7BN+oL9nfqUrynp1GDO5Fm5UwfFlHBJaX
XLBziCEcvgaA5T1KDCNAqYD9JcIiObQslrcAOL72YNliISX55dkcQhDwvo4LDBvlgzGWDq4qBugH
Pqs58tUTbL9u7Z2l6NKiY+zi2iHgRdl7irwlzx4K6ij+agnsdAlHCvP1w9pIh9tOQS9FHop3J4Gz
tZEg0FNLzAE0trLdvjiKTcLKqFnYj9q/FwpxuhZZhZJPviMxK8pzHw7t6YKU4v7T24RcQ4l1T6RU
7LLJwbK/132A+CjwfIolfRQq79iW2knakzghB3cleBLcPzQRIg6gsU6cSsbPjpZqf2l43NWZQABS
hgZgxNFQCyXGI8uVT/kwNeyIMdqVGgyiRcu4ABVRIxCeDNYqapaL3pbevcaysVfVxiZDid1LWiYM
xFZ1tb/rNA8HdBVBrdPKUui2thKcdxbmg1yqHHi0D/4TH5k5qvPXl3V1loXAxmYN6X6k2qrTeDyA
M6uQT3txqdl6HVV803eW4QmOE4rJ1D8JyxOp/xyeSFFO1XcqgUnpLykk+1/ycAcDKGI5Imm2RjYq
2I/62ywEqtp1Zcm74Bn6G2x5H19KmFUETM3hUHNOkqz6qHqqsY8KQISkdaiIQsHIOtu+4YlP2LIE
iN7oQvZ1CQKqIVzO772apVHydO+1FXQu47K/x3PwGmvLhZFnpUmJs4qxBu28GARAOvF7c7xNfDDm
LCqYmM+NT39Ry3AoCskTcI4U8OtELWfDu/bQn901EsX+6/2go9Hgn94qz51EbriLwTeJbsnnJUL1
UrVNh6qAg1NOgF4+Hfw8F5h6L8Ex+bL7DUAF968tAu9sIbifXdkOzA7oI2fw4NQkto2rNMiZCcPM
4GfhmFY/gUykmPoullyFgYbYNcYqF02l/ep19ik1iQWj4189TQ4/OVeenfJO1QMqksDGJ6P5TDwB
o17eD/B4YduffGHGvxqRX6tYGq2gxjOgSIYkW8dvOay4fEFK3XwZeUR+WfPL+D43aAG3JRUh5kWz
VXNmgimr3PX8IaG3Wqtj7GYT/kgcen41aW3eqC8OdS+/w3m4Sw5cZi206bBI7k3fVomrxH2jAEwk
vQ4nI7JL+vKE1PwXNhD7FmjrbAdxxFqGQs9aIMuwcA4t8+L3n3sfvy9UaEbSmHJ0jCCmoPL30eRW
Ll3ZTFx6Wf3qhthg0Jtpk/tfOyb8t9DrvAR2wUF4kGCTNUP5k8H8AM5fTJpxwi/Z7rklPO6judE5
nfmr1oLNRApF9+g3sYZLE3WB9IliApBW0z9FfJEDAwh44h9EWXTOkiEZXvPINWOjdLE94pMWfFWJ
0GcVCw9uHu17wfueOjdr0rbB+4TePVjKPw+HAdm7YpElYwaN+YBqSunWfy3b1sUUBWA+IGZGe7mP
rXcJamn4Q1D7ffvXiDzC50mxrJJlfB82lkOpTOB6EdIE6T9Qz4eeRzKerYemYhnvIbGwI/gC2XDT
TRe6QJdL8FuLOBKbaGKpwPp4tfHmzyQ+Ox6mwxzUI0rI7aJbn7lW6b88JtgMRcjnsXT5I6L547tt
UAELGYm6zIJBcQ3miFYqRcrfoi7RCX9MxdgHKqxx0eGmQajngMDCLlciIDdE0OG6KbphHJXewEAp
pSfz0pDinfpVyC8F+dPWqlwuKzqYQaRJYGUVk1QOOLDyzNlYZaJf/c1rykPanhu2UpoRgL2yUAWl
VPJN+8wDTWbBRkHWjbezsFEh5PFZcr4ST+ZhkR5XEGyW6KPPIipK4NvmiYc+2uj8BtdWoZnENrTy
vLPucjguW4GDLbVb9yJgFzYRTHeWUbycxLY8aTq0VjX84B5haeIXANpj/c8XV4qb0joMKoxW4er0
nhTNPWCn7xohx+gPC6V+w6L3WI7kTC+K10xGR/Q+n9S5FJNL54nNdziK5aoWo3D2+7juPTCTw+jv
xeFTvuh5M+XOCpqZ+kwfpUld3DuBlNhtOsbRCm08F4xK3zEwxQIwxCLQuzVSczb2P8ClUOAVeOZc
ezWgOe9e+lNvt5nMjgNLL0jikBjXtV1Q19FFCEDzjyA/TfthCx82olHWU7fe2xrJ5ydC2k8stl86
QBXDi/CDBtlLGJOOv4hofKBp5VE5juwp6CXZK6rrTNnwQTSB3oiaTsXZWgrLpgq6N8IsMIJgWJbp
Du0Iz8H5QxS4OWpTz2x6f6Rfndm93r1iEB43vFELh8g/n3oNzK2OO0rtbCSbF+Q7BHvbXCvoeZ0f
YX0PXSR88zWjqm0PQtGvXCqtab5owJQJatGWk+pXNOmc1coKQPOwBq6FBL+MnTcXcR2aMGSwTmLs
86oayxheMrUKIBunZN0aj/bJZxdEeCiyimFSLPVEYXJNqRb49WVX+5zkOhOJsCY2xMVgMaG9BLjJ
MqETggcxqRBc249AbIJywSAhCDgCnScggqQsbJe8EUGRxXlSQNfnDCzOnCap+srUDzKbqg+YsAsW
vT5Z31TTD/rURm9swoIyIOABa6K5NxwQ3OWZvs7W/HhC54Nxbw9U+GNimhwoq/UWNeTMV8+183hK
WLb4UEnuFmEHo9/guG6WjcFnokMCBQTxc+bUHjv9xLA+B2vyg/mooW2DcWukMai2KiRoerAsDkmB
WZ0ui/pPr83vA9TLnR7f+o3bqXT6rAH4ZhMd487ihG5GfJm3wAdifsbJg6TlvsTIJVygwwBajMOw
evUdKO8KHkuOH4OCLYru6AsKzSnqPXlaa30WvFSmoREaKhebLmQQ2+dL2rrOnF6rIxmUmA7c2Jz9
fso9lRSZ732aOMjBF7U2RHmRsR4H9OcO6yn1Y8q587lsFJnY7YsWYTYqD2iyp67iehlx7aNKKvAl
g2BA+By1ZifMuChFbhEfoRVbo5mdT9V3FuTDPDn1g+2Yb6g3wIYWDKrntVZLBcRH4qcJz7VARpYM
5+ymzRMzG7gGU23iA1HDrWpfoKWlRvYh4cYuYo5KyKNypnwma4on6lUDQDoiOXj+IzDN3lAF2TN7
z7Mvzr+Rjku6isTvuve5Wh6iOMnvm1tBYfntrjOzb00iNHAZ2EmQOaLSLRT55/cnoipH7WuPyvCA
xKfmtNGslercXvNEtiThQH8kb0/Pipp27BOXyh7FNbbH7begyNLyub2woJ/IPmGmWQT9zFAuYIsn
X8I0sVFIRjaQNdb6TXOK0d5ZDpIjjSP8LgVt5UEXRgs0KNrtJ0iETj6OM72Qh6RyhTLYcdpY1h9V
e0VzPqy8CUYRU3vvnQPk0eOLivj52KcU6rWrtDXJWQaGfXvvdkT9KO1FPnU7GiWKu6Bc4vdvljJY
852i4F0QJOxcqVYBEnCpf9ollmwuAJ2ez9T5pmYwWuFKG1ue7t2+llNwN82zpEo53F28Zem1Q6CY
iCJK6OMq91dC756v2+w1SzbAYPBJ4pSHG0jDZHbPfoNg74EVx5tXyOkViN0bVgZFhQjTki3kzNTH
/qI6rP4y+o2t49KH18DaGoCh4pz4dtv5A2HhAAAXzY+Tm4njkBYplw0z0NQERCMeQQCE8wjA6aeJ
Rt8/sA7aF2eoPVsB6AdQRmn9fNyuGDUFZBaWfK7R7/Edyb5ogyqbUVX5RPpjw8xyKMHg5WRX+rFH
zfWB81TRmxrsJ0INDjqBAiYsTMBLI3/7Io/G9BFG3o5dCTyQMW7Cb1f4bde35MOqWSh5U/IWKjBC
keZAFPA0Sd8/640DHD7fsCGOBXQmcSrJOL0JsT29ZV/q0xvOm0C8toJOqW4W+xvd0zHMoNtf+WSa
a3jxFFjrsrmycVl0GlJoCyjk9JRYAChfGhPIEcHeUW9qQEJ9bQuT0RWFKnxhe2/Q8T3ld9VTTiQy
BLw1CJH0LIrVBOwDRC4JN6dQHd9VDeWIUxchP9lU0b/8dZl6GF8syW6k4k6dHpPFGcfl3QLNhs1i
lJKbI730u+8FN+0P+DkBOu3MdY2JC51kAON/E/1PXCAjUZl5uXuAVKgeBEQ84D/Ra9kqQ8exJAZZ
Wz9m4M5hu2g0gRjG0ULoo7+S0dJdsr/NnGtd4Z8S9w50+wmwvYyxB03vRMOz1VboSWUwrYu0P+zg
TXYbmW/6PaXTqt4DqrAzGbeuLsg4rxycg3Z3Np2a1+VEmGIdW5KD02/a3PpbXc5QFvD6qV7vkh4+
80tumYkfIMgi+M1EQfLJtA4iNBhFALIHpFTSBMvPS1i+w5sQA+CPmMPfe4/fglguuwSwzjrWSQAA
1D/hPnuqI6QUdiFmQcDClzBBrLTzsAQ3sM5iqODBFgmu4XWwqOV843tNAn7EbOrt29VwXRrKvWIQ
Q3H1FYFfsSjVHc177iv56+mHCE/MbOs4ek77uLnHlp/E4TB6wcJA1AIezkXgi5SIa+Lh7XEJA9ra
JJ7gpWe28P6LZ5jB9lwCCMSmBE6/dEwzE+GqWirwX0i585ymJ7E9Gq2Z2avtBLFZspvv6/8mtEUr
0hTHDXyEHA2wUgeU5eAB3v89qegrRUtzhKE3IjXXpG+cLT3tKoYA35ykKPU1xA3csilBPXXCflpl
7EgTTqOKKp7cSfEOytcb4Hk4MlN89T5EMGnDszxjw/K5l8AkuL3o/lczTE3oUL5GTkoey1QMj1jB
VDQ4OXc8mIcIm6oYCfmejY8NRKTAh/8XwFyaLkiecxJ/CFrRJMsUNZT8nLSwyDhVBJ3a7QbrfHkh
KskHnTTHnkG5mGtTgZZ2mkL846bu4NpjzIXVJ9dX+TuyTUIZ6INvynEozM+NDBCXp2nWr4XeBC5y
HUSdU+p8OqxbM5/CVVwq2ejtTWR5TLEHmPd8Q6oSI6DHGaW8TBbWTtCh2rTyZ3Ju5MX6J3WZwSTI
dD2dPZfORQQ4//ufPV/4jHHCsnekqkaa5rDekPZ5wMgRoz6J9qtdxxnNFrN7HUqqOqQYfYPaFUL+
1VzUUTkPWIGQ0Yv1Pe95DER/JCLTm/JnQQyO3n11zvuuXJXqD2NxNCeYXCC4DhVO22AIb5nNUSS7
lNWmB5Mco0ndShwiM9gsdbXftpeTg589eIPv0Ko6D0V9+6VlBs1sEHlmdk/KjvySNWoP6OIin5Aq
Mu7cdHXuwH7CdkRJjQdUY0GI6Iyn1k6/VgB06V1riNBYHGJ19/CnJABhLkysCtO9LMjxqi/vyBBB
ccXjD+6QgQZmW4t+jCwSJ1szx8UWPP7K2doQMhchYdvkV4L6PSgu/W67WZz1rJCre3ZOj9dSupV3
2u2ZiDRiV/9iFttrRKyNzIJh5OPlodpHa1ejdWTezolL56WD08pB636oxhCpw6TEzNhXtcDP9+VM
QnglmK6NjKE/esz4+Kkl4Jz22eBktCDYLjs4SYcr/Qe727CN8Y9IWOk8NWSygeRHaDu/Q5zXrnIX
O8j/KYZ0kLjCU2pyJOfcqtyH+L0dZBfk8qyntdvgPQjJ2UNzpSjQU6V2LQz0m2oIWouVqJQZ2IfI
d2TP/UANZ5pO0inCy8LGV/jDdwZeKlSwfPY81yJY0HWk17yb0g09qKEBRKhwDA7XI0VSSNRg+AJa
XuwVAGQu0prCg7J4uEZyCUqB1UCUI+0/YLLlS5UAWR/zGukEwflikJeSHv2juvmmTIc2l6+fd1X/
ATbz2GRvQ5dXiVagsI7P7t2iuFd6r2XjnqXVsPLg7wJG0eR5T81Jw+fYBYB+7WwhbccgmhBYNkQa
dwKXMeT5YtUyaaEMwcNtmzB6onRZxl425boL1wuY1gZr0B4ch7Agt+X6VpkmmwGSn8cnoiFzx+3E
GgECJsNct19691YZWOfxsuIEceNvkOiKzB8cT8ttjmMDp0tTT4HWsWEI4VoL+7ILHBk10p/dZifr
/zWObyzMn4JQHPO3F7+ipQEtKcEf6srd+y+wuyYtozN6jt421juCmueNB2BtpujslGrH62h/duY/
RpJZhl+mFajcbbIAS80aesRpxvqceBkONRcJ5hQ8cicFTdQ7xIDADrNEVsG4l/QlOfsh3PSYazzE
KG5c7qFuyKuWr9tUJrV49v7PXT7XQWq5Wso3tgQbqLXUGUrJtxMA/ezG2lzflymCS9yijYfg9/OR
7Ect7QJHLb87vzqCJkOQNeY6Ind30Yux2u0LIhQ1CEstvdPGOnyCtzvJxIQsXwZ/JgNIwVZ1jMZu
is17sJeE0gt/kXUWN8q/8kzDyrQsHFi236pYQi7TAT92qWrW/vW+GKzRk3dTk2KRD0Xh2FACBlqb
sTphIiVadu8ZFFgfraqKmsYIuXdKvwoArsT1Q7F6gqR5tBzrpf06Q84wHuSjZHJoutWxCo57l/Ei
zvEspjPEShSXgRtyh5kPCR1+7X2fqHPrRPriFPWbyQrREXO1WvGN+imLp9/JsO1XiIPiToIO3Dj3
feA88PI3r6paPmU99c6RpNFLZNhHLYvZhP4x6tQzl4xJE0Du4AtJcqHSfid/pBIVbfn0ukonlgzv
LIsUK5PVSQgyaNPc4Z6nyQWyrSecQm1iuYsBZMO76dlazhOhrPf3Hjep+zPMo9Sbi6lEqbtYW/C1
ZINf9r0++nR5L5vANe/5pMfIhn+GS/XGJ9KyEcQsxBGQ2RjJnAkkIZox4otEXkW0LD1x/Jblx4El
SVqHH5/S8xIn+7m57NcfkZnkwZLIMp+/MUHVPoy4L5rEtf2HTGXDfvFYNmF08zMQb2jKETnDZgCl
wpI/BbPc4htOc51sXx6zqA9ntAevrHxchh+NIZbcfYbGfaX7r8MbRmbWlks2QhoEcxRba+ZhDZD/
3UMTq9zcztkmxY/nF6AaIS6z2elMFTKf7MPb9RTmdbpjDdhVmZd47mzhorlRgD+l4ssBVPc5zx+Q
EHSX64tlUT0ZWk8h49F2vnCzNQeAKpaFMy56IUs4Z4riUwaUOb0L2PYkav2mLz6rNk1nxN8CVyHk
j+vbwX3ScNRmX8j/y1QBcPd7nm6XQiIr1qc0butq1jNdoXyieZPbQTlHhgQkeGlUvRg4g+LYqDto
tf5vFajhY4Acy3Pj5h/Ey7pkt2p5eLFDAe150WPklG4CsrBGHAxAEC7dzgqdXRAGOhyBWd9T/F1t
TBl/6H+2Nl+LSfugBZxdEcnZxY82jpY2Jjvrk58adLN54o3rmMwqhCkZzfJGTUaFchwN0TN2JTWv
AcCgd1HDs9frFpD2N+CN00SgtElq1PL90mSr2h3XIsVyLCyjG+02LqWlFmzlRVRZ+NwbSLuyOn+o
UJ5ntwFVyVpETwy2JxxVGe7g8W6f5eeqdh6euPJNb4FddTin1GkJFx4x+KGaILYrLGmbmIjFts7A
4U9a6jA1Ksbu0wQp4yhUssHs5ugsQK5icZgf7PBYj7+pW8jdByx46auFrK9aiYfgEt/hAzz0358Y
N4RG8wARSEE802eqLLJ1MeTuYRUTXNDkyLoTSkZ2DQ6WiSLltmsZ++8nMVEjJwIonM0BC0ty51Ut
7pGO0cPbdHFwsfgOIS8DH+tcHYksxPZf12cb2NbKj7PkSVC51fUePTRTuhv0faZOEQXLV8K/W59+
lzI/cVh1jtnOQvf/9o+oSoYy+UD5fstxNwr5l4ILStvQ+/HqnP4SndEwiFwA99IlJIU8xEPhq5cU
6SFPfXTGSM5jn5PD7o739qM9Am+C6zB+Es4bQv291TAAIZc34Y8m1jF5scks/U336tk23KFfuWvv
Jp5jUgrQQx5b/7HGET63M3MEYsPx0S7tNqMogKoIqkV8aKNwNCFL2WD5BJnYFPFZ0t1alNJ+/wLr
95qpfpojaeiqjXZ/LTDPPHypp21ke6ydqTEkfsDsak1c6/hkKSoZyrR3xNDfekSiMWQ4XyRkZLl0
fmgXKXIB3mkBU2IrEjOk8ojTI8r9f4flATjYww/o5wbm2OHDmhsPcZ/JRe1/1KGOovbGfMV0fScI
MCPWdUqRmYThHnHjtSR4KzamX5jeiDVxIOhq+zGGVZomvqfOOfd5G6kxExl1QSzpmInEcFEw2bDR
FviwqiWFrv9iHsDg1rE3xysHfumdDciyuVQQzRm+rAHPiRKLPOkZQVIdlTGB/1JvyHrvU4ykuKV3
UP0WUnPrZWyawMbbXYnwBU5+MTDZXhrOKWpYjiDxON7ifqatgPcB0M3zMsPueNUE9OOdRKl/63XY
wHFILRLPUPAqx9AqZOXciWXAEa5tQqhGU9LpwTFppN98PgEzMDntFfa5hhnL/AIYdNraJhUWxFHw
oNvhHlTAHbAJAPkFaClomKVxHSsSQiSsWRz11mUKdsjR1dPFEVmLboc/GiPc++LJMf5CI/Y74naQ
OqpNs6Ddu81n8g9Tgqs4rnZln3dmzAbiatKcDr8ZZHiDxYhJ9P3PgSQjFKncHhRPw9MWBARkwv7L
XaFwDmsDW+Gp6AoJr01y2KCM7rooIAbg7i32ZBS4LPk7UDEvo6/fxEv8ksoD2E8wwX2MFURtyGdQ
X3wH6dleL9aoSoN+MfluLF0ZMxPdN7dOMLX3rjuMvBdAgRQABhnIBNnt7a4DmiesCEWyJ8IqJl6H
X9PMJ4bAcgfuUSTmS62+xaSkI5zwt56zFlxSHhM/QuNNnWrH7yStgUl4CNxsBNhXyLbPmnrYG+R0
BYUEENWI+2S2OfvV1lBUpb2KTt0E3naTL2EXwwz3u/rXz7AWXjfWMOPmiS3ZI7QVw0fR3jTe3MVE
m4E0/9FYQBkXbKwy5gKqNpp5aj8UafwQGvbGdlFTNHqnO9Ybi+3Uv2QRVapCUn43XVyFk6WNArsD
G4k7LRiTknxnEVZ8DbCZ5kSq6K0clULhp1IeVwyfLNfXPWK1B/Fr+jHLaNE9pIB2avuoIt+Yuj0f
8VJP4Llm9XFCKOyNLwnM19e1XkeaxF/k5Qb8t4iLmsAAog8YEWYuxhJaLTZrEKWjqgk7m+Px4apy
7Az0rA/VCeqTFC4PeB5M2va6b2sA6xYV6alFz7xueY0zecKfTyDC+JhvhkpvHVLKxXmHuyBVWcSn
CgC/Dik2GSDR3gu6RHxE9BSDnnLGPiFs7KEV161mHKmmjaLYtaSK4+FjTesvwPsfxlIhWhOmDrBQ
Reom0/r8tgkyIzrC8hsVSrshDXlUSFwSgCwkkm4AIgJvtNxGSdmdV5AzdC+zkLyA0CA49FGL8nz0
leDyPm34/e7gjGODIcdf3T52CxX37zSfRXjFOb/jt18FJkOqV6qaRM6pGpjeNQikZgu1/uKbdtdq
c09k55klUEzbor6fMpTgXZahyfG6dG1iUTuywbJn961lHhPFAXGe9VycggviA4G4oDfZaL0uVeeQ
/EBAeaBUgDIfz6R0NnrzX56/G2BbWgq1bco3+3r0i4TidVhK6z9Hyzz9kX72PoHgDikeC8WyryVK
ipRs6UZkioSocHaeQS4VxkCBff4tXkoaClDJMRQS0gz+fBTT+gjWHJT6iWogzaS0r3cfhvc5qGhy
wly/qYikLfUMiwllvFke54WU+oiXlzz1zjwCqU3tr5ZxyCAMcVh3wUn2OEho6wRcjROm/hCVYEoL
nHJtzEhJ570zut3kjfn7wgedl2yW9pUWRwC2uCeTIWtrTA4c0efoVUk1MjmgA0YpwYY+Kr6kjn9x
2+t87qKSkckeEB1P7yNcFtePY3fimQKhN1uYOBUq4hjyNSXPQR4ZizhWlNpDXak0PJFGSmDd9bEM
aaPkc3WCGi/fWHPtbaSjTA/2GrRLgPMhoOE80dqJjEgb7+F9TiiZATgW34CVsX5wZPWri2um+UIu
8VQd6EMeRWyFGqzUp7eeKYXjtgck0ZL0yuom0hmYiSqGXrz1beK9l28o33zPf0nqzYHp1VYPgN2f
YX4oYFuZy5mv3kdZYkBfKg+6IEXm43OWdgLEqS3Y6LnYrAnmtMkVNzuxnoQdFuKyfFJ9ag0ptWws
qyhUiBm8R3PqHlpyIruS8Z/YPRS2fQMd/7kZHQ531dJyidajWuxN4bRV0kqe4a3cvC+1ym22qM75
9jm3qpAR2dSku73NPNvsR2ZsByLIw+jO7BEB6IV9I4fhJgtYX7bWjO3LiMPyDGZJpj/lJDadzJO2
pYDQqja1FBwbLM70c78Pb/sRFVp+WEhFxKBOz+mnbJCxN68Ti7bSnSC/rZxkUbv6HXW6ygs86zjp
FtIiMhNZzUx9N1jRDPMckuOnDZgdh1QVuQTExO9D4iauyss3QoU5UAk9YjhOojSvXfry98qpTAJ7
365q1kCh8SsiDcMOpGma0Gs/c22lzxz7AtCR0wT9jcKVy9VTe/dAkFwS9EiJeL3gwT7Ns2h8lF8C
puh5nFdf7vqIO6Hys3dLc+0DfsKvfEEbY04b/jKYLPLw2cO4zDApFxvcltz8SjtSu9u0LeeA1jbe
FIfCWxxjjXWKV+Apd+Kz4HRMYuOZwBW3wHhXQeCsseOkg1xWSuM6tW7r93j1yahCYJRESpNsE3p6
NBB3rYctkxTJCOhVnJPIlD4HhKxyoYoi6IQ9gntwczxJZ3aT4/sirz4p35RvIaTZj8EBDXDPJ31H
/26p/O9UuIxrLUJaEKG0irHz2CT/cO5g6Vbpfl46pNJXGa3X6t7V6vE/bssMiTA4whUpuDT3g3TA
/dkDaTcDVX6QoI/jQN8YHauWrF94FK9f7V/XTJj+rod4SH8DXVPXn1ZX9H/BwSvyhA3tN3KlEAsJ
cseuyWy6MhO6O5/lkgYEGr7+Up5EbVvGNogDp9RiCCaTMX4JhAtS9/G8qIuRYuHMOffNpNaZBbtd
y9BeUBO5H7p1KPLH6baGBubD3VpYUkWoIzhNy9Tnw5ZhDUcLwyzNKWc8g7zp9ns9Pqgquu06+dSI
YpUTD+hWcu+sKrKl4Qwr94dVNPiIxq2j7fTNXLE4Uve8pcKXgJ4s3D6/LF/9AsEtw1rDWoC2s7Z5
Cu6Vyp5VaeuhjA0ZHJw9RtPKSJC1S+4L20LdasFKIfv5m//yHitv/UvSCBuYqF5W9Egt0qw+zbpD
pRkEfkZsTzgvVFFga2sqRcDdkJ61f4nQR2Zdum0jx3SrOaYKYZPRExUzUiiVo8k4+sVcklrYWSB/
5qmBhFWBZFUqLd7eMOVa7qe3YjZf2J83tjsDFP9WDNqvPAhpVK15QwGmjzJfVEXemccFSE7CisV+
t/vp3EAKBCMPEaifyiYaJ0K7jnM+3SR3z/bBFoeuSLem9U/L4dGON2y7vwUjLdgB2Bm30g2dAyhR
Enrs+T1FbdO42itIGt9eNqLxUpAtXM5awRdaBUTnZ8++TgA0Y1K9u6LvOIwkVyYj01mQztSYr8hY
may92YZepymfeLovQKiFoz2p59eCqOpDJ2cYQeuoSzZBH4clKHCAvTUX+bnnGns2F2GlzYHVCe/J
KXQx2qApnjWXmK5QG5NiZLuHS/usrAU8LIIJX44J6gWtzbpkLGH0Z8n1UdHP9URvPDNvGPisGJm2
FN8WNT/2ryRntQs0dStVA73BrEwyZGJKymyFXynfnKvIVPvyoOTqZ/hZZUMTK3bP5A94+lMITmdA
53tJMISvxijLOfsDfBVJb19q0EyjpyIFyloY1UeeuNNBGl9rvjlO4w9UiE1l+/hyXdWKoeSm/zDV
g3MHzAAHbPPHU3AAcCaZ+1zRK9XNYmQ11bJVDv5tMkhWSOV1I8iDiNVMh7joTvCahe0zemM1xzK3
87qNHYvMcFnm1kUjjf3IeiGYa5zjR73dkfXZNavpmLvk5Rc2YW2R1LlnsirNQr4oz6HotiDRNsI9
MPkIMIQ1d/aPjOaTTH3cvraL9L4Kt2CThgdIIxkaDiUhhbPLPx/mGBGfLPj37SJ5pfLnrMkZ1m9F
l2G4xixGRrNlVSaC3teSF8nF02YIbD2DSBHiprEL3LSC2mLIcIOB+wwEtDbRatgodbBKyJ8kKBXP
/cmkql7la2mTfiqH7TYsQcCYqTXNMC7nh+8LAxeYbUDhqQarak5HGv9jKctT3NkZNydwkWoAzJVv
HSNLEaggUtKZgbce3dym9F5gDLrEzRlhhFokbeymZsHla2qo4Dnnk8odkb5ybrXyhe4+4hXuah4H
LZQu+isb51miLtuKuJFd/RXINAruU/zAWTxpViaZD73tOoFSyZHiwC+IvOFLO5xinCVOEPggvRtN
Q8A33On5GlKyujueKC/F5gkJzKJQuB5z0kgXEoDJj5Rltpt2KAxWqwwYcfBdblm2qgNUUodCgAsg
Zc8pUQQFFArimiRfQKquQzZsYxcfnw54g/HzmeLS4w/b10ZP8Wo7+izi0sn7+2rUIcAX9zOUPdbM
0LZQf9jlarwQjEFYit/BVAKqyGv2xNQe9iZaSYlA2G/V4ghpa+fsdwlSYdB/iiphXKiEEQbhN+/F
852bEkO16/a+K9hSOYUNvikkGk3nOYdCWKv1lHMb1knpqEjPumS+0t4T2OUbOUR89DosNNhYgS+L
Wt1cnn/ckRFTEdHNXA7ffWWHqShQrbl0xqaQ7ZGqnjIG0CLmPZeWjxk1qFZN7p1Athp3J5KRreaG
SqlHApIdWXVlMhuIXExrHBhDcwObZXDuCL9CAcSD0+wFIbjw9/+EJ4WS24xTagg0kD0T68gy06XO
SkEzFGpMcyVxV5ynELsMXpcqzpnrSiectv0SBmLx1QxXv7FBAiFmGWKcsEsMcQwHDIpVYAqMjkG/
8dGNW/cOVpia8IaGSP/a0sb7vkB2uvWPWmchUGlIiXkpAueiKqrQAiuczOIpW1l3opSjfayovEI5
GRaenRyOE2WtSTRLn4ivjyCU1ZtUeLZru+UmK0NUEWS2i7TgYK8PtyI71x69QUC3CIKPc2qa3lW9
bpCFtCk4Fe2BEEO4/750/a0xc9D5uLUq6YPM6zv9zGUY08HgsL7Y7RtI6Gx3lHbr4RsOlppO9QZV
rfm6l/11SdtA+uPyDmza3DdnBMBAy+BBs9ifg7MUF2UqJFHiZOpXnwpMtl0S4untgZGtwEEc1jaL
1igzHX3WNICDHoZptC8Jw23h8o7fVAeHGfHJJIC5JUda6WNl4lZUxf4EDFp2mFjBvjNkS/YLR7EF
L4xGh1dnqVMQrzJZclMneHiL1dw7j+YT6NXJH6Vv+SQrTrCC4zwjy2SgzWEpdivXbTGxyAOy9b+t
DwWiFghg0Fm0KZtUsqPITgyveRF4LkZm6tNW/v95ztTbFUp0mQg0T5hr8WaYd13dzROATT/s+Mku
1yLeuNmLeJU1QYoNTy8YAaBkGWBYKpeDpYVkMLGwOTT4pYmQ7W13n73P0e+OS0wowI2ZOfm8UVBf
S+ddWU5OIrrQ/pnxJoKb/qZNnZGS+lirXTFUoD9W10MDFqO7zY+jP0DIgjxMnT8/mJc8pjQ3qwYg
krkOyWkxd8Uewm7l4kqHGN/gvLCDTFLN5un+btjhPfeWmw8H1LByEezurIuxm4I30tc2CgxHp8bv
tvsgkRC067+ls0dSLiDshCqAceBz7Mndsme414kaBpeq2vx0Uj/IxuKsyK27UjiXL9rVFMnIqJWn
c81rTL20RpCUNDYf7DakTRySaECkF+vbfW8bxn94WwuFogb76pJzzAemL77FKTpa49ZmEZ5XFnSw
ZVNyNdgJHMv0BuiiiYsaVQ+2eEnPrWhqjWAPXVQxJUdxOIwPon91n8uvhcG92bVkletFIi9mBiGr
DlZWZfYR2mLLT4p1Jqv8LBOXuQSnFQ0tSBce1OECNg/jEaUIz/rSiGBVbEgeFXWyzTqvPr1DsDbH
9YtZWJFliIED5cl4geZaLH3KG0ewvfA6Qk5oRpCEnjYhO0jwhzt/or/Qm4OosA9FDhJ+QAc3rdN8
BvsDpgf6aZ8bvSAoLGClssL3NukBdT8vdUP9QXaM57CwYKy5jpOS/waRuBHoIQIcZjQA/54ttWdy
O1I7/5d1p2FARGblfbCvZ7krmylG+NStE4HSx6lEBGXCn9svngYehfcdpqs4HDqbTaiN9oOILC+g
s3xZHLSRdwhleLP4acqCblaaVQO4+4mK2bzuVYVkq9hFWl5vODtKDgB8j0GbpNrDvJl2cKFOgiPb
o9e1TxukV+/vJqZHEB2V8a9iS1Kxqf7Hmr+7j4/Qp9ZaH4mw/eX1/NBxRTiET2IqKnnjJJgLvEaV
GudJDN9e4Ohz9+DN5eUT8fnqRma4eE+WvfxREl6pWgWhl9265JWIbqol8CRPlEAyfGBp8WbkCM+6
LRgg1wkxyIPC20pyKU77d7WaNdoRRxbC2/pE0f7UCN9rn5aQOcYhHMGLzINopQjS/CUV7lJusFwH
Z7xZeSKM82Uie6hKHQj6k1VHZ1ldEUPAVg/E1OL9uYqIrvS6pSKJL+eDUUzxCNBKT0Moz8fO5jxi
W6RntGa5guuE3aMNNitIcUkWwDoLWhOQg7G0eqbVUvdvEXzFmjoVLmGwe2T2uRJBOZ7brLHl2wud
wL8xMpzxSVKDyp8FFkoTMuJqXmRkrgCrf32UPTXUwOv1Pf6M6bjHSfHwiitSvyLP2s/UJzYM0BUR
rTtPYFPxjtLrc13UoRlZQgDNGyiudfgDZJFj1Nc2BAKVtGEI+p+MxRqaq+Lnq7mULpHc0KoJ+QbC
RSqzhE7/WKm8Y5iwF8s72E0NqSFnF0RBZW6pZT2nQu3I6jupNy2fbbPQTEgu6yAwvjGnVX0B4eTN
wi0TX+vsjJH8hiflpUOysytt46jEI46vO7ozroydkIZyJs754FWVViB960DtWA/2/HtXBBGpNI6g
psEgrQjyapPHelgAoTZ812sOdjSCZQCTucpwOoiIOxJcYhffrN9EjCN2oB7EuCUpxnvuxMhaf/YP
H3liUMoJBpvg7Ij5wJzyRF/P3cOVkTyKTY3fn4gAGFRLNSh+JgcD0dRq++h0UHK9Ur38kL2hN1fZ
elqisDDIXIbIaTSEZHkq5AQ/llTgkaZ92Kok2VJrnhueu7vaw1cANpm5YpK5j3lEQclL/J45F1D/
PYUw2qzSeij5yOnr/d/kjVXiGuf1ISYhkb8dZNCiByZFApoMcXCin5YpnwDe2NyG/vaDXF5m8BYz
j2nSBLIVy2Q/KoM7Ngs+tUkCwaKt5hikUX7gR6nlm9ZbJvS/jVur+ZABWlkoaPqOWInK172vMNY+
X8BIgM0D6bfasgxj0qyAmXvE+dJKAqafzjcVJzJmAhEfGvJWXPTdBAeCvLzid2SIDHMwY8OloExQ
ZFQTSLadANJd4N+w2etzkUIdlDUN2HEKemNOxtz7M+wpAa6jwpOFhwx7HELaNKPnYIyGfgbGl/cm
NuFJyhKQJEqQE57RdHnbKzINwooVzek8HADEZMMCxTex2oU9MJ+5Dtdk5w81rT2p4Ms4pFG7HQI6
GkjOjP76He2zVkTn4vdYOAS71Qtlq/T6nMAdbae1QHPPS/+WKwNrdZ4Sv1FrczHIkVJLquBZuzpk
Cp4JNRZY+SfK1bEx3QXlrczg3rLeLfUm9adX8uD8a4HTaFnBA2EmNZE6IyZ5zgmY31UAfd9wM09q
mPCr9i34uRSTZREzen0eAXu0U0K1/75DU7KMXDb/7LMp2RiGuwkkr4pWvcjdgToWnF7Zo1lClxG3
CDEKI1hNgHdFXBVfJqEJs2HoBDI+d5pZoPI8wgLOnfb3rdX1Vb8DWxt2xk+vxI5gQxEJGfsQbPc3
uD8qSI+NntlylIXIy62n1fgTmOXNzcnGAWinqwuS9iJ0/z+z9gukwa3hcRvP8eaKYu/hqTPQvqLd
0JoR1K3Z6lH+90fX+JRUFt57F3jtVMzepANnNFlfJNtiH98zvVbqmDNURWM/fOsyQ1Ly3o/RDUzA
Np2BtYwi8Mryk3dUbJjwvScxAy8gwF7fOj66T5WRo+yN2d78/JdSYz5xdBq5DBHr+DBQcvEvRteI
EDaGC2jbO9DgVVCqkOLPoeK2N1wDYncXuKR+2ZQdvYovFb+30oRfVWGQhTAu0xfH3IC4hm9wqa7v
fuGUZxvo3466r0v5y17WRrHrhP+fIp8Z0nX42ljo/LhvSmwIyvkc2Z+OWoxpW4ThKV/hOQ/g6PgS
8OUv/655k8tMx+/mtctwt+d5RR27UDi829s5mQ4H7ApSVIKvKj7YzQvEXMAv5U9FjQAJPxSlFAQb
SCVUp6omMBye7WSnSOyrlwVEsbKXjQbviE8awHnR+jARrrBmmgmiokuDg0CGcN29MM2f23z/dVj6
G8Revh+Lue1jf7f10aEMls7w0uZjLclZeYKZuFU0EvKp5uTsvlbKuyGCr30MekU8aDkGGxt6reeA
/Rwk2M7qrW5mbxnsm3Yc5d8LwB/9w4thei+qxi8OLqS0l52dV64CJMcFQ+ZS4KLOn8NK8lqPpWwO
1Pk93S5/mogpUn9PRLx8fTAKrcHaKffKtHwyX8C3VJLNpN/dyFzyuSfWrpR5989WN4UIw9eohtry
MVTQEGs988t3eJ+RXYMtMuFi+dpNqYsQwaLV+wHR5FtekXJiXA3smNOEVDOp12hZ9wnSWD0HfNaP
+uG9cwNCBX4Dzo0Nd32s60jBtANQMRSmXbiX1k7tvaaCTl82v9lLidFiD9y1VHRAYr5r6SYVEeVJ
y795J3fO1qXKsTa2HLGe3yVIC9Xe2L5f91OHv25eZWdDKPCBkB6xIrczx/+qXtgyET1o3nilOBUx
SKuizOxsDuyUFXNoPIJ/7T/lA36cmSD9dRPRPUDFtYcUYVUkrxbCBWzy2gGvH9sv/MUvadUx5+Dy
trqYmw8F5/Rmfdc6GnnYIgP7VrDfCjJikkm1+7CVK/Tzz1p5NHxvEYIinwH5kEiQc5yOa+0nBMKl
JmwuieZe8zoTWyHEJnkUbc73UDQYVV/5Evur5bKlZpTG8RwLQ94AOU/kQr8ai2wfZM/IK0QueY+t
yBdUdQru+B4fJfu1XM8KnC7tWC3gfmVVqb0n0Qll7WiPJvsVhe1TAR1RLWMcDGtWsPtM5G36piiT
UWgttZbX5E/b+B56FJDYcDFBxasJrrmlLWrEyBDUSkqDorANa9o9kH+ng8KOvl+0UCk4lEl/jbuh
OUFDqAojEgDtSS97xtfVVggviT//OqYqPbme5rvr2yidJ7rbwQF7k95NDlpJqtQZ7Mz1I7Q88+g9
ozWVUlJmDV8AH1sq+VJuwb1wyP04yfBjgvTaLn26zWNP687dVOF5tCXLgHJRdeDaOx1C4cGqsxQV
ln4AELRFjEuY3aLBpSREz/2CCms3GIz7WUETb34Z658Td3++6XHzQRjtjpHBbPgxCH46vHNtRd9U
v3rJeTuTLhrl/lMmqxfNXw35VM9f6QiD5vay6AjOgvusSNTEmtZCOTvXgvbHxK7kRDBCGdj/eNCO
doueixQJdxASnPxFrEp0GFMgBDDEhZCRoFwcyEmRnXE0sDFxj/DFo3i3TnlmLW3d1PJk1zPQMZuh
aXCfsFQDF77LUaDMNkWyyg0eW8myXPfXIKI8WtGnENY9o7UieaGUsWffw4znecV+2lHbj3fNg8xB
RinUSexsLc+sv5FvT9KDIwnLAl0cS6Ir5CWsvDzuBnbDN2JXenmlpdYuSxrJRix3id7R4YY7xxQ6
fCGr73elQ0aYOEHTcQh1wBLTWB3P2LuYY7AjaRAtr7DRpJuCsQDvXbCe4IsLN7hyJXaKy/xbaZaF
ENHDuUbSWWlbgj6bnp0dZPTXD1KomzBf6lAOA/oqgSsQgItGN+2oU4WrJCUyi4UuzMDc3bp74Y+K
GVaKZs9ehP6EqvrVbbpeK3miQk9Nt+ufWj2Ss1Sl2tcgs4LbnMqwCc4UnXQPdGC+8rFEq3o4nbKX
m+UzHcT+yd0k/TDibWQHc5GQXx+aZjJmzvHz+EeCF71iYO7iVq4/RJ6hg907XIE6q5Ffv7z8JBqN
6iGbMF+87p8lqO5aBkJWUoReiuINt0SSMbs7jI1qKUIk0KRzoAgjb94VzJ+ADoy1K04rQcuHCl1V
plXLP0IxFJzd6Ra4Ykf0b7Qv3aZxkuEr+G+xJ5NdbTGCcdRgORVc8rfKiC8rl+TYMO8OmLcd5jhi
I39c+kL1oRw/EqvDpwO8v0Nz8OYcQyjxg3Qi6SHG1X+K25Gr9LpVbOIM6JGbkrOkOc4MYHkZ36NI
CwuZoAs0Woz4A2r/8PeLjaHM++mie5I7oxiFT0H2RQp58X5/sX2n/BhZ+yvExqtGvNv7r8ow0KVd
iij89JU/JAN6EztqvKZje8lsrX4JeuhmMuhdTuRcR7AmDs2V8vN7Roai/w88u22ELh1iuhwkjVha
QlDdSnCkrGdexDp7ickqLx+F3pL1Ijopw2jK1InfE0z16s8VwvOoRHHTzR7NcUNcxvxgOJX9zAx+
7oBYsioOcMSmvjRXKfsVyj+NSNohVvHif6XRNvJ6z8PtBZtwe03KUqpGP7cn86HgpOtgaXWndXB/
hT5T4642uAvf5M2H8CWVCr44Kv2Z20Uey/x0O17ij218hcyjG2M0zAxcf8OtDCpBi0UPpkfpbhls
c7XCCutaOkef9EBWCkp++xX5/2t2NpkCNi3hPJHd3SQC7Ut4T2Hu7KcogtcZXZpHT84LwhyNlWZM
To9uZQ7Q8oJiLPqnkb2/4GfjWx5dAjtA7eFeDVrHQw8NwwumnUaLz1uJzZXkLFpssfHgc66+KQw2
6BuZpP80TEV0i40npdEwnSMN45PlH2SlyR/1iM24+jWA+sfeYDSf82cQo1lGZBuV+lz4tzYon0CM
UPUGp6kbd1rGQBULl49JDFYmpyi4xLkeqSb5FfztxVwY/Wf3q5sY+fpSaokHkZ09inohq5Ltkmdg
J1YHC6T4N70MqTBFQvcO3AKpniLHEgDJItfxVE6vE3/MZA4Q5QPD+OB3Ozmq0n62Fc0xBxaG0G8E
KMOoxJ6Vg+xRWyQlWrgaazmApp0ens/lpErTrkzNy6WiN8n0bF4+y6c83SG5QnQD/wXjyG79+G0u
8NicNH5pRT+VaAUzrLmovMhMEhHpwRTCltk2dzsSuu5iXCHniBh6QHkDLphu3lvLuOG7noHI2Wg3
/Pp1lblBQLpS0Q0QeE7ndpcaSCU0mxU3k8OoMIyWp0cC1TXyVVrDBmFbZePgbIiiiiE+B21HvRMR
iIhGfd77tgy0zbJKi+rRie7I3EdR/Ercq+tc8YQlHG54Pize3Xy9dVtFhwwX/OfBatc0BVTn6Els
afprxdMga9+h9E2OI/LoTqrceV1+l9OG+hXD2WiqVa5C9pKnVE9QQ9Yljx+UM4w9srpZfkRXyJLH
ibG72oduYe3h8NaavkG/bStQbcLwTS03R0QHRJgEK4l645EccG9RcuNxwWvfZ6AC74blZfLhtVj/
tBNu4YHlMDJE0HFH4DOxV0iTMqrPdRkaeSkMLESHOBzD5l3hVhxHZWhpo+t9m6NS3eWKAYNCsvpr
5cWaiiMZxQYo+MKIU4b/HRunO9GkGd0X9Bn5exGMDOLw+q7Sbp6hTkg4fsXPy74v7BO0OgAHUQBG
QJRmg5T/ROGjPPbOKE90kwbzHD5sUsDN4gR/zOPoAv7rKxYeLTwhTPoVirr3oZiV3IhxFSp9vPuP
B8rFuyr5t27PWgRk8qvTj4hdBbA6zFejcTUoIBVuIiTYa6Zok8Yu6g1vFX2prfTMXwCSv6ATuwkg
3zlInPkpooL5YP0B4sTv9lxSuBVAGWohcVkfUH5toLWXofv3iuIi89FfjMshnRo11J1o27w5f6Gb
p9H4dpkS0ExBBfQ1mZ5d5NHuliqeJBcHNWNPypU7iEK/HLO5wbP6KkGNb9HaK5aaIqSKmW7kdXck
Bm6H7BdStr1+H/4nnxdtw3EQQzsM0qdklGRzlAvfgzK5zYWfidI9vjo0/VrqI678YSwuFSPGYrHz
JOo6DoD78XaBc73Bu3mU9Ty+6G2MfvbqF2EUxqb4AMIod6OFgaAJQalK9dUNBva3EhzmrlRBW5lM
xvueW4wXRZCgw6HtVT/adRLMeySMmK6eaZk2a5FnZK37UI/g6FUkcHDevATjOuXOB/xVCPcG1/eZ
QtjrNt+ojHWz33NxkKaWi6SawNJhLfCj4DxPwo93WZTvwvetsqqJWQBYP7nHLWbD5kWRIpVfairN
lNZKxwgtU/DbLeVPalHHDHOAMPLzUomcLND60cEtDZR5ihtMPIb8aEbQ4ID0n816BtTzW58gU4aj
mMSrbHLQc0Bpevj8m6q0wZNN05yA6AwJvZnHrUinNVH6JJc8O/obPjPbNMj96ewVTjpaBdiuwpXY
ZGr23r4r8aST3zGyHpF1fvJFHC8J8OCXL7+10V1jGE7WREXqHT4O0hUYS4ZAmZYBVzXUjoaejSbv
Tc5oqiwSCFMToS66Rj0cKrmgQt6Ifav8UvEWymKz0pc7QaVDlvDZPA/nxJVhLUXWwpdWONDPiyCK
A3vp4q+fqkwK131lh0SJaK2x7EC/jSebI84tBoosX8q6LfXutkC4BZS/GNZIznKsDdaQC0qIKwZk
7i/cCqzZZTzdbsNEvEmfr36Us3i76QXBD28TMrDFcEFYiw0JkN1U3BFI1+qui90oZUF4+x5WqLak
aL40Cl21csFf2pa0HtT/e5dUXS0w1OIK0vSOa2nGYpNHf7NO0pDY6XvKUeCdI/WVDilTVLSOKcJ8
/SnpL6VYF7Z1LXaJhgsk6WHXfi9ygOu1sqOTBfdd169mk8ve1LpmRHq7QKNDfJ8uUPO2xx0dTqc1
gnJvBHaAM2OsyTa8t61BLEWOFDokBiVyeYCMc0bFMKKsmCsb3fEsw1eUAi/LZbRNnA4/mFbO8e+a
ShXNxj7Es7C+I7UAcw/BVdNaSsKjcQFLVRn5NxLHo1ecnYhCrae/1XwT4DMB/kRl10y2e3xkpDen
DbavSlIOZAib5vaRzTXzvIcbBG2N+vyvyYUstMLilpD93sx4+yAZla6P6pG/UrqbugYAtwufLjKZ
5vAL2nXLzEJr6q5M+qOReIe6Xb2C/WfQnUyPruBGSvb8e/uOjmywrXSTpmKZKm/flGADU9+q58Rl
mcuokJ6mGNu8K2iZK551IeuOii+/S4OPFFbl1DwlBTFP/HwwKvOvy5hM1dMn8GhXAHcLFVAPPooc
8/i9uyftw4AMhomMJWU4AqXjlk+YCJajw5LkOFUjDVyebeKd39oOrg3zQq/hS8FVgrQm/5PG+tFe
RS6ZR4EksQkgpC9HR6OkgXYxBXAN3hhOZKlE2uL9aIVI4C6bt+GF0THHslUiIjBkj5sKwlCFGUiX
q85b1J9X/ubnKpqi4fZL+JwZuFORyB7SG2wuPzj9/GiwF6ThRB8Yq4y7IoxqrUJLrtYdFNJde9oD
Lp6acDyJZYX9KSqDlNU89hWJRA3TSc6Mc2eR1d05lupUcEY778HPpx0lpX+viJyO5yl0He0y/kXl
Of47ioe/VswdokeX1Hd7tWLCY5PNnfrsTfSE98SkJX4vX01vbmA2P+ZFuVr3Pb95fw9oBuAUJ4Eb
fD6rfCbnwkEiDWiXc4SMz8W1Q1lIhlE1FBBARjGlP2zoqnMqgrjoh9Pb+pKgNnBELHJOV4Njrz1P
FEHDdS9H1DpyOJzwvgUNNCWfcSS4s20xdNaOVRSk3lJbdy5W/ce0DHlk3KXKLhdOcnGC0osJUj4i
Td8Jitpefw43fzXZY1gZYdfsdPA09XJSEnzR5DbXgdQsGZ6PV8CfykMhSOwYpyLeGhN3NLLjVmP4
o/LDCHLXQM1+y5Lw+cz68X3rVXJDUZZEl4agC5MEIULAtlOWDtGW6Fe1kw5lPfxXB/71fGHp6tOU
uKh0Fnn0GpF5vH+PkNATFGMBbQ6kMeZqeant7ifbRVAHqBVL1Z8Os9S+qKaYhK+70hcsza2rnVvc
5QFpD+1flpQG7Gxdho51cQXcxmA6sP8vI3NHb/Hto6nUUTkmSpaDAXSJLCvDBohIEhRuH1ceZQvz
ArswGnBPk67+POL6pUejoGLpu9mmnLn1WWMZk9t4Saupq80lXALO0f1lTBqVHFptwQPxXONwqFms
8lpx4i/6ILgS0IPjRdmH+WLXRgfunzjL0eHWqZBx7Ro+WkZWi1w+c61uzwTn2FmcqwXyM6wPXA3V
yEgowF2gOEwEAgF9vKgyzXbmIdqSgFzugB5MuVDZQNlp0QwPoapDsdi/rhIsyVI8vHATFod400Xi
pwK2xgmWkFQaMTGu0MKcv3vZdZlLB9TJCWzYIHAodg57DM/G7xi04QYhpBLndKc/rQmNeJPXrgF1
IViWrF7116vKb5MgFKnm6+hYTvR+YN2vLB9/0X0mlWoDyG6ajLOLPdQjkjMhvwiFVzNULM/NPE6C
vgT9/ZdUngSw3vgbcTGyEIW5V17bSekT+ga0FcadJjf+okVjMPYc1VMn1XW53jpSQAYp3PobqVCq
38vI3HDNYowUyAy+Ih0Ny/X52F4ffkfWYloTB3ovYfZePAJjoWbh6YorP0vxH4ce9/Bj6t4RtG72
dZQckf4C3O4uSsmpNYH04iFC8rHFId/9X1+52AgkrF6g6Yo2tawt7z0CtIoaRz/Jit5TBBy1vHqM
PzrqmSszYspbmIAJuARlu5p4h/YGjQnddIR0v7nHPZBZi7+gbSnM/r8/dPXqjawMP9E2E14VeArr
UFC27tN3gktav846j1jkoszcjIJ/EL2IddX03Uw1nDxMOJv/JbBaBW+gR9UtjG4vGYGyMKNJrdHo
8RAXL1tEtMf2A3hMRkFucvT7Gr2o2C79iAnpGNjm0up3w4VXbQSx4Wo84yWC7ikMIJYJC37E4N+B
YK7NhS3n3ELENAwPqAntl90ZnYusPHRasM5SX5YwyhpOm/v/ig7JWI8Hgj6GQFuYqsG3d0+Z5TRQ
5VQCCZUKNPy0xlmW6ZWN71+LlKJ2XZra3Pupc/5vu0kde1ML3E/BVDvTq2QDrVEuzVQoL26stI0F
CCCU9sr8fxySHaKlJa8rDQQDHOCUD5S6XUqBXx0cgaiEB3rglt8BTIpWTx1aRDlV/wtWtVTRlLyg
cQhQo9IXyd6yC4Wo1XyMpDUysznySUV0SGyOcSifI9Q3MO01AoUKblOstiyfxZ2gCmkBNQ+sZOwe
q1XZXVPUp9628NBd7Etlr8uqkD7QUubrT3aPo9KKQ2+6CG+Bvv3n7bNYI8PI+cUEZvraASD/dD3M
KPAUxN4Eehc/BI4AZl8O5W2t73p9+CXrwF5/gt7CLk2XiDaMo0cNGihT3SlaNQ8NmDkm5Jk9kksc
0wWFPXR26wQ+/7X1+4afh30GRRmMAtMojls+ThvQ0j9yqqNjKEZoGdDqGSf9Ub3mmxeR1p5SyMYF
e2u0DMmZ2nHSjG0oSBFfE42Po70/EfMyBrRGEOiKQrOgkWr3gn44FUHthuaPx/p8mlf/IfNaDQJz
BXOndQWyvVBWR1IqgJQmI4IexBWa2NCOqeYKOJOtH16SloMEexPlp/1HzUmDauT6dsGAyAttBkZB
ZU5aW6upoRVGDOPGXuVVtjNz9KA+RoUYk0PyuloQa25Wi7HwsLPj4eIVTmf316sNQZJblYwj18jS
KCPMmn/JnIoxrVAsksMwy0I+IZLiar0zyZ/6PwWjPMTr+bX+OMiuLHJsUk6RKtJ6aSFP0oTk7yMd
YHRMCwGvyaFEjODMmOcXc6zgPBE1j8VevQuhnBYJ3UZluRMrW9xE23PrMKfra6+6usOZHs1a1fPs
3q3su9so1xu1/1E5V81QzScvLZtZcGsckwpUb9r9XK+OsCJYfXsSfKjrm27Hm9W99+XPzXtH2ZOG
slGpPg2UfCnMvq/JPRJdizYO5UfTh66JDaHJX+T7GcHehKWroF73Ai3gRAkPHQnRSmWbiLGodosM
GxMD6Oou7YYnH1ivGiUNtX+q5ZfrCzyk8iZRMJJVSuSH1/XYvUhGJxBT5KdKV/muwHVywgL8RURP
V1EQmk5X9BjslmwLDKkdox7Y7B1IVE9wYGridm9eN71e7eI23jNdaFcPtxBGiDuEwvFj8bFnKQqF
3ptSjdcRsDu+a9UH5f3sNqscAVZVlk4W4bqBbSqGEgl+gQBW1dqKIPHfvHyOALFfFVmusDEvAiyv
+FQbuak/A+8PUM/SVmnpFx9q5r8nZf5SLpKnsN5k/MOQqNoSUlhnpqvyAAshhF0xEcSq45trzpkb
tRaG2SGmFqHiA15vGkt8GgDRkGkqP1VVgsTuANDqwj5lxHx7UHdnKfuZj7BCbXP2lb4xRwL4ql8Y
mJtShVJlymjQEEvxVBDr2Zi/NnL9tzEHueRJwOPqXEjsQHusemVjRD9YccXdzS/X9ehRnaxNgh85
vilWm07nhs23Ao543WRUdqK5QjT7peSI148LaW3ivv6wkVIpKCOsE/Gx10sHFwq+i+p9J3yj8GZM
9b9aApbB2Yj/aiBOlon2ivGF19HDtu1X/krRYLsEEeYTv1aZpjtLAq7M5w2VGfP7QQ/aFhcB+qlt
rFJNAlgc+SczfJlYvK9YEQxUAvMXMnoC8+SjnfL7qx4pOoOmccEciOjOcicM560DCGe8iK9FvVgE
6bSVkkf8hC937cO0xTwS+6y6RhLtAd3yO7etRsGBnSvHkhv7L36nK3uKEAhg1tTbT1w/GyOnNM6v
7eMsC2JguDwUMCM0vJnYGn44aBQ2Gar+V56oQoeyrr5IQju5bhVjR1jt2a/6puHp7rFgdOj05VL6
4QzL+PZ9n1aG9srgug1RKufL4ubA0juwxETBQP67bGfA5kGAdBxZFFLWS4BtSw0BVatiPlNY+Q6c
m4JzWpsgKLNUC2AbcVfQly5VP4r5pfameC4veZMgVb6Dj/stxdrJRPws2Zn/+tbIHbV+CfBbT1jC
F1p+yrWlAFh4aeou2iNCqOfVmQlnoLECfnCQZAQ0XJbt29drMOEGBaO3sAskbYtPd2CApP2n2dbd
xvHOLFg+JcABfMshvoTPsCH2Cu9BtAxUkGM8iVG0uYCPxuEQ5O+Y4IFvlHjoxziruDvPEZrdPaSD
//4ln+oXU0BI01kI+5Ibo+kGKPcLc+24DJugy9mgfqgOhoTGkfVtkaQgmHft1T5oNaTAsICfGtWj
YU1kihfZR8hH2tQT/IIkFz1hMo58Q5HnD6RxW86NDkkmehVlcHQoGTE0TeegkY7GBaR17tGiIuGA
kMSPaawJhQDekjq3PzHFkNIHFvE7L28Ms/xQHDkMgFVoOkp3qggpfwjhiXSoIJaqZHeU1W0bPc3S
wMmnRp9Cd4ddNtANl/of9xmBP/97LPLMpCxnV7Hs2s0yMicza+xjqls+8CHzXOOP6sYGknTzr3Ii
gJCaFsKLrdnmj3/V3LHsJbmZrKxIXgBo7aClIJWRb6vHvjgSiHbsTBCK+kYlUtxeUx8TEOGUc8pv
EtgqldG1tvJNVXcqdIhti5SGlN/oLluczjrHauMlMqvZrZs4nfArx3bY3ehdhvAu1fjFKG9RVcE4
X+p7wSMR9ukIcoLEOQMA0xzcNTBeinG5AMPIAppMli1se2Z2NP4hU3qszLDqsR0zDVDlxeUcGCdk
b8dhFhRJTJT88Sv65uP2fhxODW7XBIkqRHLij62ANPIyDZ6iapbXA5zKxq9Mbq/8lINghIw/U92m
lontbilI/lwhF8mps354gjjQLj735UEi6odtrH2UA4RktCKGMlcdSBjF/22nVQ9BM80a70CB5wl5
SR08o34sOK+tmRYJPUFmnRQoja2tK6Pm5f8XKARpYGpy57XVejeKxwSvsBblxdsNQLIHklnhL/3z
S5MxWFResA+VRm1YwOw0JjIwNNeqCuX+OM6jBOmelVYSAgBWG157f+n/hhbCzOeCheCOltkCVqX2
wHFCpX4Nv4GNv5TdAeRVtZlsA2XdaQdkRTiP1+EI+49ITKhs43WXxYrHNQG42kRm5nwvWqBECdY+
nXw9xBLqGGIPefE7Hr9Nn5cCklqgLH5ZncVXzbre7DEJigQaTe016tN15ASmQMRcp58ncKAg3LKU
nTmCkWPqW26t282OxC5XVfbQuPIec2VJ2Mi/4RfjqVWW7Wc/uSiRLWUN2eZ5/RlrwYCCbdlEk5IF
ZG3z230rNGujgIWulIraE/gmnQqALWPwaNSQMfcmd+DNR89jElW3wRWha2FAHilZCYy9o1PpcwRM
yrDLLHL2JsAbe0F8CTKAojG4+S71pHbMwGQLjO2iCR2W64xZ1YT2DR0B1lrTNNme2xZ2NDZWiMUJ
iMV2tYfaaWGmrPjiDxAa90YhhBxI58XCwMoPyLd+rsB4rD/YMOABvgkhvYeCyHc6okDXuS3vWuDl
jmjdyElOvyIhOHjTSO9onKn/qVMBwcgHVLpFUi01PXtG0QSYvIPHpjGNNfPLJPQg9E3qDiZG/EC4
6tMo4IWHDEJIEAjaL6LRDU2swpQ+TNfnW9Q5XYRgiM/CAIYYwp8GW7EK9GPvJwyqGb2+O0lno/qk
GxYZCC0N0RDSFfaHh4KJmtbE4TlSNvo1NL5RmEk60GkAl9dZKbXtfRvMpqlshyER5KPOdwy0jRgz
I0ergVpL7oFx8Pj9zY8QpFFVL7HZmw+t233/FHX1EqLmO1Uu/Z51SeSHX+j4bvJ0sSjaruHVD0IJ
zvYfHXRVtPoq2lDmCbhFhikW603/r5uf6EkcW7Je4WuQZ0AWzUuz+bEREYkDkgJ5aXjOiMGlXBHL
dKq6kHcYcLCIApDHiVKHq2WoBqGxuHPH3D0VZeiRSmX8J0Jl0rOi6lpWuOcS0CN+P9jba69EGH0y
trBJX4Yz+Mt8R3JDzR8om/MoEnx49/EZIVkOpWHcd3CGvWjw65gT/vYd1JEcTsUONgCrPpFFux7v
Tp8s7MpaR1SsdyOCsxgYjOM6DrL4KNSgJveWDnAsKw6ErjW+Z7loqIq5S48V5ly72uJ/hJ+wVFWC
ffdC9ljo0XpX4WDHjz23KYG5Eqrkz3xsKt0RMEcffGrBA8WSp5e2QlZeGWVAFun8lmDka37kGi1l
hifu0N53uHCu/CPyS3Ct3SrgJpwAr9CDdj6dlUGjWrldgd0b7o912fFGobeupPXKLlhR6w/Gx76b
bjipCkK8ZK0HFRStBVETv+dftWUcICKlH4v3FaqnCE7ADWtNTPkogPiBm5XNHWFzVItIHuUu+7q4
kXk6e3crFXb2wcWfk6NFO9kl7zTS6JJxizZhuFkAZ0Zl+lPexg2/q+TnBlCthar5m49HMtGkRJqq
IA6XaqgAFzVibgAFgTiYeySLk7vGF1d6DhAshE9U+Y+lkamoC2gOaqeLbbSnRTTah1Ce+Cwj6L9e
FMgvdhP/IiQz+xPPh20uXAYzOCEZSA6m3zos/wDTvjjjMmUjjZEg0WiFTrxn/5PZY9OghK/Dkczw
krzWmXLpxB4gaAOq0HuEyXWl9jbLPV2nnleOMTO2W3xikmgpkodaayhTbGXBXNkPxJpRuKrhtWxg
lhB2YaR4Fjp8EQ6AcCU5cadyZQONuDDDC8KtHwM3XT2PXt5ldM1NMsECFhXbtTQOWX9ZQcnBVLrJ
D7tpFdeG14oVEjPSwbvjVcq6Zzgf7EYqE5USnGTJXqXB7PCvKU9TBIVwqUMwZD8dTVAD0HKZqWXl
SqGNsJlNMR0LHC6rG2RuhFNF0FTvq5FnEIaN4skpO6nvXL7r1qcvHsq78UktGCTlObjr9Yj9r2rz
y4vAT7axIPmPQxdQM015KSBq60yvVTjP9PpwecywEHSQj4bPwwLyHUmzW7MOx7TllQuvCO7eBQql
C8fDMZ33bR0hxjskfjwUQEEusHScgQY2xItEiqEYItkW1PShIZpYVpGtgTiDVn2YcngSIKSywaGg
TPbZTrSJ1QfDgw5kX5wO7hleS+EGdFTbFr3L8R8BzW+0U3prEX1ermDFn5Gweijy3v/+dCFfiSE8
3/1UA06u11kKCPozFM1JzjF5cLVD02Fr08NuluHnDvyMNhNgau1XXeQHmCuJzjDmY6P+b9cuVZl+
4wA1yEVQ9AXRbF6w3xntps1QbWP/H9y5tP8pZ5DNLndS4WR7ZPYY/yUfng3YQrbuDPgrUwvxBYox
kqXiNyx1ce4qiLvK6ey8bBcgjs1gqPsZA4oW1idAh/GBglhNijvbfgliGdGsP8O7/YB+6MQxsCeA
M2nWCg4BOTpMWjtGxTjzuPdJQUQE6l2QdQLxvJnEmrR0xMd9nVygJixFDHTEIf95MipcI+MgyToR
S3taq/kRa9l+ylSOkYDzp74fzxySfTZ+xXBtKEO3gEyl6KjzuNbZGE4OBkWv6ilibOuTbbEXHFGi
qo57KZPQo+w5NU2E2WzFwxWV+vnb/+Lw+L1FyPDPXG/HgiCIHZ98h7V+Qj18/pYtJRWoK0y68Msd
mWdkXmBSfeDNFHZoLi7LTAqY1SzCY5dmldX9xC0rxs4EH+HO7P/tnJsSVLBnNtFooXJkNPg8PI60
bX+8u5nNPYS3nZeKKZN++bFsfWnV7b7V5KTxivuZfCGbJW8Gy4O18OX5+3KWdwSUGkKhB5qtnNzm
rViua4bo4rRH9dXBoW2nF2OXcoXcSkSOzHwoaPBw5grh5pyQ9AqoB2Dh6tn7lSI/bb5nmk5RlTRC
lGg+eVZwYlKumly4d5X+SDYLWmpunFaoNC1t8p8BbqP77ttGTyeoubFrb7hWJWsLuIeCo2LFTYjm
MQm9x66B42nIti6ZWfW+R8e1aJ0yimDScul7H91/WbIv3riPSG9sIjikIuxIuD7e6b5TooEpGP6G
JfnJdqQhUsX5uZDct2+Cn4J4qNOvtVBgXz4sMftXpqTHzemjXr4C/2754esw6aUwzFTssMAITgRq
pb3TyXxl88S0bKjIRhaViH2ilLilOPyL8bmaLP5E0SeqM5zo1c3e63Kcp5M/8BSwaQ2ch6uuWVEp
jDx8aW46rhcGPUnmZdCP4O4v7wrUkj6YIxgnfbZ2h983edYWs5bp0HJf95eb+4JNF9PBJI1XD0lV
LqDY3BumldQBGMLUFRqwRGhgc1Hhjc67/iDnvEdRxKW1MqxMa5DUrY+zLq23/QEN91RXTPJyhVxy
7G+P8wWAzNj5xaH1Ns89SHwXxhOCXdwf3J9E3+o6z8Nl2b798rTFKbtOCQl0ob7Ws6pSiuOWaXFt
5CnGikM9UpKSBtsdJWQBXz5SMZzymx7MYBY2tscv2utsT+Sm0hI+YY8TEnmNcU/SJlNfJAWi0ZK1
ZuDglPCrehLd78EFQcPZe1y3YHJvEFRvyZfXEurkLotf/WP2KSo8QCYrLHY7CrQCumrDFOgnJCoz
ncNfAd6i/9F5MmR7bMWsMibm5gFvjBVSRu2FYwFSMgK22F3M6Y0uAaqqVtC/nAHGGMuZDCj/Pyps
+vfcfXhwKoSUHsucM+er3CnNFkZk4kV44CoN2NYvUMsErPuTUWHEz6rCzEY0rtz6nJBgVE7G0qxS
5ZKjH/fBlKi3Y22wp0WObfHMNqjP3Y5V5Uu36VI0J4IafFE26cEq3OLNlyKjOb6RPFqufyw+kcl+
1OfFkbdAxrEHcuDtjJf5xJPI8XCwT3yRVRelBQRKlyiGYK+OYMBw82dGwjcRbEdaw5485SVBKS8v
1gMGEe8a30VzX3QmtoTAIO1EOYKxVsxSiNQFvUclYHpJQhgLEaz+XTc7xOKKsTIGNmDGaVSJPbyt
RbtDtEhmWokQkAyQBidfUtWma+m5J3uIjjzG24oxwWy5HRQtGnfJ7RSyqHqSsKQCblyFOEfOvX4H
Cd615+Rbq+9IRSdDABpHzWY5jwncFu1aDwW7wq6GDZ4GUFMiDV2GJ1s1PYW8K524lSgXI0a9vUlG
M8qPioKZ0es6Eff2El8XH1yBaWpLu65408SFkoFpF4tOkfNdgtmKnyMyG8XNLuaV4aB7EK1CmRD9
+FURul9nBX7bw8l1o3yuYLBDzn0CapaQQhB/jxq0eR+g20RIm43XooOfUJFgqQBItkFbbMxK1UKf
MhYRfZ+Iheel1ZViV3IULoKnxFBppoe6E5bo7MbSURNp+zd3Qc+Zs1EMmuV0vwlXJfkeAUnNZgwm
IeXnBYvBBaceF+gq1+xEl0j8SXLJO+FvOs2cAHDbS4CGMZaIp1lRItLDHf2xfX0MRECZx5ZjAxdU
FJMB9nGEw8KicrGgT2sRY+YBK6uWiVtpk8eqiVzMpz2m7gBYu7aLh4owQQROqn/ophScoj0YJYcL
a/QVPeqmLHQp4kmBQq+YmHKB5qfHOilRh03JgsO7JFTQd5Y8uRvyRt6ARSH2mbdqlpUhnauz8uDX
9XLxoIax2ovENy69pvt+vYI59eNI5oPlLdege8AvSREXfIkXXRrfmTvHClBFAfO2GF6bYJqhU+w1
uY17JeoEkVcqocF/Oem/skXk1S+NhxD1iK8ToLsjYMOnCd7sg+n5FcIgxO2Zh5M+8Mjn+zsDLh2D
e2FuK+ZnzBRFvj29vzS8/gDuT6CUXQANI2tlaSgcZL97oWZO4vOtEdZV0hjg+A421hqgq5KO/IvL
zBs8CCuMuuC+nE2lCPrFD7u/w8gUjRNLung6luhEC3MB+ir56qs0AxoyUCIPfuwmMl+TnxpMyngb
yy/Fmwe5Q/buQJXZyP6D12CHYFJQCpj1SG67VWpiskhlnJ0hGiZ+HRbA8Sm/hPSi3LYHP6yTNuYZ
LrjKt3BIh6IP6i7OsBPHs6QQXCpCerb4p8QGxfXzjpLTyki1E1x9GnYlQQdTZoR9snOd3Gz4Za77
RysPFC0UsBbYPKJbWvjEl/IGlRa7lVViq2GnOODUdZWdr6E+c/jb8RiG8UQ3A2AXZm1ONJ1kZgqT
Ebb7rIIQ5pL6CMcHOjpB/zoiwe1gRaQ2BZ34FcyLxDbJqJxgNE+HaEu59ChDfk+Il/hss3P/NSdA
LTyTNfks1fGVQVBvE6CqHSpTCRx6EVolgKgeulwI/sh3Tc5HBqnn5XbMPyWr26WL32YABCw9c4Zs
FoswbZ2S1ueKFhO9xQdzBFTq522lMFxIDZARIgwSJSG5gm2Ufy3E8/9dscw4JvTEY2IgxhNVP5zU
F4/xZb9VscfG+jd1EoSvVwxqOHJ3rJDS1MRSyEDA+bmwLHZ6RFi64d/GHJ2L7uelOXUn84/c0g5K
kdeLy7RTnZ2aS8MDNb1asX1y57OQ5/R8hE2n8z/4yctAZFBKKrLiMeMTKO3UqKgj3D2+Rkk1ckPx
HYguo52pP7mbjdsql9g1MEcnbyVOTVsQ5etpThDw8c0YTMR6iQ7sEm4kAS8rijAIXFXgI6b+AeZx
xHVnHsYfdKTZUxcm1cu+lUYNV7Qb8mqNxtiNxUTW1NVUUv0EwOMVUfMGNmRDv2FF/0EYWJxqzLf7
h9OhT+nAjHHtUurSXqPEx+pk1OrzUWoWIWFP29I4XCZDUcr0WAnvRgZKut6ASbBTlzXhd5/f2VCx
rxGpoNS633crdWIqfpkyp1fgx3sJsCVqFXLpLbRXMc9F6wPk5EFOQ9avdqKO4aXIcbXsZnGQxfP/
LqdjIHEoMfnhOGiNjWGm4Xd9LS3vYq37zEub+vlQA8Q8hylR3qUei29Mt/v47rD3m3Tqt1Qi2nt8
mdEjErwgwPNdxOwaij/0/Qq1/tePZPVNrihSnrQ6iWQs2HOeIu7k6muk9cpROCatJWoJYV3Ao/y/
0bS4EIjnidhhrmKjHLZdf8tq5myL5OuRPKnsGdRVY0Ae3cb8KvYUxrZL2Ro1jGqGu7y8mKinXFxW
p4Iia6E4LqSItj/gvxVeGXCrluMRJexXcm5lb+DMhb2hDrJ7dTRYS/wPn0yywIM2LtUuLWPxhMyl
gKeaOgHQP4b48ptAmZeLV4Yw39CJ/nX0mKHwBMqFKaiwQ1bUrqXlW3Oh6wmDNxo2yDu+je6CxL7b
/lkfDD7HOG1jCgFE6BWLC5ihTM8Nvx3lQogVN7stKv9yP0isMGmBaPKtNd7p4/mdNzEcM8gr4dWQ
45JtjIMgo3EdvVMxWRLYwrvFZ4VdeFNsGXKPshNKQGRS/HoTNTBfXWCg6qyIDznOut/47HTA3MUr
FXFl2OaPkw+rM1ipSfa2RGYwvSw6Xq9QMDeuYZXkQB1GoTvZ5pmFMJV7hNmW1cKXSSkz1rNfVkoU
TIcEZNmOjMyXwSHzM7K7C6QcyMQDIRb0KNCfdaAeSZwttkvsM7s5NE2rNZXN7VWd/7rhrKp+7jK8
7P/cnNC1HLuvQDVZqgcLYXlGI5I56+roHxyMzn1R3ISzK37tFIS72ECaId265/9g//Z1K3/YVHtq
Efb9X1epkShH5770AvLw846NERSG7Bk64/YKL3cp7D6v9Tv0x06vuiTXcbGMiEK77ZqmO4tlGwDd
+Va4KoNDDfUEF82n7O+8+kNgKEG8J7dxT8NrGn/td6dlgD8fLKtMxjSKn0t4D9sZKUSuvPWS1+4S
X/PinYASheyYjiKZpLzUx/E9uyn6T9gkjDY7jWxUBjDHlGssKnc6NvRalCsUQnWQ54j4DGGjVzpF
XtawCirnnusqMhd0DTfBi5VYiBSF4WNYiaLvSZVPuLfY9/5vF/XSJ2SKiKz+BoQfC3C8ely/ClrE
fUvAmvALxV+iJBOJGiKKmO7ZkJNBHpepFoFp6LlNUC+Qn6bLcqt9YdLO8ukO2ySOHechfTOFvgLO
WFPtSA3kPN1svPsG9hajZXEGhktoHoF6va2aKDBbWzE7ow2Gu+In5qfwi06WWfYuqg+4Oecd+nPW
rozhgkwY+MBCkLeiA40gky9qhxERtwAovRVKgU0OOU5TaAfXLDcDzB98bXpZ94h3FFnTfRHq/9Eg
1FR5J2z2K8afQtbBCs0VnmjIGmgs/hohGp8WMK7UKvhfWwfdFEOIJMiCN2mQm35EA4X+yPDjbAX3
4m6CX1x1HoTavvALQpDrkLB+w+cE4uo7XytNumyEnx7QftytWngGBcUD2c0xpVAjZdGZMjBDUBD2
u+xHFYPH6Gbd7h7lTjHoji6S1LcchLWRFg8+gSqHe8TwO5Tu9nljxO/BWU74f0hI9o1i8pwAGFPj
c2TVYRX8+Nyk3SfB1/8s7oobMA1PvwkqlbNvyvmnbx08+0JABmR3A+7CZjuqFs0ne4eMtOO+l+QC
9Z2Zs6T8hYzpcKtPzZk6XjquweGKoIpmOIvjjwGDrP8TxUU6E1vQ1h27SyGh9fLC3/eLhL9mHXLa
7kaLFB5H1agVKsDN1aJ+yewollzoKOzHXWuDo0cyCKr3FIGKn1f2IO4LAxKdqSlLJdbjCPKmxUOA
x3DcVrVBaLFQSIqdUlDFtqQ1fbhIyJ3O6i+ZEnoa6H/xt/pVSlLyog22ccylto+nZXg1q0GnFd2k
2WXFFdN6U5ARfBURtwlibwFz3E84qmcRWy/F/8MJnweaf723ktiJPfHlXWyBeLqHxIdYLFMEXGk0
dT5dNrcYLq/VYZTn81kbcRbNR2z16nk+S4i01JHGl3JvTdUv/O90kwXTyP3xpkg3uK2SceY4cSmR
z/vMgQKi+Ta/s6uz7DInF30F919fHBh2jSa28qYxytuGu/Ia3BI+Wn/zxgxNAx3nxP0Otof0VYu1
R51LZSiU1mgFxSAXpNI4KCmJc3ojKDq2T2opKQAB6Lm7k5NrrgcEhW4GIoEWXMSScGuc378iq+Ca
pl+66vRYHR4Lratn6MupFhgAHzu3KvVmUjbGNkVWN2nr1O9KSAn4E1NS8wSdFz3dz3vraJhbJ3D8
YhplDqvmFrq6K6svHRmvPeWTti8AxK+ZRA0Wk1NNkmXRRU/x4IbCIugh3KqueI3GZPvui/qsfZy5
pMxA9yfifi46VE4ODlUEse6pIx1pv12+DD29vNP+IJmg40nElClWcWOoV1l9Qgpn3cDS2U7hKUST
8qNflpR7KFwEOI48xE7KGiMPcOtuC64hY3iRwwUr6izJmLHLvk9INdfDzxTv99nMI8V9O2wEsY9T
v0DuOvmGp5H1DC/LkoyPdORCUFKM/VWXQy/7XW2QVv+45J10wxDUT9GP922qSnCyd85RuUsGWVPc
a6GWrX27dEpbq6kIqjYNelONqR1ykzPlQAjIbQq08kM8+b0GhXQUB76LXQeDmAO45MgZTGgaw48E
JPCmc5gOtOWAOJzl1Pi9jPD3ObB2PRGXxVmLGB3GEuIQG3ymuBwBH0LYZpxHwZqdK925vfHiLWJf
6POxDHrsYBSuVwbAqURn3zyz+NHig87OTG1idh8EOSxyU38Zgcic2jAwMwX3shOUuM+CJFWStwP3
QuhM1dV59eGqe7Vm/mC0HCy2uobMz+FGlEXcvWlkllta1RZRlchjsEeAKOthoX/SrbpCopFPHI1A
Uk/Dtkb0c+HzFCAZ2JMDqZoZLGK4VcvCYADTJiUgQc3HuXwX/3/uETHKcd1H/mxt8T41WlAJjaiH
EkNJNla10CmlKuwqUQZK0sM6+n/HC86bYsh4oaHqxnNHbEMShd5AO75De4+b2Y7BDQ0UE5eXpK2/
qSWcVGG8Um0w2Xj6SN8DlegMaoVe48iaphmWNidzf11C/zs7ABcRfnBfSe2OaP4sDzkeR1eJU9Xe
D57SAAIu3RNcwEJwOL/xCW0Ce34TUB7DAxJg9FX1LMmsKBqq/GzllLQS+Ljst2h3KB+PpxPOa2B2
H4SQLBFceg/T9jPwe+zco3ENtKFZrSkEbsN3yzDHfNTyhIlVcZ5YDwlT56kutoQtt0wlF8uappWA
xAmDgmgn3+3YHUwmYfCalKIEKR2ER8ndbxlCu3Qu3bLI3KsPTMqwpKY7EGp4Xq7X5HE798tnHwwF
QO7tJHKKvEWn75EzobHgfGcmyWP1QlLZg96/GfQn5EBEcETwqjru5u9Lz0xFnRsrpv8UN5zAULPt
W9KLTKoeFiA2FrohgR9C4rKDUJzutcVN9nooeE/qwbtPx1JvM3Dt8dhuTYbS1ucmyUX/qYTyoVhc
OmvqivcGvVTLTZsohwS1g2BeSYKBK7pklIutAvnyUuD6Az0icj2AGkb8NZ/tjqER1bwwhcUsNTDC
VSMBQ+s9zOiXhgL9aHtXbPgHe07nnicQeHwrsyjpgO1P2aO7Y95T/HA3ZaQz97l1t3fM3VcG7qzN
Xxed5U7mtU76YykPq1cEmhRG3MUPUIdcrR+DHc9np3kRFL+oTzLQxLD6HvabX41QxnbFo20SJJ2b
UbrSaE1oBiBw/XpAqG3mocr0eUjNUsJEHiFJj7yxrfDXJUF0hRxSxSCVTSLE+SiXA5rsFHEGt+Ov
zIaoZ8LPw0/CWa/rjW9fvAFH6k/s5PXJzncxgdRtE8bwpUnDIbYbiYdt7oGa+pIlcChkau99z61Z
DomnmZIG8nGV3UKMuqoj2ZPjmWPb5iP/0skNZBH9u3C88qs7HwWSlFnVKKykU/edhAtjU0uSaheQ
qxBbmLdBhzW9ZVD9+gePOKwewktfYAZyCRzG7RjQz0SGB3dZ6Javuot5ALFq3UaGye4Zw7ip2Tf0
cerx15XWwKqlxkq/sKzaRErjJq3mMCIYDXvsxGrWfaMlkjY6+qA35b2fhJTtDfDHzowTsi7IYXhJ
dOfSJ9CAxhL3+OWGcgBdyY6rcaC9Se+NkuCLtrOR7KKrLEAfuyCFwzuYLs1VqMduz3D1I7X4QSVB
i+D0lwkvl9nXEtcwomPMIaVkhIm/KBOCAhYBZ9G4TqB74dH6p6XhhE14xZ4BWIYJ9sq2Fvv0LdAl
aSsMkAPZ/+fp/QB0UwOyRAP+VET/DEo0zGjzcJRJbX5iR1ks4MLvYlnbJ3RpaFzU1CHyVqyt1CgR
fhu6cTc0p94FNTp0vKpRBcizGGVVWPfwjU5ekNijIuyeH/ExlrV+XcuxVUPYSFJPmcsljNIVhFDg
aTPGObyZ7d1Rbx9rz8IN26ohbRlvoXeZKIt5f6JRFhr2A/7RVnwE/Pa3xyViUFskEBbDOK4BfOp0
7U75xkh8WEEuJcUsWqb/42uTBApF9uIUiGtrTcwjOPwgWYRhvcUFfvPMRwTwt4G6NL0MgXn3wMoT
Z6MAwxNLZw2VIuBxgupQZ8Xo53m05qryEWTt2my/opFxIZDcGssvner+tsosImd9fc0uHYec9HoT
aosNBJOcIuiljA0REzhW+npxT7nN5fm/lPAOXST89IMu/bBOpvahVHTEycdAUuhcoXXsC1P05wmL
yADrvfHilqWZTOe7Gq5md9tMqIkyTsPcTYuoxapTK8bvw91z1W5aLjP0PSrxWNcQBrDx0JTr3omG
xetUQwuMXUBULzV9oUZixD4BOwp0/YtorDOXciWZZSWmAEbLqaINfeKiJbnaag2yvIoMKkKSy09X
++DOcqyotPeFVF1EWEq0TA3RtCxnKkHOJHuIu0OI1HfUI8bsMVE0KVVfbCU71ijaigmMYllYSNJz
nuUdYPg4ERI3BIzeY9envpKU/io9UthDEktCLZXDPAuX2cS7Iu3jHSA2etClMJ5NG+rRzoGcwGQW
uOp4Q5FKU1/e6UqpbNohqQGvywpDwcH1OOJcNJMfAtleSx++EIYjIY89VcP64f2M0xpmJ0gj9B7w
rc7542cA1vph5xxHS4T4XQEazmBXB1lIBjH5h47Git6LgXFtVHkraZCTVU0QS943etCaNAnmVDEo
K5FM1cS5dnQaroFq/mgX0ALJF0dZCYOGbohogExCWYdWxkIPd1aR0UJcAvl3Yzi1Dyu1Bp8vCN7r
+TMDYOa7BQV0UwLwQ8UrSLku/oOzHkHegzt8h3GdzAf8EDCsVF5YNn5mKmFERQ7+Bhgj39FVJSDX
/rtLmCShxPeZDTMbCSMw+Xnw4mrferxQF/pZ/ZWLLHD0/qWm44xE6bfM6DIll1KFCYzlwzjPI4td
fui5J+iVrOiz+xKpqwawtTwOgyUj6xcPhH+bBPsSbd7+ckcQgAYfD5lppThw1xFgx0+JI9szr5EP
i1ykmZFYljxVDd/XgNzEoo/MNZHkCwAV7CkDRH/9qY0BBAqjEYrUGze8zZnPWb5uzXJMP1pDRxkP
ayso+/5Lwm/eD6gmeHje5eu4Wc2yQ3OPCeKf8/xMilkqb9lPwKUI+X2yG+66fxk4FPFo3x40s1BV
qYRWkutitwkBTZ42V4+Jow3BYnPt6ctfEeDGkuUoVpKero+UnJ69imQNU07i8Rv3uGHGj6Ag2SR5
Tn/nBxnu+C6nlo5wHofAgQKme82UBToXSbBkBdmrbMa7+s/VclS+Qo/yiYab2CdECLm+akGhX3z6
ohWolycNVYooYyLjLjd1o1hjGuR0hkAuLkDBuqJc0znmAhD6GSIGHeFz5YI+eoOVwrEz2dXFrkHN
SxVIPd8HmLuYHKPS6T6CTbLbEuiCd74NWRKdaatsl5EvzR/voVmZiHRZRYbcEXBhMIsGfqdN+WWo
Db2q65iplzlU2S+HlZQZqi3st45idWwWGHZV2wcf/EgssrpN2ednKigD5ob4hd4NPgTIoaXSKaX7
+rHPNNaeoIT91P7strxp5r0rjLFAOh4TSHhDqB5bhdNZZrO4fSN5+pqnCYEN/kaB/G74/541racp
grnd2TYO50TDY8U8yBbq5b5UwiQsOz3dSqV9TEvSd8Eyv6I/HCQ+pewvFbAJSMhn/Eb0Roo/DHoh
SKAycLaZI5km/8IIeaKIlZmgo0S/VNS2BD1tcMxgRxmZudCO6y/fS5LMzCdDd7I8BqBJvj7UnDKU
waEnMo7esY2DOniKLzPnZ6OZI9cPBp0sfYLWf6nO2dhHdzG7qUdnYf1kzdGCojaLL0Y8PLvB1WQ7
gGKseJr01Y2+u7HlMVY2M8TMov38VFChi8Zr0Al5eRCRn0HBuxa9waPi6+8Pge9gQr09FfspWAeC
Ii1DGjiin6EaVgoWMM6l+KuYaov+a2BRatenP4c932xPdBA8dcGkg3wxTCQsXv15M5E2uqyyEVjk
2M/hqrV0YtrQ7+NbLbN+Do3nYHfXJDBhFUj4QNGyAj4l3mRlbblxfgVy63/EJcsTEgkiNQrD9gDw
YZJkRt0AUOp2fBWUsao7BjNE9beuUrGzBQ7LOZX/VGLFlcWyDICQS0iGzk+ZIISg4TpeUGA3oJaB
wRlbvG8dXLGs8FI7DllHmyr+Z7wocWDGIsWurl9Tr4tLFtNnxFG1Tybcr5xDtYpbY7j6/7xl4ldm
8Tjz9A1yW97jyyUC9XvvvnZ83nTm474wUJ4OIU/ykAI630aJwLCNEbI/32xsgyoqJs9hPG72PquJ
LWSLrk2y3AJIKnFEBTNVWB9t65E8/xcbENe0ziPEePT0LZb/SBlKhamBOV9Tn49GWVgyBA4jZifU
LMiu4mdWhQMIhFSS85lE6koXc0DdyTQeEthFybC32W8Nexct4HPi5QpJfk5K013+GzFZzdVmUAnT
EX3BKcx8WyxMofhqIuu7yGuSUSssqx2xmXyxjeSaVBaW+emjkz3TWbba0qQ2SYVP1DyzfPw4YKMi
vjFVpURbKscz6WQNNeflwrLVp067es9EcAH1p2ra8lKt+zTHcZfEP/hLp2LJSE7TeE9DbTQWV2mC
dfMAPHGF8FMI97zOvu2Edp3r6ZFVVaRsYjVGmy0eo7R26/Nh5ld8UgEvFd9YaTuYvgwzrQffqMRA
U17TsqBSNL192HOoIUTjUz3trV7RXf0X8A4iMWg25uLEXATWX/LH19SgKyIZmseEymt3VFRI1wcz
ruu4xnk5u3XaKvZTegU3WSW75ucqvhL8GaVxqCVrqEwSAmjhW3M415c+mHJKPHEXxVmbsHoX0gFB
BPWIcYM+SJ8krxnpvD3yTOY6RM2MdtjFH/cH+yQlkxXV3A4f/MDfkEt3HP5hOhafEpdzDDOTuT7C
dy9C7o7W6SyG8Tj50wyV3XvDLHNWOWuEE+NEha1bkhjVMd4+0u59b6EyHHVVUW42q2/wvjCv9SJW
K/NH7dscGlkR8pUt3Y4DOrusC6glVIRYrWdGetbZolBEFFQOs+hy0ZO5jkiggrQdxAvJBLVW+Axv
C8CCy6bvCXY6lUjC7y3eoW805dNKkL7+22hWRllDGu1IGr1u+hlspz30Zr37Nuo/pWi/uCFQSSjU
a6qLgD2nmh5Vd2oHbJp4l1cWnZrppe3zdG7w1SVecOJ0n3pq1enwyO+kks84BfJ86nKQG6aJMPju
ttGW7aRujt3QHtmQSiSQGUlfSdwK+eNdx0ICjiySZ2mJrOQxb1Mdc+spy6bUemocK2/S3GXQelkG
ksWFVgSL2hDOJizo7cjEyO17PEJ+PtA0BgxRagcidXFZgY7CFBKWDq8mt0God6O6vCKR0NP1vVsd
SBr6+1E7u0IuvfFeJheWDa9kTFReVMX34VHupacydq6auwIS/qD3xuKmmCpsExEazY2xDscpTTum
G1cMn6pikpBNEbcG5M/QZ7m4MQG6bMXkMStXT/J/iWBJ5CYIiS1jQarDekCqGAnL4g0DaJ7DlYQu
hYcyEaCR+Jh+6T+AhKsz7F/fOt9OO4Th8y/3wcUob4zYnsPJDnXHNl3Cus9Oj+s9T0i0d8zUsjVl
8PPCWcuv1GNzxoVbJqf1msndO8EPAXFR52N2N72oU/SmKvQnQTJF+qCBOPtdj411Vgjj66gWrWDu
OAcz2BIcYiqANS4HdrdY+n0DyarETJZjI7AoG2Wo7W3QQzxxUQXkjAIwVbUR/kiUNi28b5+cTpZH
1P/3hiep5btW8H3SQNlQ7BzyjVBC6ryvgPVDjXR/n4Q4mkdLY/HzBT9B6MdVRI356gnqakq7zk76
ZYQdwml4vz5vUv7hPvNrL1vAv/fm41jiE9Ag722WtlC4MxvpOykks+usMieESzifA7aM/u6JOBhn
UHJKr2tod7Tv+EjlnyDB9d/KDq6QZ9yw3FDzXJ/xUOzvRRjz0xd3hlpGFYzBDxOCJjKI2XTti6ca
nxmpkq6FMtJ/TYunIUW8arOv/r5MUbx6C1tF7qdpUV6ugkLMtoV7+JHSsUAJ7x2/cuxavPTesrAO
cKzeu5w7cbfHXImEjESxtRqqD8w3eoyZ5J8Oe+w2hLn7BqsaDcINxpvcl9Bl1Hnhb+i8zhAIoC4e
+0J4k5mtLsBgLJFwrpNyy/jHwHn3SOy6YFv1DkYul03PkCYZDjyILB5arIp7rwsw46k1mXDZTkT/
F2H4WT7q21Ss4Onu0V0QBjkgYDv6TL5FLeqZq3AYj7tSDKDLLoD2qBHng6/RAS2IoP4ylQhRbTNs
f7M5idgcYRJMXDhAo9R6p5qShrxyHk/eu1Xa53RvaqRoPe6ejY/1UYQbJou8jM3tThGP6uPi7RhB
XpoNlRhyOe+Spz9NlkLlCeNCKXEYib9LIQWcjVjOLK1Ad7xCsMTL1HJ66Lxv4hIctE9NuqHqNlQc
1N9DuWMDNAuyX1bcRO8wULUZt0NfUbh0fNd8D2928GcBefk/3tHLKaj/4q00OAe0RWjybCL6KfxV
SGKnVx/VP0wxTvMdEQuSddtS0IVF6DxYF62kz34S2fCvYx+Wg6yYQ7u7zcrnSJe0RtgqZewenrjB
ucltGDGilyExuk+TDO6awlEHb5cOQKOfHyMcPk8U+qKhvko1NUqgtaxZF6LS+kq9UpDA/gr0iTuS
8zMYPn77Kr6Wq8azaitn9yNWytOxZlf+SzO3HIz3EDn/6hGLoVzEsMBhzpNyGLWKYu0fDooeaZUX
pF6IQSVzdoO8TBaAFzqJ9Cg5KdXlt+XWaK6Ke435W+aVUzh3f4IA0LrTzlL4RtKLKKrO+5NeOxro
p+0UYQztmXl84rL2Y8SV0+QAIqBxtY33nvgtpjUThFG/0gdYzzVtYD6lPUKJmoFXJ1kldLHdfGOf
jAwPytoojmLKk3lgsWXvAPoxFOlZSWPtnxaqnfIju1DDyhsCQudQ40zfWgj5fRi2YahisNMoqTax
DFr5bEUW+E46xr2/COtAwpgXR7whB9gVCzIQgNztJEZ8TcAOiSJx+GFllvh7ZtKy0DJ1LbsFr8uo
GNmmvSkdZGwH5vj0Wn0PDSW8Oyob91alhGA8TTcdInBcnFdiGMCAOnMcfI4jz1JJ/F8rMbtTOCao
X5ZjURgePSEukYhDjfqgVXlUy1Bk4mdJKQhWRvJAh1GSsE6hM6Mk94TW1Y97oLVRDeYXL/TrNnph
wl2Oeq5SAqh23jWopjZH6sKjAtCS0PeWazEchFcMUyA/VuzzZiMXxqpAt6f0CjNjlLzAhjOs8FbT
OEPPQ3//XH/Hvof1U1F5hzQgvKgNeyYsDIDtBGOM8yzokZcHrdmSQkWQhDLm3vEj8ha/0Wyh/naS
ERpwX6VWM5p052TF7JnxM5mQiaBHsqS+LYsESC0shqakgzyl5YePhGR5vydEm3HPX4EN/lWS/t1C
yYmrYemqzpgEz0+eyE92fX2Tou18Sjjfvk3CUFhiwJMAcjBJS+6XUQf3osfJSaz+UdBnO3h4Nneu
tUFDUjKWiuq15esLfDoZJTEgtR6JG+QYJkBdgT0D4SHRlFNGHA2lsIYeiHPGd7IgMT71LEM6E55F
lH9+11pFwjw8y6nmwicFp4l6GN87cM1GW25oid2kuRpimROwIH59RsikcguY+FD5rPljjTStYU1i
HM4HdpF1ZaWmhjoxPkV4ensH76lBTuPmGObJXMVvFNPcCgSwH1FpLg1Oe/lztFEgcFZFLcOaVrKN
pddq2rgv3DgXSRjkMplDqVJw/LoZqaktdrYq/Ngt2s35kAjUNk10pjUZ+u5joQHBAPJkmttijB4T
TTOhkvzN2l3e16OPCxlF3H4g1mtia9W+1FslN9ddHGcbe4SS25iTW0ClPpNeQPKKITyk29AKvu8a
a3KSCsff7+uHTRLZnBNqGSYTrJvUMSL+QJIhDg9sEf5ifgFVhldPfKxeoaV3/1nDzWDRXwTvGBmE
PZwudqBC2sTZCSKysR0G01nN8lu6FWCWK118ad5/tupbseeGHS/0Qb2jWLw1zZ0R+qx/mbNKwp0g
Nh6Ud3QaiIVYyzTQ+e3XFGy7PozWv/oYw51Hboq22CJeWb6eutmO81xCpyAcIWC7kq/pSKEbito7
8hhPOpdQ1j2cYduaZ+nCY6wJneCJFvUj3sWaXiqca1j7MLjbE0uSPYxkFSv7M6eKib/m4tvfQ3QL
YMKC+K8R+Wb97sSWMuvgU+xfYNP/P5nvUAh1iAk2TXlU7tkJAk6FDFAnFIQbQQ3sEQGsiAF/UwIi
eC3mIX1uEkbx+xndXXy2SZDTkJT3sUBf129y6jezuMDY3FEnfJZJCN+3+BUI24uiqchcxeHb9uEu
E2Eob/13cAs7Pf054hmCuNSLdSW98amjoL85CchN/wNMO4pDH5kzJ3JOSpgPRXp7WJZo3VH7wcLw
9HumUcKSMQqF/BVWMznXf/S2tN+1bMfl7GRkyj6gdg4cU2QlT+FvdPUloXqSGniq7nJenCe+WDEz
PI5z08/nEcH3LV6dNsagxx83ZObSpBrWajd8HmSBPKTu9fCmlJjOn6zdR9AiXs9F2c4PMpAq1xoZ
pm/SarCWeL4v6XG5LpudHvQQRYbuhvvz0yHKU8eQyisuLfrjP7SznK2B+9DeyVGKnnDedLhLzox+
CUKxfN7V8lJXP+EN2FD5onHl5I5VHdykh+hp6iEpv/y2Ad+hi6DeGBnHkvwrBM4aybAjgGCNZ42g
c320uXS9/qdonMshEGFiwZXSrpqsgJZn4K0Ktjw5CoI9VH0lo2soOhHShiGremmPZ2yCDiuZT4Ve
FT2r9W7iqY8myQG05o+gR3Ek61doDv5PhPsYq1xFLenZqHJ2cspR5GrQTAiYJU6+pq9LliPphNLC
SGSa0CRGA8SKGZVkkrW4d/KgnImSYB+YlT+Zvx7yTY+cvzmVIrZWaJOlW9R0HbTgx4hNODC2Pj1o
8ZHduk4WMPEC6AeHU0NU8N0PkKNNAbxczlbXhIJiCXvTSqeMSXFgan7yCRNkuNvkpg5FZrlMWoPP
zSMebNjNtJ070ngVv3KPMbMvVgKiC6VUlZFn2+JSZ0zKCM3MWgTa3F1pCqlstCygNAOdCyViuvRU
2cFatHyB8pwvDGmoqIF4UPGARexdjyEIDuSAYikvh2s5NISyO0A9mt4AapcMSDLHlBYzJGoJMjvb
Pln/sly9Lvy9N7unr2fTb17iLs5uuXe1Ff2QN4RdlfmxqN2SFfiBVm25Xn8CWUc32UytlFmNpqFx
KYxBiSkaXloP4Jyphti7GJnNkALWfmVzgpPvkMibx0hW+7N0u+Qy16WAqmJ5hynQcPK7PSqRdo+m
Y8NxhR1WI/03vddx55IRjhMOFejIH4oyRAPcbfgoHJ/2sWXc7MlhYqa/oqK7jqEx387S4JWUrBEV
j+ZP2b/+aOqnkwjS13c8xslEIHRU3E47WHOkOU2Vuz+Lf3n3+kHgA8+KhncwKMW8BAwYV+MJqEf3
c/4kNhLwmjWgYF7dYwL4shf/zlqgWujma886HV5/SLwInrG3t9z8pmFqyAhSZJond2Q4Pm68ouyS
hf8RRKWODbh3A7+4NGxQOd4ye+XArur5kN4M1rzY60lrU0DRgf0I8ej9qRnI3nANxHjK9j3AWyxk
oloSFpLq/I2eEKAlM8Aojgw8Q75OtAnWkQL+QstM7MeY9CLa/C+ZSKzKCA9ChlAgi32oQD+LIJy4
rEEaNg7jwkhFaBrSMzjBytuSuCF4rLfefRfVQXGuZRKv3ZE60N0BiRWgmaVLSYuHaQ9qbtsfqQDK
1rnRv4Z4jA7xP3kZ4a7270FR2EbWxqnzWVmHE1DDa+9gbYNC33N/1ng3c4dAsM7QzW3d5cL645qz
/fWN2HW5gN8n1YWUMFzDjBBIRBOKNKxV2Xu0FfYRrOKJpCiaL8D57oyJQrU3zVEbJ6ga0ltpqtp1
3KS5FFVy5EopRlIyHAtIkTuIHb5pzQw9qafO61xMlUl98n2oKt/YJ5NXEMy/8wYRHXp+JDTf1qs3
agzfy4eaefoxfcL9QBvoo/5iYq5g57TPQLtCoV9pv/XllZgcpWOLxJh44JR2Id+dEog9Mhs+T1NL
hxTBQdSs4l2mvkhjrQXlDTS8fjQizY1xPdWFZkpnukrDk7ENXTu29BpUcga8jtVOfpyVgS0xPQa0
d+Tqh3ryTnkJQytoMNigvXicp96EeD1tDt9E+iGVLEiE0HHJChmUQOdiUqarbDEgzk5QRaFs51rD
Z9RMowWpdfAhOmJ1H2RTpSFaoYWp3MOmwP5AES0mgF8zOTlEFdI9vmRD51GyuTwgJQdHZO4iaWQp
J1T3Q3UJEOjrz58405IZXN17OgOJ/WmnCtbcUAmZiysn96JPDR8fsvxGkhsEFNrQ2DsLioVSfj9f
UOPEpP5b+XMyfq15vUg4j8DoJtAdgvVIT6gWjwmshzFMVeqhplhPSC/d1o2Old21QoSjQtiW/LyW
7oBENKYm8U2UAjOrTO8MT6LQ4xNFBBGkL0FrKV6ubQJr7l7OCNLucaqK9YCmv/aWolpC34D+uRhM
zqYiQ3H4cmvtDTLYDrJGVZxNVR/JWMk5R+W4TEv44x8rLiBbZTig25pC1ZpTa4ipnUJ8GKgNsLao
L8DWqS2rc2SQK4ZUdJF2x+POYieDMHKRSE2uUxEgjj3myADUdAEVUP1CAQVaYGoGVsgPNk/XCwKu
0761+6A+3WSVOwg/idEQiK8PsngMwjtaIyJiO4D91bhgQ/fUXcbCoYMxgluGgnPXlJ1NwFZeMBgK
Xyc5KYDFzm+2rynPgxF4AqgSWHg6xVttclSRXyr62HAW+GffEaVtR9EKrUAblnNU4sCXQGBO42gq
uaR/Wnx29bcohEHhUPjd8cE7fK92pr2Mz6/8K2ni1gXVqsjJ0dqufWf4gKXg7XWLVszswrOOq8+i
orBZDnRKHcPt0n3E6J5pdCQEFOwtH4PAGo8bKDaUbq5lvKLO4n73j7C30qZ8f8feEqPMflRBY8Dq
mRsBZH6Gpt69r+DTHcE/jlzcmvsghi10OPzwT0BTEhzd346pmTeTqcLlx2HxKtQwlCFQt8PZDnoi
K3p0nJuZkMRlkYXtdxg/3LbShosL5+d67pENzNwjJS9Nhm5bEIKAQ6nXXpOoSOBXIE0fLIIu9hc9
47COePL3o5OJcC8Y96N7Kvh8Rb4vlHFgwGkcgeQC9rIRWEBUodwzgOnw16dufz36RFFLRFf++p5J
d7HhYPWn8k5tXCC2vVfF23pM9HzCxnTCdD4VSpHxMYA71XzrYZta0U1I48yT2EPlOincE9zXCIY+
zvhNDX/6h/gsVSDG+WP5DNTj0amEfCsAZVLueb+JuzVU1a/V7R3Qj5Obc46CVsu9DbImsl6F52Nr
N1p44eRUgUKAJgzC5gHDFYYRMFYJXElmbhSU6eadl7Uy0VjBJwI3nAlkU/BoFrRHvIlHUYaF1EDb
op54NLffVOqQ3ZxyzEqWYqXzWnM/ZOsjcMDHVL9SmN1Y2VQBbzTAWQ7+ccI8+5IxLdwHM9Tw7Y/T
Bk4eB0y4kquvdKdRf86nTgezi/4grS4g23WQK2UrJxJ18rlbafI5zDEG43XDIgx8kCtjFtzpqvF9
03cm3C39I1BkS0d/gfygmxMbOsP/lfvAkJfBxi6IVbmTIwbWjN3MEVbuqFLx+NnDlmeJxa/jJlQh
7mIr6IhMC/VRBDdAliUBupnvEalDm/EdS4dMNhtt4Y+9Q8mI1mcWdY3YcMSHaqii8JpDTZ8L1LgD
a/Lx1ifzi9594oJGweGein1uXiP41OI1NbujFJCSZ5kpr42Gz5uGvKEWQbKej9j4/PiPNfGZfXDJ
sHvogEsxECAN4qMaK46iEy5jDAlaSnrGBwvW0jc6+fdd14G/6vXY8+hj5y/ZjhSdugNNSLzw9Ehz
sL/JDUurshzLknw98GFED0UdXn8AG3SSy2A19KMOTogdd+yjowNo9xMqZoY++R39nCB8sPs5drch
Tx+qNX4/20Rjv3QvgLU6KdcxAKTzjxZkujatGy4oVqRRjj3fxDTWpJ+plsqvRhrAXVfGsa9YMvLe
CQRC6N50yFihev1W4FpA6xwjU0PryK2v5aiglcqKlwt1GrkW4Oq/LI2hsEyEqZByStU2mxPgF+k+
2Myl/LX5NwkNNmsInAi5sngszhFCpkpR5HbVvK7LvaPbuE0SUng/aYuAT/9JDCjvnKhRUPfh5YmQ
bc01GMU8ijkXA+97nNme6wnspYGRw0eoxdA1syZcZcuS8EWexqMSwly+OoCVt5iCvgcFPEck2bfa
WXb8/E/ZYw0F2AateHNApCBacPYW1hPJrBpR/NZQFJS0ocH7EPygaY74jGLz8w4MDrDv7lLwZLmB
E6r+R7ejJiqkKyoR+BsMUxyCLlwZ+iE7oqsXzQz1OGIeCLLx0RP0qgS9nbX94QWEbMZnuSsmrDN0
EBCf6iJqsyzFQHVdH3ktW3myUD3mdpLdSW5IhAKBVOrno1RvHfn9sBSf7OGy4KHpxcQrrDJLqIDI
SToVj8sCM6rg67p63u8HBzpo6HjEpMeRNUXO+MWLbzIz2oZlrcSn2orvs9SfF86FtM4lm4sihZRD
aDmsKIuj+hK3Axdc9ZwJ9f9k9UoHnfCN6YMoer/9Zzuh8zEC1QrTqMQEbCrYIJNIj4avlp5MUusq
b14AkYiMcHwbMMg+oZYs49YGePJOxdd7OaONEBueYN8yUvdARZmduxUWSseXI6G3LXZVnWcKB/VL
IXXrEjVRud8FI4su7kByh7A7MRDNgg7qNZz4C7txtOM2iYConFFJQ4A+60d8S2zLermwzW8nNGOr
/BYwLxYrhV5UrRqvirzgHBk=
`pragma protect end_protected


endmodule
