// Amazon FPGA Hardware Development Kit
//
// Copyright 2016 Amazon.com, Inc. or its affiliates. All Rights Reserved.
//
// Licensed under the Amazon Software License (the "License"). You may not use
// this file except in compliance with the License. A copy of the License is
// located at
//
// http://aws.amazon.com/asl/
//
// or in the "license" file accompanying this file. This file is distributed on
// an "AS IS" BASIS, WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, express or
// implied. See the License for the specific language governing permissions and
// limitations under the License.

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
cvbXGwIUDpzqkCnsIYDB4C+VQV5n7pq2Dw7G3h1UV2xWKaJB7FemfXwKK7DdHZ223rv9fqOcp+7+
z1vatlC9Mo0SM0t7ms3e7exOMxK2bqPoaK5MOjt4PpW2OePqRvzjMlRvCjqswFP0wYu2PEwdreTl
wGVnD/wrj0rJ9XOuk1NbN76030MvnSEMsw+abC5ior1ZoxYogE76EWaab3FWk4H303gweApvp4lf
f0oS5j1Xn6tmViLEsj7D3C8+aQca8G9rMM/Yp6+xsTIKMyu3qpKFbxuVGRXUbymwIEJQ+j/pY6uF
D+4NQLsNxM+mCq5tNNOIKS1hvBGqodQqIVT6JA==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
QLpmkGdkR7RgL7vp6Mz3TR9QxWKgNxujaRjBG6ltKTDydZJZWaydKwj49578xVIqb2JnzPQTFTwQ
HMOgjqc/BTHvTk6JI4KqpXMnB+pu5ssCqIhtx7zd/YJC4GpWR50tuFOUcodWuPpgbtqrS97ywbgY
ZP0U7CwbwqcJbZUtGT4=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
YFsCJttmyIAtD6l0g4WvSbqCBj7YhOaSUglb8QTx8UVh7m/UjHOXk9Y3jXM99CatGmdJc57d4ZC5
KPevWq1Ko3k623Zd6p9oz8Ak9iIM0jfh2yHVem064WUnaIShsv51BHH+Q5lg6UCUlQXWcx5vilNh
nwQkuRkqBLWspHBuwec=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1600)
`pragma protect data_block
jrrCz81hlR5dUfVR25qLeOvT0SFkNbl17+TI9xBQcX0r23xBtqwWDTYyjxQUPf5HiuJLHFxFTw8Q
+PpNi1R3hsn2lAmjLgvnkrfydRbBaXjDm76beLOlh3y+QrfxXimF6BzTjqs5yZYWjf6ENWjB1qlQ
t42R2ryiYEj+HYlLNzIf6UAQftMwkfW3DN5lyNIapJPTjqiZ/xwtdCxEQD9EiN9bo1dqio/LqenD
dZWwKCHKX3gZJRYVmWMvwD5xUIdfxFiQu0uZnqxQ/4brqkI8DOKBd9BuUsrNBob1dSDaEat401DR
FL3qWBWWpSMvzba5+UNpLNeH/DsQO955F8LLTIqW6KMBKZ8zu8sIiOjTxx6cPAe73WIUxQhWo9Yf
YxM7VsIS7/n0ugUXvn0iaxtynXV4/+XjRfGFSfh4rBU0cGhq88gH3SsYuVLv553Fy3b6HDchKutY
k4geDPfHI7HveeMdShY8+HsBfM8iTD7cyL51Jw30kH/Qjr9oXSo/E+/rOtqaqKY3VXKh81Uy1qwZ
rGXvEp3gTQsM0ef8+DjOPmpc6oKfvyBaF4nP1EPNxt1EoeS/ECA7wqo2KhvAxON72QOzlPMRzzUS
tmLRUdyZTlVcgOjaFS7My60aVYa6RKtj+V0be5ACXl478E9DNeNlrWRrmr0q29Czsfvdqqav1w38
8crt+Io6iyvRVUHURvqVi3q5f5lFH2WD54ywV5SgqTEbsBk1NLYxaANomNlR5Kucnr/K+a2FFVR+
+aOPEyBl44yjB57ciOSUb44j/1QeLuwH9FX0FSkmR8pjsiOVOdJttJUZx8ypZQiwUvIHTRfRXCLp
hmfA2rrCMDRVemMf+Ddtfo38+fVZtpJpniJnbPb7TAGQcBN04nyrj8G6yXu71YSWqw/dV3aB+J8w
YvjnhVWPeOC4z8Pm+l5vS/ZglWT17KxKHzhb51vkoGwxXWC5UpZWq8+HNpyxPVWdAE0tXI0yMGRG
rwyCNFS27FbVCMeRR9CAmHPQW9NNBCHYfpNT/x8lary5hAfqHoT/lJPGTH1/Y4U4bzLUC3FFmxuV
ZOSyFz/rgmOILa55o5em2A63N3FnCMfzvr0iJVODMT7+SXw2Qa9R7oHjHHbQ42mgL75YuSyL1oQw
9SeXv4iDD8XFJyC2qMt9dckT4L9bxkfXcJa2qw3MH5osFiOQ7/Vwq6Kc4ibriaafNymnMlix9yqI
bi6x50Fc3nO7zQSu5dteBAXDTXb2yFcFy768f/KemR7GHgVxnp6teRG/C6PLKPdgWPglrZuVzti1
BNe9ZwNPGb1cSH9/JiezEbX1bk2GrdJAb/Zgpv5w8zJBv5dNgLgyFQITtGNtUvM8feJT1Azfiy+U
GJGVAQcId0YSS1TgGOnQBLOCuhLNy/vDlDXL67EKfwgWDzxIQggx6d+uaqjvRdqnxRgoWnlrvlBi
Kit3pQuDY9W+2oMV4TazPPdIj0aaUlNT3LPPiLTDCF/jdhONSedThdR1cocXxxzztk5OSX9BSXdS
kCPAxf0Ga10whiA79flrYx2g5Khdg63EuCZ8VfX80DzdzN3DVwZ4re9LIPLtngX0Gn/K0Y7niRX2
FXXzWMdwm0puGCSoJTL1wMu4qysdZx3jKVCAWJT4x5JlQdRqE6a0uuHk95IMKD6yJmH6TbFWNZ2J
MrRlvNrm6n+8fiRwmUNDdn0J1WM2sApY3o000qFUwiMdTcpGTpWd7q6aXUlSFdrwWe0oqbBjJv3E
zSqk+idhe6sKX3KiAky30W+wfUweyuDWljbW5FCoNuxd9SsBlOA3zaRvDox6kKI2AlL/Cm9x8oDd
T78EPs0tjI8aN2fbHPOAGDt+qcCg0auRVmyymzTawr2XvllQlSpvcLDcTXMIJGQEbcoUE7g2SlBk
3vcoss4qvq83S7QlKu6Kdo+NAXHEW4/RtTN5M9UpfmMdtS8pUAGruOThCkiFQCQo0GWC46svh+3k
WO5EdZaqL0lCOnFZtEOHZtDbkB8+fBbSkK3ott1rCFdySm9xPtf7cB7EmnSejjufVsr0WVlVqrK+
X/SeCBJdLh5Caa+hVKIuVeWZyPwdt6AguK354yjAwOBmcrIVF6sUwaq+BuwXwr24LY/86PMBBPzE
fuCoJA==
`pragma protect end_protected
