// =============================================================================
// Copyright 2016 Amazon.com, Inc. or its affiliates.
// All Rights Reserved Worldwide.
// Amazon Confidential information
// Restricted NDA Material
// =============================================================================


//FIXME -- Need to do the clocking correctly:
//    - Async Stream between PCIe cores and User logic

module sh #(
                     parameter NUM_HMC = 4,
                     parameter NUM_QSFP = 4,
                     parameter NUM_PCIE = 1,
                     parameter NUM_GTY = 4,
                     parameter NUM_I2C = 2,
                     parameter NUM_POWER = 4,
                     parameter DDR_C_PRESENT = 0
                  )

   (
   //--------------------
   // Main input clock
   //--------------------
//   input clk_in_n,
//   input clk_in_p,
//
//   input rst_n,
//

   input                       clk_xtra_p,
   input                       clk_xtra_n,

   input [31:0]                cl_sh_status0,
   input [31:0]                cl_sh_status1,
   input [31:0]                cl_sh_id0,
   input [31:0]                cl_sh_id1,

   output logic[31:0]          sh_cl_ctl0,
   output logic[31:0]          sh_cl_ctl1,
   output logic                clk_xtra,
   output logic                rst_xtra_n,
   output logic[1:0]           sh_cl_pwr_state,

   //------------------------
   // PCI Express
   //------------------------
   output logic [15:0]         pci_txp,
   output logic [15:0]         pci_txn,
   input [15:0]                pci_rxp,
   input [15:0]                pci_rxn,

   input                       pci_clk_p,
   input                       pci_clk_n,
   input                       pci_rst_n,

    
   output logic                clk_out,
   output logic                rst_out_n,

   output logic                sh_cl_flr_assert,
   input                       cl_sh_flr_done

   //-------------------------------   
   // HMC
   //-------------------------------   
   ,
   output logic               hmc_iic_scl_i,
   input                      hmc_iic_scl_o,
   input                      hmc_iic_scl_t,
   output logic               hmc_iic_sda_i,
   input                      hmc_iic_sda_o,
   input                      hmc_iic_sda_t,

   output[7:0]                 sh_hmc_stat_addr,
   output                      sh_hmc_stat_wr,
   output                      sh_hmc_stat_rd,
   output[31:0]                sh_hmc_stat_wdata,

   input                       hmc_sh_stat_ack,
   input [31:0]                hmc_sh_stat_rdata,

   input[7:0]                  hmc_sh_stat_int

    
   ,
   //-------------------------------------
   // PCIe Interface from CL (AXI-4) (CL is PCI-master)
   //-------------------------------------
   input [4:0]                 cl_sh_pcim_awid[NUM_PCIE-1:0],
   input [63:0]                cl_sh_pcim_awaddr[NUM_PCIE-1:0],
   input [7:0]                 cl_sh_pcim_awlen[NUM_PCIE-1:0],
   input [18:0]                cl_sh_pcim_awuser[NUM_PCIE-1:0], //DW length of transfer
   input [NUM_PCIE-1:0]        cl_sh_pcim_awvalid,
   output logic [NUM_PCIE-1:0] sh_cl_pcim_awready,

//Not used   input [4:0]                 cl_sh_pcim_wid[NUM_PCIE-1:0],
   input [511:0]               cl_sh_pcim_wdata[NUM_PCIE-1:0],
   input [63:0]                cl_sh_pcim_wstrb[NUM_PCIE-1:0],
   input [NUM_PCIE-1:0]        cl_sh_pcim_wlast,
   input [NUM_PCIE-1:0]        cl_sh_pcim_wvalid,
   output logic [NUM_PCIE-1:0] sh_cl_pcim_wready,

   output logic [4:0]          sh_cl_pcim_bid[NUM_PCIE-1:0],
   output logic [1:0]          sh_cl_pcim_bresp[NUM_PCIE-1:0],
   output logic [NUM_PCIE-1:0] sh_cl_pcim_bvalid,
   input [NUM_PCIE-1:0]        cl_sh_pcim_bready,

   input [4:0]                 cl_sh_pcim_arid[NUM_PCIE-1:0],
   input [63:0]                cl_sh_pcim_araddr[NUM_PCIE-1:0],
   input [7:0]                 cl_sh_pcim_arlen[NUM_PCIE-1:0],
   input [18:0]                cl_sh_pcim_aruser[NUM_PCIE-1:0], //DW length of transfer
   input [NUM_PCIE-1:0]        cl_sh_pcim_arvalid,
   output logic [NUM_PCIE-1:0] sh_cl_pcim_arready,

   output logic [4:0]          sh_cl_pcim_rid[NUM_PCIE-1:0],
   output logic [511:0]        sh_cl_pcim_rdata[NUM_PCIE-1:0],
   output logic [1:0]          sh_cl_pcim_rresp[NUM_PCIE-1:0],
   output logic [NUM_PCIE-1:0] sh_cl_pcim_rlast,
   output logic [NUM_PCIE-1:0] sh_cl_pcim_rvalid,
   input [NUM_PCIE-1:0]        cl_sh_pcim_rready,

   output logic[1:0] cfg_max_payload[NUM_PCIE-1:0],               //Max payload size - 00:128B, 01:256B, 10:512B
   output logic[2:0] cfg_max_read_req[NUM_PCIE-1:0],              //Max read requst size - 000b:128B, 001b:256B, 010b:512B, 011b:1024B
                                                                  // 100b-2048B, 101b:4096B


   //-------------------------------------
   // PCIe Interface to CL (AXI-4) (CL is PCI-slave)
   //-------------------------------------
   output [63:0]               sh_cl_pcis_awaddr[NUM_PCIE-1:0],
   output [4:0]                sh_cl_pcis_awid[NUM_PCIE-1:0],
   output [7:0]                sh_cl_pcis_awlen[NUM_PCIE-1:0],
//   output [7:0]                sh_cl_pcis_awuser[NUM_PCIE-1:0],
   output [NUM_PCIE-1:0]       sh_cl_pcis_awvalid,
   input [NUM_PCIE-1:0]        cl_sh_pcis_awready,

   output [511:0]              sh_cl_pcis_wdata[NUM_PCIE-1:0],
   output [63:0]               sh_cl_pcis_wstrb[NUM_PCIE-1:0],
   output [NUM_PCIE-1:0]       sh_cl_pcis_wvalid,
   output [NUM_PCIE-1:0]       sh_cl_pcis_wlast,
   input [NUM_PCIE-1:0]        cl_sh_pcis_wready,

   input [1:0]                 cl_sh_pcis_bresp[NUM_PCIE-1:0],
   input [NUM_PCIE-1:0]        cl_sh_pcis_bvalid,
   input [4:0]                 cl_sh_pcis_bid[NUM_PCIE-1:0],
   output [NUM_PCIE-1:0]       sh_cl_pcis_bready,

   output [63:0]               sh_cl_pcis_araddr[NUM_PCIE-1:0],
   output [4:0]                sh_cl_pcis_arid[NUM_PCIE-1:0],
   output [7:0]                sh_cl_pcis_arlen[NUM_PCIE-1:0],
//   output [7:0]                sh_cl_pcis_aruser[NUM_PCIE-1:0],
   output [NUM_PCIE-1:0]       sh_cl_pcis_arvalid,
   input [NUM_PCIE-1:0]        cl_sh_pcis_arready,

   input [4:0]                 cl_sh_pcis_rid[NUM_PCIE-1:0],
   input [511:0]               cl_sh_pcis_rdata[NUM_PCIE-1:0],
   input [1:0]                 cl_sh_pcis_rresp[NUM_PCIE-1:0],
   input [NUM_PCIE-1:0]        cl_sh_pcis_rlast,
   input [NUM_PCIE-1:0]        cl_sh_pcis_rvalid,
   output [NUM_PCIE-1:0]       sh_cl_pcis_rready

`ifndef NO_XDMA
    ,
    input [15:0] cl_sh_irq_req,
    output [15:0] sh_cl_irq_ack
`else
    
`ifndef VU190    

`ifdef MSIX_PRESENT
   ,
   //-----------------------------------------
   // CL MSIX
   //-----------------------------------------
    input               cl_sh_msix_int,
    input [7:0]         cl_sh_msix_vec,
    output logic        sh_cl_msix_int_sent,
    output logic        sh_cl_msix_int_ack
`endif //  `ifdef MSIX_PRESENT

`endif //  `ifndef VU190
         
`endif // !`ifndef NO_XDMA
    
   ,
   input [NUM_GTY-1:0]        cl_sh_aurora_channel_up,
   output[7:0]                 sh_aurora_stat_addr,
   output                      sh_aurora_stat_wr,
   output                      sh_aurora_stat_rd,
   output[31:0]                sh_aurora_stat_wdata,

   input                       aurora_sh_stat_ack,
   input [31:0]                aurora_sh_stat_rdata,
   input[7:0]                 aurora_sh_stat_int

   //--------------------------------------------------------------
   // DDR[3] (M_C_) interface 
   //--------------------------------------------------------------
   ,
   // ------------------- DDR4 x72 RDIMM 2100 Interface C ----------------------------------
   input                       CLK_300M_DIMM2_DP,
   input                       CLK_300M_DIMM2_DN,
   output logic                M_C_ACT_N,
   output logic [16:0]         M_C_MA,
   output logic [1:0]          M_C_BA,
   output logic [1:0]          M_C_BG,
   output logic [0:0]          M_C_CKE,
   output logic [0:0]          M_C_ODT,
   output logic [0:0]          M_C_CS_N,
   output logic [0:0]          M_C_CLK_DN,
   output logic [0:0]          M_C_CLK_DP,
   output logic                RST_DIMM_C_N,
   output logic                M_C_PAR,
   inout [63:0]                M_C_DQ,
   inout [7:0]                 M_C_ECC,
   inout [17:0]                M_C_DQS_DP,
   inout [17:0]                M_C_DQS_DN,



   //----------------------------------------------
   // DDR stats
   //----------------------------------------------
   output logic[7:0]           sh_ddr_stat_addr[2:0],
   output logic[2:0]           sh_ddr_stat_wr,
   output logic[2:0]           sh_ddr_stat_rd,
   output logic[31:0]          sh_ddr_stat_wdata[2:0],

   input [2:0]                 ddr_sh_stat_ack,
   input [31:0]                ddr_sh_stat_rdata[2:0],
   input[7:0]                  ddr_sh_stat_int[2:0],

   input [5:0]                 cl_sh_ddr_awid,
   input [63:0]                cl_sh_ddr_awaddr,
   input [7:0]                 cl_sh_ddr_awlen,
   input                       cl_sh_ddr_awvalid,
   output logic                sh_cl_ddr_awready,

   input [5:0]                 cl_sh_ddr_wid,
   input [511:0]               cl_sh_ddr_wdata,
   input [63:0]                cl_sh_ddr_wstrb,
   input                       cl_sh_ddr_wlast,
   input                       cl_sh_ddr_wvalid,
   output logic                sh_cl_ddr_wready,

   output logic [5:0]          sh_cl_ddr_bid,
   output logic [1:0]          sh_cl_ddr_bresp,
   output logic                sh_cl_ddr_bvalid,
   input                       cl_sh_ddr_bready,

   input [5:0]                 cl_sh_ddr_arid,
   input [63:0]                cl_sh_ddr_araddr,
   input [7:0]                 cl_sh_ddr_arlen,
   input                       cl_sh_ddr_arvalid,
   output logic                sh_cl_ddr_arready,

   output logic [5:0]          sh_cl_ddr_rid,
   output logic [511:0]        sh_cl_ddr_rdata,
   output logic [1:0]          sh_cl_ddr_rresp,
   output logic                sh_cl_ddr_rlast,
   output logic                sh_cl_ddr_rvalid,
   input                       cl_sh_ddr_rready,

   output logic                sh_cl_ddr_is_ready,

   inout                       SYSMON_SCL,
   inout                       SYSMON_SDA,

   inout[3:0]                 fpga_uctrl_gpio

   //--------------------------------
   // Debug bridge
   //--------------------------------
`ifdef ENABLE_CHIPSCOPE_DEBUG
   ,
   output drck,
   output shift,
   output tdi,
   output update,
   output sel,
   input logic tdo,
   output tms,
   output tck,
   output runtest,
   output reset,
   output capture,
   input logic[31:0] bscanid
`endif


`ifndef NO_CL_DDR
   ,
   output              sh_RST_DIMM_A_N,
   output              sh_RST_DIMM_B_N,
   output              sh_RST_DIMM_D_N
`endif  
                               
`ifdef I2C_SPI
   ,
   //--------------------------------------------------------  
   // I2C
   //--------------------------------------------------------  
   output logic [NUM_I2C-1:0]  i2c_scl_o,
   output logic [NUM_I2C-1:0]  i2c_scl_oe,
   input [NUM_I2C-1:0]         i2c_scl_i,

   output logic [NUM_I2C-1:0]  i2c_sda_o,
   output logic [NUM_I2C-1:0]  i2c_sda_oe,
   input [NUM_I2C-1:0]         i2c_sda_i,

   //--------------------------------------------------------  
   // SPI
   //--------------------------------------------------------  
   input                       spi_sck,
   output                      spi_miso,
   input                       spi_mosi,
   input                       spi_cs_n,
   output                      spi_int_n

`endif //  `ifdef I2C_SPI

`ifndef NO_XDMA
   ,

   //-----------------------------------------------
   // AXI-L interface to access XDMA configuration
   //-----------------------------------------------
   input [31:0] cl_sh_xdcfg_awaddr,

   input cl_sh_xdcfg_awvalid,
   output logic sh_cl_xdcfg_awready,
   input[31:0] cl_sh_xdcfg_wdata,
   input[3:0] cl_sh_xdcfg_wstrb,
   input cl_sh_xdcfg_wvalid,
   output logic sh_cl_xdcfg_wready,
   output logic sh_cl_xdcfg_bvalid,
   output logic[1:0] sh_cl_xdcfg_bresp,
   input cl_sh_xdcfg_bready,

   input[31:0] cl_sh_xdcfg_araddr,
   input cl_sh_xdcfg_arvalid,
   output logic sh_cl_xdcfg_arready,
   output logic[31:0] sh_cl_xdcfg_rdata,
   output logic[1:0] sh_cl_xdcfg_rresp,
   output logic sh_cl_xdcfg_rvalid,
   input cl_sh_xdcfg_rready,

   //----------------------------------------------------
   // XDMA AXI-4 interface to master cycles to CL
   //----------------------------------------------------
   output logic[4:0] sh_cl_xdma_awid,
   output logic[63:0] sh_cl_xdma_awaddr,
   output logic[7:0] sh_cl_xdma_awlen,
   output logic sh_cl_xdma_awvalid,
   input cl_sh_xdma_awready,

   output logic[511:0] sh_cl_xdma_wdata,
   output logic[63:0] sh_cl_xdma_wstrb,
   output logic sh_cl_xdma_wlast,
   output logic sh_cl_xdma_wvalid,
   input cl_sh_xdma_wready,

   input[4:0] cl_sh_xdma_bid,
   input[1:0] cl_sh_xdma_bresp,
   input cl_sh_xdma_bvalid,
   output logic sh_cl_xdma_bready,

   output logic[4:0] sh_cl_xdma_arid,
   output logic[63:0] sh_cl_xdma_araddr,
   output logic[7:0] sh_cl_xdma_arlen,
   output logic sh_cl_xdma_arvalid,
   input cl_sh_xdma_arready,

   input[4:0] cl_sh_xdma_rid,
   input[511:0] cl_sh_xdma_rdata,
   input[1:0] cl_sh_xdma_rresp,
   input cl_sh_xdma_rlast,
   input cl_sh_xdma_rvalid,
   output logic sh_cl_xdma_rready
`endif
    
  
   );


`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
X3+x/zLAvBl3AfFUnKJlfXo9S/FLDfQj06ga2K1mv2mmEz9whyq7E9Gkt0hm2k8fGg8I+brOHLL0
HrusKmVVh4mZwscWsXrf7g5b7VgYVO1FPt3E9puWUNDFAA9FRblM8/ITFoH8aU/W0XZhwTa41iYZ
80brmbGmVpCeCib1OqbtZjDeLnII0V3+XY7HkZbeAGR8w+8FnDJwXxnjR+cYzvAL2b1jRk6PnP2u
025SkPH2x7yk+pOtKGX0YORMfnpbXL1ENtolW5mP0SyYOBXthGV/yUtNKga0Hw0IUMTt/qSBqY6+
d/YWIplVeitljeJhJ5ur0Khd27bTIdXxf4i+OA==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
bEs7rhLaPQTtAfLBeEGbmaBDeCe7vebYbsyZ7G4GvLZI9X5IskOUjgHLBynNBwJBM8MhYg0+Zxuc
oaLoW1AwZ1qzjnkU+xFOJpdhUIlQkSHCwdI53pzanF7Ke/aqwXRTo3O6qhO8xP9z9AXmv9ZWutTJ
4dHmi6Li0XovLZO0iqI=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
KQV0JQQ3Wba5xnxW7AzIf6TUqaXvCAoI0W8SXSCOivHdGCvoauX5HCJDzKt/zY4jmZ/Araat1KPO
Ql4jcaEDC8GxAv1evguZTTZU0xfgdTugr+0+6kqOWezhGfU/MPXlFBpgR2A9wGrKruy/XXeKOInh
UDS15RNBrnZ5WFVrEac=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 118416)
`pragma protect data_block
4dDFjwbH5EgfuI7O73Q3+H5G86Cvn1A/0KIKwdOWi0dtyhk9OIIulBeERYW7KfavjYenlafPoIpp
GmAjzhZik/otklVuyeoaBz1JO9B8qQCbtd8KIo4QMWjW5m2SKowwAjJauzyNCw96Xc4iuR/kQgyl
4Es6g2JT8UwPET/6wTiEkvnwnHtlkWjEDkhM3sOOXH9FtmxWhUoe7+n6pjMzMlL179fVWRcXdNCB
krEFmMDyvG2odIzvcROoUdJ5H+YGiqoq3YecqeK9RXUbSmJ7dYYdhd+JCSHE51gYPXp7tFh6C7lF
QMwaedKMy6ny47fKtFQLGyU99J5bH7Irc7vo4+SzPlr12kSD0qFP4YQGzcee+ghgQiXkWr8UK7qR
D92skxM5HTkKxdqiDbDLXXdOqcjc85W1nqNukFPLQiPgbwy9EyJKzs3gDL+I+PeWrXteH7raIWgw
udlv8gEkTF+OzGWuaKKTQ8QMkwKPNzNqpusY7Il5liC1fiY+SkhvSAEckcplm2iLEQ384J6CgXWL
AKqxliv/vO1EGHAT+0HMW3k5AZrp9hL3p0EhQP8Dqo192QUPq+w6NQBzj8veUxI/6g/kQBOcJ5BI
9wTl6oJOfFMRfbbgg/SzIgwy850+ePOcU+LtN4FreCaetDiDvbMBG6XhvHcpiDjUYMbc2afl5WD0
gpTRRCCYiV2WIReeSOeOFpqN0193WDNnsOj8Kcp1jVNfFnfoKkdzh0Ug9z01TZi5D1dvcVDWPumI
saoNStajldISAy5wuIM+MeE8LW9ZCUE2sHWULAyKf8ABiKjb0Sh3JsDWkC47lh5pUxAtZGpwbw71
fugL9k7YhlynMUx2ydRezND3QsNSHjvvFCS0PsKZ7kqp0Wbg/W62AeDrtaXry/I5TAtNVd6/AvTC
FQUxDMdQWuRq4zKetP9QGomhNWrlxKVExPMwpakp4XYJcQDg6Vugy0I1uafKVw+mSw5yAOViU8NY
GAyT7k7rJlS4TIEkwcJ33KfoBB0v4Xkht0OUwQgf+ytT3RBTKrQ8IeRvmFUrmQKBRPZ03814h97s
haPLii1+I+Jvc/vaxC3pmIfAhIbws1TociES7zXY5Tyjg/Tu6xLQOAX0c2tiwEMelrlHmHokqFN2
34iJwbsQcCEVlYMz0bpMHWgir7XRwd4suqadIprNFY0datRQpJn38OjXLdAdWBvqDzED0rvr7oDC
VJFs5nORvaxqYpY17cmWXN7Hsadmfza75OJOtgHfgPVleYI7LGEPLgwmW7byW5vzEZxUCnmgofD5
bMUXmGGV8UMi1+wG4/dsyTP/YP10qtxy5oIw+xbS2RIBPfNXT2ub/XW5K8Jt6HuMgN3BCgbn6fWR
LXUc4fXeLHYju5vgyyZsj6vfALa9vdUUIGVrDH/e4xkkOB/gCb97SZAAUwgLfUYNH/Dv0toHgnbC
uTWP+gyhNaAZ5T/1voRVf0+huC02wa8lemd/Wrucw8GUmBiK0nzDg7o5jRHtGPIAzGNSNgSVAH4L
QDzZ6Sd91+2rixexc6XWdcAM1O0rJGrtxxiwwR4DjgeT63qtWzRyjzzmycqs4g3NT/Gdr0dtCl/6
b3mgv4l9upHlb1zSUElF9YiSwwYIHjhqJsyhZy3ibZenNbVr9EtFQXGoZxZI0hajZmIkywCb2u8o
tWhyGg8ORt6pK+1AOXt0dh8QLEeToCPOHsTh5m4WEGhuyCQi/lxN+OyPZABZfdPGyIfGDqPlKdTl
sSt7wqKDEO1r2KH9vnt1E1CqWMT1W1bsW+yQmeYrM26tJlUEV7qwfJyszukIwTzZHSeqcUXD2Htk
YRF7q4lQXkAm/IKA4oYeD5P86PpWzq74dqRGuss80tXWP+jGMuagzxnAUaWnujZ031k788xuPLpk
qU3DM0CaygZMn18Z/0artm3nN9s4Ey6/xuX9i55IdCFzbTYZ/6lGss7WppeLBF98YIxsufwhtGCl
kumyPCSEq2T2+TueYSIVO71hx4q5lX6Dz1PCDCw8O91TPWHNWAlNNZHNjISQQZ2cW9IU1+4TRn57
RuZB770u8RWoamG7iRQzk5a5L95+Z6nb5dbc/HrsHR7Skx17/frPoFzyfO8h8zu9I751alFSUhQX
JGZMoAWkmjsAuwacBACHEdUna8K1ePyCmJs9WzuhTIlxpFe2L6EBos4HrirIsvyxqCNnLwf3E3Cz
fTEYw1AEHI7q65JA47/dtBuofLzW1iPpc7Fu5HrOBT8ipL4hom96hWZx35hYxbxLHIQM1/dxDBQx
S9PxpI4rak4lUTs2mFL1IL7IwqJzVJnKlACGIBYRUHW4+H78UURdqWtOW28K2LZWi+HpkdUm65uc
ZDmSEwP3WKccybVdsNFqfk+L7O3mxLycIGeOi93V5VM+RtrwTpXApxi+JG6o4NLyRPZGspAMH3Ph
0wExJU8mReVVcvCSXiMxQLGDQIrqI+Bu7srSM2bQ/Xu1EfhJXOvHvu/tcFhG23otn8Mo27iVaxUp
1bE2Zd1u3juE8bhdgKfwtuUtvRXQ5JNSvVMPSVeHTBgsqzxekSr7Z0NMXF88s9Zij4rGqJHfyLdW
LVMZBux5CX0cUbbNvlMG1o80PDnmnBThr/vxo29Hd4fIZw3OGqx/nOgkuS2O5ezYGLnmqkkwf1Yf
uxa1r/mjWJav7ALY/iYPM4J0GLGdSdCLLu/QbX6exgiazetYI16kj7xchO22sRA0alLLuc4Kvi36
L0F2d/NBzfg6zVaZF6rKSOcF2iCkIUYpJWzvilT4k6g7Wi+dKOcHFKbqXXOsgxTybi5F6NfQvSVP
NPyLpqm09M6HvsAk1pzWkodTyeKH5R40wrJ2INX0fbHMKDtAMU3UZtSd9uO90pS+he4I3TlkxbPP
XeHickRTN2L5E/W0Gm86LTBCWsDY3pTVuTmSxKoOyC15xl9jHeqNp4QfjkxP9ffCv3CEURJkHTOu
JAlLW1L486v8dGpwWF1Dwir5tcdSjLA3C0nTDRRN+sECr5ifdXjDcM41bmBl58hWpQGvPLLOWslf
POT5Gw1mCHsJpsdLN9CxIg9OECuNAXXr4YxfgB5p7Nnx/jELnOQSK37PQBdXlllTNDqoJ5J0yDZb
gxGrrq6UWfF8GyrQL9J6YhlP1hAy42LG7ur1kqfxXU7xwC+T0zsfN4exjhPDyU1Qv8JrTyUxwlX/
nYOPgC0ahVpbFsS5EQlY7L/d1EKBH6CUct0sb1x+CSGEEc11wVxVuAtIxcFGAtFQhxoMcdGuEYn6
MirsiuSz0fmziTZbVoe/ZOm+X7zf17CYEE1V2e3enwEYJz0ZmSAbDFd4sImC7pCQ5JWBPs4vh6a5
2IYFMgm3Dmf6WjngL30l2pgKYZ2CLO6Yf1wH4y1DjaRNRsPleAY8UVaH6jMbu9KLYEwW86a3kKrS
zgFlRqgzdI1fsHr9SgsxSL0Zm8bf+fjeKk2rqdO4F2dwRbROdCIsZk3v2fDI4oqLrw6El8l9U8o2
VChlUA8sVtYkkG3cWcFSgrnC9qaZc83AsrALxOO3cEQQ/sxA+8uwL6VQ4axvqWaGB9092LEVmUSo
Qk0pd7opLOMXIrnkTtmsdSl6PRwFT/vf8QZthxQMQNbIt63mCY+8vISKr5GRARba1+XQ8n+vfBPC
Sr6/GXq8RWLmsDBwDiEG3cWDnaMDXqMBwiEn8i/HhvUXnf+v09KdDSH8Co9ul0+uvBBs70RUtIYW
tYo8TbplPBr9BgO0d+8y/mYo7YSLUrot4XcpSQvyySXFb8ncxg0ZX6DED70E8Rl42JiVYUqgwU0k
eJfAKBhIqaTQPHASRNu5yaTWLt/oHR2x16b82ZhTHyIoJmxAyfh/EKIor19FHG9Ryxn71EIfIPM1
hWZLmN++vXcQZGLEDbBFoOQerbELZ88aDb2IbAejynS9JnRa56uljL8SCiX0W8l/mpNXYMZzjlIo
7Q9GFki2DnliflaO9NS4JAZtjR+Mgg26YS8xH1O0RBDmp7NL0WoeeRzbFqAprAci3LCycG/TkZIu
8smKxd0Wc9gck75zrwx2184MmUfGd8ytH0+4REEscmdhsYmicVoTFqhva2HxDc7nrckTe7sNV2rY
imUueMjGd9da+xRXSq2yRTnUdu+LTAQAOIwLxSok225qo9CWqUJuFMpm1IJlzK7n8zZ2E65YQcEZ
DwQR+v8SAvPRKfh1vhVn2b+tRUF4HBhk1cr/BcRGhMqKWcKLz+1Gfd4moJmA9xNpmCKbzGwIFl8m
Oo7d1KHbuH0kAP0TpkPQx987OUjTaqI+jmCIE0He5q6peJSO2OFwPrdDtuvCAQoOO7hX68NY+re/
zFNy7hM2/I/mCp6Rmn1XxZwLhW7MTMonSxqsu2MQ5GK+pcz7KkoOEF7pBIZ0l12BKwxkq0GBuP/x
q832dQT2dq4fNkowBb9wbuHl/4pqO4d7ZBLWqlwpoiWIyYN7KibHYdXsMNNGO9KOD/fWnhI4vqbF
V5XRLeVLUg7HSLIpMM0LdsDPDTtP9CTm3cXjMn65kj4LuAomB1HDdUY0XWA8GE7fgEiIt5S+F2Tq
87F6Of7gSaJDVS34ASxZ4ffjINB7cFxV0KYPxGhK0Mpgj9k5OwKJOK4qjPT3dLShCKc/1wkm6GbZ
VGs6xNhNsMz0b2OjkdtapaSBJ7sysHiom2IvpzEQh/YueFY5hzx18FzV3P/wp/xQyN6DW0bvP83L
GFyV0CXVLn66gmgzQrDnWLccrykhG3D45pN7VT3K8/KH7lD1Q/IIUSR6hfIdxkdwWVyju7ZDuy88
51K0RySWcYc3C15hctX8cZYheoT4CN7rp4gfATaoaCfg5z69PXw7mVE7YdZpBvAsxk85Ys4KdzzA
wYmZ+hzc/AEViqg2SLZKeBkJfqEd3daGj4llIvyfmjt8oV3xX632yBQpYnbrjsL0jFqemg01QIN+
cRULomiD9gy0vZ8JoMPXz7pzu8bo6RMV4zSDjoxwvYV0MijHuZ64+5+8ckjPv91c2g87JAnjNKx0
phjW8tFz9DB05552xxsPr37smXy49WrOdAzvxXJip0v5tzzKfMupiLYfl0FUToIbMpINmDnmz2bB
mC9pw/Kznk7bpjz2cZoLldZrshH8eiTnVLolHiEzXZ/qBPjAC50GXqBPq2MZvOYqSay0X3dcbyPa
hHfQOH89M9lZQBpzZ5f4yopTGgxpZGFqABZgFXehk9PwOvfaSmsWEbEF7bW1O8Z23KCSgbsyk0/Q
ee6GUyqWYw2CWUXmkwlxOQWslK8OXsRqE4yOnOWJ5NgmZug16FsY6NJoyomV57nihGEEXYdZ4uDs
QSVV48S+lhlxIXb/n8SGpUx9ftYaF7KV9RZuUEj334vbAH7WZQnhCq7L8oXbFLhq7FSls1T0L1j/
Cia1z3E8duYg+DSO61kckL4mYtm9oFJ0k1Sa/kxfJ7JAzXP8oXUWYYOwKctd+OCHLXUtNoEnmYtF
FKOT+NBtjhummWCF+UcmdlGmTaz802Wz72enzGk/6qCuRI8qQOVVj/q4qRldJf4zyXd+mXAkbIs3
uzM8ILkVHVavHkavNQHL6goiMte+ggF+QKKH1FwO8+jEUBrrbAywt2E6TJ4MkE6D3VRRbovRkxLf
lCRR4NVKGg8gmXuJBnGuSBctp7pe9zSsB7OxejjIA9pEfqDb7xNSGUm01PESvgJ1+F44IyEpgG1Q
bjhlqjIJp171yMHkGyRlz+C+yONmrdpVYYcyoQBs9jCyc5wJ7bk8FO9Lyw+NZKvykAJIn2qp4fj0
xz31Br+GZhNvgMEI5zZyr7ryu64Drc5pCiyLT2ARP/oV8fLf2YIzOfCyzS1bKprstowLmjBHkAoB
yMfAKD4I3SrPMnxmjRLMx1sopc2Wm/dmJFqKLzdoLMHDYMKBpSL1iSGtycFZMAHJiIVuq4zxqFTV
zcpsAUrEHNF9FhzR0mPxguC49vpVIUZumPdf0ffA3TN6QFT2RUGaGHrThXG03IHLD0ekBcBcKFgZ
qRR35uvUCin6pTwM5dJL2M2f1lqG+lZKtoQfMhiDG9tH2jEHYSPVPUvB1oRzPFnvs6otKA9HhYTD
Rd40dTFMQohDUstMSSYXj0kjr6v59h/rzc1cv4h5r7RNj7HENKWCxmuMffkNsPjIV7Mfde4xM2S2
xZDsSp5vvJpN2nsZjZUMoe1c8Wi8YTfQszADaLJIaKK5UIYBMcSxw78d5F6CuOc/cJc9mlS2ZNZU
pd2+tmYdMWEeuaC8VRl3LTFI+JKbV+HTbH5OHE90fJlqJ+N2kbL5te+liPcq4TXTgmworc6w+i1P
aLJhyYAn+tGiIaKQob+e0EhqXXZJL40dAXg+VYBbnW85xL9YEGA3UeMDT8YXC7I3iON/hjmdfDVo
8uE3cIuBvZlnLlnPmLQTWH1fkMB8CkettNHBB1c/EvPeXENdnrWzY5QzduQwzPFeC0kxlFPyA20K
jIjfezBc+r6qIEzr04XcFEFqT34HFUb0DOLyCIZriQv6E1A4Vke3nYtq5GkMmwGn4Fx/sd1+KhKS
tUqVEbOfmlR4GDnvbmSt7f/it6gGXIfdOBxwmr4wW5r8CV+zj8amcZfGq9jlAftJ0P1PEt2t7xYc
lFBO4A9cETYdx/phoe2IoItUIqe3HG2H356m+GIQEkWATeD1pDSTndsnez0I7wb5n4irOYrtYxlI
HCX8w+RTqeQs0VOqKnnb1tlafG24emkjk+ufoddLWV1EQ2RqwR6tslsljqhlxsLiaaNvgl9VMb7r
UnIfcZka89XbXe1csH2GFe+74+Tpv/UhUpvnbh3oSVfVpH86gWa9vuETHieugtHCUSq87Fzi4ONE
Z2Kp5DBPSzcX40KULWwWWm+vi6YBgOyW8ypN0h90YwDnHd0bpY5OrbB8CajK0XE4FBwxjsNiqZy+
iFVOzR1w8HSEquWA17MNjFwExmB/GZBbefJoEfQhABBRbwQG/GFMYPmADm66EYX/VUupSgeFvWW2
o5IA2AJrd+dtDPwwrYx9XAop/LqoFo8Jz+2YOJiYifFgphG9k6QCHNWK7XOjjJM075AAYlYzQrPF
CkzRszkRJpt1V169kDBx+7Df4Ylh8MfWEMKeZ0ib9ESzFyRaRcgB5j6ieTTuVGiGR+a+HovUz5Rl
RcHhkOCj4l67Ym0+/Bv3enRJFAdK8ng2jeotbtZUmDCf0tVMsy0m07wpmOESxcNTRYLawUNX9//O
c7yTg1yf6fNyYE//GRuAWCjiorZpPEJFLY/kYA3pkfo2S0SLY4MUyDzQaHC4F34Vge2GEdykN9X0
sLusSdKFjnDxgVJqxtkPwIBfVniTY57lWLcpis5KqrmR9EDmZpLDlTskAEhE8Jerbc6faGQRgZA0
dVElfX2Io6Dj+7Wfq4UQ5mHV5x7FeprqAP4yVRVNe8psRlm+XruFcNIj4NdM9Abz5FBBbra4Apti
hB3Nz3C1pjyQhosKbbCwTIR/f2CdbgRmpKFGhjmiJV5K6+5jXldGLjXCa2dqf9CfI7CneWfgGL40
EsFy6t1wuHtEqBSBGB1fQ0zB2XO3pHiHXdvaoBFsKVlIBYvI2+CliEzKY+/+CHw7Dlp/8UrSGjFE
OIzY8H31lJtB2uM4+3TSRDdHoDkxXfiqij57AjCPA0J/TILV0ilmwF3LAUMBSOfcOmatX+KXDrPF
/KtdQ4kDe5/v5iNhmYsrx3XhxCqoR5BN8oXm0FbSSJ7eqyH+zVgO/JTAJG9MK4JWM7gaYJcxS8Df
hyX1tXBlgZhxIVMKyUjFsbp5nJlTjl30CLqxrVCHbJOYBrA9VRVDXybVDW4y+HZXWttEsVtT7o09
r3EQsTIYlN5IHnlZhjn26UiTYzUFFn7iqCQl461WaRD/WRew20j25uaVj9/rAMlb8KQXjoksdzX5
rAi3KNznfxvQrQ2fUA7eFF58sRZ08uDa2i+JPAe5qFai+OSXfAFXtybFNSM5hDdSL1XXP7+xW5Sx
wFkyWgWo+HuTVdE2eaAY9s/fUZKWwsnUYR/Ix7YqmyoFM3rBqHgW06TQ/0ihmLZPqQvDYsrj1KIk
LP71M3rULlCAIMBkQDAFsY0StQPqcbSBiY91ALTePNoBN8UTWSA3TaR+lTswnrOw3Q1AJO+CMJDy
63P6YQSzRpmX96xPqtASIy6pFzm7M5GqASJaSz9fLY+eXe4gA0ftnkObg7aZhJjS08jqOS1aqS9X
NqmQ0k2ACVnyUSECWY0cM4i7Y82aDXuXvVkK7S4/ldJ+KVLspMyRg0EsHEBypXfDiQZ/tRf8f12C
IDHn18NS3fgInwt10Ay9rNcpJvm8UzgRPfuMEv9PF6pth7b9RzZ6B+yNHqyNhyW0ZiVn0bfiVBsc
CrC+Z/VBUsknRqLvxQ7IwUmiZOE0DuIJzGRGbQHj4HXwdsOOmUNwDcgtlTaZrEg2bnhYDdYrIZjX
ZbsP9yZEsKrnlgyyHAxL+ZD3XEDJhK+4oHOlhvTlu1JTXgb6dlimTsGb6EF0mZjfxs54h4zwr8zY
7/qebNcWet7VjTgzNjTc7h0LqnQaVzWp+klXoUSWaok9lfn+U/WUOCzKjcoNuNl6C+crtnuNM9PU
3kyM3K6KeiHTs0NKZBrdzt/ue+7WpLtZheN6LMLbpAB/QuuDE2OhmKL5A94datdiP/SeJoNpafB+
lS1vP8rLOu4+nFf+AGxDIm8AuakFZq+kUb0UkddZi9cvXQh5yqk8wkJVKBI7VF32tZP6hhA67lRT
1u+eKuOXkPobNKXaH+t49p+KWiVe/pDarP3+U/wRpbPRLyj4ODSlBfxBMkVg+E/Yx7kpIvnrazs6
whgCygnFfk4Tc+2u+DdGu4NXHxWMVUBPJ+RBhHquEKNhRctgeZnG3rAf+pGTpk4SNRxYAX/z4brk
5/EDYDM4Z6nOMjpUFyrHcJbwxxsdGhQz7074BT8epcwHL4/WWciSI8jsCRse1p/wYMgZOam8QRUZ
p69ETWp73NBPWYZS9o0IBUW3ZgVh1Zho1fyPJbNPKvBsStU7Rjrjq6/SpyOT5vyH0P1+QuOP6h31
IP0ubKj2KbzweTKVnz1Q8xOtBpRii8OhzhCOgYkdqoEL8jeh2WBRMuQxKwe5xwFMGqEgjGQqRw+p
HDDCZh7Lg83+xJX5yBOwYRiw27bTPJfegvVWs46kLrSmfurtxY2h93quORram0okgAPOMpeWWWYg
0iDPn4XrILWxdMEga3D9SaOV8M6gmIGDlgXcBvbUwH5+YmMaQt8hBzV9lx9+osNV44fmX0t2zh1T
IF9Of2KX98CjIFLb92sPG0OKIFIiQaRt8kUyfnLh8EmRMk5tXGqoOBlpE6UUKAR02aIF4w4CxusR
rlQZOCQLwFlL5h8QSByVi86YuuGk0iS8+6KGW5GnvRouW1C/BxXdPpB/tFfSGuIyASRkHdgEsNIC
EwXsSbm22v6i5IPTiMjlJ54FLyOhpW5jlyjpIYIUgc+WzEDQBVPHBFQaFjEv314DAQOAzH1FAWCG
C6MjOq9mpL1OhlLXneZdfW7iEFhTYcdFRSCzt9R1nzmGqf2JAOG1BaYJHLWMnF84y/31eV0RjB2z
bAHV4hLsH+a+VUnOc+etuTADajvpXvfcUgzayYIFIV+cBIG/n9gESC4kQ+JqDkSZCaFQS7tofk57
+ahCnszMCaVOUS6faxciSvmVe4hSsXM+YcD8p+90vuS48U4b0QZ5WjZIgRu1eB779SJ6/XFfBNgb
AttA29D8Ss/fN7VG3nki9QeYGgpC5o315qv+sRqtWI+5J1C2e5NHmoS01Ux9354DyHHyyEsCjhie
4I4/jR3t0crkhy8ZArT3ix8Od6VVRAdcxniB6iQwM3smi9NzycWY2lVoYN5eYUKTeVGHaINOYZmi
kd+9zbMHr7HlLXrJSWdDAJwcZd3Q48Vs4dXWAPBc1fU4Rl07VDzSM8K1MQazxogODVx0lPf8Bs1/
c1qk/NsnAE6EPc63q73u0liDcIFhtt/5ps6pGa666yGDjofcfx6boUk/LNL/3r5UfmCXYSCEifhQ
XlSerbiEU6aZFHLcr82J6qEMoFZydK0N+N7STaYj4VC8fK+vlXvxIn7QPOX/nzl7fEvdQ/nytrYK
6ch87UGhZZNJRpAZeV/PjD+sWNH77ZRdmicmeTBHaUYuONWGEp6wBJViShq5qtjAQGCPQxjfY+Mk
2toHn1SdVE26mEh/+2P5n4v+ICcZkzq2oBuUnsZvksVlwbziHxzPT5IasLgtJTVdKkxmzwDxNeUw
7fp9aag1Q7dwVnklW8GcbHk6d1Ik1cECx2r/arl3V2LdZwhb6gu02yRxZzek2JAscsvchE1XCZKz
hEd22SIrESZo67pygvWZuzD+2ngnlZmsXozK4m2fCctZADOaFtPNEv1zecAul7Dmx7jK2tsIbWU4
86bpzkCYAj+t58/1/IiYLxQb9UvHotNZgUypLEKcadTc9gRXhijmByvPN/+QKDOfjbnuLOGQjT1R
XXHrUY7RtqKthouhezKTant54DEw7Q8s45INv3qr6nZGvgbu5uRHEqluB4kDs+dqNbsUjb00iU1K
ope8L+e5blUCIC3Pc8zX65o/clEfIbosdiWX5al4Sw83tUdWAKTgx5L/SBOwAbq1lp5oDFsK/Xpu
StHjaH0QBMGW/K7H8iLAh1zj5y/vKpamV/EpTnixF1z50FRRWP/SQ+x830YkaBb81JLKy6fjJB9z
IJ/SygwT51H0khS3BlQjuS2zKA8cB99GV6ZzHtbfSTcGLU1J434qUZAbnrJeDqWyaNWk/gO191CD
tIHrD91KIxZU5Ek+wk7L1j7fNVobNyMjA/j2RrVTZ3a7qNlfBZ/WFgIzgJst4qpE9SZvIt3NXEYF
Nqzhab37WWhF8n7Pvy/3M1p8IpkAbYav//jk3mDFuwUQWWI5IJx3hl17YGEKrGovu7cCoAeC1whq
yw4LBolFCVk+WuBuOICpjSPjkbYuiOinVbWjyWrK4kazFchGEet9G9P93vdZu5NNvtoG+bEzW96Y
5Dcg21tAnk6Xg2Xp68awqrcffk3Ril0qq7cOGaraOYUZvXRPe3xtMzuzrWco4eO6w6leWJkh34ZN
OtyaooInye4wvAcv6tEyEdZLdOUhI5/xoZojzKmlJimaO5AEUbLBSk5RUwDaMfRizV7FBvuZb8++
fwQQOc1fbdem4ZBkPHpEo54pYvmGp4pj9GhB2v4xpQcX3qwr759Wr0Q3AbiGRC7N2r8HXOg0X2Oc
Pd+LijLNQ9bSrIR+7643uG2j9XZ3ZcoGWRW/oY0ryGtn5q4G5AirNcqiaxKJahq/Jr3qTu6ZYK5v
0zejOzoRU/RCxoQ5cNAeYofAp+4K47UZBXnqfeDqW+aXMSpeo+z7qEsdk7ukYvwFBw+0GYmxlkaf
+7LwJzNse+/H4Csscc3GiG1ZIN2JHqpEPnpI7Wq48rfgSEgthrbGTpOyJWJJJQE36fVWOX6DUceM
PnWvjSnaQJ134UA5Ds/NodiLCoe4xMLDyBIVboy46XN04HKZBaqz9SsJMZoB/wkhy4nqNEsR0scT
0ew4fthfR99vYj9Ur+jYlfSesPb+HdfVw7emUh2DMiiiLYv0e7BX4aySd2tXjKTqH2U4xc3bdV88
YZ3m0/H9D21kIEEdpqs2W/wB+mVwrcnjVUUGjAoiZgJF+QyHornC82YuFMuf4dxgHsw5VU9M3PIr
QFOJiomlDGotd2lkMZ7+uXqu/vZYTsHE6Ce7cZcq7kHK8JqiYGMxqRvpWDTfElF2tKh4Dv2NtdfN
Ukuv8nyhwag7lgo/4W3xxivXMxgS5HwMi6+UV45NNqA5d9fAx26Nmu0HkeH2a3vp05JXMGmcLhUE
KiBNFn3Ko+zJKpDNx463Kfxeod8040OmHyQGB7MQDIrR3p4HD/zSRaAD6op9ygyMtXcid2I4Yvxq
PlIRZnvi8Xix7GMoh0AqqubCkNCa0LnGc3YV/ayKO4gHWxnYpLemNsVHVgrx9YvKM0W7aA3J2o4b
j5TfJaTOWlzK5qWt5kPDf2Es3+2tn0FfpSL3+q+BADb8Q7BP6zbK/lBEQb4+r+DWcTUwYeUK4vvE
WWuCZLJnE//FxIDxJixscJDyOODVmzjzhk2FYuoO2LdQCog9XzMgEMkydDSzdNTIe/lai57UU0C2
rdhYW1dDdoqqK6eO+bXtLj+a8Ikg9JMMZn5sqVB/XYCFSOCVwTroCNqf+nTjD0Cad97UG5kAzclL
kY6V53vJvgaVBSCV3cj+Nztf3wDz9OtFMceoubw8vU0T5lhwMrZ+ViYseMijoapYBFfIf8i0sG3Q
fL5H3HJZXiZVGf2HcKYrEMGLV6vim24GVDufCnaGp5rZD5fbZri7h4Rf84PEKHk56Da/3iDl5nuB
HPTTAli8rGh7l1ZxvXiZNMPRehHZKqT57hiOzORHPySGFoiMl431yxO3I7GESQbadhhk2g3L5Ecv
0eJ6peztvKBzxqOu3YDIHpC9yiIxdf+j8h6nyafXi6Z/R54TomHtU+0INTfCY4zZpFb7kV8z0xx/
1RFFGxgPGcjcGzQ+QQ/xbZQoiniqh2DHr0hXkUrrVgzT2fUkJSmY0zAtErLfboLW0U62Hm2ZDHkd
Hl+i7mG2Qee8N/4Dygz7dgt0++SG9ug9hC6w5pH+KrDLnNf+zKjeQgC4joKC1AQLnIk1xEG+CBh/
E57Tz7GAXTA8Qjtmn0xiO3Z7dQAuiUI6HCD5zaJMhcf9QMYL+zDmkZTGK0j2HtRgmp+dwS+PoLdR
pgn41kksUODd1RN0A4o6/uO1STbp9ctgmHeS0XjQhIiOABESnoCe7tfEb8C0uFAX5k2BU67eBvO0
NrAsIwvfjbX13rE94uvo8lCBufntoDL/fvx3AfWRjjcOn6zohCR7VGH6KTbjeFpfSENybf0yXuML
TAyu+HVhHkunYhLN0LH6RdFyBg1Kplgce+V20eMBjgvFu0bvnSAAnVg56lOiEjD1/SylLbN8KGBc
bUmgISK1dLsJJHU0YPuaA+sYN2FX35T/RxD2zHEiF5DhN+2vQtktwz036vdGT0tH4Hyl+Lxf7NZK
E67V9qnDnx5pwb+C+9BdEZ0RyL8WlrN86C/HaltfuWy2+isXVA53u1u3MqtdWM5UqRdybb9WvbvJ
b8+9/ABNYgz1mg95kspolgVDW+T5cnLALeSYMetkGAX8z+lxWKF0fkDyKfMP87123q/KHIg8+RRy
l6czlYLqQzVrZZbpoV1Ln4cOaQ4f96gNqmHZGiqOUFCRMGAFKbZFvJ10QMwnz39a1O6HTG+YJh1E
94LXCp5AB/MYuKPKDDtc1fsOetF2L9eQ1+qQcJ6HC1HcP1nSu1FxXYbAhyC0J9/twCbDeAA+Z9Qm
AfhrpOmqvrHK7VkoNg/i+JGsCIndKgul7VdW9QphFo3QdCjoTPhBIb9lrSE55ozjsrwqtozoizO2
RQ48+0bgV9BCQlGD5Yz3nw6h2uO8cm6cPXcE7lP8wZrzwcFZCU33bQLejten3VPNSkE+CeILzSdz
5kr14GEZBqCKCN6zIzurZpIEKSCdB4rTaOtXiOz/jG1UXc3Hk1xmHNIb+v9xpJAcH198v+Uzi07o
on+hGGuv586PkOdvWi3D5Hq0cJxPCxyo7iOd2QK4MDkDa8aW0r3ioY7hw7QOBna1Oo5C3Ol5sJYl
7fp6yIZX0RovSaAw3B+YVk/aHZohpP22+Hmzt3s/TQxIIJJQHX/jhJ8+fjxDTPZngCCft0q54DRx
NMBwWOZx9fsHsSmb6tTHFf0hCNH0tT5yJeWywp+4wlfaUv3sxq85goUxP89YAQR208W2wtKqpwIa
LlhFcWOz4d7NmNk2iMbsSLM06CqV32e3vJb4zx+Q9JmyhpcRXfLN4kwUETCStv9IDpeAE40mMXMf
fNKu4uFA0lcQEVpohQceyG9MKHbxObSFpm1n8+Sj2ZspOPuwxClohOFemnrZyPSoVuSfffQG9m3S
T7YHFIwlxlCJ0Zx+ql3xmdYmuDK43nZf2YcHph4v2tAWUbsIU2hu6nxXj/6QTAJPIf0ehEdbqmO7
8vUro8cfuXw3NO97ZdAt2vZbo4djuhtALejFWfkVJkU95cLjvWKOkwTM2GuzNrtb6plHciFQKwCs
cujyabOOPB4vF7Gl8C6svuxVcymp2HMTcIR+s+sIoi5sHP0ng1AchfAzRK+jY9bS205usGVLMPDb
RX4+PCZSXYsZz9QEwIYaMcUwsOmXT/xbGErggxR6ASXsLqEkHtNR7cmizDa/jtQ+xf0xomkQl3Vh
2S0hPmH2DrMugwmjGMeyZA0Ah5Vr8SgEEu118LTO0eDMc4dKdZhZTXrHyzU1b++ujIC84f8zNdqZ
SblW1ffdOqlQ3NAs+7E2RsTmGHlfkBcaWq0ivIsUMRfHgcbPVajd0FpSkuwnM25NpGtuHs924+2J
t91hMb/dTB1stPaEj4rbiBPOe2XxymyyQ0c6ZulZoMTo8kagmRJkMASgmBDw0OcoGyyeUl9NPzaI
8ADWgqEBTi+Fn8SfEmpzFE8iGbXif8Sf3GYCdf8ERM/fkbhlpwaoDrki34tAOP2RiFGjE0bmmPuM
u7CVcxv0aX+zKWny5/xRTrFrPGZXIj7zhnubXH/zbi9bDAqBi/stUB4DnhblOf52GcLOC1XsbPJy
RgcKSOIaCA1vQg5cXN3vmKjytAPJ8OO8p6XTkWA62xtv5/M6XFQVsnMr0+CHmEgT9K58wtBar0CG
CGlZVAZR0attG28DhFwwGUk/DL+mvdQPdKYN5+83GwlFCx1sU9MvJWlhWqQyPDaG9Z0TmTKWKGma
EzH9MpLFGqQWdr4SzyDGG6uB0e2oRaCHe33oLrMIr08GRJEO2ttygzBjHzYK8sWNv+Dnjvb75zKv
Dhy/OfZCuNOaIz5DAKxol+4L9V7vWKjMXWpOyuKl0Emozrw7mdK18SU/W93IlKQZmBCvVafyRwuy
DR6OdDouzui2j1CAWjiDThx6RiprxtjD2X3NJvwopM/knbCbVnubdcnFq2Yd6D7gWgsKkMLLSpg7
50z4Ntecvb+2XQxqR+i/Bo8i3lr45AKjWCGz/liAysQc19GxiFkNQgHzidqZXiVspIo7F68JX3yX
yBWf9erMg3kzUNoyGOi0++mT1X1Y/2R3Zk+zUXy6ckLFZgaZbnteFsOZC9GAIk22GMozl0jiG5QD
WgXLJcRygr182bemh3tMg7BxNKTfCvFQgVPP0Nv/SeGBzAu9oR//LpT94ijJXOPGsGQBDqsMjeRO
f5mhjEsqYFpvdlWLD3LOEONqpJVLmjYi6RNT1B17WhWaKoFn+nACFP7K205ctwLo9sXpHI8xOMe2
aVQ9y2WT41AMIAH12mC5zhEazaFC3/htHLSAbrY6EJ5n9fldVkViFlV2dy5Q7K7VCZdvGWTGGp9t
rwLfnwOZGkw6iO5F541eX04V+m8cR3E4MAEMfYi5toVbM3fP+zgwmPSVA3gfzQwrA3xQtkfJVSok
vkmc22HRrNwQEXWXoB0XtlSqmRDtbjUu5tiwCfR1Kykc6bIjQk0kp+tUFCfqwuaQsyyvIfDEMezq
9tZC4Yz5dPO7k61fOKV+XcaU2FWY/rN/H5+hmbpqCJ2c7KW0+ijn3TvKC7uLS3GsNBbUuAgT1mM7
EGUq/cARKar9JQrmeiIPT2jWX+75V6RkdLf3AJrQynMFSJCN5FPS49IJ0IcRZ4VWkACyOCohCOyX
sGBQz0ofJpwJQ+TU/OP5Yv/vjaZWdiNOg2B2hbw0KB10MoTQcYTJGBymCfRYdNmulPj6QJVoT+U5
FgYjqBr1ET/eZDYwn7m0dKyHA3ihUjYo8qjGhxIckZ1SErILnobfdbmQ9hCebzkRF8al8Y1Tqc/S
UBWyQ4Nt4EP6sZKxWGUNOlJ7YVploNLO1aFs6gFNZr8oiqO/YhQTC/bVPzpge+GE9kEJuBl5GdzR
MwcmIEFyzFfHI3rN7sryEz5QbMsnaChabCmUAe4w/eR//Z7VFD2xOyUExJD4Q5xglsccl7YGRAWi
LbC3dPi5XK+nqka2gGHPzF4zMDvBSGd1MoBhSAZ/U+p5Mp5gAd0pEk7G9xb3Jl2RqBhJouwyyPIY
Dy13znQtzfXkik/v29nrcLM8xwQd/HCTHPGdsNg93CEiMILWwrtCdpFexgmrPqnqwWw/WHU5aU+X
EKNnsmkbrorWgzHcjPyK1aV0hGvM/fW0IaCTfgEJHlHDK6W17jsNR38vbhr2P8aXIq+T4MxP5rBV
KxTvka/PxVAtUzLonZsB3M2UE7NTqSlmqBvCBPgefj9KbGMRTIlCblRUNFBiowTxfzEHWlZ5cOeO
KwGqgGkWDUBiA4/wsbRoJtM4wBoEXXgMGf1l+o8GZ650xTKWUVmGpWt65F87A1XCgUMMjZOXt5VD
QFbSBQ/EOL7nHPA8UYf6xF4q4fOv/9H0Bcohccn4QvwsNauPnzRh5B4gw4lqzJ1EuV+Ovsv+To9S
zNnApB4gbSMo3kIqdsz3uJbTrSRSTQxLAXoAFA8hwfcTP/ci9lRzGdTnax9e74jByvjeqMKjvdG3
KmcWyhl6fJRZogGIqQVoTp/s0QPaVzmxrHSC2sPykrElZsSea1s8t+5vlEoeIbYnONu6x7Yd8wJz
2nHUn4b5FsIf5lX8NEnZKpsMDPl1K0n47QIofFDMS6sm7LFJJ5ZX+3/zBEPmPAsUIonu3t9gdUC0
nfui/ZLKE6HMALymmCjbE3j0n4/hPRZgYB123cVpUKOuPKMyhVqXo/g7QmCnTpZUr2dd13wNZPbE
IdeY6pdF2CsfKUFE7sWDSs6hBiEfbsVbUOfo++ngk/8B3i9B8zMfVM+doZ71haO89+K4d0Dp49+Q
/WbgtsfWCPzF5YSe+f3EYDTQrgsXAttToKkNVqzRm/GI0Up9xasDvc1uVj2E9L0lS+RKtifnvkMn
MYqr9FiHW5LLFzOwnOyNXxIY2uzcqRAug5Ng+1wH0lUQxYDEDqgCty1PUs631hHPZOCvjZkXN0GB
i29fQAhGTX/guhMNnuQTbhERlqLymQ1FZncSm3MzY+cHgJkKKd6gwVaYO+WM54q5sIA+FI8AxqIS
1lY3T1xRqyXcMvWyYw6fciLMFLgFgcLYw3ao7QryO9Hm3tFmwYCGHbiguevf3UUrfWZVSBchVxhd
Uz7P6TuJFQeIXFFu0IlIhhi9JTWVBRS+E0Yo6FSVKyM/2ae0nCdOy3CpdoRfDcOSVXFNaa1Ti/UN
4I4c4rpgK2CS9G43bK56FkfoHvZbB3tAAtRHq2HC7RXWbn2SjvFjI5lY+/Z7BHUKXlpxjzIESnBB
f7sqaZedn8lpk8WMqZ8vcnNEZ/EMVXShcHymW8DuUblG6fN/QZCQ5ykDi+WNNu/sEJGXiJj6cYuS
mgaTLgz84eBv+CUN/oaS8o79LdEDxyJkE4GaLxmycxH0/UNEHwRbS8uMqSwH2COt0KNnO8Is+Y2P
mvfqhMaDzv/TmvWEqF+4rz5kwLMfN3YbBDHdLX8fVpz8G+LUk+rCdUQDQg+rYeMe2frHDiGB36Sj
cj8e96WC9ZQae0IPun0Vod8Kvhz6G8OXMeTZPknpx6R90cJ2pdkYU6DuMA/tBnHAB8tc5Knzbw4C
oF5t/E6jpRVfWfLp4g3HM6+yaVfbHHpxqTdVHc7jQoQxd/1mE4f1Co+Q7BiLK8jKq+4VRK8oSevg
fVGuNVcGXo1WK1Hi0xyOK6uvcIU0sPXsQ6VsYggArWUnqAFo3Svu7IMN/MMoVk9W1DL0Tt7QicBc
6/O2jhgNGgWZmj3O+oCCm/4yD0hVSRWzI5KQC+vk7IUCz9LVi+BApmWcyVnPAZqT2+qAYZCVaZHM
SaZXo5hxQQ3oTwMdVmknQ2eu97dWCVrEU8VJprJIoMzlgi8bdhiuzhfeYqtJYoDnIzxCI/9ZNt/a
cOBZVYeLoycOCbN3NsLppJEQ5dI4haXSYLS3lfRhUHd6nAy/pnoum/X0lXYKZJtj0K34f4Bld5AM
YqykfcsfAV+dSQjFxFbQEvs3KEsYVARTKIOKavPmcsT4YzOY/fdBrfeXdp/chdwmE4pLC6MxuxDS
hbz8VvRirIgVJpnfGuY1ynR82Smex4rEiP8k7dCmkfnwtp3+nxTmFQ14Dzs+pNrWZIhKp0XadHB2
uw3SghJNWPWjezE4mYMUaTsT6tN+R7E+oBLdMvxEQX3QmMz0Nd2/4tuFEor+Gx4NucmPnsn76Yeh
EYiGipISYj2dqdlK7Fz6CmCyZvFMlGJoFKLoLBgIJ7xsuSTCtkTlPuw4RxyDOFWlVxaN8QU+OsvW
Oqj6QH7bnOJ16IKXgsajOeHpFlQefPOSeecTludPemMdq+Oso+E6l9MmC/GN4kPT/Vh2H8bg3014
8ZkqNYAw6WY1dOqPJS1xuIIj8t1jb5bGQy74YV3GyJFWuE+byk8QjqKkbeLm4tOO09aIFi+V9ffQ
sKi44HXvEYA1nInyqtjX7E73qfd5YE1FnDNfQmkaZNIa7qya2t8heSQwBs/BIhQ4dXXOyU7+3ROr
+HtUUQfC54XkUpJDnBR5DSkl4UZAJLcCbSDXevMVONtVLcHPpY48d4T4H37Ye3NUFuNOkcCPwbdC
TGQgwYnOgwlZWshahUOrPV3o08CmWL9XvTW3rD7edzVZy3l1Dx5ARh4q3fJjSLyJvkCAPC1m+Oun
pX/v+S2/tKYmBMhzGLXFZm3TKAN82NIE+v5R5xmMUp+4CvUBq2XSCbrnJjKRiCFAXyfXck4Xrnzp
CIKWi4gNatuzSn6o0Pp3V2xf2aYGY8IfVgvAHf8oIKJLOaADNXwVFwjiPl9D3pxR6f8zsXhxoCp6
kHpVIQ+0sy0Afoy3U3Cjw1FAjk9FuZ6M9BPB3/ao4ZP/FNyFstu4HZVZxpfD07ttBEDdwMRGKCnT
hPDLsPc3p7AYsEynR/nvtdg0HP6yXBCiS31fF51y/hQhDl93Gd/G49hdn4qkZau6UuNhYItpXyi+
47D8F7d3YyezxNnJqPPLVXRBGZXsshalIrPCSrCrtXqAufzliqN+iPXt6pOlfvy4vURSqubfyM9q
GLNHrbJH9vmRFuNasYzRRwF8BNWlqXp5z9GJDolQnVM6X/weMSY5Rri8pnH6LsO2Yk1smiY0Q1vx
iNuaZV2g1yw911UO+jswv+qJEn1FUxSyBtDoomDYoEP9IUPshaC1mcUrdS+kz4huLrCcaTf9sQGZ
Obh8Bsv2BvMv41ZCA7Vp8mlFz5Z69hQ++IIcqNZ8VpeBoOfrz5Y8FJA2qppqvviziLwpaDkO37G1
nikLyIQQanjXPmysZUr0DY7dYZrmZXlj4g7DtHrx/xMOYjjsZIylTjp0IIQs2/HIaTVT3Ujak+2u
uxKexzrClwP3/aXwMNI/o3crpkiwrG9AVtz5mmkLo7F0Olw3iTn4/vwbqHn3t0zSIgmta/hqOXsk
BefPUIhJSKYp+sM0Rb94oDSVQeqgQ+U0b+Ypz3+kazFRGNyTFRCQX+smmAuOQst6daktOwNQb0wN
3RLN82/T3qJx0C4d3IfTo2Y0m/lRNV3BCuq2SDkCdexT65a1u3gKpfXhRbwC24ApvddvWWyFsK6w
M9VFtKiVa3Qwf9WMisnv8oC1KTWsQSW0h3phQCNDQU85eVoenlyxALvmze4MPAbFYp3OkNz3kpM5
o84XRQh+NUaSSw+CcA7V9cslYkEHorInWMLzh4RFEPGmNd4ouiiwOFfuU4xZaXs72MRR5Jnb4Vy7
wWMTpQFfpGeHcWP/0cvWRtl8DI/uvFGkBy+XnNSbEI2dtOXs0oq2NPK7MNwsK1V9N2B2Fo+jYl2Q
qXHMbhS84wy97r9bFpWh4KLcRjYrf8XSW9QzeOvaz4UnXXP0H3uBnObcBSNbhGNo1IoKQuw2el0W
RIm/9K0pQWnD/0htlAM/yP6GDCHnsLe2T60FgUeh/D1Qtq4kiejirB05itCq0dKrDOinZZFcAhT9
aXS/nJbfIBwNqzoio0Q9EjfdglG4xHT0x7LMq1OcBwoUW8Q8lywDVBKWArPAB1OLD9nwNGkZiqDI
WCiGzFlWMrGn0NOMeWYB84SUDbomErnzxYPgZJ8YkwbZuTiyPkJN2N7H+IRl5iwuejssHITUB1k5
GjorkRaRpXTIfwNijg21r6rEIShZsxi2w/3Yf01tlsgLVLu8mUXFowpe93h7NhYGFE9TFpoTuic8
TyAraJ5MI75NqKvIWYQpLYnDGPJMmbt7rukDe1Qk95JgZGJNH8lRZO1HHyxVLx+NNPSXs5p4aj97
qbCuNvfAu5znAU60JYKCEbU1cfOSWoH+86uUtwIX9Kakd34hXo1EiCOedpEx7eYeyyyMah12Xyzl
BTm1DFrqSI7c2oX9XMJ8v+aqJj74ltHoD7UwcIG9OO7es445UBhM+dlPgz1arBndMgGm3VwvJmgD
4Xlfv3TKUeUTo2ppK67+ogSdBqB1gtia6ab3KkEexrdvfCtXLJgtzPvm6vS7WAR4/urHQBSVmTz1
+wi9fSBp7yYFPBkNlz+m7ojBzQQGuXMD+EzMTfJlkFuBrsgVaXshnKOAq8KCw2S0ifhbb2vTclHp
os15zT7RqXWcy9FzAzlFyuHYCasON7b+DuA7J94wdEL2wm26El6r7J7q7Mxv4w+CgRmXDBPy806U
NwUAcVUx3R514zhU2UO6Rd7DOejR74ot7NSa78CYco8eB79bySY5ge4NCF6z27qCVxj6USCNLFJM
dGGvjdmjm3cQP9Sy6r7fPA2bNKP2MAtn5WG28lCECkCHhIs9hQri+qwTL6yP8DZLRbZPwoSG9yNK
fIU4TtBIPDGgDwBD1nHSC5qj8dh12V4dnuq29vBLyYHLJ48ll6MBVR6ITuj2Xzexm98jPiu5AzJD
reiYwzEzpUtRqiKnPJh4ihVI8vcY1AXiSLSeCj6N7Em1tDWIPxNxs7d4lCoI56W4aCpc/AP2V0eX
/HL6j3kMPMCQ0xmAFK82rbfOcb94o3vI2/YEzL6kHUbs0vqo27PhdpPQYyRPhiECgzIT0TorPOlQ
bachukaFoyAbAXLEksBpjaniN/+h+Vxf9xfYgvijV8FdDgRJ1YhrHOxaElXN0aLcUmCDChZANFEh
JPE8Dg4q4GRVvOPL6nbF+Owav8dXYN+RYlcan2tnVEEtuxXdQpRa5XcymCn8ULu/sG1Apx1Y1uCX
MDNXX/DoJTU0Or0sxgc+HPVJql6UiPWS1ygkCD2vynZC7ym5AnudbDkH3VDtcGmx02NuYh3xXRBe
xWR3BQKbLckqy2fMT3i8r74/PErnv7KYOhqD9Nm/t6GnG1qFx1DU2XJ7U3VUDDRJ6A+anzaLFj9i
ZGQttoBl0bwq0w90ARYrVoQXF3jTWY3KkbEtlHvjsPa9aLyWg9D+zqnAXoOuqwE20q93FR1zXLm4
OXfF/TSZYJOalFDpWJ0b7lr4JUqlT2EDUhSoVAP+R7SEckVo5PgFNlx0ZzUoMLLX5LDUBjrZpm41
Q6PDIYvFdUvY0hRcsIIUZr7fzOwBjj/g6f/iqZkU53bVfq8kpLmlKZWi0hgY+qEEyoxrwFjx8vva
LnrHwXmpOnVaCj4aE8neSUpDllS/UBR1Tf94rkLpANPcwtCwiaU+8m8cRf9erP2A8zQvYaXPhrZ4
3uoLtnc4bh2FJen5tFY4NQIpksksC8i6LZJP9NL9f0qWMVNTPh0QnAPt62kl5g05cxVHZfcFMsEh
PjMKQBWHJvb/I4F+eN3B3nSe/RMdqy+B2bMJm7ACoPx+c/8haCGO/3apZWEDwKYp/AneUej2kgah
MLcu+7CaZPN7UbFgEfY50k+eWzDeBfB6Gb4RGF5LfbcksR4M8D337BwDW/JvwlGbh0sP5mgV0BS7
U6+KcQ1XuniCkKRzQ1tF0ralXTr0NoKvHtynSSLWSRBYYA3sizgoC33Hsvbf+bbg2eGG0RjGKoGs
3oHIByYjRkDP4u1AtoOHLyg/cvdFY3MsBUil9584JlAQtdElmNq4DWFeuncHKbCWOK4U9/qFHbEa
xljaXx9WTeD7hrvF6iBLlchYtbJjUsKrrDF9KquO4KXvFJUAZuv6B1zNj7Uj03Jyr0yWGuoS+XMB
lW+aH5a8ChqyUG/6u74xU59vIqzJZ2lwyCzJOUQ72GmZwmu4tXjduccj5Zrp9ESJGqLYV0EMLOqM
oqCATZYEtnkcv6qRgKxcVCRQZW3HeKwS/C7MxEiCssHjn1B5Q5WlKRXBNIR2X+HUkRMi8iQBpNGo
2W+lM8dP5R9V8qy9ffpknEUFKsumiwzeJcgBWL9clHQWQNWQvFtoP0C/YE2wxXE+jmz0TBB4LDdj
KlpPzuPn89Xl63YsBo69fa/AJGDzutffR1E6qBSyA8ZIY3ePPzpJ/P9hSou5T9gCX2bSWia+WIbX
iim+hG488/PrlFpkKo4gBxOYbsklbJKZD+/qSF3Pcrx/ru4en8YO3B8AjW+RWQ+KuhyKGeU9/M1L
R9M2XnEI1ucCLl00wsW13X6Tw2TAGfl1c3TeKy3zClFm//Qbo2rl3eX9mfkvjx10Ek0i89MQ0QG7
t5GkDrSWD32TX9TxSCoNutMNkgRak8yBcSLOk31Yg2n4H0Gd8wYT4+ZwbP0q7Vr1nQaVknAi3kXA
JoRuwiwTTa0rRP87defr9glVM6H9jC3dWkFZvRyhMq1vGgQNc46f4j1LL4w9Bc90BkKzVRm5m27c
fhG9WiYr1xohh9odMMyMJs+l+zS5F7yA1ff9psiGY06/u0zaK8ljFpkJikaErpHcKIBchP2ENOSm
NSM1Q5mYgc9mL2Zt0tajvgnJJPLk1qowMbOYk1vAkYLdvsEwBtTlo31oJTcF41VmCphxlodUV4U1
N4Apg0lK9abnGY/qHvOkY4IUBmixzDhBL2q+wZY0294VGl5MgIYt9p3BJH75IE+ZohWHbGQeAk5/
LOwgkS6dvGjTMIuaIv2qJblckpabuZO5DvXXVyQkCD6loK3nwJTawZos7YUc0g30bOGWi0DIpm0M
wyuCVSVdAk09XAivWhFe3RTwEAsgWiXgJm8GiHiMrLxjCDFOF5YMoWUeqUWeNZoRMXSGONbpXlHo
6vGZI+6KS4tTCaIUhu6eyIQuCn9MOGwGKoTXKl2cR/fLOH5XNPXrTCeOpdb461UZquzLE/hlrnV1
UA5uq0ye9Xv4BuXhaQxQ9gr0Xp1M8yBwz/AS+O6PE1F7YSGHD5rZNorqbJ41T3qQOsf72566Vi89
FngZea3vD8Gjf5zlDTumxrCwVjbkBofPdK2A+YYx9cKqEdKrRcbrACI+iGN4vib/GLrru0W2f0po
MEtyKHWxEgtyG2mkkq4Gn0uR6p3UwnE5tCOIBo2+nu+mRKeDqsgYkBGEz1tRp+vsKB8Hg3eKRNX4
jMXQm8hqs5dn7iCHpS73/ZmhAXcQvrpq5CmDNNDClgPBaX8wO5OeNwduGHQcF/6VLtC+v/dZ+D3b
6Xoqk/JIndPJAc6XVm7CMc6OLC0eWgoItNDU9tDYF5xBIn2lEyv1FHUyXnMMK73gT9H4dMl6z9Hk
D/QLI6IcSR7+TI34sUFD+8/RZ65EH87E8S3HxWOeO54A4quPuIST13uWiKi2YadzULvpKCjMatYP
EmERer2cm7/nLo9d4Fm0PPz0XF74rZQFwaTpvr8nC7DHUmaewSuOFDnLDDYRGZAqZXvwv+OEK/tM
heQz6wsXOBJsM8Wd9olSGOE8zEDPhfJgwaj+BjRTamkxqR6CEgPei/SdunIxA5qTaY3sXRzT6gTG
CdRKMmG8qAmPAXgTEYbnExWyCUhbcGedmrSnuIwgHHKf7WDGMVUeDx/Cy4VNOLobKntkKpTcLEFV
NAnwjLzK9oNmwXbW6UuOvpgeSUmWvm6/mzKamnj5Fn/5OChwU2JkGg3wlGUU7hI5hO1goQ+e2OYv
lNmfLIwSxAO60wvzGFkhJP31uPzGd+vec+CM/o6QQTe3Xh6NG0cqG4FRnsdeqwdBDZhr4CNWoD4z
grystRbj7V9gx5nPZqLDNgFZnfpjQ0yBYREF4pulsUoJi4SaVUkB+cP6wfC7HJ/34kAYTnwgszRh
rJ9yPlh21ecg6IMVpKcdCfY9VUeshGZN3kJltZmwPwGr24ULLI04NY72cs19TpicTfPfPAGVFnuQ
hF4fThKExw3pR4iw+QofSrg5lRj3wuj/5fHG92HfUcqC0FXB/Btb79mZPWy/Irhj0LEayODoG7ow
jMdIOeFDb8GzaTK2Uw0lwJE54AJZJkykm+NxLGEnsZAEV0lEHGsaBlkKYT0iN2a7791oU4B/iwhp
QjK4zM7NxeCb2tltMAh01mTYsnxCnokVKMk8nLsfIlhJ3FA/LlFCPrMAEeGWuymxY3AFLilR7av/
gdWvgeJRsUvi4MJxilefVXg0LFt3rGRBlGgis57XA1Cmb0XZzBUcGz0vlftRNfxKV9XeIdHwmdKI
sBUOE5+tVocbUnvAZgpikwZROr30E9PhHFEYnEDED1gWYiafpgt8b+dc5uzmhP4Wclsc1DJ+/Gm8
UsarvJ4vKonGVthnRYbWCzioZRdCWJIIULs+/0uFnuPRKu3RBuRm30HxOq2ri28c8ajAgtFYwuCM
MDH3ib4VTkcc0eKNmtTB8VM6IQed+yQ6ty8HqW887U2+ATel3GK9ZWsPWqTIiklS3gn2QcaAlXaS
UYfsd98NnSoiqfJQRfiQ8TB80JlpOwFPQ2+PIVAmvYBpmvLUGVnZWkYEeoWV7LXzCkn/L7f6C0RO
vSRPQiZ13jHmaaxCDMa4uJKg/I6FzOBHa8VWpZpRSPrwKfjx3xW426JNv3DQ/FZf8uGFLxuuQBm3
qfaYiL+p/5dhCBVsa8l37rtCvF8C57E2Lz5P3CGvlmQrm38J7SjDi+a+BKp94+kHBx43okuiqIpK
3wbjRlIgpDHtPM0SK8d0QgFiWksRvdxr9njCVub0IKQucdCRJ1sBYvrsvj7JOKgQv/gULK1aClPI
ZKQK/c2ZW24yrlTK1k3hawPVZNynRvf3LP7cgRvGpzLDRsFyZlYBLNGUe3UlyAkFllevx+RnN/lP
bTAT3vKdthpOrs7KbiIxNjQruBvNcCXjsVRLQ6tVtt9XbLOqq28km2KEP6euCSMgT2NQbwgjgwHh
574DV+FvtojPLWwZwlhS0UfmRATHfAHeqJO3N/4l20TGrk7A0BcDlG73Rd8928Lxr2Cj9OPKJjsJ
voVamnRyBG/zuND4EmnqkZef8qI3tRjbGnrqmMZMI/vGNwqfSOFpLq9Is3dSZPT7E0pfj5MwAuj4
WeVNImvVzKs32TJktA0hX0BvWPsmQIZMXFxhBwQsI9WQRTQKpUJy7hnaAs38lf7dXI5h38AfEdL9
VfijI/zi/DAdKXR4+WbiZ3YRW9U7pmfLzzWma8hU5O9X36UZO9TItPv5ZItrehmGdgGiR/WlXTNI
/bbqGwuJQXPFZRrwpy1WsecgquX6k82mgAkIM2YwIT7C6OooA3Q63jdL1HJzkTvaG4+L4XS9p0qY
37nzWeuCfwhj5fVnr/6d/qR64pgXJRPy+PEFV02Ho45u2MltWqLMJaEEpI6XexL0930kUvbPeJWk
IGsgyP/PHZOzObiKgN5hcSMcYpX0C2oq5a+gH9dYB9Pou9O/pohP9iy4ss9TqBOERGjILYn8JPUR
CCTbcKf5K0n01C7/7sIUtum1MdrIiiaMyQrBoRLKE68JBwaa032YRELcQqjDpOKfEsSB4RZXor9K
AW1V7tooL9FSmnPsw3GCOTPwcZHfX6qoxQaALg4nUT0OZ3u7nTLRoTf2R/YUmjtMn8utDxTkKvsG
elIIEWmneGGf3oUL9qCe5hsFa2U1sVWKJK6xAV73CHI99scH0dbR9UynT2rn2xCLtPw5GmS3w4PJ
eCOlRPxcpuYgXNEmramMcftDcGWso5/sJyBkUhCl3iakvFK8ZT6EQDTL0IlghoaLJKQSgS+mLLbm
aQUp5ZEGybxoC3Myy54+psjxN0z/okUrjNavsD2ejtGWyKfdTgGs3yJ6BgEpqipuNGZpDwF1Dw2t
SYEHLyox2joE/kjKrspQVY4ta9vT8LG/bagMAghiOV+Y82j+r+RaNX+s452y5lo16kjSYu948RMF
KcQdRsOJBdm9IoXdTqiGGJnUuSkqf7J66izAdjMjiH9wESe5e+4Dz7xSWmXwObr96hYjDPsBfa3r
Iah5SoM8pI+CZ6U7EEEpC7NKvuKGWY/7FtAnWnXuLREpmh6WdKy5wyxMKNYrUjCrF7T6LOVTjf6J
1a9xhvNc+SKFlHMnCRMDhRbnkcWT79Ljlx+VnwCfIpSV8s1Pqvd0v/6WRGkte6uK4aKskq6sSSQJ
yOSha8uZXGdABWCyOk5K/31aDpLX0xqP5SsHJerLoaFi5VH13prf4HyrQIkuYBcPC2jw4CIWRowV
+lNVxPwnsI2Dz8FNBjw55mCdGiLnZL36PWwNXj3e27bb3GD8IeHUF4ZCdoxHZ9vNXfI6c2zkmL7o
h8ttmQ8net1ONsfBHRGzY1bbikeo/a0qzG8xOA8r3QjY0Itd8qNVYJG28Io+g726CNOJgX1m5nGB
EU0jStZznfMUAMyVtFxCjxPlc3YmzNcIaKRMznM2cAo5AjtTpMZ5GbF1kU/q2iqBfRGMvm6V1wQ1
oFkqQXNZMZu4sLSy4dHWPiDbgJPL8cZON6Ifmwa1UVDIE/IWh7xk649GIe+9pG7UkRDJsPE+KFLF
LegmIuO/28+sqKK0qQUMZmSJ6y2ao72lbNl13Dw85nWZmp3diX1oM2322ahWcwvDIpQ6CB8Ys5RF
SDujZZh7Ha4GEC5+I6/KYoFQOn+4mKy4EEJsAvouASR3SpDScqfaNoDbB6Yk9dkOoTWcK4YyRSRM
rtN+kbZo0zZGoThJrZgeQUyIf+YDl3dBq1bYcj6KMLWz/9lQL6aCC2Z4EnQ2EXN+toC9L1ZhBVFx
GdkKt92sfZIaVxBpfxmAdER5J/ki+Lj43SdI1sfF5t1SgiaVr3rbHNdpMOhZHQgZ0pJ6peijIIZT
LKpTZwSYwzS/gWRCC3lcaLnscN5my2PR951iLY5kNnAJEDJj455TffN4rMjl0Ea2kWW+v7YPqkUJ
ky8JNDoc7nMj0KvnAOKpDrflT9zF79fGJM+ueyBUWqbJi1PBlEXCDG4MefynzaW9A/ysp7MUHhXJ
hDJ2HePNL+VarVMoDQ1Qipi9ObItZlSmxnePyInv3tRU2YusiYkcu8h6kCmykoid9kaxQ/xxhz9f
0S1bmQKmCxIj9DsMFZGjw9SNOj1dvfxQH8h/NFbRozakqxiiLGcyiOi7P6WFbYKGrtSoSshiImHO
dDSZq5p4i+f1HiWgZ/kb/b6Gob+lsW8XgfW+f09q5cyEj3ti5XQ/0/fjWdn7s819O8ZO6nTexDEO
YbFLxng3IW4/Z7N5t9t6ttaukdYX/W0k2mWQkZyZoAC5z/SPecoQWFCPsU1Q4FnU1bJ3zY1aS0oU
/JnqsohnKttZa7zQ1OiNs+jQRstJs7Bd55kdCL/RBCEO2uwPZmqdVkvysJt2zzNtuGICLo7tdQH/
VecdJJ83dqTLZOmoYKzl7Ab/ottOyOFKq38l1uS2oiVIq0p0+vKD//UlwVsaNqqkn6hkIcTqIeb+
fGKOFslAnZ9lOmtcTevyTiApT9W3TPJnmjthmnK6+POjL4ly3CO4voyR10rp4dGaLzP3pqdP9Xv0
7Z0dFRIum4QRSffDFm+lagSE+xIlU54YTcgZ/nB6mctKRt4KBfk8qFoq+2+3o6DjadR9RuQGynY+
SGlZDrEqLjwzwZyFp4P2Og4ndfhXWnBrvziKF+xuCFmjoeCXNz18GSJwoKhEKboiS8Ec4BJqiNog
yCFXiXJbFfzJ6O5sO49TWEnicKqYW7LYQeURN+NdJ0pVDOimEC7B88NRxv2VYDMq9dU1KQgN7Sjf
io3RjMgw6spuFvr2aABD8Jars6k14kjKcqEQGxAgclTLCPs53RAwLA3CJPTIMOpQmn7BExG81wmj
akTx9q3MF+2Ek4HsidDdtd9pvN23Y/tTfVn0/2n6kdtE+Wd9QUAzY2TDI1HHmOlw8cwgzCW/VWNW
ec1AhvWYh51IS3vsdCrtxSmGi8KhTROWHz28mMCuCOMjPFNMhPrci0Iu6/646aL1dyHwUKs3PLTM
6rD9n3FyKsbjKy0EXJ+3iLTj/TDa6/rsHzTylkYHPBiSv5N+DMSc7b6laadUOuSUaIEM+5PvYk4B
wmpc12M3j97Ngdxa89DyOCM9ou7Xezwp6gT1UPcA+AmJ3l2JmMjtk6NV75Iy78lrCncu0ZsIE12O
KmI1at7RIkE25lNk3MzxgW1eCBuAeRSX68QLm++pIC1cl/5KqvcMdjedC/pcEsvqMvIUOqHSP2Pg
040PKZ20QQZEJFKZeAOI0MPCgglwR/svOu/7Dq43wALjc3PskBeUi4hNuQeKlskA+SzJ5wX8ii4/
IP0vXDYoXjIx/rRRFjqE4+JCMRTfecbYvFYuSXqRPxF0+GpoxDsaRlfNiZ08DkbExDBn2G5iuNBK
3dcdy7v5MpUorQH73cmFOfWpr2EWJ1pHp0tlqIWlX4oNp10M5AocTzsbn0V2tuB9UWTDDXt9aI/z
MwK0ZgTZ9FTWTAcTKO1VtENep7hQxnBBvudOjWwULbznBTkqR83Ss0GZpQKTxdQ+fl+A/WAj2Zru
yqh/PZu8XnBmRvfLla/EnxxqJpxYY9qifRplkc9WC5JmZqEkQMGkS1TyYL0b4V2WtsUxVa4jbOgQ
XHadQGkCgEXWBGGkXjuYKEVJyRWSmFJGq3r7//DXZCyAzVGr8TlyFsQRbh/PeIW8UUVSHLBpARMn
ATf6c+i61vFzra8rd75wY7Tc8s+SLok+KmvEHGr3xRXBG5TYhxVS0FWvhMKQBvLzqDsPcIffI28y
zL29br/xMc4RcsSX1HRRLHyWTRX3mgF+9+H4kzlUAQvfKgqRXKY5mT2vrG/kQNbxLKpaYpb5ltYs
LUx4yPzQFBWUj/l5slin0+GzIpkc0Ww9i1ngdtVWd969Xo5ryAZm05RU9/QVAKVIl5OJ2ni43Gfv
DhrlAkLUAV4oD/jbPdXEO0dHWR67n9+H+df8Y7G6ftrLM4wn9HVUwJHRniIFdrGw1acI+d5+jcXe
rSlPCw8uFopLwFMkrz9tXg4IDM9y3NtY8Kukt59jCEYUfV5OFeVTnUizUf/RM5utZ+LZvnCSwB6s
+OXY1LgBJYeM6LOdat9dzpxLwONmRZHPH/5v1t7PeilUhMykxlAuGrgh81TxmtYBlRVtqXLj8C/z
9/0mdyPC55a6zDGzID71Fv41hwjWiI1vxBoO0UomvEtTzf0RNXzw3RJ80Uh/uG1uqMCmJ68swoR+
0wog+HbYHOW6S+rDUU/fHy5ou1orvPM07+GYavcBF6Ds2ySOEdkwXRvr4vCivNGDXKKws/HHdOH2
T6qz0VnHfOXVEnFVGQZBF+b2Uu+mrC9FhVHFgkd4DUSNEgVE+OlM9iKljpIeaqiGHIOF7PqLjU2X
RfkOe/hx7n5EmLs93m/AwwaelSClwNUsOC8NiU2G/7rO095QNxtEkJJXE89gFYtTnY26vkaB+dyS
ZnLTAymrcQ3qN+S0nYsK/QIYk5xrb6yVuZSPliF245vpm2OF+MGRaRIzF4pcf7QQG4hdrSLoLzop
XsXwrrMysY7Vw7UNm7jpv8uNMWU3VSDGOSDz2GQwN0LU28OlGudiANnalJ3eTRN6M5PQowTiPIeo
fKODyUdbNBvW+XNJtSWLaXgeC+hV9md6AXsUPt1vhLNkEFHVl6xjfyoYytOvqCotDL1UCo3FKYPl
AcAPwwZUyonwKDKmuN4e+q74qZKKXQLTi8rEHmtgWvMjjQVqlJ7+fNuuDvR1IRyC2NZ673PGj370
zYusIVvbmslnjcvbeRGOUJk9jR+M6K1Uoyn0cJDZKmb1j/N+3Ofo+o/EdTNX6sKROxbIyz3143aR
9qPeP81Rx5qJZh6hC34E+0j24iL2aao/uqR0rnfY5paIHhvRDTHwlvy6OQynzJIObxSyiS2BvfHV
4BhKR3C2WQmDFpLFC7Ykc5iOr11gm5gf9PqpgktvAQGMDGWRvxZTxBXms3KutQOPUsmCphbCztLo
0aoHFWHJ4YcjagmU//gH8Bkcu2HNq/CYzq8nnpfgxTReab8Dvfqn359Nbo7H5Bh/u6qDjBRXm/ce
sX71cVtZuOjXOxqHgW/bZRDpblJayBO8g6ZjCshZF1qu1m7VHHnmANLHbZ7KQpuHQcJc+MXiYpP9
n9hO1hxqFTC20VlVH+WiUqmWoe2DiBmPpU8y4I7Bk9NztJQQx95vyX/OTeXwcMWYQ4KxOwTS79lM
2hB4AVuimRD2cCnOfkA/qVf7umsrqcSzCcmrPicOYpmsc5gFeOcgZrPkjsETeaM6O818NzKtdC9U
pW9Ss2QXV/3S5u2ZioqvRXtdi3LhCc7H6gsB+lTpFBL9qFrfLVLbgvLZOWp134MSQ7R2RYGjCB+m
wQNQocsyEWCo0mPPft8pfefFl0//DfA3mvZmgef2FECn3D54qMPBumPruG8Dn0VBUIXmdGfzgykN
hz0W247cmumbMvgAI226ZkJfNu3DwJmpa87PYTysjDhAlJCjmoH33qcrUeB2KeWLAyMo0Hbn4syD
DWfBUs1vVDWk9JSTey05NYZIjauHgqiRrw7p6ciXsANuoEfr6QzST4Wkm1M2Ddxvf/eS7gqlsnkX
iXAzByZH1+MJSaLa7pqz87H+u5sUXDuG4T7bhwEaU07+yBOWm0XPCvFPMBrDQiwqaarkXFRxWpvb
xfk8y05/dKlkRm2/GImvrxzoBFpN62OHye6+Nn+k58PdMMf4czxciXN1DfTusq645TaKaTHsAXm/
WpzxwdTq2cz78sZ6UvN1dmh7RjxLGOonM6yt/UBPtgqgMgqcbOTf4Jc+TY52R2nDvbRV56LkWTL7
06fxTcF5bfVvpck4vQlkZQnIDYCyr/8SnJW6ZK47+Vx623kuzIOqtgIdNEkCp929qrv8kvAXrE2T
OMkfdQaptcfJFEf9Hn4Z9B48xAUhs7kAxIPT3Ec+VH4Wt4nwBK35NVvNQC10JUBff3jbH9caBgnq
21eZXZDYPaJ46B0QSiQeuQC1Wfav7BOnIUQ9nRwgZKtEm604m+oYSzZSJWAdNzYfnBZ/JvlD/4YG
vceN1imUv21Z1RMIjDI8TGr59DnmphqQM8abRhdOm2PaVYRZyJko2qinoJw3kHlgQaEUx2By7nXW
k0d84NPpluNIoAghuXWrvtIPt/aJL8DG8yftmmInIy+8YgriuLSHeinb94yrhOiKCBnD1lGCTQ2W
v+RxfCXBaOzX9ZwkKrB/WoFY+QdLHgvTdvr9scLySKfSCUBXRql/c9ZHXcDlzkJbOzMlEmtvMXfH
VqzLcECKgJ6wSt9bcEk6VWRQwOHDW1yqsswpSrEnQiBj7e7Z6GrBkrJ0HLRHrBPqIrgto66frldg
wiO50tkBGM88ueugK0VOVkn/RLYkMhwnVdo1f2g1B6qYwldRVcNenwiLSl75re0sacw3F/PrllKs
yQ44AYtFB+HCKeJxsyGdu8zSsIzAVtpUT1vuWiJsd0aH9J2PN8U4O5lbndBBPnYdrBP+5TiGKBff
SdNMQDrsxPgxkzTlY6FulZ4wOHbVqftRh8sz4mynXjiTG91YKg/msxfZN5e4azTOIMiSEG72GNNV
WdIoONg+kF7PT8ipVSDhhVnkWBtJpwk2MwnpNB/pPpxGzZhBmTfR23ayA2HFBodzn1UsDqBiIjni
JLInxIXshVPyXuqrQTVY8KNXJYz6/QBk3s3tZJnw2SWOuZIRvbkTVrOeqjzY16P1vXhUDs7x3gIu
XkAy41qV899ud54OZIHEwSlzJlRu4vHaLg4K9Sd4SaVUnyXzBOFgiO82lwtYMlL3wM/udJB+4AdE
2qgIFjzX2k+iE0byOkWTixvPVIzAZeeEjaEHgyfBYqipWsfOm8cS79lzwFxCJHzfmXI6BquMo+ba
FRBPWkutgdjENvyMKDxOM8dSiv6YGvzH723W9Q2s/+euU1aCAhy9yBE2dPVxtuBud8Z84uWNQjN6
pE4zpg/8I8ZBrU3FwHDgWodHHIxfG8ImoEyZtNf+YZSJDRi+hOfkXf0yr0gY2WcMeqddhYHOWCJf
eYLqfyTgGOHZ/L79P4frk6P1TBfGGC/L89mK74XwQzldLangexOacBvby1MM6OMDlImtgbo1ucnN
9jqnrdJjHK5/blFV/Y79PYn34ffD88jOpY+GMl77HGQnxGh+1dJky/EeaHTopx1VFHH+oRbxQcA7
QdD82iVhlbQxS3g7D0/MHOFif82boiWYcvmQh+dDAawylmZ4iSNHV1NjWqs29OBVTbAtM7A3BSD1
3K+J9SMsjY8oKA1X2qGcv2SL3PU0tGeCWIl6H1feNi+d08uLmaZQTwt0RX7GINXksRoNX0OlHc4S
x8d7X1yLYFs7Avtkm44/x/0UlDoMXo9S3nB+xzrsUobz2QPZLs0ypmb9payKdpw0Q6VujWBwOZ5d
wTIgaiLbFvVL0eVEO33DWp/QLMy/eTbB1DsvQY4vEaYzs7ih8xiJLInkXGJo6neDC8KEP2qoutl1
lV9Oqk6oOM0OSEzc9318uI2LEKBfRY6be/tLA3/3O3S6rJojkZlDBKBy3qBmzLE8cD45oCLL3JXy
IgkMp0mMMhE8HZSiyBOY7BgKzDDFAQZvK5p57nr4eHOglQeXeE8p12C25Mn/p1X4UTGXpmi/De20
9/UBkI2xatgojiJniCUogjFNIE0SM2/1VXEZiigsRPbswrNK2hTaKx4IrzcHRyWVLhg1kpFYeXF4
/vyqkHiOaRTcMJVpRY2kEzoniY3paIGgNbxZIk4zdrYB84wEFaOvjLhplstRlkc/3PIAUvyd1Fhh
pe0rHqaSwhFfeWSOHaac3Fdtz1Tf+WZCYUsxrKIBweHULITxNKK5+M1o3NywF2QAJtSgni0OjF0d
J+GWlVWIltFa9XZmBTR+cr6uQfZJSoZKZhg1Q0FqxNNqY15Es9heiXTGCqc7TQ8cxhZbtvPwstIg
fvUDpNi7cEkGI68bCtUXT9xPbyDWe+tnV3edrj//AdHreO2XRa6q/V69u2qgqEPIY07xJWfwN449
9ASeagPDQ0VxhdhCtmIXD3TxC5oR+ucVQBftwA4dQvW8ws2xSRGnBc0WYM1OGkYnHolDlPrjo0DJ
RtRpFIv7kiEPjdHG+5IfxEJ9FXjZuUwcHOEpDW4sgfqpPkmOGCsCFKA7jP26l2uz/kh5KlwibqCL
bNXcCmApP8kEYowjleRz26yergQE7lo1bxiMmzdwo33uW2B8geK5xkjPK0TF85QS1WhPsaimYve/
KLQHIskgGesVmBhWfIgLfLV/j1lKgoB2fyYv01i/hQUwHPwFkhV08SCgqvcZV/ChNba01KbDOTuH
AKI+c8QIyZzo0hVU5Z5Ng5jNXTZ8/zyHfc6agki1W6RpEcEWr4WXnl2STuczvkXOMFtRH4H0lEgT
l/BWPiSj8OyLIyCMZADXGRPPr7oXpVql7yCWGVZZxhEx84HXmtFXJNbSRS/hAkNQllZV1J7Bt7Wg
7krw/PPSG4FhC8YnVdY9Zdk09vSrizAd2mZOJC4mnHD1gVcBirl0m2o/gqeWA7wr4kGbkxhB4nW3
JVG0naqv0SX1ICJiV+v341KdB/am6rGMLZPN+Nf9wmb5Yoxw/XMzalWoD3CF2xCT0IxQiDa9kBqV
Ue+yGsPaQU3fEFvQbzsAmpNY1IgoLvJODY7LF7f8EpXUocVzBwZtc+ZfZgjdputhjXI8VUxPbNob
eYCwRRUy/ihB08QKKQMwrdzuzG/7gBsD3rrzgWRScq1wph5pfCWBHJ8pjhCldYxIBkt0j0XD2O3E
TS93fAVcNvMHAAfUG/jqcTXAI9Qw0fD2lMP0RixPUHuD3vUkwqyCq65rmqoHTKpMx1V79ZqKl6pj
8cihs5DiS4B5ciPdsYPDdmPSBiHb7cAFKsvVd+n/c+52NcqqxpgLaQlSF5YdyXbpqj7ej9K5g6zY
ojgHcjcyK26EiNQHiVqln2DEnr7xdoTfK6o/uSPPAfuXoCLOWxbzAS1fKQAYOHPNKKKuXfOmopUr
tlnQlLb05gh+Z9YhnXnc/4xjU3JAEcsHxI+fSDPa8CWf7me/hF+UhxLOGvjv/o6fIPOu7O8Krg2c
dgdpZC/KNSY2583e2xr3rEGVyIj6bYh+ZGgQ9Vz/3yBPP83PdgLZbc/ZeKdg6yY87HSyQL0aUP4x
zuf80IcSpCGTrzltVgciqKpRNON7WARH5UyZMQ1OZ9R2A9MCN3HGZWutYRKiyXoggUmFfTo+2DR4
T9A2T+Lf7FUlsXnH1gc8Nd4eCbkYyz36a/3a1MZyfwCcdK0Hb1lUofHYoZA+asO0kyqP7hpGYgOk
o523rUsxHjzlW/k3WWdKdbYU/wsLC2MNn+RO9jd2JKdtn09sX7SkvtUhi5iHUaXJH+LbGwLqeH3A
XwDLiZzgp0yHtoeqIfXSgYPffMpCy7TncvZY4eh1G1TyS9DZZHgE7khGp/9JX98BskO9lamOvAzB
pQvA58Cunlr/v8V8EeKNbnbzv7KLVrsFTJ/A5kJKDe3iB7bUsUHL+UK4dNyP7rHPu7YrWlwkr/uv
r3/P2RKgtf7HsfNBBNGQWOiYmMwUvZIc06u/yhgbLzIEIAA5Ftby0STBmUZ50oT+PEE8BQCygsbf
y6O23Z13booU0oBrqvj2ezsEpNk5OpzEOzoRLYcwf9tq+ytv7CbDTXFZ1x+9RhdOljtYcVzueTUT
K+bvQMiRwAJ4bJkqB6YCyHhJ6agZ85iavGQ6u/2+pmkH+pO3K9qioKV5ltvnPrhdAEKPGnUXHLN4
TsfeTKA764XjsYJSMK3JP2raBO2BT384gAgyipSOPgsBXZN2lR+aDRIIUuTzS6f7McNcHHVgspAW
ueGZ1FqeMZfDV4u3WGNYqRTSUv0EOoE6uG4obmUIVKNl5ofxQOqYuSCQUyowLWaJKh3rn8cHYsMv
nkzKxuPLpWtUR83u+MMYa7/GioQFdHuwEkJPGdrbBl2XexAbwfJDHvt9KzdvFHfe5BYbTE6LDIn+
HQ3bFRcm9AEyhvFGatp22vvullFDm8NPXR9uC1Z+W3yF2EsRo26XbSmjQzAou1itRNwyT0OTMAfp
Fu6rMOJdAVcefpHN7L2m2wBWRi6IK0D/fwz1TIJp+/g8pj41Yhx7lBLe0pl2PYbrqjksTNj1iUUg
88/IBa5LGzKZZkmugSEIOttPvTdWBgIBdYVmlapBRSPKNRUtdAk8wyTt7bzIG93N3x8CD77sIk+Z
uU4vEzuSkX6SAkN3VEvJtg7vYSOTqyzvT/NlImrqMNxaomJEqeioRTb1gOl9XU3GmtFS3NlacEjZ
vKvABzcPkeaHTB96a3uUU2pWjXV/pqnKSrbWJgIO9oa3vf1llHffR6nilmaYRPysmMz6W3tMnJgm
Qc087jOK8RcHvSixDC5G69wCce0/XKHjleTai3tYktkTg4mNSSuS9E8QqQRWB+e+yX0e5vRGsf6i
PsboyITgbohg7gwQ9dA9TYVtMD3SxtiM5a06Ke5xEFnPowOeuWNWQ7MbC+bZADv+JsrhVK4wQVoq
8g2YQY6BGvGm6HjhcJIB2rnjCzHJpqc96XlkK6Ze5kXjWki4HMhXgd0d4NEROibgMzAwhgEMrvso
p7uhMyrrkWj6qp/IxBSZjsDq/qh3Ii2HLVsRjy9YoV6Y/9DA5mu6pGni6OxQtjym5Ql4gXdTvNDd
1zaP9mz3LaVDhm0l4eu7DfpqsaNL18o1bYLLkm6mKaEnS3uhqCTTJ5cXyagQMGNl7RM8pKtQLb5R
mSNTzjM8cACcy0Tp4aBrVZovPWUxfc1cIh9U2djIOvnr/QgqP9yAbfLcEY1/Klhq4nAm2w3DUd0Q
1OYoVQu0boEQWlL5wPpe1Xang2SgzOS20lcMMXM4Gs4RittB/RyF+yPodyTvCR5IngUFWXNUQCy8
gqPF2aHLv8xmWVOHjk+b59drTef8MqroVePnIXAvwvwRJWzzt+e7XzyMQsmycjXIArFp++o9gDk4
GY+C0DPEfRywxd2T9w2/P49+1kOT35YJWRUsgCZQKufFVGKjt9ZafYFqkKq2x4wh2wWgSQ+2uMu2
XFMms6Zp9WZ31R5XCaA3Mtm5TetdzZCgx2e8qjGOhTV4LZArp/bX42q9TXI2RUaxQGh9ZlVvqGPj
X/rMJZnMvEY6cGeqPIU6Bh70giTOX00g+Vy2dgS4SOHIxRpmBBu2bqaJW/kR7Fhjz/QnqOG6Wb8T
Y6VqpBMSjnTsQDYP3oWLyD7aYd7QPC2j3sLWfEObg5OCEgKdJuFQ6W2/qBXHHF50pXfJE70pq1RR
anXA7pXM5kYYzlg4jt1vC+NMzjhAAI4Gg/LfyYNgbWh0TwCQcg8+JKq6rgpAAHEPucjxmRixF/L0
6QX0tLDvT9S3rLEMhxThNyuNGT5y7Ju6Mn33OVfAMYbbjY9ohI+0WFOTaQzP7PMkMtWeq9IaBetU
KFODYkenaYy2D5+Fi7xJN0OM2uB6nO4CJmqnjG8rZC6KzmQM/5IzA4als2a4zv+b2zmqy1S8gss7
2N0Bn11TstfAS0XROYZFWoxgzLqa4j9JTrHvzt1D+rUnXOFFAiz25GdCV6h6mLm834TimjA/EJGN
aR6Y4YUGPEjJa9n2C5x3+NSBHXlC5V8pHb+XmtNl9Y0A4hK5BPHMRmEnufecYDYC58OoUy4R1wXb
8+Aj+yLdncezuqbuG7FlSam7kLf81DLMLqEe4QLhEcDWobiR8jlIoO4YOzyY8CqaOZyB0CULBsKy
PY83CU4MQm1Y310NwKF2EBm5kcPr40/GXkUMUis04BmSJwqfweiAVSSYKZJsUP6iVAc0ZJ4w9fhQ
LdQTmF05mPuSc8LxUd7SOq0TnbvnHgn5M7QfIxyvrvR7tkj1qwXUEKWiRDicEp59UIbwba18U/80
Kl+UKPV89VnHzyqP1l3gegAo/c7sVa+SyO89ow9+IaJ7IBwPAz9DClFSHFvHiP02lkOkx3Qman3X
YPy/JpPiSy7GtwAZ8aUuo6wZQ/Jsr0Pr39xULCL4Qt4KPw4YKaLSyDCaIX5Z4DSjPz9HfvR83250
ix+4fZD7o+cOiREp9vGX92uhPPPd6gNSsHF4grW1zSJOQ4z5rcvVc4AfgK0Hb02U2Fuz9Y6HM/nd
Pqm1x6YnjthfgewbyNq8lMV4ntBRmSXEv0cLRIbvV4ovb3Fpe20T++GnCCJmx5TFkm0qZB5JWJfA
2c+SS3d5Jr+ThLRJjOW5Fbb0laJdvHJwd9CM/0+TEZ//wp6Mt6R/kvMAHZmhg4Hu512oXPgy+/AX
Y2BpdrGtGoRY6PtI/SKUgPwzAWgiboVDnCIPb08V0zL1NPCq4isRVPqW4ByiaiaMtjP35im9FwGk
jT4x0qMXU4t7DsI+ml3NfN6R7Sby96IatH+pijE2/WyYSYaOWOyrampLhaBCPZI6SNWoKiabYCcf
C3RwIZViKaZrHn9213btOAi4CgIearfQn1KYwagJPepLYF3VyAw5TYGYle+Wk/q58rXq0ZZpSFf7
R5/cdBs7fibqMIuvgb4INZhlfqBpHv3eO5UGKzxknDOMZObLApH7ZQIg+7BGBtQMZbAcu03j1A8k
Nv6EnzrPjWOZCNH5py687SsqoDKw/Psn4tPHLd484j8GKb3Ku8uH6uuajjkncWSkoYotY+c//I54
JvNUhHATL0bVXidjyQDzIpPuqBfekarKjs0bZtupFWfItg4+4Imz8AtObWW7x1okm2tD9pKTsBTj
xq8urtJy9NnuaQq4llpkUqt7KB0SsPgh6MqOiLRevNUmbm11BI2jZ1U2MP8nG6uEgGAqmheQ7G78
BBjmSYnNCn/YkkZyT05Tk7mqsgUemI6Y4VhXUVUhX0ThI7GaisKItiz3rEZndPGL1a/nbJwsqnDy
2L75dB4w1qK8gN/UHEX4+idIEFCQuedo32rTxkIAgKsV5Mcfi5K+YpascOyLIMGbb+7Qp24KYSbA
u+WCUWdD3EkrJuFAK28RsRQJlRjW9uJyrIWxmGwcvBiZpOxCH8Z+RChwXsQo5OVOHtxRDC4klj+a
JoA/9EAyncnF5zmus3AeJ7iGqNGzjbUG3vSDd09fJndKzYPQtTIG3Xd4bsx/ROB6NRUaht5rZTQC
MPl7cLDVP+C2c1Q7qgfKPq6HdfVjkkaLxf6MeDRNyfDta9lT1vKcy0k5Qsfbjo8PZl9N2aQlbARw
Omc6s3OLECWJXY6EhRprf0SwUpopc7TwfdMZVgY2HHDPIp/m0yK2BRORv7shbc4T0WRGLOaFmist
EfW+4SWRs25eD2ypzx10HaIA+P+dLGbL2xHBYYiasdRCBSyBEvwGsGixJp8bbiNo5KICdcp0puqt
XXRAsZHejmQzf1DW7BydODKDKHvDb18qO/5GloWW8ymHOxP/IBU5+GJmmtxf6GtJUj+GYXJv9bgD
2fnHUdeoOX4+B4rJeBSCIbDwXtFjhKyK8PtC0w8YswaZTn9wxtZ1v93brkraoYTkNl4i+mmrR3xO
2nYEslOUQKwyu0asClQSD4t8zzKa/wGgJlQkH9ob7dbYXnXJrrJfHt6VYcymfUF0Sl8t3dhM1Ile
maoSwEM3Hw0O6HAkhgRxnMNPIh+CskhsyBar6YFasNDGREyu9QdGixxMcU7hwxQjMxF25UEsWnba
QTFYpjjz/94mkEX+rptQxHMqsyS9FxzBMxMMGkWDsvHJZ/8e78BIGcAEWkmFjT8Af7RKdfjrr7C0
KUUjrY77UVGMtcgpV4sfypDoDFigRnkWWFea4YiBNuwUeZQOPHQCr1TvOM8yHcGEON3tUkqJwDDh
+UpoU06wmy0UfMfoGl+HUa79pFR8QSN17ioDCKDkR0zYMf1c+AD4DE6WTFf43VMdITheGegUkbf7
gEjuvwdR44ZwRlZoEOQ+7F4FL/lPIpssB89sHY5Nd7+SbM/zcNo+6dKF/93GtqspsxULLnJw964u
1kvi/c1dPokTACE0NdHkE3Np0O8suV38KywUXwB0V28J/LfBF0B/WKMjmrvn6RnFca66babn/U1Q
4g0EhFKRyT8wRC7+qm77NVd4169H6ofrqfQh9Tz5CzZIOj2vk91zqGIJpdhkgmmnq0VUzBv37qPF
T+/C1xj9DE9gwOOToqiORwPzbjV9k4E4XyHs+1ZBh8lok4QGx8FdVxgYGT/C0coU66GSZtuU5tUL
PejUc9zgkemtrbKMe/pJBkyteIu8o4Hg80zEdLTL82VfwTaqQV2pE5shhhukigJQppMq73WWsO6F
4Dp/NNxvx+i1jLyruW4f3FjYEMmLBuqEsogTBDfrnV+ah+8iC0rnOzVo+Ah16/BbfBYwrt1lOdGS
Wk33jPRRPzy6YFpEbRB0A+SAeOODxy70FsLYvh4HdoXt9dqRdTISQIc1XVTzQSzl7Hfz1sLjppb2
VwfNfD4zAM1lCSuZHiSRNtRwucsOcvc+hD8O9LW2HGZhcW41Z2KZ+MzKjyVDicnAibUJ8MeXKMhU
nGRfn34wTPw0o2CftnoB1iBjhepshd0GYQ3Q0eEhw1RHCEh3hHAMjc1ZNdD2G/xRmT69UwA7c8Uv
tEvAdaHE+7nbaSZwmU778LF2Uh/AnOLQ4DLfwU2RGkXGI9shcNdT1rqYvMMaSTF7znnCaxl32a3D
e2yz4l8atDrfoAnEjB1lSL7dZLN3uK9594WBQtlZCQUNvSNENeNayLv+lMNze6+7eFeta2CCDjC3
gCnsD6+k2KiQ6hMYkrevTKz8U4nocZ67C9CQW6aqbBu6+MooLWi33zg9+6zpf6pb7h2nUMw+gvZV
YbJxZ9/qZTeEFMPjBIFGmQipRpBxaJjVTbCwn/6SFRS7JL5VcvK/nJf4xJwSaeZETmbjG712iQbX
NzW72FtuGcQmVeOG781OojlUWaJIhxLJO72m01ykrn21vDX29hz90cswVmbFQmx+IOAFNIeP2yhG
pY1vt4C5ZtPBb1FYRdHyCHI1aiJUnOdESMkf6QjghzDza7MLAl33q5UGKDTJbWeIueyQA2VQO1k4
2m8PUKonygAGgBFYinhiKC/LDsc33D+EyrttmkjOJPd/3CI9eJS37a12Kwf0IR4FZmhlkAGPx9qx
rff289hzKbcO2t38DZqsKre2cLy/Y4BCjgAaH7//J8BL8M9DZ8nSvMW+SZexVv42VErWqTz1UaYI
LEQzS70z1vu7I9dmTWbzoGFxUgGAWLYSSJvU42Qt3x5jbaGdWTbDfP248wyG6wVjEXwY71mCMAfe
BgU9bCskKbMbeYxVpOJnwIkB5WBO7e9/SpqhqO7WYK5KNeKJA0+4MSbtBtHwH8cajquOr/5DY0OP
9FWmAs5ilyJvXshQUV+cjdO9znVK7IDph5MU+p166fLUKtWrUh4Eegfx7kGlU1Ab5b9rovyx2VA6
WKMhDxbcMjgO1hVf2haKiuIYOhDRq74LjaIU6dSI6986e1J+XSnIMMiLFxVqKYVo+SJfe/GMLMU0
Fw/Y30ewIK8ou/AEijpko+GeFkeJ0h5kUptVMTaKIqDGspc9vEDVL0rF/9bX0FqghKrqvx3k7LFd
GIgJZkPraqMXw6i4W/rCjLuKH79f1xs+yqlVeP4zWRFj04W9kAxqthwVDKl6IrK/Z/kEuDHKyR8F
rltT0hfu9ebSJ4B0Xm4cS+UlTe9Mknhh3ZT3m7ety/LfLAeBgL8xHfiigEOs10LWBp60Eg2716Je
1/ZT3pACXQcL+6Ng2w2EZmGr9y3cLpRee2i207zxJFOqMj/ITAUdKaPAvRFVrDrLfk5OjUpISUvB
n4uIjj5x0x8omvqQQk0jiCOJGCwCOXVgdnPfSNBY8LvtYpFKLjUKdBMVUoWD0ks1oK78QIhovmSz
vbUtZ3rfmRtxm5zq6MLZmg83XVDvkbTYLDR04kLtaP1MO+t5b7T37xzEF9FKh4nyPPXykWmtOcK0
4K67FfUglksQDoDdKbdbG6AH5cCPeNuIki9zfH2xco2Rkk8g6l/d/1eaf6UyGF1mDjznatplK54R
fkwS2D6VyWO8FprJrScpZr462VnUUQw+WHNG7PaP4f94GL57DjCbVjMl0KabAsBuqQFmV2/zCq+h
wpZgGz1WbQyCEqXwPlVZlUmkw1JcigsRhCX2wQsWhDlDd92rjpKwZ9HWzUTPm1sAHxU9XlzpMAQN
UvTgKkAcoiDGwHyNseo7rZF/7xM+SP5ZxyOIvyyg6Wxkq8rbO/ZPyK3qOXpvFoj41AWR5I7VrAm6
62HxFYCpAaZc1Obx3f2Uenp3al6SnurIVqOMjhDc4Nfqjm1hRGVbLEzMjwCGDIcheektVX2wLxKi
+wjWbZqxRCU1312qu58+FxdQN+RNxej3LKIdimU2DiQL6ODZ7lPT+uEMNFfHcAo9bP+qLmAZyHp6
LohomQoSqZAFOQO/Tu9pn/R6+zMGoMfYRJ6d4/JGeZprTFoBtqP8cnjHSUylBHzr0tmmOoasv5pN
Mw9Qde3ngBSqT4Uw+3E4lmJVNAlQkuQYGMRr9vitq/xIJBhaWjXngHBRu+iMdYdNVVr16gmPogYc
CjmbTzP0OeA1RJhyumf1JUqak65O4VtW6VAxff89ctMZFVvV/Q+eA/lkx8k+TU1hAFApC9q8P6+9
+uipMMSWziKDaTzst58MEjckO4d3Lhb8hjLDUMMSRdWfrvbuYtsaMEsHIbYkZT5mfWsssAj36Iy9
WWZgd5Zq3V2zHbrC/VFLHsPyh+N7Xe9PD/CMjQnyERIBN3EMmM6NB3jQcCP67+cmc3e9cav/lB2c
77bx5UVTZz5GUcxrwbfSB45In5YJZNwxOhMI1DKLBoef0mW6qV5We5EKnFSNW75I10jTlDwhN5g7
I+p+Fpt/NLG75HN5RfIeCg/ARR5HFOa86zWJtNjrmxYBKPCM7n1fEb9IzLANfA61LN4lRcuEl8N+
kgGbk0VxA2x4MtiYUwS5CceYjZDVqdGTkcoU3dba9TurEQr0qlGknc3zXB6PAsDMb/NPs8uyVP/T
x7YRi48EaVrW+msKthfz+UEdHxRSV1ygMaS0YuDmuO30RIo4Ei1D8FNkrINCFZFo2JLRUCQLd1IA
uxso9Asxvvc8KNFquNSc00bW0wWiPF6ItO8/uL2sEWRYXl8McO5h6ra72gTwV9ycXNdY+TyMX9Pj
W8xNQ284fRgCYRc+U4X0iPYq+AGEHQ9PLjVb1y0Ii42eQ8GnMdg8ivoaimOuiQJ0Sjsrg8Xb0HlC
jAYxDYmxTMiYqTJGb66Fvd+HKeju9Lp7fRlcqltabrT2Bv6c+Yhn6vJJBfQ+hPlthA+2piS4AOQj
R52IWRxOsBl93YSM/xh9a8tExFONTgoErQ3wLWqkUt4TVdtufwPlh6irPQHPVqMsny/eRLy3ezsz
u0aBSTAxbceKPUBF2dFN9CmK2YY7JA/IoCWllVq2SLP08XXmtj3cS932gyDl6ekdG04Q7Aya8XK8
4yDkSto6AUFUaDfy12/siNdh4eX8GF1uDiSFXD//PeaQaN8hOBsSGumAQVnKlSnozwHZqeI9gRLV
YWiP+6TauJ6lmGXfkHx8YwtcgsbULA3Im7CSrZiBFrzAPbfuY+U0Jo10rRCkpaCy2g6n1aJp0+zw
/ayXxdJzHbcSZmEJxGVAV7QB27IIZLhQyRowdDZdNiok2Qt9T/WCJ77ylE5yeK49QqWLSO5dYIOd
aaQXobRcKE//Fxo+uJ4iwD64N29Sv7Ux312OaGegAmuFiTah9wgXjaDfQd7rcuZS+ESl9Q5AcSAa
/03BALR0RZ85SueVVA4CIk0Lvv+mvqVIpiGcPSLu9Uqjwvt8IbUtGJmO6qcxcZjUNv9wE4qkcVhF
nygcPlCRx0OItA9NWv+68Ihk2HN/2ItQdSJJwtU+Z4tKDh+cqb8r32AmHjdEemLocjahqQQBqyFX
/hwBgtoEY5rN3pMiZl2ZCdvsGLXe3WKO1njH/nKmXU/vrfLH5YkzLdBCxPpydRpaHB1tF4yLCa9V
5XRH1qrgzC2QVdtuAsGp/iHwvMgISlmJ6ib03qADKdFbzTMJ99RgvpmojLA+5J0rzjxphkKRe8Zs
h3DwIevyPmimsR7MkZbV8Paq2FtEq5oS0QNqRpYilYXKdoOSmFsBSo1Fa6dk8QLjIBBJ57S8VdTn
UbflTQO1m4g+a1TNosNHaSkvdbuFDTTjGVBirUt1KixgHD086RNZZNjrGBNvRRWbVpirUQrjmhgw
074kxVcvBmLm9vROa3vMBMYy37f9sjqXidfNz915TcFwjx5zJb6Fd2FYVtEXnNGFEvYw6EhbwF9o
hStR4MNOTcBNoTxicMFTzsSu82qUZXiz7kUTYzxCPiN2EBIONu9CvdkGizr3M6ipvNrBT13az1cP
g3QkD/aqRI9fktbHG6CYovO70yym8P/QNZ7Q8KiUSvlqXI9H0f1IUmJaGPtgcVQVqNUmgEVh8zu1
G97yY8fXoh2lzdh7BIhv/8k1EhWvsPi+n+xADRFNOQOGrz+sp+JAIMJbhIcSxoAZhFmPrkcrA5tC
1AuwYk4mhiFBp3VKoSIv8iqnT+WBcDlCRO0qdGLeTfmp2US7OnAP5yJ4LjJ4MhVua3sHlEgZ5hQy
I87TCEpbn9K2JVf/uCxw6GHK6K+yRw/qlkuFksEdcc8fnk12YjQGWH/YbBkpUslVl+USz+bLTtfS
SChr6NvT2oK6DHVOWWCJ2ZEA65WJ1cx7S+BxO1CvVFiC8948Nf+gb08dcWGRNIvuflBK8sKkXNIt
ftiMT/1C4+C/s1jkA80JTqWRt8PrCT+cVfi3MxCiVUSK+s9LswyAQ+Pmr5LTjYqW1+n/v8yqgdFo
RUaXFxdKFZLGmc15s9cIFPth55HEznX638p3GA6VeQs3aHz030UZYKvKDlbFmmqD8taE8KLnII92
t0BOJq3ZX5P0JEloh5FtIZAcNqzfGHNpZmzfIuYdo4XpjLYLr9S0yRSBirfTTrrl5om0/ysfS545
dB3+l3XmJuJwsKqYGyElwR/syMnJF/D5WJAPWk5Ju4PQ+R6KThY4BxBE06nvnOt2Nef1mEFq3wNA
3ffnT/k9XK3fbEHR/Mhxu2AEe64glcgYMVTruzD9xq4wmW0gOHB6Cn0eXgXE8z4L77u5sGIsNaFk
acrJi2DaMFc7C2GhQ+3EX1iVbLBmFri3M6woTwCjuVhXHP1tN9vbUqefb8Ho6n260Zrf7kwnSAUP
0k68KGp1Af1kAP7oqcy9uSIQ2g5kMkoCbvF//KsEo4Bzc5mJMW+LeespJcJbcMNlxfujs1+4fc5S
6iCLHG3HkxyASgbuSWiGYUpTTHVJdxW9hnmKMWFMIGQOfllz1xC593qIuvilaD37qCmt3m9GN4SI
ornNibs4FRYoJoh/co1g10kBMgT15gTKYFgf3engEA4uOE4n2u8581hMhwU49qOSMCCRhi7/yEmo
XVfMkrmeHDYLa1Ur0RsqT8Vdt50pgSHQqnMy6RF073oQCL7YICDv5QKP6BhPRCynYi5p5j1pWw+p
AEst6GkhV8ig1aSgzaX344KYfeycBwLprqHES4tSHRdMJsOSnofdzbW+NCUPofe5IY4LHaf2vMbf
BwTTC9lFYNjCDQOHENEW1oI34p1LzC1LIoSIsDzwUplzI3xwl2TIY8oxci7LfrIOgGfp8eXi99Js
MAZLfJ6eWM2Nwu2OcDu/2yWr1BxgNaGB1BP+MEWsKkhTPQyjoJY76wpxKd7DRHMA0VYz846NhpTY
gLgTx9i2iF0hL9CMxZrrfP2pS9MPah2EoRvI90DQDOj5gTJfvc3XFqmcTOAt80Xv6o+Ty2A7n8V3
HxgULrRaB4cIJLbj7cFNed7uPfTjW/5kQtC3uQyJ+rbACBuCsjbunKG8XBWgcbaa762z1WP8uFYt
7Slu9g6LmlzpvMExf1rwqCI4ifzFb8RzOSbBBhbHm2/vf5Rp3Lv6uxshFVZFksWU0QwPvYM7r3zV
5EsoznLeMbZyi3Y4xXnxshs4URvyxecBv2qcRf0RQVqnn7PYh57+ak5ZythOPUv3kV/Xb66ByFSG
F1r963pIxranAMRe9PX3PQWuodM5w1n0muITTUdBDy+cw854ieRFKckenUyO/+aEbGNRfjZoQqlw
6NBD7DXkdsBeR2zXyz4FkdBgZo6H7keD9AA0V+EfNYavaw2SDl4ecd2lt7c/PDf+vwMMWIFxeyNn
uTeLttxya/zPw7Pm3Vh7t6wkbOgYzKRP2ESsPyAothb9+5IDjtHB0D+EFp/yF6nnoFa3en+PQGrV
hKNEYQxreXq4evPaNRcbb8bKucvpMVYLYrb7AhaEyKe13H3SUjooVJphvMLNvbgZLCe6wtFLfrL8
ipVnLR1OHvxuvSr+8bdDX7HxDVl0r2v0KX29bUYaIb2Ge2O/TfFm+cOXggJfkmQUDZJM2/7IUHEK
TKxwJUx+BHyFIjbPqFx2DdycKriTU66BiOVuHHSvTAFN0+rQSrSC3vtM2VRcP1orlId9GUxaglLW
5IkAWlEPnFUj5J90gxTyYhs9q1Kb1s/71vvMlZETfibb2Iyk/FQT1QaY4gJwaxRGuPDfmKulVLJU
YJrgROj3UxxZ9siF8c7qeBBeRb8ss9XwgMIK0FpeFYBtp/skNhE8IS9uVbLWB2mLS0ya+7DiMZeJ
0ExHyH5vlyCzYvHPeJjgdEVNfRWtlnPRd3HD1F+oyNA5KsbkHhzoFnu2OEENVXyJWvK1bST+pU4F
QypU+W38ve8LXl3EQ5uLEXVN7Rg1WyD2ky+JG0K51EtzOJD2YeepWaWwSAMHZBybqF1Sq9NaKdU0
VDM+LdeUxNHw42fNKEokSns9B4kE80yMXCEhMcb1GDZBYcqtYGn+R3kpbKamhH7fwxhq3izZz6ZQ
lCrfpRvRTWVlSthYL7c5S+T+p5G0oVHgiLb8DGNeBvl6cEkdmkNSLgV0SiqT8vW1nubn2j0i6GB6
mUeyseNH2auqEmMxQmU755w4lPxfhY62puhEzOK5pqd2ldKrOp6d7Tq7IaAQsbCH2g7lAMVKyzkg
zg11FVf6YYdBJRyshAMey5J7p9xAOOh5DMUdQcS6e/VEkQ6C77IsmQpjlUWlxjABYkf1QxpE7pgD
8POEXNCMsqqjBtEwU3f5FvqrbNU8kpClC0p6RrmVG6NHKSNoUbWmPdVqRB6xRRAtK5X1aKLGkXpT
scLjC7yXorUu3ThyfrFlkROfqVmZ3WB1tA9AZWi9HxhgTH3Kb0+faMi+mrcZZftMj28GuJCbDOtY
4QxnajcwlQTuL/KDj9/5+ZXwWn6xIlTIwNvoUI/TNIVmZUubMlUgPCSyW7zX2tvVuATerVvCI6tF
rIU/smSS1sYhtE9+GVIVNq/G1ySGL9O6PpM+nv8y3yuXQ3sA0RgPfyHV+dhUj5SxQqPWPbiv/RMJ
05JMnayTSGm6IZPpvqnsaEKHwTngVecL4t3Z8I1+IzGq0hRkSqw6eQ8uhKCo6eQX+YE3cP+4Zljc
mXTtVdz5NKXLe4EFFCuSAoCinwCGVlbmNCCcIx2o8VA1voRO0AHkpfJdnXwImJo/SEOm5ho9vwVm
ul4GDaNsDWGnRdOXrMXrgFuj+6XM8Ape3l599hJzgz9Mkk1qt3MMCX9KpoJlmiJL0u+eI043m8aF
CXjh1fZG972Q2rzHJxNfzMEpua2YlC3teq7TAU/3zD3hQ9x1/w+g7leirEnJcKHWaPeCAxnKvTq8
Zx9Jc2qlEnbOVUpz2COoQ4MsuVfID3k8GEwbBu885mt0fYNuC0bUQMxl4hCroy5leMjxkbkyvEC7
zS7V+DFoNxFgAogY62BCl+NzZfMXnfbgzy1DEBlF5Q4Ir7t466vgvUGG/GgzNbNtS8mXD3sZh/sQ
zkX30d5EtWV/UqmJzF0JcT3uALV13UKw/+vUBftqYjjiFdhBaMZa2xgEnZ1E2JnF77N1LhMr9cZ2
IyaPt+xVQHDxDT/jJVu3Dxbh3UlEidclH/YksfM7ry/yCsIBH+QU1k3Le69mX0oOZoQapAHJ4MCO
vInqRA81Cl4r5VZ8fZMKapEya3HmDL67s/aAGaGL0+TJ6/6CKfIyxeNZKwJVNyF64IHlupHUSFFl
Ar+RH8nfx6CVE0kA0kBDTjMwsM7iMqtgi4WtxWt3PSdeXnLibZMvit1hG04Zr3gs2R82uMq+14pI
PCgNjl5yJ1GPHFz7rFrRgh+QOUd0MlepIo+H0LeQf1uns7xQJ2SPrsCDWL0UJ0q8WGrvMTXRcGTk
YlzzfCiZ6ByFLa4cyJ8Zx0LfMoKC8sSTuZOyvHqRcXdFdPywVGdNVH+MdQpsdatuKpu/i3uqtd5Z
WzSXOC2Ig7uQOprjTwdpGKd0idpjiVMYH2CnXppIHVuA51VfEASZ+ogu9B3c5y9ncj0bCacVVdD3
Xbtr+JvJlYa/YCy+r4FYrIA0lthJKgL39ikkjFxgWNdy4y/EkvtLni3S05c9pqQQv2uBAHGGuGc1
qZ4zfHU/byZUPYwf58z52ayc3tHh+gkkrc4DBvl3WDDTSFB/i89b3D0GdjURt0ah3y37EHnOWaUk
JVTJyVoRKYMmhkeCdCGPIlCjapIUmo5FkRBiaNoomyp+4aZ5h3FwaCxfJRrUY2+4aV/qFU39BTbx
yy/S0lE+ErhJTu90DHdBmHhVawaZB9GXe1f6NxCLQWvASKgELmdUXErR/I17CgdN+yKBGr7xyOWY
BLrKr/TehzWiuSacWU068S9rpCV99mdoJFFX/UT3a5VhkaNcjXYYCVcijL8Vqz0q6wC8Y/946M54
1aveUnnyIkR90G19lVk5ZJFNTtS9qtYLpZgp1rLZ03ZBhQ46idgLRvH91YL6v0mi2JWfQ49OWwHb
39l+sEmtPIOtZflvbVCpb/Xze9nnFpU6IULpPj02ZcrB1V8H6NsSgdcdRIlM8WwviDqrMBLn7mRU
FJXG2Ge3UxPDAEJxo3yg83DAaiOZ9/BwCYdDY2XNANEHxSBm+GgAKKRiW2e6tJu7UoR1XQUI9VUW
v8ExO503waaB2xUfsG3RTScejLIQsuiDsStXMwguMh6DfpxNaZjU7VjuUpEjjeC3bW1PtzEJMHrl
bAL0hqbUXicHCO4Pn8XwGfvtfARivH5NsFhAZR1O5d126unh213B/bq775FVDX7wNnYOtyFoA2Yz
CWOjVe2kps7bJ2E7JELj1o16clzNlAfqVmOodyVXGqLIRtlIkBs5+VC3UZGez/wud3CeCpwFmsp1
sZ/C5SCJfMBHUVpUPbdWxGJj/xqJP9E9FjTHWziAqM+947e+j6kYipc75jClnyAs/+eWJbr2U7IA
UR2lB58tcXvDmS1yAgz6ERf66YinHIgnnnQ16HiOkE+p5YhU0krEs4ZUczlM1bf5Yp5/mt9o0kju
s9IRIhW7a66sPQHMQf3MwO56qFzwZVX/MkbOXxF0OS6ltTSSjjSfp56WcnSeZaQ1WjIsljKpd2DC
R7BVScZ2hIjrHLZlzgYqOFrBwwadJVlblhkbUA8xNBexGc3j0w409ET7F6/e1ZvGoLChJ83UgGbB
lM2S5QfoSK5r3KAaOERMi/uCf4EGaC7/0uS0eIKl0YujvpgLbl4hwHa2EJjfLMlkxBppni7BV2Y4
L96xqy51MSGJbzgxKyNwE/kTma0AIGwrNa5R4i910OcI+AiXk0lIoldsOVyAl1Vg9/SCWmtyFFwK
/buOK7NYcr6uPKvsVVR51hG1GI3rgeFUfPatqQnzKMp8x0kNQFA0kDRGjqIK4twYgvMCEKLminXJ
Sye6lF8xbaNn4DUu9W09tWgxKov9mn8lq3ojKhhQUtCeyOWzAOrf7uWEY7nGcWbjtxoOMN2aLG/Y
3j0ZYtGVrrYYz5iMnC3n3Z4zsO/V6EJFp9Io9nRqYnFrm3Pwj/I7hOCd82IHk0kXHfSXrXt/kO2t
TU7i1UN9Dua1YZbSB5t3wmJPU6b0ANv8hWoqZbGV/hJnV+tzwfq7TrTpW/N3Cilu7+ysj4URIHMl
WgwOt5lyHvBdBpNsVgtJesApcVydLfXt8+Qq1L6AobNDBF5ZktKGXyJLR3yPj2GlaXLrxb+fWnND
7/93VG5SoGxFauAfCATuCvk1faJ5bW1iXOnVpYbma5pzjYS45m0yr19mDJXY8AWc+nZX6iGURPNA
fF0VOIEDR6qqcZMnShF2VWssXW+L4jRDvDgPN9OCkT2O/hLU1lKfusJL2IciqRm9xRghX5LETYwt
iiRwJ/kX+83m/QFn/DOLYECfXa6Svb06sIiEJIn5L5lpILt8xM0JhN3PMqMb/KGlXH3gyJLg7C42
FScyIHmao6NyQrYD2EOgTDIjcOuepVbAPb1cGUmgnMJTflhJadIpDw4y/9Fgo33yi2+DJy96uCux
Rm4kYpkEVTewf+eVARVqjWS10bIpKOZs65hq52NLdZZDtNHE5p52W36sqX6U9Nmu5VtGRxZP6/bR
fv7jiHggTQ4bokHx6wCYRJOhpp54pTA8tuGhQe+82GJlhT5PXIvrnKBHSpWicYaZFCSN+3v2QFlu
G1Cn1N+ccXsEUE5CAYSKbKiElkOcgi2KT7q1ZoMisa+4Ozxtm1l5qlKIMqbTsGOSOoigIFzzhQAB
icStBDzENjvs9pVZ+d/xo70nO/wV58GgBWVC1PLLQGiwJDp/g8+ZAdXkARoSDhKUuHH61PUXdtXV
nahUuHud4iWr2ZHs2ZoCg1umzk3vT+VFek1em/wNLD2n+1y5OMfMXh0/zH9fqceert7vVzaJHHL7
fqvxCzpAyt5dekrYG5Ov3ZcDktA9sbGJGmCtg2GvzrhNL+Ni0zRS98BVWyjTpXoFFT9sQeMheCPZ
8/N1Cnr5OPlZJJCB+tyJMhNWPFYL7bGpV9JA5+S/sJ7lmvs46XA3d3JREGyiUe3hFAGfIQoZ94/Z
zEotyFO2vtg0XYNDO6COBWHsf4Xzt+3cSexGSZ//vFIJ5zDW+oFWLWabb1qMuQVy8M9ensG6pDOX
zqUzjn8+hGnjFlLI3CyQmwo1mXU7VUc3B0boTRB/hlMyJZeZdm1GJJykcGAvIiIOEwRbkss8gxDV
kXkdKoQEWaJ5U1dmJjMusWUTtVb+3pegn3hU37/pdcaoPwQUknf1+SjrCRhq4askaIJRRIOlRL44
V+Nvc0C972c8s/a5AZMJaP3weu7cHey69ECWKdo0ljN8xb91ziSJTxN6VRwV8Se8BTlx7mAUEhTh
otuLtcF1umPsX9OYN/GiGp0pUU1YEP7RnidkpCtk457QChiZ1CoAojpR8IAuCot0ZBySOQp5PO/6
fsQTULAAxeU+91pd2MTCvfFlreb5OD2ICZU8VXV0lc8MncJjAah26y8c02I0xWfL1NhN1v9kwoFw
gp3gubh+xrSkyl71riUA9kn1smaw6DGq+J+ssD7niLk8AKRr3LLf6vOtw97+gkFpZW2HeftZq4Lj
xTtHGoWenSFc2PHlwlHCGIe3EcLwfQ8+06q5VBbc/fd8Uig0XxN1KYkoEbVOiwHobZKRbb1rHcvz
bFQUcFQ0U71uX+KombVxryzn5UDVTl/jMUljxEQSxcspQJ/paPyxWy1RbFZLCZI0vR/Kli6aA85V
dl/qbdqBTkZmF5IEPrKvTgf6Wun9YCOrQHlX5tvjmboz3VSHHwddJkJsAAoTQ1NYz+sw1xglOw5n
HcadNMA+XC59yvrVZNlGSx5JHlaqcwT6OuEhq8Rzpnf902GRL6WUgiGVY8ynNo9P2/lwAW+M+oof
CDAX+EM4+TVtp+wISEkEbVLJY/RUqg2l9m7s30Z9hmqfSSEaJrxTIZygZbp05XGZvh5RIpyEy3dW
uWLB0KWnDcwNAGEzQKIzVsT/58QcEF+YodXm2QZ2F+ffilwADv8d2WdnCCDlUOtyCLsa+8KEGTST
kteXYUDXvZh33JfMk83q1vM7IqLpvODsVKcp9AJg6gMbGVHk/VpzakFPLECtTEZLMTJAbWWpfCv4
aBQxT8Iz7TNO3jZ5cFunvoPtn0l3FE3WxzxE2yXnDjeDwDzoLPKsK6NfziqmO6T0Fgp64ZMH1GcK
uN6FPgdKt72N+qXLbIRGF/4QHa7VPBjV2c50/IuFQ38IHC7BImo3ROc9W8prBQYQevubnJuvKXMq
iDkv0/S1Viw4dYoJiA/nSWl6ngSqDOdS91wsrukSh+kRL0gNPozhRBiuZ6HvwLo2nqQ4v8BFlVHB
b8FfGFA+Y0guzrHzxSTlMLzQF5NcSCyKHB5jkTllr3qz4gRizgd288P9bXuGCOuGT2Q8XgVJiAC2
N8tKzz2zVOBpLcrnKB3JLPs87WrAEch9QbA+aG4eNNkKrbWOCNz54r3kGGdz6zTmXoaZ2Ti3FZ8J
044PmmMfPsAhkaVJzbrfLR20NchbgH4W1mcy/U8OH3AvKTkix7khf3zpU/LJg4ZwSbtbeU1VVxZA
aZ2eNuILEfrNvVUj6xcFIQbrF5iXZVhiQaV2OYX8bLTk4kWB4W+qRuSW3nMAwpMrjoUSzNYEmN08
EbirLbOwTKa7lhAYBAPx4VU+7nIGUMlA8q+SVjCQU2yFhiiaOmgMCgF10H1rcG3C3C0AWXXh5fc1
kroF6ytj7jo7A11qAxR+dhAbsGxV8OFsBgK/yMMR7KWHjZkxWVOpSweATYJUVRHoUBwqiRKLR9wN
O5iVGSsQ+IYMEOp1PohSkSU6N+wsfEgSzgqrYr3DCY1vsiu9HG3aqXNdOdLmeMmsRXy9t+KgAh6S
qZ4RM97SZTG1gvmRRnSzCdesOCkniTuaFk5LhZfZettrIIcXvjBEn/gzdf2YBkd+aDc3VOkSutch
d2JsZb5aURj66VuAGWKDC0iUl+gfKa2Ab9clyftY18KoLohB+DDzEX87Fj1ql3UsCHNxAFj2NYFY
qHcLjvzMoRiFxPktnHo4luPiVLz4rkK+oio3E3jP+yPuewu83tMOQZxukkFLB6RvSiUkpdwNNbI/
x6xQzPfaPa/1MLzeh/C/N6QQVq0UAxq0a7rFRyEVlx3/9wycqGXTO0kUOzZ/FEZM+uYzDpNLpNVG
U7pOzAwa59dA9DNWAF97T8Jfjx1eIVfB2t1eQmNDo5C41P70fqJrtRJWoRqvHu4UdiLFKYMGa39k
r/yq9tFR3X9VoVzDVdruFY3Cii9Vm22CVmdNTlh4Svwrvx587EqgyivPcgFYqLdckuQBjP68Npf+
JFtqmuqgsjM3f63jfszZZ7HPdoZX2Bhhc5jYzEXXJgb3svwO79zbFSgqwX/hUe3A+/17ijUJUJ0v
rvAYjY5XPuHaFCYMf3Z6l/x1+D9aRW/rg4FvdMO7IBN23dw5cUKD2bLcj2VGQBmeziKpxQjtVpEs
IP1tRR2RlbsEbLsSFr20LJZJjW004qCVnuSRkqyv097d8aZL7bVbOH/fQWp8DBr1AVwMv5QkJbtu
TT3FlXV65PDk6mBoK5PtEK+w6UyTn6PN/fmMesDarkfgYbjecAWKEkWZ8WKXEcWoj8obymwKEiqk
V3uAQL6yhvDpTTOaYrNl22MCL/dBoyo3QUy59jcysV5iUhDi5gdwCY0OoaJ9aRcRCIB4wry/Wb0C
denfkn9YTAQziWEDcSSHuDgg/giyfCfdJyo86uzPLJSQu+AjYWACqO82i0bJqyC65w+pmOLHBEUm
CcB2u0DjBeLYFrrDrNWRH6ciQpDUG7fsckQ2LOBuUPo0AZOT1v8wO3QxwokCzhca2hsogR3Kh6UQ
Rtz4BHnC2P/E1B0k3ZSdz7RDkpTGR1XfyTveJPa33fQYMPH+jON5prPJ2BROqbqemOuHt9hGe7Ak
r9+pWkcm9Wb8iSlJnKxmBqNXu5PzH+99qtb0diPGQG0oiTChNER//pbf2sQaNkrb+B3iATYTXLVx
MofoQA360JL2hYdpLasrcZ0+Bhp5PIWG6tNYxwNIHmQ8hXejrmmWZDD5gZGxuF82dM5DoQdpUfp4
iwB2yQ6eB3O9fqU56YOHZcsBLgKUdhGHhls74lcT5e1H06ERmjO8r4bMr44pnDY7eYURTd4VSgyA
VhJVXKNfnTjY132px2dYDq+iKHlfeLDtJkoG6bVgCS4cC/onjZuO1EAAF1h/8n+0HqlKydLEqnEo
4UHfIHlAVKNBuugGUzdbsw/yOtMTeM4GqnegY/+cyGNgpMNaqmwlAdEgHtltJHRhcOvFQ7ZaLU1I
/JcbfiaaT9r41FO+oAWUhmZWPtFQs3pGwI81Upiu3mwRZ/O6V1XHUgvrzoPup/3r69yJ8JqGpOC+
eLKik5D939lh8CbGJfaiuxlilxz8oVdESVjJk9G55BermrdET2a/O6FTsB8VvrCa4t17/zbr+6ik
uRPBGVN3FgqlJUQSxtDVWtMnyDZguwGeB7Y5hD51o2NToP96zAT49yW5Yye22/h7epdMKvlWW5LO
3bfk6/Mij//fF8C6UdEtRXjkG+s5TQjcUFfBeG7YlYVaK8FVzlGNXDU+IEUznpJ5uhpxJbH4QddL
lQS9C1vYlh4JNNKc3lm7E8P7v7wQUzJLe3FyD2INPsMJdPzNQ5KxySN3w17im24bbfgHVQOAhhM4
GhGy9XEb7O0hFtmh7TEbC5L57Gk6si2mkAXo2cYwwChOjQseHUnYlXGjs1j46ukzAFoix0iY1+XI
+edyDoQO+D7IJfNW/lOSsvjaVcLe5gWuJ2eMPW72/YgDUfEPuj8lcY1li5XHTRll+LXE19dI/UgJ
Vy6nO72RQnbyikYWsqiZnX+skLLhDX4geh0srMWYoG457GNxeM7Mtk4QuB9zCXboFjZm3OvWGpqo
wgGfpkL+ilMcgpL2i0gd5sSQ1Z4oR3Dt7NKbcayptO/gxlDJWpbk6AwzOOwCB2DP2rO9K0dsLU7w
2FIEVpFCL+1Wd670CGLmem0RKCT8+dk5GWTTy1GmhaKgPGzEnTF3oP/0pepI9DFzXF0Dg3LlN4Xd
glv7hBtNdFKB+uzytOq9oyN7Xmi7/UAfuAVab7S6XeMqaZBtbo7/LaRM7zLcyoKXscV0L41xfVqU
0kdg26F+yOhehxktyCNhZdIy86mWToBQwgEmQCTSnh/j3da3LDLe8PbGdPuOuGucTcqjVNNrtjAe
r5pFlBO9GTgkwH2IQ/db5hzGyInmJQL9cTnVNr9bKGOl0Zwc7BGpIaGCJhg2osCk8ipXWvLtMWhZ
OIy1c7EnOcmJUxQSimPW8nsFXEfKqU48b3NPiG3qBpZbHbOi4I6CO9TSIE1Xq3imbuGtslHsSvj0
KADdVKhCUGbiCdKgulKdmzYwwdqJxPj9EB+dUTTC4ivdSqwfKP4WhDe9RwPJIMZAAMiJ4+hA0XUS
QxNAoYhn1yBcFGxeD9tpzJgkRH97XCbnuzQVRwlpeslRIFe3dI3YiiLnG63Rjspjx7w7jKVHjLZt
r+2LgfMqBJVljKMYjamaRMbwZ5vXW/CB+CN+l201dVbwOpTStMayaFI9huXkixoAZfLwp0s6FHsv
Z2eqNT0hoebDEIsTMiOMmDOaTLZwiBw4O19HymqrMw4WbUAWJZmmWic9E2K5+UoW1tq/bTw51Blw
rmZHvNOVx//1Q5YGPl57b9jH5/mT1wG2Xvkhuweoc7J6pa7Fi4zJkPeggY/Ja50tevpGa9zPaXP7
xUtrfj1uiseGTKdcADoCwKg0jkOmYj5CQ6t9Yxxv/A/1l8CmwcIENmZOpwruL7vAAvsMpkpKKxTi
bzUNwamvGnBfN/WGqdcBe4DsbXXVmoujAmUIaSD601JdfXQW2Iyc0OuuK3CVrGC2sTBZJZHD1FNd
Rhth68iKyTgXBZzb1PsABAeNKRuZujjPW0a3lj87jbgZZeeBcVpUgBhQSkuzJs+cZf3hwQ99HG91
qCGxal+7+FyNwt3RN53FNlVLJiBMHvwc+//nuEe4evxCgEL5TX2mfh5WzFi/R1mhoxHOnuabIH+J
Lymg5mqwSP9ogBfo9qf6WzpRy40HSxsWP5gpTb011mFDMc0KZsQ7AyCXo/iO8jqLsIRldaA9QWlP
g8PENH//7iPWtjTi5E/ZpObjus6TkraI3u5a30vPnUWD7LVmgMUMU8rqxbRwsV+6H9hkswnS2OSG
tZ0MZg8awYcADbFx4VfrGmHrrHXz/NYa7qdRfQMGjQIMKHlb3s+uLXKZpy64zn1ztKkDLvhr6LEe
50nVRg9IxxnsfA2nVF5U96gLSj6PPKn0CBDWRSTSV4PVGSVPwQI4CTb1szKocYfqI67F+h37vClH
yJBBHQdOn9SASssLIQWh9Hrl8Z4tkjesLw3Kjd9ed1CO0h5xvBDpClGrZXwydUV7CqIcbWpqULB3
8zvIunPtnPD7IQ72O/5v8tYEgPNhOp3i6ywEoU/N7NCB13e/VSgvm4RFHqblyE7smtQpTBevmCFn
X+smzD7AbRrNy2KPNfwzxnbfciU8ctsW/MDne0uDoCRGxMQyld2LrYJFC6p1yLUHzLCQhOjd4Tl6
pBc9UyujivNtLhS51U1ePUt9Ksz9XSOBSOJKgWy6ui1ytN8xgfNAsxUR9n4+CKYw8KTOdAzfwqbD
JfF883pxm81lJvMPYwx2HUSwVQnIMD/gvsaQ4GZP5d2DSfdZ6hGXsWy9BU9VpWhzlF3Ej24FyDV5
17yh3r8uh7cBfFmgoFelokk6kKnwlkveDksDOsLtmo2sETlhVx6kgM/sjhHbUzrRuxu2AyU3ZiVX
U3uVkP+Jb4rw6skqT80t9tBepGJOoYZ1ihKtMZmsfryjVfnoBIAtkbWdq3PHfYebYMozwcljs1GS
lE9uvsbPv62coQvYqcEL+bdJtHQ3g2J3AYaaSu4RZVLbYWkg9EJQhflFZVrjTQcXA32eFSeIXN+8
/SUReNMoR26zw7dzqsw3B3oGXrd2UkccNBil9l9VkfbKBtRCRnOtcYqVnGGbY1HUOgGLqotaInVJ
s2fWbYUloV2HnibDa5hH1e1oBAhj1euEr5KdqZTmGCb8Zwo7jTNxOFPMiqo5UpzgyKiBtABZApyB
Srtymf8hqsN2IbJWGx8mG0OcEYErwKDGPijzcF2Zvar5SGYP76rM8WtYx9546iODgngzV/26W+TQ
7EfsGd2AVphQ0xy9Hm8mMzdm+G8zg47l8leLejD3php7+tkwOJKRw+h8lU23qr4EEFLbXX21lxL4
YormTYfU4WW/74Ez8A3cjmmu2m7qdQ6TFWzvOAu8mAnPU9uk8yuC9EHAMWopd0xl2F5phHbALSH7
xeRG5r6ue0qkc/d55/3yrrK8nwCuNak0FupVGFI/D2sMqMAuz2epwrUq5iMcV+SlgnO5C/ELfXSr
Riw4m3rZWgFtlOwugYM6lvMYuvr3R3O5ofzn/lrBbyZ066YwgGifYmrD0/foTSn++Txk+5Wk0aKB
0rJe0Lp1XHcof7LDSeOyDP3FoCZkaOSKKYmOcDODZc60S9fjXw+bzTorsYgL6ZhYIpAzz9YtNQjH
A6OnSLdZkgP3+xmzsfOtsehVMigjyCcKj26lbaRSEUHHO5X+q7OE51717wMPmTM2LOrDfN/TePY6
Cju8HgoaiDUqM+d/woJRUuYdA7RJEyDjDgeu0NvatDEznTLwBtj1n9Iy2IXUqVKBJIqOtXMP2KGc
cXiHHf5RqSGTdTMbfxqUopB6jZaZHFDFFkiuvTShGpx+KhlxPuyXpSG5fWb38rtvdwAovC9esW6d
DAODF/9CFj/FPbq00TyPP6P8oChVzaPC2Evc5cdwsVoHw9aCFSOC9c1aakXSgwVa63/wIZD+aJAD
UnJV1Ky4ardFz53qqP1Yq405FO7yA/gBpSimoxZ6PT3gLw2/sDqsbqF2DkiQYb/GNiioneppFe7B
GEkKZSXWRM9XFWNAkO1N4pYDacsiQ0KltDO4Al0apd+v0jvas8aFGw05fOQMhd5lChW1wGxeL7fI
Vq2Bo0UgJnyQD8bW/nTIX6IA3D4G69VyVdUx5iUpkX2vSSaavwrXC3RcvVYQoySFXnAh0YI/RaNA
WW1Va2BHIv71seE8khlj4DAevNFhl7FgWCLD4+hnPhZO+QELqjW8vql1STd5mbeZKWIUFW4WWxm5
cEECRhcPXP5kT80mkWj2JcSmcWKLpf1hGVJiWnLLN9QuHzpqNL0zPt7S80l2c/oPGnXgjckkdoGN
KCXLpgwQ7Mrz+v7px1dSZ/vfKlh/IQ5dpAZDGFcHvX3GLrqoOOsgYv9c1sn1kZxXQA5bo6T8Wz2Y
W0V6Qpu34COyClWT/sQop1txxrzV24dDft+A0Nz0UXgHJ5hWR3ufy1FPeBdEswEMoVAJ4m9L96h5
IZBA7wFeykM0VZzXAeVLXco2y4e5OofqdzcDRh3Rwn4pl/G5JCh+ALgP20DZ/4UEfeO4kKNN96Ig
GCOawILQIWlKzkVArySG8cDDR9GeIcJ3w2BUxk9MittxUY+kCCK4SGpJTdc2fCCwr9Or/TkxpWIC
DdM0avmoQDPHhmBMCddrEV9WyPsmlpYzWLFAGh5yENTc5CG2jjb0siyThr4/x0ndXEmAAM875v6x
9+p5xKshJ/6KCeyW31dBfpqz0CLHXlAZiesgrGTgzYKRXJK2IBOJlhQlSX3CGN/R44gXjm1wEFBT
YOd+4h8KdhZvexFmah1ZEg0gGZ7DtXUwGE7P6fJTNIpH9/0aqry2i6fGACxS17fvNUvu08t8pW3s
hw6PCyu86Q6GWueV0upPwzpcPikMW6LH3r8M60oaoSlLV7aK/YlabiXcIX53+lD83sxX9zAIDMnh
HdO8ROc0DAE6R0JAq5MR1ohosxDXL++IzxbwIWnHyCG8xjFkjanscapG9oGSZmch/fTyEXmBA5V3
8EKlYXUhNdO1/xqHnS0vhnz1SqzkzWdzzfN1Fd+2CNZy8+EbvucSoIN3O7tMXYO4RSlFa+G/msWn
WAZrjxJaq7NwPFL5A5Y0xb7M1ZvSzvWZk6T2c3VxG4UODCtk55TSAKbAWRo1SFdv5y6Kft7Vv8Ak
ASJ+8kSJiFvDJTiHl9ymgI9ekGfFaIJfK1yQUyGTPRJezuxbPqLUfqgmSoDCkV/QDzQwb6dEEldj
+uJU2nVhOaolYRsBa6X6X39xRmxNYe1m0C6CMI2jhMicytKPMWmIEsXVk17yEwbVODYumK33oZJO
HcXqFsVnIK/8I4Zbv/JYfsnAfS4zoXbGx2UKywvmF2wNJjYwI5h9T9SDjaGG9+cCFvw0WbCiXS76
nS1BJZifezfWeAgmVhFLiF0qFLY5YqD3VjS/e8qUzroI7eWQM53OBaD+ePFqzHPo04doDaWp6dND
I3IC+rFSB1D+v9u+2kyHAXW4WS26lijEErc8dlmQFS6lzWcrrpWYgx06rMuAsHMtmEMZTSz9oOb2
YgAKeaHQEcdoW5xUcXmdPYyWgbbPKrUCqb25xpl4IdnZal8sTg7qXbpHwCH5eH5e1Ueo0Zjrp7OX
Krp4YpT977yNpftokU62cs5+3V3QK7W3H/7d3hmTE2jcCLCBmThWq7yqjIQr6r5kyZfuoHGR/nxw
/Q5Bhnm2SpJF418x832bF2EDOuV42SDoZZb1YqmgAngy5wM9Sko9cvcIBCztwH8Ch+n3kjugDuf6
/SVNkviEigYbCRBC1O4i7Z9oMkHPuYeWjSnMzIRfb4c61F9k6MWOAlAZdcxKG5//eBvj2y+rUKGr
1EbMnJ1axtzJ+nBXqHX4OLspqtPVCWMKTV9s6y5i+UkS1+I4TqkiOXt3YD5lobFD/6HbhoxJAfZo
WNj+KX3hLpV5VIXHmoQqE2LzNOouf8ULtkvkH2eQAXdeKsWcYHtWJC3D8sgFyKYJ00pM/0hnQkTY
oQOcM5YLFEmlD8phOOy7Q3YH/DYJhPsXIutkN51INrp+zc5bo2g1xF++qaHHzQ1klG9e6oRnLEyS
G8+J3EyPtxMuvcl1RjDJwExiEcas1sgd/sMrhF2StKZ61kwEwoQ0bs2mDpWLdgZKUh3Nj38xRF+8
EfMGLHZiPQqDuoJtKct5C0CuNCYgWw8khTtD5qzz6HLZij2dzwODxBoFf5CSEKU724mayJvtA3Pz
A2u29LdenR5GQsCPo6b9WlqBG3Qz2atqLBX0/OHBcUqz+RYCmazacIGe2xYYWWhE8BuELsRotml0
/zIZxCOGNNVMmbmAuxfLMu9mS2vYYVn1SKsIoHpJSQB9nWUd0gbZXDVfjlIvolKR9TurbNbaJsHR
gZeUu3fGj8j/bMGPUCGnxJsbBQqfP0OS28m+RHXY5fipV72C4MYislG+q/GQQEmhdHwcg3roJEaW
Ae+4aCyhZ31Rbo9PjoOxLV8ojh/QPvFuZ7KaPLad4YwvPExtODIRydr7PrFNdrpEPfzpcBSxWS0E
YqYPMl79yhrqtjE06JmoPiJUp1QbzqQB4Ws4e04syF7YIrOjLV4irpvtwKi028kPAIjumhjr/CF+
RsfalH59yKhxN2R4ZeNXE4hEwpA+HPy9BDuKk8/v8lktMth/S2fUwT5wgDDl1WWdhwazrVXpBamo
h2Q19LDeqZkCk2AKGNPotYitlhMIuGUulnIXxBYDy9lR5qTzmyGTvbXyDpQB1c6gbs7D3i/Yg/eW
TRpANbqGO3VHxnT38kQxDUc1K3n6HXjgbBP31HlffuoSB3XDMMBN9LpGkC83OE7mp3eOhcHZqn7l
Knd3OxIj/Ln1jUhIIgMrk4NbJ0viQihBc2I65siFRX1IkyN+iq+ps7SUPaNP+hi+/x7KYM3ZqLga
0PEahyuElNezT6MtFdCSMUbfU1oUuOjs7JhiMpRH0v27odMWhaeXjSs+pMKjiZljpfLwfUUbxmuT
9rR1skTFIQ1PKO63XMtrH2BMD853TyYt658C4KX5mMCbYgVwNif5IZTRUxaD46ocpY5HyhYEJ4Cn
rQXuHo7qvLK2gdYXXGOgyi72YkigMOAFyYyz0S9qtCPp0gSG5bWl5NGS945Bsv3BCMnIaQyZTTVP
ZnUo7QUzcokFccEjxWZAdJUK9soZwG+Ff1DWwGu2Fy73e/Bdqlc3SP9wbUuMLadtWuUpzrGl47FX
ZCS7hdON7a9mQCUKSQwJ3/TVu132+BIdC4LeGEr7uDl/+7KKcwJXxMV5yAwQsHWyz7jk0g4uclol
O/l1qpS55TVUStlQnFAkcRFOHF8xTJSTgxwXML4tcH5PtN8YAzyGLZOu0zs5h45mCYtwAGM66qhW
QCV+elSNa5uM3GB7rcgavEYRTasNmYdjJoDcs6K8UgWifF98cvJWXXTFUQ/PR76z1rtYLugp6C1U
PPCmYLp7m3bfsiUuuREU+8QQY5es6FrKBp7TNMG2Czsag0ANpZMrqSzvJjGISap4BbKVT1KiBoyh
GXy1xxMqF1edgkaCVgu4hxMOVf6qH0a7cQJEHpyiesw+GzXXIB24SpBdp19xjBRSjn2bFkb6fLUi
NroXoryyq/XC2vzBtDbWxz3AgEPeo2CqJC9kqgbnoTGmKZZ4BOUa+F6J7ZhaPqQG0sTE7OVxEoE5
ihrn1+Z9ggYJn9nRtlhAj+ns+Ijywh8W/APSVfV0rJXVmaQfjk0nZRHe8S8iZlLrjXMbHn9Yz8kk
ys+Hmd+wzNvEpYElcPgeb6G6cKn8qI0QCa6UBApn3Q2j+G0xYacqDvTXxkVQLLLYbDFEOmz/pOKu
MrpwXVl+4oPfItJUJsJa7MunpUlAqJFsoW9Ez11SKcO6qnII+hV0f5sKU7GEq/CcQWpMEejaaWpQ
bac4Rox8Qe810Dq9CzEvx1eTGDJbfnaGf7xiiRkp/I1m6BHNB7gY9NbsLWTrGME++q9kqrw8+zbC
Q/VuRAcKiA8xM11TFpyLnKJw9TFUXhDDiAqzoqA6lxdL3G3e5gCamXGkOPEWAoFJivrmG1AgtYDM
Fi6c+23NWUBufIUodMN4BNLmYzoyQgkdpQutICAIFtlFS0SanaGAjKs9kSGNrfIfGkQ5cYbqCJ8Z
C/E65uVct4IswcHkN+e9wKVT6tGkUbfZ5+2CE9nTG+mu9mhKCrnkwGDIH++F7p1uR69l2H8k7nzB
gjBHrs7XeJDMBoh0XuKRtMSOTi/9/jD9wWyepgqsp6LxWxhAaAxqebt2Qkbv/0/OtUpw1lr858FG
Aeqeq/tHOI0UybsrSTcedg7wgNeDx3LeFGqCBlunYHOCZlF/yb2GfNrgzn69vxR/pGuDsm3AxGsT
t1w4ILUhzA6FVtIqRGZlfD3ijwbPtgCays5D8bLTT6Fd1jYVJI3MX4NG/V7ZE5O8tKfA0tZ030nf
BAH0E3ibvCUhgP0A95M5n16mfmfHli03HcQOp2GYLHoWvGrIQ6HNo4BRr/airySj9tg+GdTtgS8B
rxe+nrDqEWgZHXcyEf07P20g3ZuezSLwM8Qx7eV3YrmwXGPXGvyH93rTL1XKvyi7XRoOUoiA3A4s
UqHx9js17RGgCZJV4WKEQHFE6tl/ZP2+k5udA4KyK2v+rhBU/eN3GCvUgn3fjV5ymKIXtNl05Fao
abyCuqpNs4SnyS/3S+tzrfTHaIcGnuJNQ04dgYKA8nQ7SwQhcCg6kPniWR8ahaVafkXFxbjqg7t6
XHKKxtQssLF7F9qFxoOb8TEKRYUtKFXTHrZpjmJmH0QjhEZ7ljOmKyCQv3wzdRLhEbmZbcWskMEc
6ZuSiFFA1Ci6aEtA+zBUgf1HITVd9J+d6sYJNb5io7eebx/B1HKxLFLjlD5m+flMupU0YGI0VBCu
/PEEpVrR1rtHK2wEXOhht+u8GvsNDWoQwriM8d40uAR/TvWrQWPSKy1G7cDO8VWOQ7BTxIlQstst
g9kWIYqAk5LijM6ZcsblYNYGefXdSVxnhGWmQbvvDrfes1LQ8zlCfxcSLpJ5Db1Us2PBPw25RyJW
PW4/yHBrvW6Nj1L4i7nS+Cl+NPHyO+ED/B6b+qDaGzieVOlX1urJnfx9Gfhwj0MdhV2w6mZM1Ltm
q0wAfsfrKsKtxzqwE1sfY5p7YTmCjrOwEW2OT6TIxnKqTVjx9SykqSitevSfwt3xKxKOL07v7Mip
ovStza95MFXOIAMm1TTKbQ4OpUzBgTQCXoHcaTaKp3EdXo5+vI5qZxXtEAJct1nGCzIM0pXMl+vw
OyDlqTBS+8zIuiPBjYJvJVOfLUSSBFTnKb6OIval9h7ZQBz4M7hhAQ8KUzH7DBLE2pgZdTnMJSd6
uL4WSpMKfXZUMQS/h6iTHzpERtdlfpe+n2WVM60KsPG18TCnFokm8rRLgGHF7IBUO4DcWeD7CauK
738H3jsKazL95RSJtwd+xZI0KJTWcJr5QA7PkwXyQINBO+Qg7mCX0cZdaHx8V3i6vL9c9pW9s1D4
ZyWFzhYp0/j0s8qbPvzUcQ5uJS1UfJUYPXMalXUd2yB+U6JPFyEG6QF7su+D5aLWWikdsXiypnw/
/QKCezXYGhdN2jY1yFpc92zelg92Wzn8QL9rFuZHDNgwHpFmhk0xcUTrMa6hs4JBNH/UyulCMnTK
RAY75XptIW4nCXSo6i2x68pYTXF+Aqn6euGP7xuYy8+BmNj9Z660VJMkP/CSNkCslw8WzaE/ked/
J7gcx12ceIz7JPpUva+tRnqoteQL9oITbB+8zYvnkeCEOcr8+LjOkUs2cJ4cGkkhMjQmUjkclWSP
3Q289EhAscyLqMV7B3A4bzmIVAR0Ee78MUKnFI++Rov6xphoc6T5K7WW0jOT/r8qU6paSKgRoAJN
5uRIs85kwE1HeRx3yUgZ2zKtHwjrNK9ZqFYVQ3aF/CMhVEnPK2jYXAkT3FIeyDjCkGXbo8p6FsGv
Lu8oRFrnHZ1Y5F9P0OlSirMbJnmQ2jAGEUI18G/820Sb8x4Y8qF5mGnAH23rkgqtE2spILvU27ze
66F9WX3ykRf9xWTL6YNUUeuNoqPwul8eOFfw30B4pgCw/toCk1EtQPMyVnhUchulMG4Je3ILWknu
m/lK+qYk0BfMuUgTODFKJdVHaE0caDHaX5WJz9lW899wU7o8ALTfLrcTZyQoUh853OJW9in+buLI
pjKnH1GYt2YAxm6N3V/XDCit5SyYhxpjLi60xdoDd2CETyvjKlCHGmzzemmVimI7oE1spXTMz8md
OqmQkmw90G5aE8IzgbMh6r0gyWvmQ2X5MmASVeMoAwKrg+l36Vh+z6F8nGWll7TvtPFLX5ZgxQT9
gExoqu/WRy9tWASXm8jFYZzk/XcHpaMJKx6fwRYLdSnFZwvxV4ItuyVG/Cm5RJ04nkgPz3vU28+O
jb4tf6ZH795HfTSJbsTjtmSi5WgofmpCK69uzYLy5o6V1jiXkehdC1WLI7FyFlAvM9zSoNrKoo3C
hniHp9iwlPSRC7Uiwz0Wm75CgP8alDxUOM8d2Ssj4acB1v0E7c7q+fv0JcLGau5jjvx97u6NmDQh
J/u9MgoUJKWyma+BNMGmJ/mnVkT5YLh7JuokfdrLEvSTzbxOpvMJ2u6wZYPAXIwYw+pXqn/lsJDz
BofX6kSxupacS5UuEfdgB1XeejEEBra+wmop2ARyL4+YFPBGsJposMcIs5jc1owA0mZoMbGLHEJh
xwH8WHf3sjcrltLqCy66TzNp7n+lY42p2CXjj1DAxurXxJCICmUQ0LM2umjYHhSelwJaicF4FVjd
EtXqT755x14c8/LeCMBCWFb15qundHWr52i0TDk11EQSgHaVvFfTfB+/+4/YZDvkbPMQnu4EkDqX
Hjc2O+gHpLiLiOdYFPs+fP65RuIqPPMDrj22vDrBwdyi/KMDKmc6CvzR7Gb5SzhfnKVyR104IzFi
md9h8c+3FDrC1b/vfi74S/L+2OqCxnfxYzViMT3RRl95+ov0LkfpC69YAZuLrtWcikPYg5hQMRFF
f47dHiTHQQPWARxsjLFG/jxqEB7aWak3BnJEKSTvbk27+DGGXgNZOK39H+2KiYJrdSrqke6NWzTN
TbvqCDAGdWgsFY/i0zAqfVDXAtNMepEYTJX7+enKfCsQxGPS8Sw4L+ggqoWdlZM2DEF59zANE67V
B55xattF4oLNOCqtR2oncmypryhCLPXZ2fhHXBFbqUAwLRDEUpvk/NzrOk1Whpxr+FyHfFHhHnUN
JeBpxFxJ2RJbbSmTTp5wpKiiV5TTiWn85MxRrRRpdLY2Jxi4orIfWXskTflXdtLpYKg3Cdm1zXbx
NxxYvYC7OMojpjZDeCfa8mSUelfYD/hNZge+YoFM/lBNGLRxz6wPANnQsqRryb4FxF5DdEHvjJa/
EkNTckGDNTbnOis5kC04qf/xbIfFcpagZ11bkApMTM6cRP5kAoo2qFRpBCYEV0xNION4Q+O6UCmv
FlpuxMRJaRSJLkNuCh5KncnHrNecDGOFznyXAc7rP5z/RGxxWuAmlK4+CPwZbwKMk7HU3QzFWRak
G9opLJwcYKngDsaAfDVCfcCw2gzPFVjmHhiN2HUbL5I/KoiBnRgw85P94K753i6fJ8AD9fIgB4s5
ZkabmTNNrYw87wfyW6HAUA5YRRAx24mIFkXt4faVnBuENEw3fNq8LWIqcxJ9HlXAqhfHwsOTs3oq
5PnX9NSsyy9uVVVfXBtTpdznzLlF4ilylGNQlhaSR6vcCh626j1QdCi9cQJMnm6XBx3/eYvtWLAT
8G4irZaA8lcBRYDUu+t9VCdnMg855gBheczj7Yok8MHUl2seqqkzJ7hwuw8FPqRUs2tplMzzqhjk
4nqhK3GYMwgzO5Nhz468BWb4muwNTTLiBqi+G8G/jMQSzIVoIXO6wx23G1O1gel0qoNAvjkiBRKx
91nGC9pwwdVn2tzcylgOywSLhwIib3h7/VjUlQNwMBJxYdWcaOdVNGvNkTRyw9Z+h94XPiFGoTqL
2aM4HXkFl9KiIL1FgFI2A1y3iHALIVlpjVe6od+7t9CUu52DFSPFPmswA4ah3oKmaVHBWs8jZDmk
CpqCmQFi4CzFxxDrEXyeKS85GNO/lOdWK2v3hLj5MsNwgbK+I4EYKPK9LMMzh6I9W5VVGxUSEU1B
SfWo/8PpWJWQElRyPtP1i5fTEXRIyN7vcBY045yKurjlbUg6zpfo3mNrBH9LwA+ZQoBV10K8EGHP
UwmI63O+g+ZTIB2VjpkeOO7zHTqudKL4SZxlWaJR+tI9+ahuzaGmckafoATwX+rSIc1jOc+bnSiM
QEur5NyRYyqRQ6ETnWktjgWaHMOmWSdGtRJ9b+d7bZWHUEyaHDTGg+JgelxFqIh3fAmJ88mpex+h
chp0gM+H8KdTiKBg190ZKe09PtmuF/yitHjX+o6ViHKO+AoCPjn3L/aD3auLxNMbXlhIL3Y9WjHO
XF3qaMtxGxr0gKVLiNXq5NwWEBA1g9wD50fwDEt3Ugfyewa7F1vM3tYL5UfocSEaG6g6/Yoq1ceo
3fRb3XZzQSAQHkdjKyjrz6mo67o5ioaw3YsASI6+DPXOkb5vKbjJmflSqzjsrzF2sWe2tJOnw9aD
tBTasLANeveWUPxR3olXJx0OlAuGnwIPeczoJs8bp7YMerfRg/5NckyZpTjZSU4XcftiEq+BzTXv
hmegN7VmHToHsVneaGzTy+fvwOaJvNEjyggf2G5pbCExzOC80ibIOfiLoHqSGfRA55Qbnm1WXOuL
Atl6xtWplb6PgHsn5RF6PX13ckHVwfVXjqKJ2aKc93pXNZNucrhCrbNmSN1Wz3dUhyu5v3eNGlIh
lWrgWQTFxCAfjH3eLKp1myHbUCC01QkC7sApVCX+/e/MqUDoejm7RG2Y3pXwsB4TbyXIl0fQbaEu
VM92jcIUoGNNcOMj8urF6bEe7TqPpcm/inkro9S2fIXHrztJS/1jvu0h2PE4kNQoqKShpRYgx6Z2
YlYsWcb4d1U7HDmA6+vrOT9hY4ePZvh0as1SRs1TRNsCo6yOJexyHMkbq36TFWSoNTZ9Gwwg20kq
Qsf1/JHUv9pE/jb+tnB4Cnh6iCTqZ/2C59TNX6MKcforB0sPM+HUlK2iRuW6pWyFEI7PALX9l0gi
3cvhQ4/rqV2rMm9lnTRFzX4YclF9Ud8oGHIw2cvyo39LRcsVefgmRUyTOy0R/SsS0TrI6jYkFoNp
jU3P8i59uTnCsBi0zJ/hcUuCVY5kCRRo+FJhLY8CQNA/PGY+9ySW1DUKu6imkG7fxB16eQ5dAtU7
JuddIvbrxFrjZY1PkorWlrA69llLj93YLDEji7LRKZA0G8Wf5qMUPFE3JWn/yrhVy9bprYu1gTur
MmCilnujWusiUfgrKSEQY0qNxtrxR+ccEb5WDrLJ8DFlImK6M1oDEd/xyV1mCZkmHxQQTVxumcbV
oumfZGiwwyIZUbdio2pEGVR1yJ1AaEAJ2jxuhHkuTXsudwYDbVJzTk1yeU3yLknH2l1jH9zsaXCE
NZ+Qeshz72yArpGfKP+EvJAu6+5FvNoycb2Q0sgl0+Hj6tCgvwirycOk7028eCK7APx0esQUarER
72ZvI1PD7p6pLibB9gEOvtlC48+fQy/Ke2aKxU1uCDXYY94MqAnSqBSCGTTCb3FdbkU/lcY5Pye3
sxqUOEVyhVa53ANWQ74HXmqGwsJnmZbu9+uhoblhr8oPAgCV4SkSvPn9CUJj1JRk91AlnI5PQjHZ
YepxVNflGr8OwGBW7Mukf9C+E45WTFjYo1tAKeASLOdz8gu4vfXPnRmwkgXDoHvqVi1IpZXE7fY5
hgoEk7gUPreytBAjyvyFVWVrqinmdzbhMjQisQXgCmIYvIvgRqH7PAU4MzRpb9sW314W0OIitbQr
tOZ0TzjpnBKwMDEsOcw+uS59YLRKmEUrMHVjuwNzrEW7FIFsrVzSxdmLKpW3NHJJxzUoftgTtoDc
BwrVdxASoNG2q4Tg3zUyZ04WA7dr1el2AsPwZ3PzEJo81pJNe0OBGko36Ns7bWQrxpaBTY0ndTjg
yqb5EEETa1lVJIt7m4vveM8tuxKb1vZ/joIWFhCk3Lh0Z1fi12MUDO7BPz7bEHlP+a/jgGZYcUbE
BvxfE7S7jJstqdrV6An/DTWNe71OtSP5IhkvkC+cbhpaLLeeqGVbaYzylkPou3xVewDmEoy8f/Rh
mIAykaNjWbJi3FXvKbLoY2AdHj5BhWiNLgyMgxfd5AuJUN6VjRl5pA2PS/Qzkc2CkO6/ftNrjzHQ
T8wL8T/4/khUmlL4FqWWBeE3Zn8LE2pcI8z3u/26adICE0MnmL1+YanuPxxqTHTvIVRbBLx0efSx
wqCWXfdFM0v1VisWVxzvS6G5qLohVb9ULET7/F/fMdtlMygaV22fnkYeZpv9USJ/Aik00hjnS4v4
h4CyVhf/HdDi/vPam4R7gQwT3DY5aJENIOX4l8oGJZY2vxD3jMQC+CnlNGy8/tXXLlMEghudh63/
kyd3gpsol42hgviRW4N4NWGf+a/MbiImR/hHuoOwhKZShdLcYEdNUYMjejjNXs/uzS960oaH68YK
NV2/hhBwNUhSE+7s4f9GTlcebcv6ZDtQUH4+/0aXjeWVtNUGUGEMh0mhkAdCKNrbyUMx5SvGXcL/
xIHjs66fFJ6QtQ3w6fBr5ecVC/oSyn6EGP+yhyrlHwKkR2yEaNmenCacf/exzzEYy+sQc4ainVZi
diYgnUkEKBi52ZnPhcPKkbSl+s1WW/Toilm/q+mXkltgs3jQfM+2HtYz7lqxVpWNgdutCsOmNPRb
jMgqFumFsAxnSNPGQ1ljWD152Px+aNcL7xdM/Q9WkCKzMMaOVCFw4CDTddD9Jkc0AlxUdZQpNTyD
zmQp5jPOtxs4F65HhqTo0Muax6XdfHASwp6COy5buN2UXuCKZnBl2QI4zaL76cRP2X/v4q7F5tkP
XYSTwx1mXi7sOSQaTHrXU8jbD7X63AXaMmi/4iYJ4i/6Sh1/t+SmgmAnhM0hi4L3a+m099/eh9Ce
4oNsxju4wzUevFg+ENJcL14xaf1e00l9ei6/mtISGZx9+21X/HDY+XhFlpTzZt05eUynNoRid4hE
CvoKcOfExYIqAPq5xYD5HTDZ1EnqFJLh6x22VfCH/D29ir11rSkKcMRPBhInFSfe4x/rUro0+Gxd
1xXTHP13hQHLpC8ZLPUePbDtewg635m+1vZGEINBUf+X/kQnSqDt0fNKh5hUJ6wO27ETdw/73O7n
xwnoVNnfEv82VOMypkDRa+0xVO1cVe6iMGkA9ClDGCtoJm8xMlp6LK8gOq2moVBRVkv2yhr0/0Qe
gtE2jlY+LKLpFpPXa64yN0igyZl/ELADbkPb5hzK+k8FxdCBgqiWt9baPdR+jyAuq0xd/eg4OJrX
Syuk1Xdm78YKo4M5Y/M30z4iVDlYbGxqsWYXPDO1Chz4e5uUR8xLrRp/9b6NzyOqS8Aj4d6nkbxq
+63berPHeOaEooJJx2WrIy2If2CVB+mQjyRRlCsbkLDUajDd7GLMOFTkUOL0nGR1B/Mxcw1ci/3H
PPjTq9Nm2rwaWUZVVUb5vqrX4Pz4r37Pur1UEjyrtd35+1o5tWHeRmwUFz6fDT1qwnFiF/5xlwyU
soM9ZWa2+FyLEfmVlcVu0LudZrRMUBdGkO+WxOZ5eNTtn7Zav9O1lDBErAYnIof4ggj11LrWi6BR
kdLoN/aGtdzzGjCAwhrgpX+jv94FblP0o7rG67o1fsAgyzp9S/YFYZtz8SIcua4pbCnvTNVHRPGj
F+75ZxPNYvnJ5wK8IbvrRbc3pne3706rZHTtawtMXJLngtp7gJdmqVNB1oUVNS5nTEkLLMc2qk8r
RB2im0b5bBae4Kah7Dft0Pan12jyIKQVplcJoiN3HVI1lPcrCOcyXaCrt3fxJzJl2IAkRWwYsgmR
p5Imguw8ogkkhwy79CCkLud9ljJd/EwvbYiZtSr3k5m4z5VgXMit2D4cYf2r19T5bjfOANIxNc6a
9cdS4dF4xIKlS7zLcfJmoQPeM197HSUzYjyfGUyXxQvC7SU10DDDkmfp3S2sFm8b7Q40LZujnCMF
fxYIg+GMWYVesjHJtWNqAG0Rnt6mMOwkCW5sGFQNqatdbeXzw2hIo34RxmQozsmYjOdL47eEeTfg
TmbU3dKfpFP85cBzV8uoN/Ku2Geq3KuEmaRfC4dT9P2VdxeLHJU3bhNiqYVA1is+sOtl2gq8YgSI
Ki5zncMjwzpHkPXxIwVPH5sxbeliCOfcI5G1ykH30ShMoa+5MqqjDDlMiQ8xbSTuCnnM5qPsYEcv
h7QUc3wGYE3+arx3vKG7enwoic1/XdcZUeL8FykgPRYht3Kjc0l/TGjqbraaCDEi5hlalg2NysPr
y6StBzOmAzfdEZ8Nycyd0jbdCrP5lee8SJhaqIAXU+DFLkhelyuJVmK3BUZkHak90nYjLdPMltfZ
BdQeawE9BUXO1HOk0coRPFk8A7saMUWxUTgUUfYPJn7IIv7erbnZYsYTYCy1tV9+zzt2V4/A3tGI
zWDrP1csXknvb0Pt2zjNFv5mg3K4sunKDXuookzazCJQF3t/bURKbV3wEciys3tLhWUeYfXMHFb4
MbWoUzkByb5CUfywIfCG4LfDhBEsZRkMJ4i6+ZfoMP941ujWbZw4yaDAzrFCbdN4GaTjcNezlizn
TkGs2raI2eB3y8miXA/Vdy6etP/eDEkAemttnYggp/bDDo63RchvE0vb2Q9NvI/p9WLdXC9gB9pP
/xcmz7w15Fdw62oCIAgFrm9l36XAYo4BUNMIFqcQrZgD5IqZcH21mYnhtxsPUO2nGTBPhEk2s1Tm
vc3sFZkG4NllPAYw9RKBwO8sg3xpYulfqa7I2G7KQrqmDrB2+EPeCon8C1LDSsiXr/QWMNdM34s5
DGPt3/6fmINLpeKz0d+Ysm9twzPu7dpJCwsf942ObniCcKOGfhcVugwRq70gu4zHrfQuHxZTFwd8
SGVOgwTlfH/OKR8B1FnSDEYgxiPKIggk4zynE3bSu2OxRKdny6Eo8FIP1Xau5HKvxY9tGsqZHRgC
NFjSCiR+uVl1NxC1AV8QT4y+xjzzFKik0+STZMTkC71wLd6C1s6sOJfjU9FAKyRZ1HDlgBeJ90Oq
8TQUqr4OtdVjgry1csN1qMonXexBkvljS4DWu74/Z2RolEUBiaBl1ZRJO5aGPSAL/w+12LPt+EL1
9EkoTeTHKETB++xQk+vmpBGSlmrif4IQ5xkyM0bMcsM+qlT8f04MUf1pxZdco/ns64WQNW5HhePM
mobgNAG7AzCo8gOQNx0XqnkcIYtCQjMlJ7b2zOfv7ahUdMkjLjV4XX8LM0ztmTY7LC35grA9LkbP
sz4BYSO/wvvtX3Z1tujxfj8bf6UfrLvZ5JrMgYBSavSx68pJj8Pi04nwrmpYjnJY2WwMYx+IyfgV
MdEJGJTR3Zs34KqjbIt8TsAaIbKANyoqCkDxSZX5V8JwmyVV3Yg4+e5HSJajEhEOGSpjrg4HW23e
GZeSLtiwMs9WNLfT9RFcilheXgIFWlARyT5g/csW7c5DxQsvcKQ5Ccsr0BaIc1a2iAJStw8xTy7A
QQ8eNcb2f600Y1VqvGsIWmSoYVkY3LXh8KddSsfbNIfGpDDcINAbQIWa8XP36WEd/6bHmAGKMTnT
vDkliHgAqtrYqFZ5N75U1t58e+ipSDJFqqTkOd2ZSxkQDmyk5EM1PVr5yGPKbV8UaX4cAYezn8q/
JcrgoL6PdHSCYbHW31Z1POhITDy/TnLCJPDdQfZcIlwQf+rXAmu3Fm0wBLxIsaY1/uXaU6w8qEyN
Nk7N8l6bSz9f4ZpnLcQFFYnzLZoAY37i0iOLDvbY6s0mMIEM2Z1xjCYCxWVp3dzIyRbbHuzAcgpI
/xyRgiNGjPHX32RLFFpx4Wwn8ak3Ezo66vOm+Mw+o51TidHTK4zEfhv6f45mEksTpo+M1uqnBRuF
TWppseQoeZA+IQg3ljKCqPT3h+G+4VAgvfxaO8Xr5LqAcsvC+glIA2+lTmqEljKFFMi4+FGaCtzM
CQ8CMZfC7frN4u3joMP6puP9/LZiXbQwNHmky8j6+G/06Jw/eF81tS8bfE10rUJuS5GBcX9Mo2mi
lykKDEZrEWMGPxxq0N9X6paHBeqBi0wr1Y8N/gxF0ox29s6jJ0OQDVtI4vlf1q1Uz4AsDoBKL5jr
fzwGuyvC0QLif5BFIFUsRhvzP4ka0knRc1AijZRq87jF6IIX+i7tprz3ebY8NCw2pE+3Xh4WZ5Gg
v7d3ZIv/NCoj/BT2we81TXktB86mwU9JpxtXA8ui4r8hofkhxWtVpaGeWzRnZeBcailkpeMzgx+i
cd7b6awODtDxWWMXD6dB2lPv6BLWPxDOOlmLFB3SnTzoyx/RCX5jVCjMq7txoCurfzj1ZI8KTEAN
tVaxEwxj4IJr/++FrwRPgyITycSKKQLjgnL54GAZt3P/IFK3oRiCbFld2pLDDoYzHN+Zn+mMqD6G
pcBegT2lV154JjqNQ66wD7VzbirA7fOFRhNJ7OtXscPPOEmmxKnK4j3xJwKY3LH2GlBLGTEVnNCI
A0Gjbk1XPi+kiVGq+GDPmAMxDCIiL+y7tVrOQ1bH2CFn9MKdyVxw1YUA1lmP9HJ9r67mARMaOcKD
reP+hVU6aA8z7aalCJgj6Bm1w56MWixuTrY2C+DEO1cr2WJJppNOaWrIBWSAwHbal3TcLjDCTTQb
p4WksADeAcIwpPjhgXf/Ut/YwZP/ks0juvkcIgEkOTi2y9Uy8YjgsUSL4SpgoT6yUwiTvbmc6cTT
v12WgYBN3PQ6RARdeX43K1Bq2xVhBG7sh311ysw7ptT5r3IZS30yKprEoJKigyU4gtBOQE++m7dA
i1KkW5nIDstBRaaBspkdsqEyT9sCMHZKLleCW194cy4tIgGGrE2Cd93uByFQMMAZ7BsFXFpV1WVK
xcPVFlFxDUfXwvMKKxtTEIiG8fhIyniUOsb/zcMqoPYV48+nhk3s3D38q1rUtfAIlDiwDIU9eRzO
U5lz61bunIgdm2WuUpko377BtOBlQlYA0Peq2VPgCt3jYwlRqLHRby45mFjVikMiNY86o4E8Gex8
FtcGFRvMo372SWv/tZGTbkffSuXpw28J2L6y4qa6jDFI4Kzjg26C3pwZLCuGaqnJIVwrnd5I7eS0
LL4jDy6AqWiUHOQm2JAgsGoXVNlLo+UwPGMDzPOB8vFgbWLcP0ga6adejn2oA4JGKrI4CH3PRaDr
QoKNeEZ9irEIudkSaXAdq82D2VtqK64fSdSOZ3u3PD6FK90PlAal0UEFnu8MHfFOTrzVDOqKv4mL
zfUhQCVIENvLL35dcLpc7D6ZR1kjHvfC1l6ch86AoTN7Q1zwwR7NFN5udYFc8nSmdGtiO0SeksL8
2n8U6MHhMwd6o24BY43015+2f/cBqu+WC6F2LGNN21P62GTHsXLmUryyC2M8TLOh8444oRHS3UDO
ShYONHl8q1zzRAUR+Ks3UtvzGHEl4wDFNyyTOBV1dgorR4C9IgjAB+JPffRa72ns5XwVGH1+gsA3
B/gDUweKNsja1CTvEPt7Dv+mLd1qD4xFblp38W5D9gXw+LAHigI/vsvjvyY/jyKoC+cPyQibDxTC
qvQR/Q3yUeyY+jjf68C5sXHHYNC0JU8/t42uNnmcRgAbncw4GVJiiaBca1V8a4vHuRKiWYYUo+pe
sYfKfhcSDpoVDXwdj1hZs0D+ybAsYKCQmtyNQgYoTG64SzFq1pjqVHM/oeQI52Jae5WpliepVrKI
S1L033QwNdcrkKLo7L8UV9uTTiKUY3I7Bnl8kiawsVXHFw5sktbdnLE2tL4dFRuOL1RcEC69fjmK
KyQlkoyk3WuoBeUlbVSmX8283SfXkRZkJQrXxdeqZcAK7VDwWHqatRfMB3AafbwOar4qabkZIGrw
QAunbi3lNMZLYXqeq0OJdinQy4Hn+ZEUgNEOvt9WyIls9MVsXb+/RKkraKRTfZiF7qSL6cFXhwAA
L2qbZkIsTHHzayhTK728xxxvJPutbXVNT7NlFKnYI6FnxlT9aGFLDt21P/69fhrS1UfWE6XZYLkZ
2Y+MBZVe9MlWJ1Z5BYeFzEIovj+bt+I1BkXZ9gQtpuac8CZM9w8tsgfxqWvgVIZ+OrtlZN66cmM7
z3YSK6rdglDarfTpNWcOzsganZk4NxMsWWRBqGtDaXmLgzRWXT8AuGrzUgopM6U3jGYg3aGslCW2
P5N8NsbNXu6TYBuw17mp2lG4yjAw+fD2c/UCNwtcIQ/eOd5Mu8L7VPmvnFzeziAHmI+bhbtaeF/l
/0BVao0fQQxDACMdVkOzbvUf9gJzK9Dea2JyrI24P3oCw0+RZuzIzauLszr7xUmMteTGW5sTNx0B
n+UQ5+3TlpbMM8woSofX5Tkl/XNAHcs8XKZbZyKtcKw7x0VzUZ85/GYxy+/IoNBxtFVslI6DmVDA
cQWUEnsSa2ionRV2xGzkMM92LggR8JUKgZ2Y5T4rf9FjLVsjzcxDbNPAF22+1qWnkyRuUdnfmwNg
SiROhg++CpU5n0dyfbTKLkADbnu+/5Gp2JrE/i0Io2rrMXV8Nxi3Duw4Eh30+RA8ae+XtL08nW24
Tnzu8yw9JW7mOM3v4EygsjFp7y6bIR5hdnQvMtk+eBdP0bqybyuYeXRVUecLAiJPeZAD+ikXxBEG
yrikARjg6I4b9h1Xlbpg1Zg3AFpbznieW4IglNuSdKZdua7wi2kbk+DG9SBX2khsBPkEtxHUYbit
Vqm933a3qud+1jHwmC/Dd4IXCBBYPHShB3Tq/AOOKvdR9Ro1uQWtQLIpojzNJ6JbGBH0aChhIbcG
+YMB74QXZNVn/eW8MY17LmY85PYXnj6/hd7Vq8smEwi4nVOId2oVMxu1FnzTxhSmYB4foxN07JEh
LksUdnyY6BLQVKLXqZMHy78rbFEzPyWwB83kGS4+0cXmpKIxyesyDG1VeK80UAJNw19900T/5YFH
uw19/LSmN2uE/mlgxVIQJCDuKBsMTvY+sIUdz3PtHQ/WNJZ0g6QvH84EPEQi7/aFMdSvFMYDOqBk
ap1QA+sPiwnxH3jgsxhN0H3JL2YXTJ6s/WtzjdSiCtEpw2xg60aJS2BsoXAJCYj5qn8TuNs565Yy
EOyGh7bpGQtv12RABX6WiYheJZ3QTj6MQdk1KuQc3IQM0gFWqRUUV+wzreRG667zvTZnZoErS8g+
dZq57QrnLaFMxnCGQgGAUZcxoRkj/oNXmrVaZH8eSRjAIp7mJTQdrGk8jfgFRJwsd0iwMOv7HoUB
0W5zH67Uh2qHJzXUXvbvKifL/Mo0rD/vvM3NjK+/a/Px7aMvsblY0rmRXezDxHSvdKubt18iUmbr
2zE9BxiutgLd9BjTprXviKUElhxg71V4izSeL+6WhSozSR+oqsDCe2Wtw2H90AKV36Trl797jk+5
nkqGfyiBwv6WL9iHXx2BepVaTBkVCvX3wX2koBaMFrzsQ54KSf94eVOIJTI1WfAOsww5wA0vP9pP
rqJL3T9RrJSujgp6GFBirT6A/qesskn/v7DKUHWrRSadzk0XaIkpN46v9xst59U1YqbCbfQcMYvi
7DyvlYMAL73fGkATWaySoZtoRgHPIt3RZPmSCJUC7EELfWZYKotqeWKRi/VmjwOexDNwckZlPNC+
/qjWPByPPTGvX9OHJSjiSUiJFJyPjqAmKagJEw9udka9hP82ESHgdCE99BVWJfh0uoE3Dh4r4UHn
dNzPuUdGCrBj0DJbeEmXtdSZl6pHvIAJ1PLYQsJeNMguTdIBFWTrkmsfH8pgvc3RaNP6212lir7v
jMOHAa3LrtE4vbvL8acx9zpjVftaiYXADdhTAybXoknIQrbLWS0SA7QK3AqithvtFGKCIjzxx6Z6
cio8Uo+eVUYrqQb6L26+/sOVWauuaaFSvTj4Hm2I0/wi7EmjWt0JKeI8KMZx6qm+/oPYtz21mW6G
lvZaM6WyL/m5HZDh72fCY13GLxfQkhPW9ABa2x57YqWWc0wvo/JQxrmGtP9tacg4aNO7HtcnUj5a
MtL7j/BvsDAI+rRkxLTO6WaWhvmjjAWDfRoOyvlfypLY6S1BsXqTb/CBc8jm/9ApTVTFNFnGcmpz
9FbQ+xAzLbhnZDX8LI9Xg+C1IJZ7Lra/WCmubpFb0CkDOlKCoFjjgD6xye+/4Mvq8vRwbxCVJVQF
NJn03UKCJR8sbw6/QDhm7k0uRvprvnMK7mgeyqVg/IrPBaj+NJ6e78KtWEz97ua1+19Bzl/7lXn4
DKV7JRacgLyxGF76/Ng1y9SJLmXBDbI9mwKMu8elIWVIi4W1z92cbYEaUSznHAPvUigiM0bV+ECW
MOZeTgN+OGNGtRbrpWqn7TCBi2kDkZsqHjXL3z/qV5kmKXb+ZBzSyGbjRFpq00frvWk11nScjFMg
xqn6Lm+MeYjTz1Yt1mikLi0jmWXvz8iFi8RtJrUyodg3POQX0nkGyzWfq7VLqTpwUNdkFvKh2nAb
110OqiUf/elisQ0AIW1eklrtg00oJX+TYQOuL2fcp2H2Owf0jiMoLfQU0UYdN+vbBWfSEtxqB3QY
EwOXtSMRsMqnqbPXX/0UgPcdLbK/bt5+RLmwqK6KGFqdi8IMcSEJI1/k9STMnZfhphCQKeXljeJe
KmO6LXybJe6vGZxYIzO10zuVNoKaBPGMukf/JvfluA4GKGsOMPX1vSsx4pNhS+a8O3BOB7vPD+eZ
rdrHPUJRjFJlMJfHVKESiDxNgSNOlH5URSJuATofmruTSrkUySCaBVYs/OSp1komvy7a5QpJdX5r
TKTzQUEH2Nvy5TlVBSTnCZryiw0hC9ObUDNG9qaoemseWKhN6KZMgNKnpKvJ0yb40iShTTHvOsoC
sZLA3GRk7Rl70OBTMTpeqzM2RoeXsGTuk5OMjYQSMH9bfTPLKVrlXiRmyAi6eTCejOldK4dX9xwW
+DDsvHTddpK7SfBRbcZaZE+pvgO9ydGFDRHC6Qe+88IITCCbi8706dDxkWw0aJySTZ4tW61ZeJKh
TWpi3kkketuQLKR3qBGWgB9IpUSI9jGORvBh1nJVqZsqSy71Tg1HH82kTqptHdaOjnPddcd+sMR2
l/jUpsR1R4qwRnY0hgsveJRIV/d1FNsd/Y4fvgrExBSUTrAkMw2ne8djRPWLCzfCnA+vewP7k/SS
SLkP1xI/hxaN8rogG7BSiGAxQvcK14YNZ1KYpmfI8d8XSoiHCjg/SnruOpgA+BlgnAXKd+GBMd/t
m687srfawgb+vSuOFUKJatUqFCz2DwVirhed5lTjajsqk+E6JuRbfa1kv3iTxJozt1KjfTPEwoWj
tD5bGF++BigXBQFr/1A6bTdsUybPrlpYv0nraDHSaZznXGRJcjCEf42Oek3oO70aDefqRSBUdtog
wO09LSTV0qI8VOd1Dwy6B1AHHmQMyjXcjkrSr0inJA3x8ripkMV4Bt7DumVyJ1mDogS3XAAXOEt8
nEb8D1atS6+DAENLvksDJANO+0JFqhbP5bttjUACaK0Y8WiwwtmXH3QsXGM7OlyNPozjxQ4WPggJ
Avs/GaK2HlWeImZrpcjh8iwGHlVh+0FdmmsPyFKzFz0wzbBNWaeyrRMNSobq2QQbAY3gWQYODPEd
/h4wpb+/FJePNr4uwfdInsTieczIOLvQEedlvWqBRb5jE6zgnsMcqybmPhys7KmnwOmQiI3b2xeG
eC3Ye7HqgEpsh/iPUkWBvi3G7t64XZlhGFWUP4UoiqzJLB2icNR8D+wPFRZD1ER1WDWhG1A2JeKu
A56qQ/Jq5PaWgwPKhsOrGtOedXvSAEHcqjUmWPNTHI0lvi38Zged3YDQI41Q8eBbmKHSHmUu6WiT
lXWicCBjNw3AI+SnSyKpKBYSzJbduky409HTSlqJ9OQUH6JWgNIYSEeQv31SHNV6DNvkdqy8Smsx
842re1wl507TxAT1W/4ncVMCK+WIyQvr1a3f14/0gXCgkFGL6nOAkou1mwbddDYbLBorE7h6xANI
K4nT2b+ZhQTpJW9pJOZx2eU1461ZdZHH23vXfrDEt7s0AHP+WJeXYEh4LE6h5eUOBfLe2wSL5w0b
nRJxc9ZJedo5VDG7M8KqRKFz93yPZrEHF7dRic6tuBmmfPeCRKSIr6wxaeaOTT/4stePXpghi5wl
jIHYInlfy8qttV0pcFSoP4TsdiH0yCaZZBykLB+6KlQD1BwZgE3nUz+7HXQVhtyIEB4GlfI146bs
8LaCXYS/b2Wg0Qm0u/Y2QvJ2mmzjPQyi2i9xtbHxYK/Kj6FwNTZdGupRlu3kSwJZbnWqbNKjpmLg
1qMujMBRoDWW53J4+zGFSXjp2ZvMOEfn+6fxM/HUrYo4+2E3B8eF6jAVcOx3/hGIGlF91U4C5ZnL
RzXzF/MnTziSonXLVlvacEA2752/w06v4VzWXhQYO+4o0qRgviNGB6vldDuTYbXoY3rQMFWPdn78
6qeCk7wcXUDKXtkFtUuLZJ3pNrFns6YJvxN+OSjMjqnYBwqiNB1J1T4YaOZWF8f1pvNrypwXarQJ
popLzgw8nsFnRRp8dR2D+XC5XoyZLPx5oyUK4g7lmSb9aAnC+fUriqCAa1L6as//PDS69RtLe+Y0
Ql+BdUFGrCk7Fhx2k/GW59WVPMmuUuF+GXrD0cuxqTHeV3hzqphFAF7UVXAJbtAHUAiWF58eQTsK
JuGmmsoEn7/khO/QGXi8l6e3IUawUyp8c7Az9awFUIuntGsxh7ZDPc/6tWUlxcoMD9ld7HND57sT
uxKnC5Eovp7x3tnxq+2t01GKLhH5YCc5RDf8n0ll64l/TuIwLerjoj5t1dhNvJ9Voau73ikNOplx
8s0UHVz/UG62CmEfCG6lOKJ+4pRCnW7UVKiE3nWsKfObJGjOPZm7Pvdzny3Az5IOBWCpN+o+/jIa
doszUDgqYawSzfssgm8BivK3jGxvDTr2LV3JFTlMGERuH8pP67//01ZZ0k5slIAHh8aPOpszQ9CI
7U83S2VV4Hrmzum5kw2qm0c5/Akuuw4N3oB+UqgjMNdjb8VOA1pnEygTw2GE9w/HMLe4iPBDBZFD
JtPfvTtuTHA8WltSuoi/x1piLXNnu4LFIXiJvXSZ1M4z5F4n7K3M9AlT0uy4nK6TKQ+DSXfsqGa3
jSs57SdePDTyYpg9qmfmcvweUgTS79rUxbXe6r8DRffCOpUln+/toElirN/5FffN8EN9Q2SFkRpo
1L5tEMTSP72SD+9tu3xgasITjRFMUPKGr3By4vCbCIsSTXViGDhIlQ0hRUy85VuoBVE1VWSRIgR2
RKr62NZjmnAlylwRksymjWXOXJX6AfnQJk8QLixL7MkC4vMJcQ3Ybt49Gv93gM9aem7TicqrPxIB
OqBpw68DTQEZzdW6XSQm9qGjKPwWPJIZuLye4lXuQIE1QK5zLhSFo+zrNWKQOZGaa0rBjulPsyGh
wWn4T9STEKjYNsMM9GWG7BhGX4hUWwMh8qd9fz6BlUA5fYml1dYTnOqpTPuSZYR0Wcf7+e973Oeo
xLXwJcUTf/5eq1Wn6cqf0c+INEYsRaJKk6ajqEBLInrQwu6qZhmM8T4Py+Q6y1cVC2tCmj9WiTG4
qsEOSKcamgGM4YwcqVSeQ54ehzu4Kieqg2Hce9a1Dp0k/PxATf97dhRRKXSCzedxVHl4yWrjPXWX
kwpj8TWmxqVhbwhdFDcmp5JtGvU4BMtYIXkihnaP61lI5uTjraNcj9X8usV2jB2Sw7GYrvdqwjLE
Hd1Cl8zFYp9nfaBFb5gbHBfrVn7lUgBLkO/3lFDA2Th87UDIYEaLmpksPFOmptqFcd8QL0NQlq3n
Ai/F89ZHcRyr2UqgFXXk/2Mp0o5d3sg1x22+qTd1o2S/NBkVyIc+zoG2MiFA2s7GMPLU7NdJ2vRO
4ATc9kEVvRoH5/3Id/dgX6nWBrMdCkaH/wOSiy02pZWBWuqgjq08F0JW1fMpWG0/7QX6My13Cgtb
pRb9czRZ6okRZj0/HRTTi7F2bsZbcosJXqs/+A/HwAduSw1O3ZQkxtkCeEviCGaiNKOHRbsGubNi
nqkCTXehUVASrKRNeLtuhA7qq9ZIHyHtqIIt8a07YRoNh9atbJ2+RkO711V2t5KACXCnRfc1FhTZ
g/cYBTarFDJ5kd0QWeenoJcyLxAsBp/5/4V7h82Zz5OzlguWpJmXYkNZsD93W8v9j/2fjRO/ngiE
ssn5BqQr+ui/6yZyxs3deYfGKjI1ti/3yTaMpjKRUQ8OlZB3y0AXDorfoB7nKUbQpdTqrU1v0VW4
o//1V1RG7FFrDihE+vEB+quD6xXYZWqwCigxTncBnHiqKIlBDmeORy1wmAxvBdSgOjIu5Pg8I65o
5h7x5dnHPEffwZjuArovsuQ72zKgnjIEyq0WUs7jii/JQKWQ8vunjx4iMwdQrf5pO/ztof4pw1mc
6CMd1+SyKkJ+weRK6R+d7d7l1KbH2I0nU23yVfCzH+zJZQabjPMVpoVkQHtzA8gmE1oTAV5wYbXO
J4BOLYUZNnIPkzv/3kxF9aW61E49DJk1YlWVYJkox6y694qTCaHMp+vVwIIUcqpuv/qsKMQcbP5y
rBb8awsIphmnn3PLBtuxnZ8LxHQ0RkMh/0AkK+Jke58NSxS6AtItYKesgA/srCaCCtfvKIjhwCTQ
HxqbFKD3uS/5r4fvN+A6xp9B4fkBgWjkwP3MeXdzf+LrnlI+Zi53dfX7x31Ig3osB2TvSkGejVGv
7YeupgMcYa9S4hkxeMADh9UjCSe2Yh/RtPmdQlwIHnXgpxFcm4eiCQg8MDuu1vqhvLlkHpW3PLF+
LDEKWgSmZOu/YfZKvJyPGrDl+G5pwxnrVRBfJMgp836UtqamNZSYs01o7KYXpOaaJN+7477FhoWN
AiGcrBf5INTA9277ZU/YVD8JnnmN/JfGEkyZleIDSQaYAzsjs6AOc1pWsx2EiAmg3wNW996hipEw
APycnwhN5gclkDyhm10cVnQHQG+IXkCttfnrBoJ3fq4FGHlZEqoewIxpM+2ZMe+43Qh/U+sbOARq
AzzG53TVMo07bM3Al7pIxe+OTJi8DDj9F0wgt7gE+G0RqkuWll1pAnQHayUWL96lEFlcfVPbwu1a
kjvgCSyv1NCnMLQq3uqLg4fytsATWOaCYPIurYnW47YxGMHsz/bCoqunabpwBy0CPmMyaL7s7p/p
WUK60swxQ2VNMmcdAg3rN3gwnuLob9ZgmwvdQpd/HfbQdDDzf2+WhQgHQ+VJRkQXiB3OcmCRiO+X
0oCG/NiMF8gpKzHNon37WN7trrDNJX5cBquWovpG9WsSDSjxM+L0nh4pbGGVjrp9aeWarshy0OT7
JoWxQr8rDvveDjkgreptW5bl/BAQIQ2Cdbq6EFyu53c11UsOR+6pzsPV3Mgdnq+XsvRe++49o4sy
+r1mIjmDlkz66rKP6D8V4tt6vszHeF1O8eUuX0+nJLhNoYu+rmTXWiUOlAwvklPWsfm9qHAJ/aaT
t5/EreNqWYp5Frdds52JXil2kTMuYizxRh5Xp+R4Yld0TQHivprv46mRPMuUxJ8yxePrLwfx2c3W
pSYhkhGndD1/maqHWiFZ2yAFhCdAtqGwGFf8QS7DrWVCKft/QkcjlRjfKL+K8szEHeqlFS5WJosZ
Hk+9S0c8YsPA3DDZn/duGO+Ewm7U0T+fgFtVwAADkkqPc1a13W/9U2lMoDRPsGAwV0UzCwweVPLV
pd6ZeqYSgC7YUBRnCCiZik33XtPtFM2yOQHF44WdOOg++uei2buCQIoT50eYg8OTmFXIcJ7jk5fu
FCpvgp6/oTX0wp5jJiPaMYLFjMC+Vgu7hJ4pciQwbaavlv3FL8WjpE7yVPqG8n5ZyZiL00gMrhmZ
Qjy7o+lzVdnJuwcBfn4BclRRC3RdAljlH+gEqTfotNyCGjxkcwBwxwiyAhe3t1dd0rxahEgBxO4Q
B4LMZzcxXD1BVKVikvRvDt3hXEzPElnjQVNPpmWUf6Umv6RA6Y88h+VWRw4JzCoHhBQ8j0BzBJbs
qudvJSoVGI2eJf6uSO1zmVVfLgCJn0k3w3affl9JFN4O2p/LrEMttAsHEVdW0A1NM08BL9h4mX5c
mMTiGzhkDZUNegWwyoWAFp4Hg/+ue4V9u7h6XNxrk5RJ8N8aDPcJM3byZ/j5HG6LpTJ6OvK7bgHa
lBX/04zWznjpMNb/BEiEfYgbvNzrxRFbDgaqszBXC5SxtqUeqou1QaawClCdS8cfJGuI5KPF/qMs
ZjH7IoqP+7HJLXd7pi2zOkHRYThK71M790LAjHb3ATB9JCndTUZJa8cHOsJtgl1YkTwFF6WxTFxT
TFFoEZRrlN01A1/G34yiDmNVOXQf7E1zvvUXOuiXTIgbg/vEsSzhKoNpPrKAEqLvzknpluYYBlev
i/KU049P9ciOt6iptjF4DDRjF1RO3OZQXJ+MXhefrojy3z2xjYMfsnTRj0/f9YjCePgiWY5blZGA
X2/plAmDzCc3z3XqZ8KOjRpBcLoieKFm37ta9ao3/STL1H3fiEeQuBBS5pCda8s/Ke/9lscm+mWw
L6fhYj1l2iee7Q1KyJVigMAvwZYNbV8UTUR/M7xmjTB3qHqzO0TsJZbm2QeqDoNufpFkzS4EXg+i
vBSxXBucUQ1MAh2BrkuaLTaz9TkeB35PGlZlq04qx76ZNwEbTMgEENxs4TIS9AW8vKk/YYCUM0fb
5EQVIr+D+q1Jav7qq/0aqeovnVGVDu/m7mEg9cIvRoqxlz2EdvJ4BXu9R6qGwHbAS7hCOsTF3U0P
5jMlWhyVPZFNAT3qn+SWXySoFIN0iwTr+535sKNAe+UY4+Il+HSAQEUzQ6S8CrnIDbnfm5fsv3fY
XAURbm9yKKRh5bRrhzlEE6HHytPKS80/taVbm8SFTWEao4EEHTXy0Gmwsq9itIwkYWsfApaXlfto
bptq7AgnkjXUCakMdMZjPBnTc/bo0SdZRWHvXtu2sEdZilqDylC472oGAR88yMV7PGaeSvPI6YSG
C5VJ9MKj0DuBx11SOuhrnMwg9Ve1p9TqI5pq4jbGPdvP5S8D1UiD3+sQmwxuijBE+islXZ5fnVzZ
Q1QYk/9W3yn+OZYGdc6Wh0x8Rl/ZKTLTzulDUMpqIjyB2hw7o1cHcxl+D9STcMCbI4k1vuRU8UNz
20zu/l0Wp5j9Z1b1znsxZcQW8p0hQ+EbcSTsGIHK1iEXp9Vvqh/cTD71/L/rNBh4gXl6dJaznI8+
oEdgYQVBBzqx7X9WlcaPPn6p9/GhvXDuW2ckH2BZH0rBNcTpEJh+9Oc7lmlLEwksbISl3rAhFrOk
2IKDiQgRoXdeUQEBEBDOjTVTbJ3sUzlfwZ11iswp1UEz80btq7V0mkgTv7ZR7u+i8/dSlfpRp4+S
AtXv/L+TDbsDUFYUSKwyEg51Rmnuoy0HxMlzFHkl+ctJc01+HpjAdebl9J2QmbbRzOFfzaJh6LjZ
9wsQvCmDhYgnb2WLTY3RejtI7YgjYLKazQm2sK1WIMp+tVkt5o1y1p9Ff+/GGDJqCeDLGbt9aXww
yKp3wE7HCAdViBjBVXxwzXidkjGv3WA0JkFJYaRuB8KRPejchWM5AqOe1SNfLIX+XEw7nRP3idk4
cvmaYgBTNDqJqxGQVYhMurOhuJI5sLV0K7O8DaYvpMxaDLP24WsdlWETHD8N9//1XQgxI7pA2QC4
LofXoR+SJsUH/l3FwesJpVBsSIdj7h2Kq/PqFnO6jC52IbrKazphgChnHQJ3Amxs7DeAoor/sBDk
NIODzwQNk91lmmOXbn7VZImNXi1u43UtkkfPaPrXHtejzhKZvBBHjvBOw34BtOllOfGcMn0dcO2Y
1xipKapnWujJ8f/goLArWqEXGzlxhuSzm8Pqyi1ZEBk+YMXoGENLJpMApcnXuOOycNiiJw1FLeEc
gUiuDvcfXUCbdHfmKHsTE4TRS43DAPRJtwDmouDLNxNlcTGaDt6zXxLROmSH6SlfmOgXRAuqf7vg
kUnDOsOTGOeSmY6LgIE/3YejWMaPjHo/Oo3Mhd1sTJXLNkoAGkaqQuh4e3EBMVFfFXLR3IWnCRGQ
TtTnyVLb16fFwwhbW4GXYkxfjUDkdcGwkNRzkIModJn+RbSo9dLBS1IVgelPHrU4HhGZRd3xj37p
OArEq9T5lZZZ8z14pmzsufywlCbMtuLHIPz/UJI++6TwXIziCjbd7LN3Jzk+bUe31PBchEYYgWDa
nwvuez116/Wkwkv8os5AR7fo4XRIhCIY0niLtXQkD9c+qWhVKJuWgNnJ0ic9DcxWYGvRSAn9fl/M
8QuhZbayZieWVjUSyblUH+9xGItUkVnCwxC+nadkOYMjnfsCgRv3EPp+464uzftdMgPPJvxvcmCh
U2m6U5BypaUlpUBMjFkwpVtzxFxabDd5eew0SU4UBwh/tCMYaT9E6WLBAeIKnTqYboi2MpDfrvJ5
Xh+dO6381u2Nkzg0doKJrSq8fyXnjZ/yyQ9EGqQaRKMO9+58LUfHKcvuX6ULU0l2Hc8aoOBNRaGp
jTgwqGcKyV2rUyjbrhCIHvbEphVrv5g/KYvRf3XmmwhA0UU8uPIudeNJK+nZNVT4wIYbS6TQfS+x
0Jf3rpClGuuuIbDVqzRJuEtyctyt0WNjjcwUGB3RHbnLQWY3Pxt75A9LfZ9ThNI6pzAgAL0JWXxB
JaCrGR65MFgrQEQPVrTF31kG1JFFyhMlqo9q2zs58JmMKs7fFbXp+/TRlPN3Modx48ITGGZjWgJn
QrQ/1rKQcpJqzK8HOa0H4XtDrWdExxtV0Y3x+MrMhrXEhbFS8Tm+Ll/uNDsKFmp+WbpOU9xe9RjG
eNIE6hD6bQ4S6KQ2IjjeFsHAqxzySqdDQ/NmqqmYwPTK2FUTZpIO3T65FsNZ3pn826yLFgTQUndu
Gj8z0ZW/2CC4RQrnX7Xq1b8Jx+Iu0b0BBvJG/qG7poK7j9Y6SMTBBg9TTfql9MLy6MU3HDXsz1J8
X4XMio6Cyb8wiTzMvTD9v97POYuzeS2VcdEDJHmfrxDFNrY8Rzd+EYN36Kg+pzFfOQSCxkt1CdEM
S92r1wD446Eqo5FddHSTVo2qttjdpQ7Hf+PSr4qitmac+oZTa3BTtW7+SvpS5z3v0BS245OvN67q
MO/0X8zxmJWGaxPtTu31GpQYigwABryomSIBO8DogrSEycG+WGRc9hUzDHImcy9GFryxdynxAaWi
Ex6fgqdSLq9OXoks4162ClLYItm1aIlKOgrM92ZS9lR1IdbsTd3j87TcTLc/QBUvaE3HvyDbqGdf
ro28fvPpLRa9eT6AOroQER3LW6O6uHimkIKlotsNkGHuA2BsCqSndQXOcdMemgD4g6p0OeooVggx
JE6cHYZi2ufi23awa5e1QqxAN+fG6PqBPEyCtqGBfyIfqfWaIc55KTR0o87FE59n75AUOfhx7zEk
F9OTXkoJiw33suR0i2kTzD/41FAWv1rw1zM7hVHqCHokzCaK3PU9rseXYyC2g6iCZ9SV7J80yjMV
jJ8BDr4c4qVw+9RsXBsXqWGliCwj7uN8/aZxaJrBLA6z5kvb1Dxyw64K6VtS/9vEq6LbjtuM8m7B
yuqNIilDFoTxsyxtyhBwQxmfpC0BN9I9L7kaZmKhB/akR/lSqaPzV8AqmwDyn9WjTw4DyScHuPot
Kjc7L5kZgfP7xg8V8oeSyAx+yrop4By1d9Kl6e66xiy3SXtnv4sbupJDYqns7mdDx0LaI6JTc/g2
N2Ti6VBbeCD0WtbguCVWNfq1n4Nwebg3F1ME3ekT1vBHMRvCal0+ftJJWdIJlLlSxB2WGEWIc2sI
m7n1apOsoMvOs5mhVuBFh1KnwbKFmL0NbAzKLKcOQ/wgQa3annYYTR1e7LmECy4mgf69BpAPmRD2
EtoDFKgd3tvN11NiFzRznsnAQsoZtG58emmt4lOVipiaERkUj3xTae1QCeQyFGHwR71Ep5jK10OY
Al/SCkhUTz1rFq5MOZfH2z2+hmDNyOT36zpvuQpZ40X+gEUtakvLrf5HmJBLoBpGUVDxq6qVyZS1
70q5GKu4EEFkiiND4bRxkxin4wgO6ZKiA7DHM5C8fLE90F0PfljKAjryIiW19vCjvl4MKt+i9Sg6
dcFuCwlwyGQPxa9yNB+B7FqF2wTuIRDbAgDQd1LXst/WHDmMwBaYJmYzrciwiLRqEApPzs+Dsz4r
UYyPidHKuSNk8lI84zCQxj8/AX+aIKJxf+mvUDZbeZ3FcRpGSB9n7Vrcydw0IVMxvDSIH59P8827
q28J+bNaJKMoN4c8xYc+XCVtw6OtU2SOd7T5YOqrwvxo9Jms0ou8bHMD3kyGTJxBOn/L2u703f9y
ElaEeoLZeygehABllegoOzKvcE2qzNM7qS7F7Y6GzM6lncNgtMj5675WMHEA2cgyDfoUbu4VncY2
wFo4Q09LsrAv/ZuysYKccJMH/zCzeZqygowOvjrP/55tAZ0fDZPHb7m44Zw4JxlUHVoIa11344sy
N+IVrDL2kcrgJHXfV0WMAAeCAYR1jrvNXBvi0sZ9la71GFmAMqtM2BVmtuvInOJc1drs2THTrNXJ
z8BgAHORcCCQv4tS71WXQrg/APKAEU0TWliqWbpzL7UVNeC8Tb6Dw9mz9elXOw6BtQQO/cTcjFnZ
kJ7E7paOXoatVqEIPVLxC0ibxwT7c3ZciMgFVZpcp77c1sK9uiGVcO9NVw6SjEX623MgCReR0MWT
eGAY3J1xVRimcpYZNP4+LzEzDGJgzx1nBzzkL9V80tGRJUmDS2fHliWtJazLtSJw78mRAc5gWcG8
QZxto/tCdNGmY5FoGGi1kh8GrALhPvnh9n5iEHe0oul/vWlYM8cyzYNTbVgjaFllUeMPTyHsSwOx
mam3ozYL0I8113Wl5OdDCaSUkiGSfWG2yR0qzCrNHQABfXOQE0xHkDGpMyPArjwZxca0S/zKnZ8h
PdRCX3N/INM50YIh6+oPcZe2t0HeF+aI3P7LRwu/cJMjHu7xCuXoVbLmM9BcpUpQXn1izgapajYs
tUSpackBa1GI2WCVds6/0c2D84tZf7UL4/mPiobWFnCW953z59VUALzp5C+zTA+iOyzWXSW1foyb
XEUTNKeztevLAPAtCraJnIZ8a7BmgykEz37dAqs9KnBNnM2rNVwqOrQyAiTcLd6KJKXIJCpS8iVs
GqpfElqvjFJ0WkCcgQQPfzdR35LSnMe8aqx/8kGE+FiskqMpw6p7B92tZWvut/KMlnRFSyd45k/q
dDclWq6i6x7N7AJMFl/gtV/nD9fhrrGf6X+gq3+nt4GVNwi557z1vGZicWXyHqVdxQvv44oDQRKR
R+WYonDLGrxCpOohNsYT+Bkdi/RZDjDUeWZB2N9YIUUtdV1/ruF2E/hTLPMhVXLmS4dTsGyboTnj
LjlQkXh9gVeHK4DNDQhoXr4wYZO+tI7IN5+3rGT3IyaxQALD5hX0TcJ9RuoBfz8JZFTJeys7K1dc
2JT+mO4Kr76k9KR5VxepiNAVgMPtL5PbCKNTUrq9zMD2Ke2xPpLJklkn4tVqcqFf/trZRn0BBJ5y
dr5gtyt0KN0TucSqPKUd9EwkLmp9+ti9AMclWCQw0QxWXwNWibl2rAPzLsdli8kwegyPwS3h7lJt
NjsXUHWalpGOfY0I5ACEnLJFowSE2hpfB0idjQLzIENtoLGOCFGXWWT0zZRWhDDVkGbXyGv4y+pp
hMGv0pymqp10iIolfiOd1y8YxDafCPR9WzyDKB6Q5Xtna6sfFoVvJwZFWr31CHqSZRd/KZpsrhsy
xgF9WyLEh0gEdPLrSVfLewrqqPYXTUE6IoJbAdvFg96FjlUyV+MEREkFctf8F0RqNRh0Y/B486fl
x3syX2mtYqjdCNiyboayktPEZwyTwd5LvNcvtjQXJVqWXUW7tUlv/N0GiL3yZWO1VA1KRfi9Dofh
fmxuJuaFX7hcS57yjH4Ih+02A/p89EcA+/wNFHxM4t4TnTv1G/EPvB1vQIospCMM/Qk1BXmrsC5N
tt7BsGv+AQYR2A1i14flgsYXQwCkx+W0YxDVlPNFh4z5Mmgux4VyG5rJob3KoHZOnHjkvQJoLqi+
nXSrxCMIBV89qToacSZraV5Cy9gueceI07s4hyDbYEdYvHVFA+6VuyNArOdr3UKqMcDfJZLK16PP
MaqliiZITkoYewN9RDV9Nz2Sgszcickl0yuKBiD0B80lg8esULko5Isi/kEhEgUsuPrz4KKqZomf
okTCRve+b3cHT/aVCsQXVzmp/5dAcyof9V3K3qpIxxjvIWvt4JjRq8pq6SbVfKMA8r0TQVOsyxdw
JYObIeRVFAp1/X0HZ9aQeN2PsOyG6oVhDdyeT21pEPT+XhPeYd8nvvpUDmWoAWam2Qaj/ZeTIvNC
Rf3QZfbQhbOZJu2rtPo7lUyquIDb0xQPrcEJwOMImfmQ+2pRbkFpNQcAtBbbAi19HD0VEmpbmizK
1YIfvJivFEVrWZPKDbIkylGBk4L2OtLMm0jSZ4wA2H6az3cciMUcMw2TSQg3CSfSZXWx7SRKQWO5
28TOSCkSz4pzXc8A+RoJZIE3lnobYnmxp+t1LoJuBBSvWbI6q7HxoQL00a8ov+u+d8j7rf+4ysBn
6MV3GSsY/ja/SlAIC2a6xSpPRMJmLLRxsH+CgzVh9YZw3Mn4lGn7ACDFdYO6Z3gO9rznYs8Thzec
VSNualz6lE4pScVCrb0f2xlbzAncwTZeUsqe5WM2prKgm6UfG1v1TOUbvayLeaQJQWNOi7OlYqOJ
ZNqPSr3oEVJZeNyf3jlVQ5D2GSX/QW9CXB0PdAQKHm8nliirjeIOjA55778W3mOlPOxvyHcw4Gce
0LAlqFuikVAMn7QAcF4esIqBQ5Wd4YiE+1NvCNQS/ruV25X7kA4Yv2OrQXDF6i8Jda7liz4J76Zx
noPZPKqk0E37Ho2YRMlSQ3KbklfZ4g/a/c5RLJGIX+r/irnLrGy+jx/OvQLp2AXuVUpcGsX0I//0
ny2CUReZMDdNfqNASJd2t7GlSDxBP2PNh+kkt9I4oUK4Z1uYEHc4iFTnfXBaCttUUJaf9395d36u
ifzQrmQpNLN9qgoit6nGy5i0WHyKYe2uYIgucbSNwtjZC+Y3v9qEERu1GysrqkyQHjggiIx66cin
G9z0g+eQ9L9luuVzTkaJ0idORThcWo2XZ84HQ9SxVeCX489KNBh7cG8srYt8gNhWyxjYFSE6i6EA
HpeYDZ1bLKa7ueLU6N90gDbj9Aa5okPVHaSrLUFdRmQnbMKgY1TLxHriFzZDFRYk/8EOQ1sniCJd
f8x2Frm0+h5V0zs09Updac/SuszEYFSBx7t7xrDwn59CKwSKPqAoG42ROQbwNH/XvwVOA0IbYIek
K1wvaAX3VnVsdpfnArl6lB4Nm53IjosqqUUDtQ00+kSibHBp2pDnAjsTEoDlFL48mKRt7axLd+lw
7M8AocqlDUIK7aRVj2QsClw/+6zeELB+GZMtKMZaCsuZGUsa/Nil5EKpRLwPoQxuAOhXa4Nc2Fol
JYyxXQtVNj7UTrgmZWqY+gGYP85amCJ3d5wV+MjMZJLtPcaorzG/aUNpWP5GowIb8+ogJmNgoxLs
G85jJIRN3RDiY6KMW9WzVGwl7TLE4o80v4rbs28z4f7jWT6lbXkvJg8hI1cJHSkjN9C61D/i1EPA
U6+5qfFFmhOcmJfTh19eQLvcMrOC/BjO5zgEdtwGXaL2sYUDXoPZtHB/Mn576+XJ5mNAsF3xICbV
HVcM7XTTAGOQF782QQ8LVzUQ8zKqN0zu8qios0vvmQMvJhd24eBqM4MiTR1DYNlBIcdjONvN5z4Q
SSjFH9i1JJrZ+zvUyzRjFUhQEoqmwegIkgP/BAB/H9tBGVfQjlzfuKZb/qxc6Br8H0RHBU+04wKu
QQGH2W4DVZFZhE6pk1Cg6dqY10ZBaUTmFMygq6uNRH6pkjSSi0ZHw5ZM5Uez+kcpPATLJKZiODxW
LT/0Ut20DbJ1o3GDXXrwo9LcyN7Aq2xAaoRSs3ZINFsvv02ibRc/uat10BYwJguPEVim3yMCOXBF
PiQI2PB+aCGA8AkNqRGZB7VrN9m0KXO88pyjVUjdum5aWuQ1VR7tS7/+rzPkP9dr61dWvOAwmmNg
VeV1fV60D0HGU3cOjG1yLJX2xX6CfuNc/KxTiCf+OSQE3fXiJodP/Fq0FCQYNbaHqub18IQjWb3t
W2g/2EdR8Uq2ADJo8/IANJR46A/b7qWpTh2eo72AlCiaq1gHjgnePlYZRP9+NETMq6sm1RsPXbFH
txXoC++BBfZJUc6t+x3Syj5F3pnNgJIbySiSylK93NXgZ3s5y9gUaKMZqkpQPZcruqbLrg47V5Ha
oQzSb6QLGYu/wk48oLPreBEoUnSrp1krekZmbE5No8Evji5eYIRq9EuAwfx0ztfTOVQgw7SW82D4
vHvbBLqvB74yHgv8DK2f+6yrk+yA7wvOoccbx2F7PyRyaYF1/gKZSDFnJGLp/piBA66DzS5Ll54p
BNoi9v4QPaWcBPpGF1DqEgdLTEpAbXYbXrBq+2kTw9d4LwzLL8reXXrUCaTT0/LlnH1nQ04+mHDH
7aC35SKxiueMIOS7biRhrJ/Nf0AT86lx3pQDfPjFLAdMjiz7I3LeIFQDNA7rugbrsnuZ70RUTs6m
9jgSdDOxhr548A5LtVrlbVsOyjqF74cnAvjwkfIqHuK5vUIJP3lMDqemBWo+XGyokiyy7hX8wSCk
TQ9g+lIBD3aDN+ywhopYhMjpQyHzOXHcNs44AZG3ybajvLTICTJn6xS5tcm2+aCyNq5kd1QOYPtk
xjFXFW1NZA+4jjtMSS3cK9XkSLglFTyNJRowTe8ZlBuXkGY2/3nQ7UXEUYH+QV1TWCHtny9V1ZfM
DGJeSKMuT+t7BSTjAi+XjkxtQt8rMSgXBP6tbSTcZWMUxGbBJkYvj0nleNrNcbukktfmNwWrxr8v
PsXASsjuiN/p51ZTJ9pyQMpa6I/4dS6ySxOJmf4gnPbpc3BIB4IcwitJ8c+hoXVroepzXOZk+0Mv
ebJ7EcJpfU/dVw0EgzIahW6FDdazIYNikppJKDc5Z/iOinuRjqECoU9Fd7nUow+RaY73fnNqhXlp
wCsfEk7xgYZmK85somPtmeK82SbDla/TQ/caEjuHyLAK0teoMx1e94JyDyeO1+SOsUA5vLAVOWNK
oItVwdrA08MycUkR1VaNU4iAKzTZcFWO49D1Kg3sfAWSMUAKR9kI6udVNQ8bhzi4Uwj81kKVc2Af
VUWWq7mo+z1zXvf0CZG9HCa/2FPk9NqfSw182zOv1dmMspzmDNnUIt94XQFwrdyWJnv0AoX8mfRN
/SULUG3pd4EN6qWht2B5Z4POBAQ0hbKZQhrLDZYfYOGKbH4/UErhietu3XJkcohDRbv8r+zQ6itu
4fdEEsgcuU1g7X9dFJ2rJpgCP/hLfaaXK35mxzm99vPtUV9aHhZ87WcRKKwsVCguCbKzVOKfE3yk
skBxRXxRJAr+llEM/f/1CMh5cg3tzUSCLvpw9R0QgSWRDGimCeluP1gt7UhY0xsMTTzZJzQyIqcD
0tstF9w/cDf1AYzKHuo4A0DB4Qc1wIUAWswaIho/4Is1NOBP8lxKpXylqssJfmphF9dJ92ZG/aQr
Sjz5kN1OWkItY2AsFDrJmPDKOabCWlKRpF/hozITp7TsEm0G/vzvs9UVzApHDNdG3ZqO8THRqEpx
76+DKQzKTm/LJlLdioqb7fmAXlOyXf6BHYEKC8AlZz1hGBZOZPuqppONCmFKT6wZcwjawf5XCJ89
4dVVwWvPkqok3C6RoejqlYWhFBKg+KqDV6iPi7WC0kFfpYBD/iTB6KF92GojM6V+H1GqWZn7PoNP
u6Hmnoz0W83dAgfrbxA3EmwR1GdEwtC0N352LC0oDzN/ve5hvDohQrjm2Zlz2pghC4jKgnadCCFN
FVxCDZdllcnxPiyRBf2YIBRTS1zebLvN5PiuUokLqmhgDlz4HKBvl+W2T2x76sibODQdom1H1Kh2
D3oRb9EG5heKDdVRDklPjgX5oW+vlc1/UpHZyoFV0tr7MjUEgu63OEsQzH3NtXMQigBW1JQ5UR8e
1EBsundAm87d/0MnBTphCn6vEgI0cdUj/w4IFFMyTH7VvKGNhw9Cm2kGSUyvE1/+KUtZu/6E4/6B
mVDV0ZOg4qJXdgDh/V+QDf6FDmkvHT66CZaf/Jbge+fv1bqRb8aOVs5rwGPd47tKGz5AWFSMm3Le
BL63H9P8R58zt9Qc+dTc5GINw+z9HMrhnn1lHgAiyO70tz6tRMml4CDUBl1ViyY63uXlm6dpA3FF
+tKtBoWXnczyiTe/c8uEe9LS+KUZGa3pEWjfyWWcacM/SeBXtKpym74CRLjtlICROeGfQyqPcDps
GDF/sHU2b+YfOwPs8JKO70TKM/eUecTJpSWSc1Yrg+RNGoKspo6ESRH3Z4lRozlx4aTOpYM7opco
js9Mhu419UgcS9FkxGZv+n89xBEIm97zlP5IU4XwLQNCepcxjncL+aON4Hjad4c9/rPK4xwEHcGZ
K5d65uk/N8ide7GqiFhMJD81HgzjpaXXcYwdHM8b3DGKtfvbb4EIEp+QudVcs3GcW9fjqMfDWive
sjVr6c2acO/n2zFZcDxUx7IjnzHapF5JVr6H/E8fNQynwknUUAxUV+2jH8RtNFhXLVNigkm1qyDC
NVbBMOt3AdzfbstxxgRHYaRao4V1m4i7sG22KxOuEu71zOfBjZdDDiJ4jDjvNVf7w7qV/ObYitrt
iblsXA8XCQZb3FXfHsc4puY6HGVZ9x0YtGK5+NnUOs62F60pnyBZkL02b0EkckyUGE+8BZ0adx+G
SycO346FRLn+jhIXKLv+ubz+pTgrXgQCR4ItLXu1HdaLBeWmMpGafq5x0zl5U15UzzUAfkSTKyTC
5nWhxoN9JZIHjnw2UAfeL4Zv5ShrzyxviCOEUww8BIlgbdnJIREUue3Ijqj+z1Wp8j3Fgu19rZmH
kVxQt3TnQtZXuAfjVtcpFlsBtp8GtX2mOuJmZGDdejAeKT1bZmPvg0YZ5zexeOAV6IND+nv5qerK
O3uJ8acgte1FOgtVvd//fbFZe227C1yuf2kKXnin5GPMGwR8LdlmFJ3hkR7DXjxGXRcRsDSUknp9
uFSKfBn/stbNyn9/kLSJ0zaGSSK0PCIazfTkrRcYEl3psarbbMizgcpOCNp5xC8fv4bH+Ysqewl3
wkU/S+VEniMwAWNdzsEgZ7VwV17c8Ul2j9BYu3oVaWIEPiUMt4SULhbxnaArhRQHpLDmEps+ZT0S
B9BDgr64NPs7Q9yQ6mhu63UvNxSkSH1AWSmarzPP/fDV8zzJeT66TLQiISJuaOBRZGIFjktyPSwP
f+KrGNFRLtpPdcrov7OzrHfO2a760jA1QCCzbed9teOxGHkhiBdkcbGJbHSNlUF+YLRxZ1jDpewc
8JN48dSQC+0GqLqNngZt60s06AewCPDe1xOPC8Nwaadplv3shu/L+WsRNvUHleWdHxl1jJrnpRx2
Lsij53O6a5jYonA0lZuLI2mTt82viZjqRu/Cp2vuiIfXX9b66C9Ht1/c3zm1TgCy5dZq7DopJltf
WnDOfTPPsX5sRAfdk3XHESUZglvt7febc8COQNQI58qTO9QyquOuR90lOOShttdvgn74F11N4Zvg
V19mKsafb+Lc7qi2YVYoUse47B8vxr2LsHTd2xETP1jRv4rDhBcPw3hz0btnW/7xrzoxt/7NJw8l
X2K8K/0PncCTLzToFs/hwG2Xv6KiqOeeWuLcN4/nFCKW8gWKjPfeJfvQh0vXwflpCgE4HBqj0QNI
IVkBxBp2VfzNXT360q4WbMbYrhRtZD7r8tkFG05bWIXhYndkWkFduTffoB2DUDQ+7nqsg62G+1Og
BiI3d+IuDdL3Onqv+ORtywW32irhWDfo6Nw3t4uSXH1Axz57F1hDrXo2jvjNb2N4x0mY/Usp5e06
PoWR3BrM87t60SMzp/PEFjH0nS6ODkP3Wty6immhQeOLRHVaDCFUbjSR+gtpBZzLyF6H8JJvAH2g
Z/8roeEGMMWmaPpcpm9oTnE/TJfrh19J0Fm6WoktZFaBDgNdOqhIfnFZlJQ2QhXuphU2yiPFh4zj
52BDIAtlyliH6LBNbNdZFHggTfO/1ZMKstAUzi665ry9TsZsx4xxnRmAMUd1F+z4wgI8PJCpwrdd
yWkPgAossEuAWbTR3VyDLkemep8vn0CH7GVR7sN10dmJR1wHxPudJr/R1B9JekvmtWBtv7w5ARuL
1elaQT1zdwB0mQMOy8TxsB6kcG57PbULe+pxmNpHbuKdMdlJ7wQT/vVhdbX2w5DM44sczBonloLv
sBjIG0KO4fyEFtPzqDtPStkcuIQ7Cj/l1oEwaDXHKdrid9lIwtSLJF0G/V3uHBTrtGZM88e58Mg2
lHHlPcxdHycXHAq0YutSTYw1G+rtlHzB1vkOCpLldZp4ex2eYkJVop/RgE5WatjCHO4M36Fjq60m
uKwbpKgofkvoa/ALd5aQ3Ut59BHXXKgIdkR8ndXbS5t/EQT8TUZ7mAwXu62L4nvlSD++LfaznaXS
JcjEifjIJUuh/rYndWhXbJBsO2wKpJ+lGzZkgi3VKAv+5iPs10Jb8sfnz8woGJvlR6lDjEZj21TY
rs5ECOYLo3bE8V+fLZvZkK+riUruHJFoKhxD+6zaOWYpd+W7VgHNC1+cP8mLKoGB+EzQxuUqRJGE
PwfmRAhpMOodlf7x/ZMdcn4j+lqsmPERaQJFYfZRlqL5PUd0wc5L0CEyK9ZuPW9BDCVw4fZgBmsj
nMpGfvx6alDDm3byeyzPsYt8zPZcKNpQBFKxPmpKyfsHoM/IT0h5QjhlFatV9tqKjnuDNI1rv6zc
D2wH2CMq2ZSNA6BbcbUssvGbGXHtELeW7WJA7wUnNzRrvMZdtknzKUm+N5mqO2gnoBQXn3B10d2K
eo0b15WtSH3hFG4A3WHzaUnxcYBa3JLTdVC1sj4lN6qae/3rYw+5HbMn0VlIHTH8STjmZQcptD/a
SH18uy/SeKhtDtMMIt51g2js6raUmj0LfDh5bVZ8Nd867i2Nk4AP9Kxd2hft5QDTyeqIGuER9jYv
fuxce/QIRnFtnBYUrrYnR11dVJJIekHrPIDAXsRYIxWyPkwQQkX24qQXRHc6kmbeHMPHrbIjx6im
gP3k1l4qY3gChMsB2lzCfKHWhrz6wWOrN9cUs0zm0PakVKbeINyCz4WPg/B20Xeoe2fJOYqT829x
MSqQ/rrRUVeRXqdMEDGwrsI39831MVJmQ+KL4uTHqWrNMz15xnsT3v3DGC2K095sf7wH1+sUTFTE
Qixr5s99KrjvpKah2aPyHhUCUm3Qzk7j/HOvHvCcKD1B6bgPj3n0DOzR5ZcKhNpJEioDvElHuyy9
P0/L4SlSgpJFfGXtSy9OYCvK4S5hmO7taLYiC7AUM1VV6jF61romHNiusFans88Ba7WJ3Slf0eq3
NSDFpz5M4d9naRzwnfLS4OttR3I0wZloGHbByXGSlWOF54D140oP6DcGFTuxXqZ0PFZ5G2IHUSdH
tD+1Pohsn6u0ldViCmPyUE7i0ESVlzX4Odyk0aJpaddCS3562i/WLW+yIi8nSJLrch4R/NSqKcrj
6NeFx4OJYlSw3Qj9PIcZ5WXWyQqQ3hXfCrpdXC9OCBF2fTJsc3tgt6JmFaUxMYS/hcin2cgwDstu
J0K/0Fi0u8+7SNOeM3vbpFDUBSD6p8+69jMFCh9FcP6qXooh5SfT0BTqqOABGAa0wOdI++MA7Nh1
ix7JotOnHKvYMQJd/Xoj454bdNo+mPX6yqEiZRQJ3CJh4K37f7ORxZ+U1SRLALSJh91BBnMJblfF
1v84oDAkRbRobSstThrxUSz5dJxZytxIYNWRxgluOAT/wtV5atzaCkgrI8kzehN8aHWK6mJgQJIT
v5fXPNW5ChbgJL3rnB9YhXH6gbeiQjSwwgmBJ6usb1uqh87BsJdAwjc4F7YSpyJBuAqm60JSAKso
qwR2Atv2assC4y8pgbfdXd5LxZ/Hvd+oYW8tA9P6/FE9hrDLJKXdcYMzTOOC7/zl7Zp+kixVRvS7
UgiszjIEC3yRH2H/O9q1z0kxA3ZgWNHRvXc8tVyCJZyqrNohGsVpjiuVxy328UYU9KoYftzgmVtQ
ThNfnqV71AW1LdnuRYuW+bIzdx0hiTBmjAmZneZUXF0IKap1CNoGs92i/et9EaWMIcF5tzbwFYSM
qGL521ZGcnBR5bMajN5YIKPX4MbSBqLBRfSHARqJFXJ2gWiUxnOLngXoWBdSWELwCNPn6uTAzGpt
Pm5QYAczh6LHzkOkGaVNBhADmJVPVjxDildmgGEyVFN3c1HYD0gRHkkUsMtuAGn6HOB2Xi82u10A
I0EbjjYr3BS7wKlM7g9y2dDo3FUdAv7dpV1AjHSo9k3EV7Zt7uUuC0OztrDtfpdtG+3eCiIV9L5n
tByxfRvEdJs/Teb+Jt9n4YSImNCAR90eDNmqIViCMZOKgeQpll/Q39ZGtJ9XoNSetNaXCZTucG90
qqOpDRt54DSBN8EzCYJR1h5fQwev0hYp/eb49uj4Y45jR9CNBRQpO9UlPWMleudGWqiiQgU3xQhr
luQDI4tpm8luNFkXPlsaPtrPp8LWsklpUgr0zX7YFDT0SS1rp5sq3e20hP7jk+4KRU16Qer8x0H3
0ml7FWsLLIA2k5+dMuJNpVLS/Gf1fbNvID9s+X0lEXTdocuQwTZisPYj8tCHMp3yZ30Tep+T7g5o
wWCbIvrEyb4L7DqW68+rXGduK7myWKMNqZx/awxSIf/8Kuq8wvPAATZZALOAzWC0znwGiZHjsDBI
M9pHBK4ezqtfdrmkFYuPBUBk3a2aVV5+IuBz/9CYiSGXrdsxhteFl0HgW382k0DiJvZ1f5zzzIos
nDxMlppjfZOo+A4KeIGO/Xa60BnPpKWOPhR0RMbIycPXaYYLosLr+9I8YO6fWmcvee5dD2JOCpVK
RADGHOAK0buZDD5YFdA4ZW2pBdss5K5IszYi+In7ootNsnXK3yVlWS70xQvh5xAIlLI6++Sx+jDB
sGvT5iokKIefvGxFjHLhe7Ms+hwGBoOYwNH+hzqxwQD60nRl4JvO3ELmZawWGCAgtIfn6S4Pxynm
F1yYsMkDOVnsAbz2DFR74VmMjIRPh4cFYHSE2M+PbxVl66WDEM39C0W26yQJHvbc+/n3ZCwkLac6
6nXZpx1wzt1Yv/aTVIE0n6+f+TkW7MujnJ8Iy33iR3V7VlvTHxamYFfYtnssdPp8oJNfqfDWoUA0
JoiMNUV2jtSI2cKIRaXzCpfTNCYr1tXCFEde8+WlR/9AKxzBKrIIOXh9fyjZGZEo5dScoKKZhHlS
7wZSvfRbUr9gbUL9avHfoqHVj1vcZMT8D5yK08h+IAC2drhv9tySK3cctfcce8HelbqeEgmypfKK
9OyAkh/4sMsbUmzXY/r+DPLKNqTofr+CdE8XGh7n13Nf3XLejDSv1jz60ngUyIZZiXI1IGjlbkiz
ucz6ouJYrEqqDWgjV2TzskM4AVZjhWBTvOySXlFP5X1CMSwdzfZS/QhiVqGmoIR5D5pMRmO+2/BA
7pZxuSSrrpDb56W/LgHj3YHrR6L9tyDU5EQ7Fb5X5Gs3n3okEFt9Fxon9r7icKcwYHslEtzoRKSF
v5Q8PD+nrR4c7n336cbTuNLF914NgoyOyiVKnBoC6onJKBLMr2wxNtFeeio7L+fRYPhMQHPP2rXv
awop0gClAT7IppHlZ0xts84OJwUWJdWhxDV+vqmkz9C0lMsY4Qtm1IeAOyFaosege5kNUpR17XD8
/sZWkQDblOhDF3YBsaL5JeUIISJ1PPeD+Sx0IwrJh0KHLWBmthm/mf5ddRwhXF+XxtL5WDFxYQ95
esLYOK4C9FlMzqX1RpcHAr15H9kuDMQg022t/VQo2JGJmwnBpQLU5OBQ8WnrJGeJ6hVIFh4/7CXl
WiMgoGwIoAKNg3VO8fbo/omtoswwefaphWyAZPydsFJaKX1PLDbx+lrKygTpOC+i/upBHxS3X7ps
NTR85uc+8Ub/RA1SJcTG0vVoIseMiL31G6yJAnsodRxKTQsU9x0GyRqpgiF/iDsNw04lBfPOYKl7
tbCRtn9kwQp1H64/NEThRxaRtmtnt5NAUINRdpVBguQT6FnN9MxeABR/LhMmVQib/9Jt0ucObF7s
NYAE2Ilk2W3v5KbRLQZgCQJLEcPP/b7PAqOI4Fbyv24ZixsHdMyjdaQ9z9qUDBqGUSLwa9/EnlX7
ti7CvFHeh5cv++yENw6TbT/cBLaukAyCDTozHHQyZV8wXdce9qZZHTGFvsdLLGQp2OgdBxNWUDVX
FnRXhL6j80xFvrEPzhsAqzajY67qgrnxOzMKZKdn/FwhLx/brEZc+0cFngyX/xT2bGzTzf7vAVE0
rAzkpIUeT9OuQKuN/k3nWKaLJ0J/IF7qGanJBBbsYECk2uFqEt2DtqPP6oLFDYM940tPAz+RXNi7
ScvtEVXShg2mrTCF5SEJ8ngP5YwUJV87rc2qgc91v+CBES3dWNriZIm8JSnF58xYSdG7M+u1nQ7C
Nd81zj6Pn7ydBIwkS14vPnEzxdghDM0xgzPiGHs784FRp2XW7eydAh7RJ7FIUz5yHyTHPlrYbwiO
BwuX+/7NW5WqTkhDdvja2/aj4w1bm/LRxVK3LkR3Qo2SKmerW61OJJVMxiEKMpeq9aGVk+8yi9FQ
jLt/XrsNRceHhICQ+871tHd6lS9jrH3HfpsJH1GWaEY3Akrs/YtlWzFPqfFKDqmvZs3FwckFktWe
vLx7tsXN1vw6bAB8fdTBSD1ASF/oF4PJb1jpRt5NAWf1HAkBg0yfctAZb6hg4wcf1GAxqTlPoeoB
hRJFD9PJcom2JFJfD9yYhRRVRx1MX7aI5mGR1y6Jpol3jPdbXDJcGbvj7IcEFX9DiM6/es1xlj9T
7ME88g49LYf1DArbQOsetDkDZEDKA3hIWipglevQ3R8UnZdWtTl47tajdk8OJ8dNEmjuRRCsPZaG
MeEvqw6ET550YecCphqthXc6GcujMDvEr5PWDMRWVbkWtpqEcS4RwnkaxbtT/EBAtUI34nnbNLF5
gzVpwG09le92b4GS1MZZInguV028uTaeHs1JSMn4SNhDg5Laid94vqQoDtlUD4+T2jThZ5D/vgqF
KX7f833wFfHvV3jTXT9iGGDgGgUxsG29F76dwGb459zPhfVOaZMBN7rSMfpN1ptxSXQt3i0KLBMT
SOnUVsBDBNDx/5OOBJM9YMuuVHaGSAdG/inblKCegXqlSaJJwAniRCM+AmtAxFs1AAgLceWE79bs
6WWNM8xAwF82HQSDhwsjXyIaOFymdFNBlj23lmYs3UeWQs1VEfj6Z1fZuPKfkjzx8vrTZPyuGU4G
Yj7zq6T5ZADVutxWmOtvJ6cQRzVrme455kl1Y7zrD6GdiR6bLsGLiwIDuVQtQ331xpL0jsa5Ekqn
FMIp5s177Ggu71Ko3gbNR5hFwlpM8lV48FUWf0EJIh9w6O6NZYvaqxS/WPibin23rMuclCITpHq6
NXBd/pQlQ/4H+eN1WGLXNAzqHQ6K8Mrm4D1a7H5hBZClvSdWv6IoTWHYctG9sQkpPHjEnV6QFd1u
03+jemWLRvMiJsluCFi+L3H4sXp8vpILIeU/bJizU5QKIqBk8CV9UpM9uf3ynyQqdQ2U32CIT1G/
zpwNHMmYyImFLox7uIAZN3SWh1EAom9YirvWOyZEEvg4juhg7w4ZlLZv90on2ekIaKajTUSBNwfN
6kLYK+0slaS86JacECh/iQEo6drJk/1HrzVjQLxHOuOM7hkpCSqbxA3gnpHLzeQVAB+cSg6Xnw4Q
WmGfSpERgclHUbZJX0sR2ot5Yt6d0cK2cAFR925eOvMFwGnzg/GlULtVhZf9pwO5rDVqU7QVfrsR
xAAkynPXdTyceJqRCGQpi2TmDsErZ/8xZXg5FlbaoB6Vq5SHTlzmzc1HPxXDu3CTnt6di16Z7QTJ
KemYXeVRB+EJesutI8Q++IZqi84fzx3lub2whzmdlOdGKMZL+QREFoA+aX4nCeotwiBlJ3gCJge6
aEMjamruL/LmVT4dwXPevjwxHLJP1P7rrVQfQjMneRBN+XT77XYQM7F4b6rtK8W7qMmkcMlFIj7/
oO00G13dzRWwqKNCUokrKlzDYLUVY2J7Dr9p6PRhjGW1G2WOEbIGcbBl4OTpwUyn95m/LhkVRSX2
Ks8AOlK3Nk/nYLDrze5Xd0Bh1TE0wKJAFClOWnJPwB2vg1sK0o4G2WGCsmqMZb1tjWFuA9L5oA32
m1cx37rXmE5dw4UClysHAo9F5X7mnjdpW/oaq1pVlrLWRhD33uOnTZFDY8xF/cfvsRzAZLer78dT
3MWnpodHi1Oo6CGeQSc6+QLjbjPdb7KLjP++Poa0BNSq5zPX0hHc+h5/gsYQ0CiH6ZPln/UxPTHs
7xUj9ZeIILKeoYWOZqLgvA9wKAC4mShyodUgSwrk1UMQfegIv9Bp/++/yED3tLeyJLdAZq4YxpxY
ReHXI1+Die4CPAgr3/whI6ydAfMNN1c60AHqibGbtW8zJA9jGkz2xvbqyjj2MybTd2KwgVG76UOR
HA+Nge8UnpIqOOyrWCEgcCSPMG8V/pbsHzJf+DqRcgD5U9W0vPU4Rk8aYe11q5Vh56L+/5KcfMV7
cRqHFJpUVc8qINL8hc57cVBaEk83qry7+Mzg/e4kMkRRakJzOzDGlXXSOVrHIOu+VyNy+yM/e2KW
HAwtk4vEQkS7yKbm4c97OcisM4qtrvldc8+Ch45N6XYoc2xxstGJJ5bb1otsGmkDEvqJO7u5Y3pW
s+UkAfmPplTQoEdNI1X9wGK2gLSV45lq8YEGgaeITiNASU7O0hzOmsiqJoC/txVcUZOmgHjcrl/+
tW/IHQjuCn1D3bhy5RFiojx+WBJHbL5lMUa0AwRKVoDa7MpZYZekcvwzeaoCJipplbjWcTQ7oJZG
2Z/vLyc4s53/gfgEdQYFFvCgK5ISH0b8GZTm8amoVK6cALZypkYznO0pOmb/mKwUAEN0QiRf8krb
C77rv2HMv/PfuYrqJxm7sTOxwVAC9b2u/9CqEm1dn80l8eiZV66NNNlBYSQ3GPSGWJQqmDpolpQr
YUo8pgpwXu/UrbzBkKtWZLr542h5xCnnxJbUbGWLOp5ljZuhFYDq/1mhid6S7YL1puhhBTZVS4pj
YfzcRovWQHSPH/rizVIxhZaADbsu7pR8k89Q0GqVnGuLYG6ooIzOQYYXd1ddZw+i04dud8BH1Udb
6lgjkklhz3Li6Wtcsr1zLfMdWCdUobdiZXmC1CG52kfAa8FPS7uSPVA8CtHuRvB2jxOoowg7BmYz
qTCnCjV6iRElM5puGfAJg7h0bRXLAxJH4tdGj8kj2zGQSirwd6Z2/FH2nb2ZW2EQWemQj32KRzWE
2HXjiq+ie7MXldGW7ESnvjQ2Nb545T46EJ2Bwsm1HUa00GXhEr2YOOGHhbI0WI6g1a650BNpK0yd
QYdp/d0KFTEVK8nLIDtIJTI/3kp0+vEPFXGwl5UMo3WSPX31ZuIAeyu8zpcA9BR0iyvkdaM637Mc
xNwXknDiQ58SJXU+SfhNOz9wAnarPO6p12mpDM9VSaJd616aMJ0FgQKRj9+rE0l0jWfw7ORSP159
ReS1SdNuUuzFJeFD/4Xy6gd2+l8qMa4J2SBfNzX+hBeMFUrtazQCHTxB/UdhT23f5velqJd8P+PC
xiifgSj7/+kcoCtN5wsslUFyd9FF9bYvwe0DNYY19X2v832LKg+UgSkuyZkpTnZg6AnA8pWSRkKx
PpALyq5MOCeQRQimRQoIxOndUzuzgoh0DyqDQKlZ5oAfisasukksQVGXiOJNxhLo8+k3g59BlXez
Dj4pBXaaITf8TbbXOjaWvIimP214AAuiZFYMfmV4g5uTR20qIX9thi5v7ipjr0c2MOaKUeAx7DuQ
UGt4zbtV92xTTCBc32VaSOUYHukhoYUWJhklMcgi30cBvPiv3I24I1WoGAjQrL220j6m+6ixHbgf
5IlbmQx9XfHqqb9ASa2TmLCt0v/+NJBRlJHVxpP8XPGTHg/0zOGISK1YmvnTl/Xml97y5X0pjhna
tsQrrzeqeoUk14hW5n0GeJn9SIdZNuMjZ3Ikymo61+20s/ZuSHn1NbmePXOlHiC0vc73O0TeU/JJ
JD8OjaNGR2/+RK9X1cVKd6VaeRaI/whumPSg1GdJQOW46iiT4XVh25+cp4G73VFlpkZVtBhgzTiM
QIk6cZtfQLigVVOWh17MXF0Stcd5uGCoiLJ0J6ay699xePk61/jNzgA92mHAdp7nqDz2Z3k2eSZl
6/WyDLwwiNAMrBLOBdG7gQuF+Y4pOXEd4P1blYWRsVRMfCkk0I6zRHXzohK40W4b58JcaTA0BWpS
/ObzweEwS+uLtEOnf0DoDcgwdJ/MnAt3VZwjEGAzwGX6jhgZk9Yo6ejhIngqemriBjirYI649j5P
l/3he/SkSwrkMD+d8i2c9mMXZ75UDhtZUEPNuh7qxW2bzNOLtfHzf7PzwkNhHfL+MHH1LY2dkdPH
YcKkWZY6DK8ifibwFY1fZ53aTb0GPYSqCzjNFtjko7hH3SnRQ3S/6YyX0W2L0K04KQcGrrpReWuK
FTUFdB/zd3gaJO4UIm38u/LmqzmegLTiB+coKM81J/ZooxQn8hFpDXYztaoym8ICOVfxGOk7senF
NQxdQC6ZZ17o4F1Dgyk2mqBqHawMi+igz4Ppu9Nsi6/ve0XTkU9mHNWWyTBFqp6/qibIy70BJVOt
d7+U6V3XEQYUPv7f2Xh7chduRgB+L4i8G8MQ7lojctpHr3q2EeMtcBsiXm7in7NkOhyEYJoe30M2
QHs5/SNvVO0fvwy2UcGNIG31K48gGeTt9RZfdMCpMVXHw3iv0IOUNdlf/vgQLaL/tZa867r+kv/h
Jni9PvdLcgBjyfaOfPUAva94M6BxYVMJf+1l8MAKbEtLTi+n6yLjaJOSIMsXdTlcy9G5XQ8eJDMp
tLB/zF0V5Lct0A2Q3736q8E2iZXmgdCeYrInb8Ap5LZAwBdmIp0VvwN7COxFgsGI0NkBpE18R6Gq
WhTlpfLndL5Z5K4CtSG6q+5fqjEPJ+QprdbwECH/C0ETtfi8XDerHYGQELGkG+DVXzqc8G6e0TN6
6Pa9kukJvUJQ+TjnwwGlI/u29TNq5V5D8Fb4NT8l5k5jz5DmDIryYOy8q7WQpnYqf3Wzv0qk1zWE
MY2mCIzfiLEQGl1KeOMOtMgCupAH0/XV1XOVUXfDte5Lr9fBlm39I0GA6AILsfWwH8QSL3/gyQIb
bLbmz+G8e3RAnFTnpdr4nbtI8St0nw6MTyffBac8S+5rZkV0zCiJJx/eWH2Tz9He6XCd9GV0Qu0I
WsWM1zR4q5HmStUscklPPug3v5nZGU1TQQljzR8qqRpLanSGGOIEky0C77v6bDkMaWv7JGsymGxy
L6R3hjkULGw2xiMhmkNe1XNHcHxy9BxVHN7mVq0R7YNRQqTquPIAvuvhYIg7ad8VSN9mYOsUEVtK
fW0/rJmTcIT84WYl0MiNM+odCSqLN0DB9qje9ibOZFbr0oq91xVwM3FLTU33YWgXtrvcqF5w0yuM
XFaCl8ifXvv1VSLUDl17zI511h9ekCKmcs+/Z4qHCBxyYCtnge1RFqXcLb7r/YVd0WuaYGjsBKUC
DHP6pR7NF45vejMC3+8X0p6YWe1LkrnplEajNNNMFSS9V9OcyWNN5Fv4emupWyzy3Fje4ysqT2K/
c8IcvnSObQyL5ChV5xTQjx8HFniUpN7RoibDCYs5rKM5lKEtpMs0ULVWUkQn/UKwFgHytFjLagzG
9KGYiaA2kU+mO+4y+OGpeI+0DgHfm+5Ha2IF8OY5/X07w+zQRBTf3LUb6IGEdT9c3mRI0QKEsnUU
i57btnLGaF2im3GhSvo3tGqfurTOJAzEIVrJIKf0tjIN5mKCTQjO4rOO6v43tsy6wmeZwGlngiKL
xHIdj5ii5z/StOWgMtmaMyoWJUNOn1HWFxuQXXYQAogpENlevN+K5A3WV1pNTUW5gZxxE8c1wU0+
aSH7Ot0kjxJ6so5Eh/mR19ImGiEw4PR1EhscQ2OMhgOJeIsAdYB6df83LyHI8+SD/bUXIcWc+j0j
pimprrTB+aZsCfgUPjzQRfFYBDeYKj+Wu16mbn2fxXDYq13T8tzW+DAfH6ma0NqL+I1kh0WHwz4f
Y2es07nf8D1uzuxQ5gh3mZJfK2FJKpu4ADC2+Fyua03+t5BDOoYYnEuEDaVM08n2LI2SEfeZ8u6R
Zh71JxeZkZys9haCUz8WxYid6czlSLlQiNCWH2WzNyONlke8QE+tiZ7rnGq2JnOER2A0xXgfE8Mz
tuywzHBFVl1LfUftQ1ujWJWR8bDMh5a5Z2hykf0QOdhrdL0KQe6adBS8qymqSLAc/fy2VmxVUJ2t
nWXM1vKV267r/wggfHVGaa5OdU4Ku5efJEKpUgKg/3RcPuYZmUiFhCwQNwB0AXFOcV1HiQe+mxlM
W2pi0na5DWoZxjPHkHj39C5+IUKSEhyHaQNsAkGZWLQ2RqRtSn2LYLSuyZkPE/Dx04dcpWXLmx0I
ivj8il+FaPEIeuFnesWFLozbEyRvRAoZ2qXIVmBdiLKKRLY5+0QmxZJ5+2a8k4xyyjFvBC/6rcos
UROeT6qR52JMroa4d8vzT7rsF72wut7gbgehlvQYZ6ywMRpyX4iIfIPY5pl2AFI/KpDGGyGHpMf5
eO1iA6oNXiasMite5J71RsQa6O/PXFrnCTypOZaD3bi8rR/lv1RQ0uUSmDzA4SNMDwrnQupYplC9
tjoUZSQyMOET61sDvRpC6EZbycftnmqGqhEINYmk/LFPUzfSPCJwlFiO5q0w4gKvj8kMU9u2Bvsx
8v70T9CulVMp4j2xqxLnVleqbxJ1RPgigcsljmQqdbPCHScQRrh9dQkI/s9SwiTNv0x6URmDY9aF
1zgzmsgkTAtkE8jRY0M7vMCkFPG0LxLnylJE84LrOCWYOCRCs0Mi9I4KVcGM6gaLDS/4RuxNta32
zmU6mswNMVRmPuoSXAgq9On/Hd2CzwxS+X5efrQ8u0Yb9yEY/us+TBhK4bY+564m9icPyJpsGqx+
C7e6wiDKahM3otQV7if3aQSPsgDfjlDjfYQsKfe5orD3QG2+sp8qv3rqautHYy+4egdVzfRA9yGg
E1VKGHFR6Cb2F0qTEFRz143NYV5iKvg/cvaszcJ7n6mH7iYsSUnoTLZDwcs7OM7x/SBpGYVM/K9E
s/Sj4UUN4qlAHCPoxeCswQrqKIzhOx23WACEuYMjC61av9feyEIrimuSmzi1bTqjGbr5nhExMbjK
6DMi3MBnrSBVDlqxi+2cnTnDiry4xEEgKCYqHwaCs83+gjqpe5IKIzI+1RAV+1zFC8MS8z45cn+m
ZPvp3zISbUh3jLjWwSc7WT+j0fHm7AMNW76KyStUMFRRoiOPgnRdDkW4ekBliBwJylsufdmmbA/C
UdS4zj+PhCsv2/Ues7C1atzkigTFNqzY0ZgTuWa6DWyBV02DuLxCmctyjT3wRfOoCyxqkOo/hcwI
gdewJvC20sDld3UeQbiadN+VXv5fpeylaIoM38Rf4L5TZSkF/hO/O86DxzIaCJKyzXvzlsoX2ylN
YlNREEexTEAAF7OcGuprwIvIcO5q/T+jFHwkQ/dL7OvdZ/FRMJ+u+d+q8Xw52fp+vMmE0DDvUwzF
8Z4kgV+WdiIwGE2H5/QzCnIh98zwIwR59hezlej7gIIMLAL9Q5qfSXaXiKq3GwNaz2F8d0Uvpg3r
BxC6T2ec1eJvLMpygGP6eoegIL4Q14vPE5x3I+xZJC7r5dOc159ATxY7qL0M7kc2LlBf6NIcMewn
L5le/4kvL40XsjqqPNo5xMAXeGIF6wYXZ5UbiweYI5s/za5XfJvXmy8HnyjnSk6iIA9c2uDbyVF2
CeyUDoL2/eCtrqYNySXK9AT2smCrTmWebMJmRq/hwZNmZRXsAatkFJh4S0JwM72P0TytVqNT/gIk
Sr3k7y98LsuccHp9cYSs06sGgsusF0RvC2++5CU1pgIVDquPorJ7A6XibxfCfnQrPBdWUlOSh3jR
9vnzwdeoBLCFZIA4uEFNiBpUcjDyq6aaPVxNK+F49wsNUDkM5JKELAW5/Z6X8llyZmW5pYnv3Kff
duIpw8511qRkCnQRD7yiqLW+v1KKEOfupsxKecTDm4sZc0oXKLmc2TagGN17cdL6p5pkIkyXPXQa
Krvnk6gqeImS5BChadQi4ozCPnIX+C45UYByGaEOgmGpGlF9gxQFBK0UNAymQTn7N8Ppy+2pZrs2
rYhOb0e1X3Twp1Z2qgcNb1e5cmRAdanpBOnMuxvgp7quU9hv4LzBrlOWRMTQ8R5c+sEc4qNacWbc
T9yNlwa/Wzwze6LhFKGhZ6lec4fnodQMxVhI7SjC8TDXW2g6LKwpAWh/qo2LIb14j3NcwQggTTt7
8xAlYlvmcaDRLAyL99aGRz8q/nCYL2d15+4M7y1H001VmBA82GxzycNhC2owy7id7TMTy53S5YVy
P97miaB/v7n+BE+sQGbD1dTCff0Q8VLaqd76Xu4xcsC8U6hfHcpCfVE+1okhz0PLx5j+ruLNQ3MY
dLXL0x9KX57zg8rb4QIdQL+f2N9ziq5Nr+u4AeFtCTLNQrFfRbkXofNKATpqUg9/SaoqNvYobY9r
RnbrA1XJh3JRKMJEZmWG3NBluIGuMngUPBE2xIxuSvwq3Avo6V627LFgs7pqf3tZ3yWY2IuXijo9
Azq1joky5scBsZurNJaA4JNZIy0SnzPjcEMSOsKcZkiqxBJlg0f3VVr3+WDJ8S85WpwTjjBBNf16
ea5Wct6daMceLyXGKyl8pd9IJTIcPT573HKGigoVsBIs5MpS6z8JpCujYKQgTTzvKngSvk2FM0Zj
A7fp5Hf8b9oHZPsu3Jk5mlIngANrhYauqUwXCDL2lijIUBPV4G22vpsMjaGa4vIClL/zFa0HRq9Y
GGUG91ccYAJ0LehyfkOoWL619OK74o3eeFo5VkiYwOJuvORrHlSTmS24uGjT0EmSKJZTitelzNDp
l+3mKfO7TuIhxZMeZVmulyPCp9DPoeEAGjdS3dFYUsp1geTMbB3+NhOige8Xs4tp4JMuHVhmpFLk
/Y+yF5zDe5Gd3SHXc2IDy8tcgoLDgNscCG+0JvHjvNX6ZdyHUIuDaf85/fwbSnTijKYKZTvpGcTo
sLtYLGCb7lxNzrYEieqJFiiUNC6sGdiLJetGwURxN+z866PRjc0c9V5ly4DTKI8o4CLSFxilhwv4
cS9zDJA/PwMSyPZPbIm3ezCdzfBe0TtoHKzgYd/MemM1UPERzLRRKZKPVqiF+8NegjzTOFltjus/
HceFIQUgJSJEPPHPS2ejcXUbdNoCHd7Xi3HuWVFwvOWah+B1HpD3sCDQ555HLuNE4ZcsD4Gm6PIP
b4ih/Xv2DeR1b8Jrnty8bsVovWNiB9xh98/FQlkXjx3mOigRHsS5BNiKjOFslQNeaymqAVd8rtOz
RP8TyI3djHSX0X4Y8Hzn8V/l32oRbhjm8l/Mm3S/B8DPdtID7T6A8sLnoWVaHTM/E5MxiRd1xegL
jX/e6Ld8yLoxS4xpzC80cosZ1E1N5c+igaJw3qtHqDsLJ9wtboZpQ/r3qjYNCD/pB556QGQFUS2l
7pH/llzxlLYPpq/iN1S34uaQrlbr446MuF2HkTSjIejIPZnlYsolzJUhybg11A94SngM2TKd4b/t
uBnxgc4GL81Amu4X75PPDYuFGfYnuVC66q62+2w9oZQW7kuKmhQgN5tVGkp+YyifzfyxRg7195gm
5cGm+RQa+uXGfpL9D0ab6JpREwC73tV0eAAO6+8m/QjhCr3XwItjNFARmY71Q4ImhVkE90fAKVC3
Eg0bnSffJ4pItHYlb/7AcJvnt3PayxgAwDJwdFSm16VUbExDWhg1YbAhG990jGd79nyUL/MQl9Bq
T8ol95q1jEGYBq036i7+Fyh5kJuyNPuQIV/rzrVI6XXMSJJu70gdm1gm8CXSC/D4BLiaR3MXXCKE
wghck+IAq941ntjHiVkUNl1Gnk2cXM2PGUx1gkOi7AA6YuBEw/gPH2DGHtavfIaepD+8ZzT30jgY
ME5dI7muOD6HbaEQFZScordWjc+Wng3LSVV74lmvpby5iR70kix7TibHsknfYDA2SGLlCzbC5JtM
NW4YK3/oYCYEMpXC8lSVlmvTbVwAvAJKwMMbdnXNJC9ooZSDjj8ao6hXd2RUPU7n2oBGAvsgrC4u
mMdClcNbkG/h2JhgfCWpUZlURFLam1g1HgrgVMsOv6O45+EcssqOpM6D4chR6v6C0zCYQQ7cw1Jv
HIZyiHcQLErJ5JrKu6VjBEBT5dsuMLlkEPwAsOL3w3LKHDU1zjI/MiwogySHjFj0KRtfwRlAKkVc
w5/64QXhwcTLhJjAPhZv3po7nkPm9iizlEhe24BM6GQpp6bINSsXUG2SFQcUZpAUF1/45BGD3DeE
gX+u0jA68bzcecnpQvREKzdk7nIrMH2LnqBLFjs79aKY7Gq/gHMQ8o/Fp1T/9e1CQTm9ifpoYPMs
WGs0gYKbgdagQvU+NIebgocKAEIslkgL6DF4fQbhHRRKDM//3HOU6V3pANLwd2n8ih5mLzGte87+
8AyVjNrvP+H0iq9Kprz3U9XuZECh7C5PU8qZovS6fyWoTEO+lTVN5y9XY53r7WLjK3r6O84Wm83B
zlDiDvpRRShnrTLV7qmlgFqBCBHIPRKi/Od0O2/xcN2DOyFfWvRIG5mkNtk/tPzzc3VRChyXkXwV
CK+vtSsZ++vqeDhwmJ+deCAPb6AME4ysBeyfQiY0mQ0J7PvBnzz327SoNMzx4wmj4JZwCiOSjctH
tEJgefS4AGixouGPRN2Gtri0mpgZ/7vQv40qky5lWoXpoCpjf50+SUHjJT7WFPDTdj1MIrxx/cpS
ygi57/XKbHimZK96+zmfwdaQs70ryofVLuUFqkcMVFW+K3tttJguZooJTz4NjR562ozvzWo6ias+
U6kHSOirbLrfGpoom/v1LcqYHwq7IvKNQimAnNA8e7VzZZh+RjI7H8SwlUUWAm3vtks6tBkC6j/l
jHiDrZWCeFH5TotZXAmsA5mUykNQwu4+0oIOSK4ruPA8N/tA+gwG9dhYj7DG2NSUgoj8RydRubfS
KbyqsiEth3D8CrEQ71Et8D6/SBsoBoChHOFsuQ9BmGg1pPa7SKQ9ig3JWtwXq0l1Vn0FCU9ZRD1Z
ZMtX35ex0i4Dqjv1+1GOOgTTFiCoPuv8CaPgtvT6kJ0MoH4phzJv2zX+VvV/mNiC3Xb/qWZ/n6Q1
zF4tdAv+cLKoCTJKkwVmkjBidZYK32pydeu8eMBJg8/wbRYoXAgMNhfcdZdO8+ntWr2lb+Y+dDOz
83cL5GLm/10oKQZn0Z/OCUiCn23uhDiBEAk3KvuE9k9dU4+Lww6JIRvEUtZKWccHalkf3YMHY4/g
QfNzqHszgHdMzKA+k0j7Qr0koXTJDjq0otjEiZ9Jkn4jVsRv2xBpbKZQRMsDbv7dFNlwHZAsMhQd
fLZ32Gq0UYqKqlruo/1DjU0LusIYbhNcuo13IvA+jpq+D8TyqeOxdHPU07+GbXMnpvy2Vn8W//0m
IZW4pH5UQLEJdSgHNurIRaYnEDYTJxYvzkwCOjdBW4tHweOauBtDrrnBsE8cwvghU7VGyqcyS05i
F41FyZNbzBm9rYXOr26SVMfJu34R44iY0ns0+DNnyiPvsW4E4okCNgRZXV00jNMz7i/wuORBz1Ub
KzdkQZ9WtgHusscOobcCP3BKvClgaZ0iL0sHhYqxHciVeoFihzXtb32mvGqjB2zisgA8U9k6qdpu
SoLIpiMTR6Yr7NLpN7l5TGV+QblXgQpm9AbdzTTb3zQOHUqDFQzl+nt2wR5ruypbg+vu1LFhy6h0
yeYnb/MlGM+6243UFIsW54XAwywW/Xc0+hetpVII4yICTT5HAqUasCyclU8yXHWHy4m00SiIhj2V
x/qbdd0HHQS35B1XGEq5INzEligzM5NFzimztPjYfyANWIBoXfUBZp1h49e+vXBW7MdeYEg3EG6P
qmAqcvEOiHZmpFmSr5lh6imdleFYZ0U4ywPoMyW3+x280YW8siNninmPNcdtChdWdp6g2cgQvYup
EWHmZBnX1JrpZk9LoPkDX5QJgmZ/nJj17MMXCOtf3eTM6Z9RpxLYJhUNkscpivXqcbkcUpfooLEV
C1J2EsJv6MqACsbFaoNMoHEh0SjjAOyGmF8HoGdJj3s2Znp72aMJXMKQH703y4asbktxrjkfKv3d
Xm0BjdmK8zf8QdA02EWMLeCFXoiHuzKvcv0GkdrgxQEOgUgElK0OYsqRIyaebuj8950UEbhi2Ece
+C+tXxJw+XsbNI9g8tWl4pVIfS9r+NOF0YLZECv/Cjvd0ylAcvt38/YLxfxuJDe3AO7bEqoYjWvB
TKm6WbtNCBggn+9oeAMWNnhYV+lbdE1HKWrlUTjeJpgqpjn8QAasN7x2l/mQTDNLl6Pw4rlcj3zZ
QZqEUh4+w2QFNDiSo0dSD5wrJpnk3ZPbWis/gWUUdjBo8YCqkwf+u8n7Rv58w/hh4FFOjJ3B/4Lk
PVQFelNVhdzgJB/A1eVpZfNtIxZrs52XjrgE48+OT+zqdHx5CRDZMa1caV/r+4FZ67kcj7jt1N7S
4LKG70WGgwEKlM95gEDUTfr0RRhBIgHSIMPdxRtDy5HY2Q3LaGquhT1FJsA6s41zjLTaqEvcKb7m
G+PQEsv4SVKv6VCTQTi4M/ePDjh9a4Kcplh9VzO0PxErjWM8FLPPPY+k7wrlv9VundsVR6DEnBLk
f55wiByJWsjRoHXgAVDT2Zg0RtkxSPtaXxCOZdAWMZ8GWORwB0vjbALgFYuidvwrkkDG+i4262G9
PdfG7k7ycp9BXdee7wWRjvtf9YEslsfj9C6f/QRyVf8/ozZt4l5mlfZFJ2ihXNHUB4+qoENFF6u4
AVp5TLvPFegbwG/drbfF4gWHTg4QTRChe/ae9Egw3lMiq4pKm2NIH5wWuz6TcEbEzC77MeuBUdhs
ssw75tF17ekD3Ifmcb9j5eYFcx6CA2KXdu6yr7pU2TSFQ1oSGmX3B1R+cpsluR5CIgLPApf0nr31
HQApQ1efSHVguWu6fCRDvlsEquN4oMXDB3ZXHTs240y3UetGaj4GojUX6KlORqeZQ5wsqX+m5K2H
DOyo1ojCaGW+QpxoNFIcaNjBrU1ZJHtOXV0FxKtCvZA52Gp76KrrmnqdDGLCdG/wH6Yx1sGS8FjZ
v2qVIe6yxVnrl7XZY637C4mEg1tccPPGJJ1CrhdDDkUPYDxk8V6ULVyh6igamT/xaHfaI4/bYKz1
G8zN9WDMb/PIUe54eiu4eur4eri+zKyqO5nQ5nkp2FgAc3X/od2ebH4C2USDxBeJ/dNah72ogfV0
2k4wAyAMIp8NFkmk69ttG+EWU9awb3sC9iV+idA6lMP0cttrt5K1GpaaBr2GwJs3S93S3twQYnl9
BRq5g3nffkTGGwvkW+ludBQt8S81Ioc5/1Tm17XGDbZ6tsNkG/ZogphsrjArEYNxJgiRPcG2/GHu
+suMRw635fz+WjeBaE91tgUpMCjrOQlhbLoFFn3pvq29tE3OPBqw8BBewfZIyNO5cvFDBtffa/Nf
JtgozzHrmoBN6YkhxI5WIvhPyCnudCrIPSujZD8p1zrr/nLhfsw3MY+QBSNYIadtSAR5VPMixKQW
hX9JxZ53b/o8oSyBJbNdRzd+Av27MHKd6drNHFFtubcu93FivscF60x9FyBQhXt9BZ1eiE3Q28fY
Kr2jL334OQjTWwSiG+N41PVDJOCSznUlw0sbn6aC76AUD085Hb57YHUdlrjK08C3tHmSTRX9o2LF
PN2aBy8jk0ruDePieqJ9Cr3S/AMVjYubb3SiewvYzEtgXgwkVLMxfpomeJeQecPRgRD4Lv5t38Pp
cPK5UM/S/y3U2ulz7GbGOOBGG+P0SdQv6tOsyNtX9CojZvnknWMlVVw0x1hajp/WXVBw/UBDsGq8
w+v17JGoxlZTULybX+QriqQ/kE2UcPRm/Yo0mUFOftuww1OQCvdkqYoYVFrzrh4eM6GzOy1xb5V/
+JZc52X+nuU7W0JLMZDqmc1yQyoac/ahOWrumrKa6zfRjSSz23od0KJ1nyH3UuHeu/jNjXCKYCiF
rZGnz0RK5CbCCA/XKp6Pl8Q/H+AiJ6zDq+QFpH2JY5m1+GWJw5x/0ESerg9faU4rBWh4pf7wJBqd
Uozt2fKLlTKCHruDAvdUuVCejETnuyIXZ2a2pGw00gJVBbT9U10FoP4RI9x6VsIubzzfYpQuaBXo
Ya/ZV+rUWTQh/kvfYrWEEi9gNzLZBI8k2TvR+2xs+wpHtvaduI2VaJMUOs6jppNc/qrDMsj11SBc
20kzD49a8jMUybUB94Istp8Z6U0gyMV9LyXFOOH5n3aU7KyCZZYAfF1conwGbbmh/RmySX/3fHgN
c7pdDccikmhXkSENxdALLsMuWUGrI/NUqNEjchnoyUF/hGYhYyyFrkfq+ahu7OkTGKG6Kh+5EzGs
AGsEEU1kgp7Agig73klrpmeXhXrOy3lSn9udRWVTm9DAVXYZcDirPjv1qSyJ6gR9cblXzJ2DSrfh
9SoPyJOfzAYlfx/W9RsZ7bK3kxFxc1vIhD6TY8VALHdfElrbDecWQJXTMqY0rQ/cYa7M2+f7q4Xe
ozOb9PT+J+MwOpGgTu+YXrn1jGKM5M2IWIRNcxtu177yE3UZY3q3t0f4GAagTKLBDiS5GSKH+L0t
hMtks5XSLA2PUl1JqeXjcv3sAb6KQJRGEC6fWboxp68SzSisOx4OydYN2woSLAuSb4t+5F5L5Gxr
AcXUXJXbUZlJjRfIhP1n4NR2wEmThy6wNi4exMvV0AUvEoxZwlSAvdPhL7+jPU9BIxdjyP3wRAlZ
pEj/MQSHucaEfPsga7Pf4kOBXGYs197uoHvK51Nw2GqcRudFPn8vKqt9TUugzEiwJHUlIrMB/LqU
Q7Ci+/qh8FbtKjZQwOM8Vg075YMgWL61NXiPnSHNmmwD9iVeBiJd2fpt5xUXuYSpiH7LLIWv9hTS
KK6ETbjEJmPP9G6B0GPXv257rnBH5rOrJY7MXyX79A1uyrkX4vtusgs595Zn8C1CEvw2pEkWjktJ
z50SZ3DYU+x57DrVW46jhUlsU6+15lIn3sAdxf6EcnPkGw1aHlvF0a8/yvbVh01AkCsWlzioMoHh
jh9nm9P7Mum3I35B/ZQbvRfq9B/4lQCKtg1UxRYJmo+q+BWghgMQfy2dn/B3AfvyY7C9RWF1F2Vd
VidrFknJh1YN12kqBYlV1mINtupnVZQyt6pQqCtnKFHDx5cTYiUzb7qURnHO9OwNAgs/xu9pat4F
oo9i5E7MTQ06zJOo5/Yyfrvtz7nX2W0nv0vkjZpJn1lGnfCY5CRNrhFu6k/MGNbQh0v+7rhxd66O
67MamPQ3qdjxcYnSZ2lqat694TBz92Y5nzPI+9faM61eI9XpkLN7BzvdxHSPlCTNONelX5Saxyxo
xJbRrnbdd6ZZajBgk8YHVAM1kivTlT51liUtr4FY2x/4PlwXeeA2y9W6hkZp2L+CM69Rd5J9UorZ
ukXPooODnnPD7szDArBotPYiDOEkHjcYEJGQYjcluoP3J67BTKV0ZS+amOHyo090DiALc3zuflMU
qsCy2DQ5KlWmV/u3KB0VLWJ5cq1hGzL6xQRucMOSyhkJNGlQZuDQk2SEDYWdXhqSdc2/TLXNEyVZ
Y7ec6DDNYr54qJyRpN3r77zadnoSL+oCNSQ+u7EPo1o8IX5HqTYrZaEM5WJRvcn6xZR9YAjmYqxD
joKNlQMVL20tMo4OBQ4I3SvYx3DJetogWETNm4bT2O+kGaskWxDaxDHf34+kU8PKaqWF/kpQsaQ/
6il27QpFKbFgWmFvajzWSnviJPB7zQCTwlg5D65oQ0M4J3Evr4whQrVQN53i3+ZoL84A8yYJujIE
WySt1AZ8JNfVQChEMu2eRCsdF3PJLx7xVdcfa3XWxLh/9B8i2Uwh8bN5Lmts8qCwQmqdJGfY77mF
kGSH1H/7v59uHvZ/seJaaXGJS/Ypc3m9uJ73WR3wHWHYlmfJlzml7gQ3ofDhY3HIsZUIke7uULkj
2ZxR058BqOOzDKFxrnYq38eNeTEfaPoW4+LvsBxQRNMqmLk9aoYKqZ7efFxNO0uW+gvg4pU4ltus
foVTqSAG9OteKjKRsx0oxkRPPkBrv4XjVlKUAiWgFqteYVW4V+hCroXevDHReIcXFVxV5I+HTzJO
A3AiBMnpWMM7vmDvUMcUBnBizM2rQZ8qlVC2LMJpB2jbHaHat9kZqO/liAmhHYHgoIhZOoG0foIo
uYjSv/AMbdo0tYWGjNPaqyZVwEJPNe+q86iCROVhU2aucAKn2mcIBeLPT6vPoTmC/RBoHnwaZyKu
p8dxj64NArymShdnfnQ+09QIYX/f+lLbUpuOKbpyl6FRK1jcW88OJdoOL3qP026x8LO5OLbnLZv6
ffSG39G2h6qwlze1AcNZvfeH95XY82c3ewGJb8q3YNpvVCcfGWJ5qXadQKlYCFDoma0rxPEi1v+h
ayA/hLD5wq4UYbaQEXEQsqRz0nFfUI2aIZtq1Dom+T3Q84dhbnvIQ38bosACR8TlX9lapBRDNlAg
eD0UDguVGSrdTE+VxEBRJthQHcbuyBAMFF9VQnmT7O+1Ex0/C7dsq1zENNRuyjCFDwc6BxB5UENZ
6oFRr/GCZVBUM7FkPs51SmT5BjBv5zXIvNLqKk4v4QvlrQDQeQnpHcULaZpbEf7X6H1vxLSQa0Qu
LpZINtuxnbzL83QCerJgRbbjTk0hyOOztFOIgRCqfxZXN9EXrzBhZaJj912rV/JfzGgBM8GefkX6
1VelsOobvOxUnlI5Oh1g/7zj2DW1q6Sq3of23i4NksSrsHcMZw1BTUyV0EVnjr8s6PrfcJzEwpDv
/Jw2i3zkTJscyCuCXesKGgsSB9h0j7yDYT8D8deNBu2AU47PtC0HaB6D4VF1O9Tp7LsXXXMSCprc
j+/Z+Sw5N2L7zYoMk+07d5ltDMYmMUG2gu5VEM94Eh478Fi3dLxT405pTG4PB4AaifdAB4Qivvdg
nXL5RBMJ3FFhJDIySiyetG2v6YtofY/EbydN/HLYEkBY8yizaOj9PY5rdbWAdwpCog6F1kbvgJTo
FwFiQptWbtQNq5653cijRigDrQy2/NZjU4Z2Xeiob9EbPyUUNq9AhvTX0h5BvWc/5JGsqersgmoT
PHME8xPYltRv6JOdFP4ULFpUVC/xu6KWujmPFbqhvp+vz4arX/wzDAifTvInwXXuReUb25lFeRnE
JHkUk44SZSn6m2cE8NmzPeBpzYRXkXJjaHCgRekj0uaVdHoFmZVXL3g26Cqz0KrGND7LPb38Oo6S
XVFMBOlYot5B4kg/JmivlQgbP/axmbl8LlwaQAyMiXqELv98h7HwMGDsekMLSWgsj4HkZotxp001
eTP32IKoZQDvDcDYtfuiy0akCO5u1oOPl+xpsLvlE83voqfn/rjkzj7Sx9VLd9rikMi5oEESank9
dMivkisY1vfNgyr/gvcMhMjjuQ6rXC/8Txm7f4tN4cUzTikg8xHDY1or/T7fG9nsvSQI+dR8jpDP
Qtqfyn/Ug/q2gMGvm5Z7rNDAjTDObV+PNe0DHDphJ5exTYmQJt3At2JCvWapOXHUHIW2KHbJmSgF
ir8oppkfoPYtT1B/yGd95NrjnlVouvGlnB2O+5mUKVly6xBgvv6StC6MdyGiPTLmXyhpt8CqTsUB
LL66sVdn9zk7G3tGZQxmtY6da7codVEGjcaYLiFiOWLBsCUlCa1uDcp75lI9DZSTnYBUpD//ojZ0
eY7DmGRNUpnQkYxaK8gvBIS+E58KRqw2LNpZFhFyE3u8fg3ytMp3yHrd1Nq/3BbVlNJifBmcRrRp
7Ss/H6Vij7diIklVXw3WZ38TtcG+/lnpfnfv6CibanV/Z9kx3hvOe45kyNYP+/vyr12+n6H+kxOB
yxxPop8Rcl17RbgGRfGymFenf2cPbQsurzi+XQ8ojeJSvswbJiHRVlNYq7IEL0NF67Qt39pKlBl/
ITbYijXyKp7RoURoIuQ7gGlNnTem6cY9v8y1wfRvW3MqX+oU6QNoEgHPQ6Wf8n2zeJAwNRSDepv3
FWar2hkv4vdjahUj8YIaVjp2V5ZVY32rwZMzfP9fqlcWCyEE4Ze93/aqt3Glx6697p7/Lko3fCA4
WgjLHAuI7QPnCgBQAGDQ1lJ6efFn9gdJjfEGJ6F4VYXWDIO/4Jf5Kmgx8L2Q1iGDjEeBC6VKJWm1
CbI47ybQpJ/MAmZiCBhusnjsOyENPbIsArCp3+AAwsSpbVdqb2IxVWBBBzVqbJOO8K1AKl+LNjtT
EQ+OGGSTieq7c/xXAalS7r9UTEQMFUf8IR2Rqh1l90OCwk054acvIfKY7WrC9CYcc9YV2PgprCgq
jqBU4E4CDbzxr7buxCQXPxnOegvf+9EVrCrovaAoWr073yhkMfj8+OZ+QVBG6nChigRT6TgB28Aq
p6GFmry+LH3nCARn+SeGTS9/M/K62TQdKwJAw06L2CYQe8ND3mH2PoDevVRaiYYR9YLxkOEbBw5d
HCuG6y0SHqqHk42a9fqwJQ/f1s8BZJnk9R+0BptTeSWw++KTmXHaNd+HhKK0zGATYr94+Sp1L0D4
SNm6QTszb1xgRPSa5aI7AjJwB2Z1wIK33GLjlWZTHP1wzQVbAEWgtPDwSx2gIWhcTxDfacZZCius
JnrUz6KBuGX0TZMHL1VYoFdRe5y/BbQs5qOFFabQj1wUmnn8ygHWRFvBH/2+qRuqcnl26n2V7t0C
Fb/1GhfiptbYq6NRGplfPgsQOfZKnTDCRpscSfM/wfv9oVNq/aqkmeP2uZq4Q4bldw/Nwtp71wpQ
KiXzaOP2hnUP553MBUjDDeERuNwxtz259m7OZYUiopLV1XXfQYrwViyKsRrvckviCbKc4Kzg6P4w
yuht/kCIlJ2pNbxhbKIqTMgY9ijUOxkCe6PKfN1dn50tjBzyQmKO7cwyGd20Jh0D1Oi1ieR/Vav6
phnoNQh/dty8ovrFIdgQqCiwcoOt8mVMywaJQN3bZn2CV5HkJ9RE+z6jr4tVL6SRWdFByykZk4o8
98qlgWq/gBD/P5e/ddlpPE6FFwNHX5v779WMNVTPRhyN0fLFznuVZiYBwwH1eXPViVv6/25vToJ5
WZvJ8S7+/4NsKOAv6WnN0k4QQbIE35JoBaNFsXulMckkJ0SngysKvaHfX53xQFsrwmMP0qPYT0wT
Fq5TrnrwLqKYHypIdf99AzouuL1m/ZcY/l7Fgn91idxHGTpccjmBwxyO0KdMfL5+k+jdcZ2/2xkV
NaFLwMg1bJOHp7uEk5u2VOCrc/2S7IogNwuoiuQg3PtD3wcd+j9NrfUtHWu+3byeYLzuCB0IoxRf
OZ69Rp0nwy3FU60FmSTT02rVBPbH1/7jgEoHL6IpRZU2XvkapYvGy/j0R/kKSNbNniLRh3UX7VxK
kg5+vA5J8XZNBYoKDhIOcmb2KGioRru3XH5OTZdDah9hD4OOUBjzLYwvreZWPJ0ou8PELwE3DTG4
pLkoIFEcFmJFF0/0ez3t+VP6rUTSYI/ki34c2CGvoS6WFJ4zIH/T065icQbI9Gu4PY/uivjY4Njm
K6QSiP2q7ExLHMazq8o8wIHbtbNLtL1LH983MxgOwNKC9T/w6KEv3/+R5cNF8EPNW1dTYh86ygLG
0hlsGnHVgz1sNp/LDYitJYugoXzo4dYteCIt94CmN5bN0WzjXXDbluAasZWVov/IlNMQvmFy3io2
A4CQ8lq0prCoHkcJsfclBrm8kx+BT3K25xNzIhOLZVL8JKLW/6Y1pllPmMGktb6tbYfNWtUGm+jn
OwT6bJbjy962WNim5ja9iQLW7GvcrVCAFUjQM7y6Nnn99wdxsVvdxO0rWhb38n/YO44HC5HEsLEn
hG4gKOOFnGQon+Z4NoOFwyez/QewCZYm/Sck8otxABDIFq7NWQOLfS+NkHSrhY+vN/fh7zwQb6Lj
dyqYjjv1/VAUrnEypH0AWoSOR7Gv3hWccCM9s+7bEomcDZLSA7Bma58OQin2gI/WemIgqhfamcoE
icxXa7B93T1VY6jtK9BoM8s0g3/8Lfo8e93ob+w8KY93GnjRUZ3WcsRiiLct92U8UYX9z9HSF3Tl
rx+5SF227MdPS2tEKs/5ORoltwgLQGkUN/N+zCMVJZ4XvWaBqGsk49w5yz1CaO4bhrj2MWOMrImW
k1Jvo0eo9zuJe2e3eo+zIxA8hwY0EgNiiqrvZe07jYQcItLieYlWvB29DCSQqrZq3ulB1ePFCufl
COJgsnl3vAAraFtPuun8j5Tf94XqyteFVK9qPWaW/JLP6kL20XctUvJ9ZELFTjupkd4Mb2OPEKQ1
wpgaCex53VGLnCosboCRAwPXNZB66vZPZLKvc3aZItqEkY33iwoSwaaZK4AcisQjE2SiydMAQSKS
9gU8IN5b4/3MJGRFCegaDXw71n4P6z/AedL1t4yaJko0l+/MZlhvceVpMMtvV2jMmy2F23D8SrTS
sIYUEnwaFk1M9y641jQ0A9dalwF5IyvHo8dD1vObWd7AtjtjHEmRDf566UQdKPpts/WWdkyGx/rR
Tm3Izqq4XGyH+N2SI8A7xRMxGADq4TDrgwhwNHxXHuLYGlxRCSkqyq/iwhVQt5svbsuhBicu+gY1
CTRZTSYExqIOQP47pgjAZj7BFIB7IzqCnNU4GZlX/cbYlfCElFJAZ1JGim88dt6GY6guuiTNfefQ
WmXoY40rbrUWGrEKMW4J5GnrCRRirGqBvaegWQwmwu2cLRGZzX+J5ReBVku3xIQVo47lLpxTTH9h
QmOTjNUZBtXG6Ho8pFgb1J5BVvyzG9DaReOGXckGjZ2UV1n4P1LaKZi8wgnb1aqYEntogpE6Fkhi
gmacpgr2hdUA1ZPlulNxVjjLRyv9ji67ZQBrGDOF63HEvlWFxYlCroLRgcJVDz8w7JVG8oAKYWcd
xp9rdKC/l86wxjj70egV7R7khzAkjbyYsQy6BFn9JFPCIJ062Q7LW+ZSnH5+HuMkVbN55zwZncEO
iHy3EnThmUTRBqpQHiDNkZuqJ2Yq7x3AhwdgRWYxhiia/9NxOpzAg8wIH4WVmSCL97C9W30z3mc0
X0gq8zzhaJdKAWWkMtC8nYx2S+L6QRGrPWXC2wh6lEu0Y2OAMREMHI2R2yrJ2rXdJIBH5jLxwQZX
H2K00LkN+Ti+EZmT5/xPnegzpnvTPziGXVn75o8g0cFgjYeCaGl8xrbrYAyuz0A402Z/pWNpHQiW
OWczU8z7xSZBF0/DFhSU1/1+3fJKmjaWI8lUyv25VYRmKTEbL2kXY8kX0akhZWVZFB3USAY+08dJ
ebTIBXRSHvZZVv5qRiuuVZag6v+81utBU4Z3ktpoBkYzggJbvYQQmtf0H5XLuvcKYJwTZ6ybE1lq
bA++MavfHxhYDACMlsdtStdev9w8VFp56upEDtuCUKmpcRoRGF1/B02pStcskyOcx2CwLby6Ai+m
Zz/yF39ScJrudMIj2Mp5dwV1sm0SMC/od+gt8vgy/es/ggAA/F3Xw0j38LDHvMCQie03iWo3Ogr9
DYD1Gra4Z6VavPtU7yUOW8CBqH+n5FckrYAn1Tnikcj9UHKLeUgkbhFw5x54X2yrRpRYluJTi7eX
sCJS+IiW2tjnoc1ngKLzBJ+33VldKr9uD6zManNxqKX861snx92H6COmXr8EdQfNdgu2Aeqg456X
zbbSfkwgKMkjPcgh8XzRavS5HPfuMulq3XOGmPOGSL51XfCp28l/R9HcZOYaOJzwlDDmjaRdEk/h
B0tN8t1ngGYVdtK5QQ9lOENgWh8McSt2bV//IQXJQLMaCZ3ukgBjkVusB1Nst6QbkWSbfdK3fvbm
tSueAa/OmBDZdVhXw7nAL5jqVUeLp7MMdRXn0HuntVAMXxhnquOWCnEqofO5lPztMp1Af30Ch8Jj
lBIj1jHkQiGmUkIGKs0DQQhJ0hb5MM2H4T20mWD/NZJBdY9XXJFVQDkOY5XN38oFNO/oGzRLlMWM
y3m69XPaq5hIvaoe98GEwbysLXyRm/91B4ueNRKbUt/R/hizreJxpPXnTAydrEspg4/mPVGAdz8Y
d9abLFkI9rw9Ue09kuhNa52b0NEKl2zfg+52W8e0YFWhgOBCLRkPcQya5DsteC1YNYWL5UmfIaTH
ScuVpSJCMN+3x9LLUQEa9Y/6ldDrCaOas+haX2Lrx191sua0i5QHW9t1+I50a6PlX8t3xTVTRB/6
ZlaRC2OQ+7k6/Y+oetPva3nSB7wepqTiMr1MNuy+xD/biLqcTKY2aavxpoJwNixcUDO7WzzFW0QY
+Ta5+YzzEGSSkhjTbxS/tvdZJ0nzbvZlg6Ymafsovm7PIaRf5S8PVJX8AJTXcaA71JdkJx9sGR9O
8oc1NwPSPbRLH+UUrTO1ybC3SjEc4s82F5c0n3JO/DFhulD14oeMPGfjc2PjiLErvtPX3UIBM6+B
AcAii094SH6OuhU6my1UrnSB3ls8jaXsT/XKH+wL60/U2NyycmUfRUXoRHSJm7HTbECdaalOQY0j
anen+4RSbFb4UKWCFgvJ28geOEH9WbQpDg4sBU+DcZNVVBFYu9IXzFhUWyfJ38kVQxf5AkuI9u1e
RgCuDrtPBoZWXMTKeW7MD90zYk/7l5Z47oRO/TVkb2cDHPfXtAEWg2vWhIQ5Dw5BNmzffmk+eaeV
kiLYABgLrkhKdInO4ENs1l2yC0Xl82s35ObBhQBr7UZpzBGneqsG3PkNrEMqVqwRKnoNbz0Dzbxd
ynT2nI2RGisKFFZtjcSbNQJdXnIlNPXQ1BK/aNpPRcmRnW8l9Trl12ajxpVsErz70X7/i1bIU0Fs
XEg7bbLk9cV99W7lCFMZZ/68lEJGUle1Zfdev8t3YczrxC638TRQecP0uZKAnSxbM3lUlJ8bU2Qu
4vV/WSrJjPm//k7Y6n8eb5URVLx041mcOgp+wQz6eXa0b/0ESSZ30RvUErYuW7fc8e4LBN53iZ3s
q8GaxKwWGWewp/edbvESBTZJHAqFr4Ow5lNedNg0ivyb/i5yfEa6ZRMLgTWSQNWECtle7S20ppnm
PW6/Dp/ytDXX5qqnqHiDSocEx0h4Ub+UdjvhdKbRRY4SlZ3115RNQzswPbOXk890/ixw993lqgI+
sFyymueZwo1+9y3JvTO4+c6kp/pex2eTWHLqzPlfX5aoviUMMbkgfClj4nesHHg+mi0k2RGQIy3X
3czWUm0hOMkK939mUKvoLk+1P9/QU0Yr3Cz1b6mKeP/EPW/JfdoFcMIlhcyGKS+M4tllF2XVkhN5
iR0tC37JNCt76XKJhdpmr0ihj+T2VD9cdsEkRPFUgE39QNBxiyaBpbUMkmGemSIMsw1VI03hDv2a
gECdKL6n125mXMx3isjB1iWSwLlbYKov2jXO/Rv+09FQZZWEmZmDyei2YPmFdYepGVN5vYh/6YzD
3J6Dxt6iNU5sArVk6zQ9XEiP8V2v0+p4aa7w2hnThsxvRVWmLS4dfb96+D0G/M0tM5J7A/zeS8tm
HHKeoPKcmKEeHc/xYrUh9y8xJSMXv9jlYqCPOHYMoaEws1EQaGUmdL/3sqm3+5LxFNVXI1VVy0jQ
SueMhZyE6ex2WA7mXBtKWkLhVHR8ETeMh6seU8qdEqvqHtOA1kLzmlzkgOH/Joc+4gfCLk0O8gAA
WC4RqK0B8+iEpiHXp4669AtkIYLwi2BGodOGp7ze4JNprjrX2gyQPe6ArCJWBAfBZM9ZanmIzOdS
9XzUWvfj+etwKQv5EvgNQ5hskI6HWs5kbagqJ2pQVF3qbpaeTnZdUDtSoyUfTBxqdmB+CQlX3NCD
6JRyPrl5YJTvrpxlW+6hQth2kESPt9qkMYmagbhsjJhLwSfWgUqN+uGYi35XUmWLLUdZdWzFdEiE
bxMxHWScpzqyIFuJx02CyEPwGXVWPbcMdOY5ufGxechhi/xZJYIapb8nVHw0CZwHPnm+XU8trb+6
Eqbv8Mwk/hsHzzIZrebhPX7R0V7D8mYAJBuD24dPg0a6IvlbAmuLq1LD2xgYnVlJp6aosz01EY0I
r2mVXYNJBhhTZoidKGrBdl+x01CTPC+NkIlKGofOg3hb9OiJu4zJ6PtyHIR9E0V0RsCR4EN+/K7h
+rvDKEoLjLorhPxq7LFhYGMMfEmRsh/AKbSqWkvPb3mgYPYvB1zFDTP57pW/O+i/QQ26+5ICTz3h
WbV4cMJ2nikbK7XpjqNZxfszb6TBKFrnHTPkVE67D1UjCWi38uH5WVuRxCMryAusxAV6fb7z8yvn
/ASjh8+GJ4Y4vmNzoFLD2U3uIiQGBc1/5K8R8fAzr55s6EXDqU1rOlXoSebp/XMRT1F+oD1h4lFV
a4bJeyOUQQgDSHgmRC6iLGTvZ+T4IIElhvit1lzxxr/7rKRibF8HWiORZ3U9SbF+jrGI4/aOZ5sR
5pR5+8M46IlhqMZ7b8GhWTzQ7f7uM+FyU2plWgacVEcCYSyaVRNIh3w5ku6Ckuz4GL7OzjvxCw1d
d8Ub8YYdHNmg3xnkT45jS+PkTHWdn2waanqC1Pwe6v+CI0Pr8s1Yur01KoM0VjVaQLzjCQ5KVZTh
sKdq5h7R+WqVomQeCBUQMyOd9ui52pbvUEdxNic2sHJd8GXz+gS+HBRwFIqbVC9WEM/L3uV/ITLN
vnyWhwmcFPVhdv/MGHaz9ESM8dRRneOucos+snv7rgUwiSBfEe2FVl+7XavIE0p+m4OQa2t/Qdtd
ikgO7uCy/YMoFQdRgFB0wVq8ZcjFwANhv3aWsAheHfSHUrWZxo7WDvADJFn87Q/h1qQbVJIouuNT
boh9qkW75+Q7hJqn7hya9BlUJTS2c/8G67JpJcY36UTnctt95FupQSKCkq3S98dbSHpgSZR+n3N7
OYhAhGVDf6qzaLAI5pfkgzYY4rf20+xZGug0dX/vtxqQI3uVgIGGD+/RvrO44ao6VIsEnB+GEkyP
dph9xNVGCEEHB4k5Zi1MkKFnncKVGKNTkTmfYXYcm2XT3967zE1C+4zG+9w6L+S10b2JaYZFLEdc
AgKyiwiMABBF2NRO2MWutTFuLrkfcuOm9+cBw4VVGyta0trUTtma4iroDIPawhPeo5K52IHryR6i
uM8tWIj29YejtwHyMty0vdg93c2C00t/ssiQ/by/pNm/NUQxr8DZtr8KqxgVr+s71peE+X4SupR6
noIPhI782qLJYmoQs9tymY36Q++l3DaOewHioRwXLx+uVV5QOZFaS1tO+B/dO3GTHjBt0MvxfTrJ
i01zFAl8iaUZ+KgxMlmerkUhR6jFh2S36pUSqQtZ/h1Cn8RIgS9RC5O0/bHwIQmn5mChDmQddn7D
bnNVJbRsqjBNha9jwXyB8Gal6U7D7irJ8JHeZezyv+p4aSz9uo/XPrqnNws6yTKu1h7oXK2ovUSS
KdP0j5Pzpm6dFupVvg/IVltzkf+tAPMYANn10uVQPUAR0sigUqBaDhsUJmq3w/keT5uQPthnrvSb
GGtc28SLY9ptu19pS4Pp1d0Am2c9EKhFT36gZsR4NQ8qDnttSUS4vSrWpxy366knaCY8ZO177a8Y
t2wdBjVKwhC8iCS4ZO+ne5uUBel1t4j7OhQoDO4zF7XnKDouDBpyr0ch0ySfs2TlPtAA+E50NO1X
69NufH/4GL0NKhj2xbLkbCrQ71ay6IBSIE/fgnbkXjT8d1xB3K81+sfARXG8qikSfZ43Bo8pWCbC
EzuRWTQNtMqrrXi53p5+c5YzFbS6ChP5S1qnMeuA7T88Co/Vqpwb6KjBBBCjzJ3rYi6UedbsA59y
g9kSzyuxsbrMo2xHyoiTDc0Y2uGWmLgfbtet5lGb4RhGZ88U8g52iX+zaffHz/foXwj/Y9YEPBWK
eQzgUhBDtwt0qihxNECxgTeMyTBnVdujWVz6iKYqGMohEosd2O2TbB8gPUAtTuU3BKbHWlsJmJkn
QWGjOSbGN6aW870+bh9RiGZlE8k1KIx7AtF1I+8CATX5yIH2pHaL/Md0KdndJmahIWfWBLzllbjr
0NmJFHR+zHKOJkpY3OmvmDyliIk5SltBzALEJnoPTI3KzA5YvAN5xXl4k49/9LvpD2uNQTarWnIf
QT+fpyPKx7G1RwQg5uC1RzFR7wCQuHEVvuUwmu8aoGtPRU17UNQcz7OM2Pmm/W0+6NinEdBWP7Fm
uQvfVxZcL2AEyHwP+hXeY1JcaOooMg5c32Bvj6ClO9WqpDM7RSw4tg/HJjL/Oe8nv+7lB0oAbHwZ
d29sxx7xaD7y4VkjD7h15TVGBl0k7fUhxW4c2kciD7A+kc5ociVboNSDcycI/J1Ecf4upbekK8PA
IiEzu/kMQ5nBs22YmZK/n2vEgOA7LH2cH/mh00emOCLxHg34FVup/RzU0LbQpRcKkTZazSWbLXRI
CRc5AsCK7k6krLOtFOfq+DUgKEXO7lwKkRfwjCpfUe5qjM+lQCCFJf24XcoZjdGWGcE7sBoQMgKU
VufWSirfCoYLk6qLn/ox+0VV9JhZTUcFdT0GvX8gvvEpKUZfCzDQTouejoecN1fWigjuBIjm4sYk
ESjhc/hB6WaLI+MrcWnlLt7dv1tAdPE8huCJo7f/IDPL3qKmmXLVfmPZK2GIDzMJzs/oOPKAHWUH
bh0B/hkBPnciMkj9Gh2aiAJmR1udvS6qO+uE27jQmYxymhlUv+PPt5C71WToW/zto6Ws//Z77O/K
D55hQOA7q2KZukGGNhtbwZqOWeybVfMLugkaG6TUDSiHagt7yg3cwCoSK5/p2hOKqkISHMW6gMnh
4WSZgychchG577EY1Q3eQ9ZIFLe0ftWP4dFtA8ceuKr1cDQkAF/N//I8lPDU1OGf0DRjJHWh9PSL
oTF09bWzwy18T6TRXG0WBWOMl8/j2M7O9ywBp91NHjYVWiWeRAWxQbPAPf049T9L8xkRiDYO2+CJ
RM3leaElvx29rsz31eyPH79xNcduolKdmKDNl0S848iwzSCZTh3LCndaS+d6WBboL7R60g/+PWXX
AAb132e80xVUhe/OBwvuUV1AFCDmohRtDw5BVSJFAEApxrtUJVBd7M+qDFs4qhtTmQ5Oo3RkBr7J
UlA6wc76Y/lY3jhRnVLnBIXHV8Z/SVnz2sGm0s8PTUKrPsY10ohN+sQcvYzXMK3bkftICmFGUdC9
U4e3LEQymzQPSZHRHdi9Sp0KKNv4exx4UIB+Ho9qg05DY6dFbyOR8NMcLZbuMT6Xcu12j1t2JN4/
06QAUk+dMxE45myZrp3eaCQ27xZnBeyY8e0G0gGEQVVI8cMe99qSnN3KGuEp0/uk1wUFdcLwcZnl
ZTRb23jj9RllaKLbov/tVtRk9tX3lWa2kUrTcNzukMOhp4OpoSvJab20CEOSh0lJ+ATewwblVYNu
ILufj16ksQaI2tYowOBwaB4S2LQI6lyHFeZjhKL2kzUvEHhwgMoGyplRGBDKufYE06tXc4zbp5g6
8HEAgLQH2eff3hMPAn01BILoij/iTdbJ9mCwSc5407mO46e5WPwszb6Od88wSa8jxYz0bogyoQ/V
1Ywwc4ie4anR6bdrl9fey4r1+XQNGm3qM/ldaENAsPcskXV4DOxEG78Iaovr3netUQe80FEUJ+KP
kNkFNE1nCsIbSN6wz4O9Xi5Do544JzCv3RdutJTxHUYd011FyQUdNDZLRKwzTxuO3yZkO0oCQAbN
UvrZ6hd86u1NyG5FfTFHWZpekJ8Su0QuxEogUL+VXDgbxS9pDx1nPVbo/j3fMyUWztX0ez3uhpjH
2iWxTFjDGejYnrx8IGCSAEs/7Pr/yHempW1GCBuSWCkbg6G5B/ppSUbenvYCfSiv6uO9VekBKaqv
AwIGWy+wJU/IEAsy38+FqXGCGdJfw694s18J/+ajkhB0W38cs9HFpwYB4C9CYcZPRzwqGfZ2EoFQ
vJOHoSRN0/dNiSRmf5ut7WkRSBm5eEuzJdmnlV0bzkykSs6LJT0FB7oyrWwob0cCujWZ1kpjuMll
DMfBF0R70cDWvbeIT8L1vuwKwAQhJ5n5JQsGMEGakORAzQEvEbZ2DUXBYGN73wO5hjWYY2UU0vcI
Ogi6woNhqe03gYX0Aol6X+IF4VGqU0SK+i4j+o5y1AmtpO1RimAkfs/YYQetbbiyaUvKl6Yx4gQ/
iteu+X/wlMb9Kp2j+gB59Bg5mZ2QQrVZHinNKM0VSZgSDtP22IOI6Re5aLcfR/p4iHpksoSkxMsX
E/jNOZJp6cPpZ5mHV1mX0Je5kPQbO2MTeE4n3KxBPFfmk4Tzg+bxH0skgXMpDDP0IjHuluEZijz5
3nfE0k5t2aus+pW9JetoMKHcFCBwG4lp7+fsedZ4Iq7LlfRCbTQWBjl85nTPaZ1hfQ+4uQYXaTD3
Un5y3hXDTnllDntIFKCWzQhyU+XrCP+xB1cOKgGOD4uMcteWxIEYbU43Ayg9IKDKuqqnADNCwyb+
nCdqS33P6lCJOLZPCIMapehkoXsRvdAVBLGYj7vRzflTPMpYp+IjTvzG4RMSuo/soOXsq8n3Uc6a
A7GWXJs8/gT9BKMBHWv5qmxJLsbdHtKiXnns3Uf199gAyoU3GzVvo0xK9BelVqJFEUNMXBTFTkq4
i2Tav65HmwYMwuax8woI4Z2Lp2v+amuzDsyo8bKM4zk+UiNAmaFfrlswXNQOiX/3KIZIcvD86qj+
42aY8LhJ8pDahvNINvQHAloUHCs75WTS0W87hBYb5UEXti2ySc+F9NcUJuECs/KRxyXuAUKP21zw
IlRZrq3gMpU4CG7/y4iTVwEqBkVOanCMYj6N4jX5gU3aCcw447+B3mRh3Zhbq+iwOMdvcZTVTFIM
9z6YpgVlucjHWCmk91b1nwAV/4NIEOtc6y6cLEb47Ot1POHiPodUfJ0Kfz5/u5v2smZJ5ToTnbRc
AACzPQ+FrBvNn8GH/fhmejaLIvS4IN6Fu2B1wADRrtrQwk2es3ufrjH937xaGdNLNIuMlfZgmsYA
eajRyyOMTZoEh92fhZZJ/YFjeClJpL38edsf8BpINyLORBnzeAesm8ur8/Njw37Bwb07TR88qNZL
TT/stiFYQLvTqFS4CJE4GytUwqvNs699X/Xh/IBElDPqp+lfApeQeEm6l1gIF/9gOpfMSZuPo0pv
ZVlfbGQINl6YE/SwPbZQbziEoiR0q6Q8ri4UyEf9J4hNPhelN16deyk/nE1SqGstvggdvvsIx18C
vJ3UiIadnG1OIRfqX1IhrXrxXxAhA1ziC3MZQKCBCKpwdSiWy6L5t6vcKUtrqkhxgBhWQCgAkjPg
fZtUI8Wm/LnZeAwBEer6okruv7JmzGaYMnPP4LY/l2HPb3fhiNZ2xj2PBvdyXI8a2bgiibNxC38S
b/tzL1J7e4kfXSVz9RbVS4bCZolDdAu+N+twtnnOGOz4xNrBta464d87Z38MNkSBLbvz4OeTaFQH
teoIEYYPhq4biWCTHBFd08pHXRiw/QxvmQiyly4JiiHjsRzcLRdEVf2nJayBPPZa9x+WfiYiXz1C
d2jOFh698lOY3vvC0nR2s6XBQRAv1HJqhISvJfT7T+LynXAnrE7R8N/si9FJ8+gJg/Y8NkwHQHy8
dCyvieWd6z1oYRnW6uDgOlnWATrGYlABVPp6BVUfy8pK8E2dvMRA3WdT+hP885rcSbbO3eS53Qj4
ThTgrEvg3d9DsqYX0mlSSOIJTDVTMkDTT/cw6FHvlQbp4QypUWuTqInZ18At5eajo1w4KBbOWRep
lFqp5tXpEVFV5gMfjK4YrA7H2DwqoHnbhaXn8ZlOl93VNA89geoJwJUIhnWWLEBFqpPHJMjRDtFz
UmW9zer5tT8jKOAhUvERCQ5hc7g2xr/I9Qx+Er5X/fL6B6UCEPJfy18n1dG3n9VnJszjn3yA6t6A
f9YS2uP7gc8hZorQ1lfmHcBPsfJgWI9GTaGdWkvPVAxNpo9It1ufkgD14K8g4PDmrKQ70og1b7N0
B633SNbdpxNwIhvYnYZ6BXAnsXWaFaKyxQ4x0iTFjjUTqmm0wyhnSHSQjGfTMnWpp9xReYBu5fuq
25IoKOzV9fH7wQ1o0onpizAwDuE0atY6m4Jz/ELD7TmQD5LXM2/KM7f6vApOP2pAiZ8APGpvagKj
TbOajaojoP+dHzXVewVjK57DdLpKPADja5RfmVjAK5rxFLxRrJ2Qeqn7dX6rJiSvyIAjyAYfhtSf
LRsqswtbWhP1Zz0/ptnawImq4FHsgzV34m6l8L4lZGXhqQOcpoS4Gb4GN/vQkEdDTW+s0+tPEH3S
++yKBysRYEW8ML0vEq3pTtoF50aivhTKJV+xuPGlqmPPf4ET9WWyoLtd4aY45W6HBAaD5i7G1ugf
it7+9FnxV9je0a4kORasK6TRc1vCvmBBCn+WBWA7G7yoSl4FcqSq7dV7HCQ8Ve4yUrkPdzdT/ZHf
uFXbzuLuCREwXuGp9DOJvHaYe+2qvz7DgU0BQiU9sWsIK+jJDQVRoGG9w3pJ2SJAuicOYfIqYA4c
WutjfDp0rMUsLVLuKhZdjHkVACRDeGCat1+NMJqS9EE0EQ5vgRA6fi9Dq8FNK6MhM6xtH2O7cv7w
O+q+Axux0qa/qoLWA/6l5Qpgo2hGSpNxr/pSqjCu7rhkMehp2jHsm1dNfz1Zn241SMGn9VtD6Jx5
gWM/uHcssU7jYONqMu378aMBKYEbHlXgH6J1lQICMXlsChWYw6cjqHu+bPaZ0rfNJCTRd+3Mx1p5
hyUTZ1l7BvPEQbMmca5F0oh0j3WPtUQmHHOVcHYX4zICfIUWr5tPtxs6W2dv+K+GjMZvGacqQFgH
AZguzx1cwXw0j2pV9n5yyZ0EZRebhkSLsVcWDFaDyQcTuyBD59lVk6fM5NNNEkpY28kWj8k42L/L
XMgsg9G2XHyJ45/aBEzK3mZ5EZqVaivemAZdgsjJ0o8wrIr7VoAJA3BCpuBrQEqHmGQx+xLHQUQO
O0gyRFHV40p3UPbyRvN6WfUJ4ohRojARzSuTzqzqijnZ5O629Rw8lNWC06LFQwBNhy6FtsgK1TAB
NK5NIsvUh2woK6arhVPZfbtHtKJ+TlmNmXXaBXcn4IMi2gk+27VuUa6d620xzn/Gt12hL7trMq08
Hj934WQhTMfSC/y/IiahQJeOrnmU/jMtx9zPha+bG2239t9Vgov+w2slbOAFb9Aod16s+HJVk1LC
Rp1NxsdvLhmbkySSky71vM4VT4ZvwqAEj+lnGzwL8nokxnM1TDST6hB593OFFEForNin961FImeG
p35l57Vm6JwYtq9ZRT0zC7T0vZiJhQqNCeRkYmA28rScPHWhV/WsZ0QMWiOdpC6IhPK0IgkLmdsY
gCZe/zMJdzTiCBKUS7IcBYLzb6vgzApRdJaRPk8Ge+iifJ6rMM1Iv4BMXhWrgTpcHmkit+wTPbr8
dK3o3BJO3kLbKuconlrAU6JZ09rsn4NwtnXY2DGhYpvckM9epnyQ3czLKfgoZG5SjTgB3FkjnfxN
1ALK16DoRBz/Fwj7YiVZb+WwiSFqIcA6w1p1V8l3ccDw7HvQn13vKciMOVR8U84A6mlzqrObOvWR
rmjGPbR0dbU5K8pWLcnEE5VMzOOuzxAtIiyWCGS3i2foMjX1LAybSWORMyE6HvKyK08abgFljqyu
6Psps0NSJs5O8kksGxtI534qwO1bzBJPgo1nO70AXrHQ7SEQ/ldu7PX2FP42OzPOWIGvWaNcmmNe
6xlbip7PFMNoK8N92C7KDhmRUrRRt2mR+YpL4T9cSLwJoaRhiBQb3kDI7q2evN3gXRSnuXZafa2H
oYWlUco6IE/y/hK2+8yDAjzjE6BAGcQraCBbEd1C7XL563Rap64QaIOJHxQExK90nf/Wnc8bZCch
iyHV6QbdWSYxP18bs4Ahf79Zu+2iaQmCauqn+i4BDrlbxw7uLKW6sAYqtMl0CPaaLYF82PpQF3q2
EPdcAG3JqUtNb3sCQITf2AHkEZliTYNmGGK2+JKW4QqN0LKOThvcJ9CZWXf/3JyRxi/v0cVY+A1y
+N4FUYR9uZEPdkvIkz8hGsxVg7P8qO1l0eZATzDLLA35PnQ9glGHAsmim4d70I0iOoTqBIwEUuSS
oMlmyXCVmkXeg1iVGMBLtDkcHzV3wWzchc3DpZxsG4T9K1Q2s3j8uvxSTgcbegZxWy15kWNLR4jq
5Uid7lLD2PPdRw99GASf6Zo1b84nczs1jG069whEUJ9glr2KELVt67Dh+EOsH0fGeAGv+JbE6KrY
/0hNwOqDcP48GudNLlwntJf7zmkCPDpTqt/APoz+XKr2jPR9jDco6n/nsW0cvAyA7evf0EU/6NlR
QQtS2nKzVZ877196R/9y8V8KEMZnMVdA79dCER5efif6awPQhSt4+m5PmxoJRKCtzU+X8BRrvCNX
A0wCQl9kTcIolXGzxIFHPHJynI8MeMD2F2XbEabs2WhGpMcbYBMYjNMojt57lDzYIjwLZRinhyIB
n6wuox4ltQZuO1N3DKrtMorMO8AL7UzKfwKpo8N4Sa8jqAE/K7xJY/WxwftafOpeh8TQyR0LuE4F
iiyJ/YxnFrI5EGCdAaq/JCYep+AL8Nt/HURiuyYUJr8VLl6JojJxxfjImjeZqarIDnDzCJBbYeYK
gcxhjAkgsxbhULja2Fb6yEGobLwG2xXzN5Yp/q24JkSucIcDPWQeUb80do8EQ1p6Et/oQ1/8x4+N
EZy2XIeh9+LAiSrrbWBt5XWjbMyRtG7dmiRRkE/++UHMXyzb+CmWvUBUQeY0I7D/2y62BBiP80Yy
49SqGNeEq+GnpSlgcgTU/kVMrMj2Itu0hNqdh1yKnEZK+yt0FcN4xIrUQj26XY9gX3GEbyQMIJWy
qKJhdRqZR/248l+OIilerzbxVTUpe2Dewt4tDoAxY6n9kqheWN+nJ5PZU8C9v0sj75HVmxg+t8YP
OqCi/XW82Ypw7vJXa66wVyLvOZ8UoZf0kdNv2CAkfBjJbbuNJ0WDe5HczGuzMN1wka/rfHyWADhk
kmyBN9PYrqc3fzzGhlZNWmpDgqV4ApmdbSEo+MD4AKAuTx1/lsYqw/m8hgGxiUxV6FyowGQp/QCD
LHWBa8Pxs7gA9iAex2T2rr27Hqvbyko85oJQ+vZJh0li/2QEqigu5yJHn+gGJc060K4P5M2GmgIO
BrxeMVPLkrQ04VGDnzqcbqF86rjtzYBLS0yiFzybznsWq3fsLLgIiOZGY6XWRCnZPw80ieNKAVjH
63zij7O5+Zge7fjeWld9RQ6WBWfkG2bHMxWAHXzCicyiIPzxlMGn5SwtIHsGC2BnPTTihgrLzVa7
QYHL+e5ac+zUCRLzEqJs8585g7KAtzgkvvHK8/Pvjpn/CFbwHcOzbOei+nY9p6PwnZuRBEtmGlhA
fcnGw6ezdQZxarU5Stja7yX1NeoGLAiPXJ2cQlAVwUlfjGx/km/+R7bywPSZYKG4xeZ1lV/gkUAg
Y1u8Cuo9DrZYXiI2gyHbGLpnOYMuO8eMYNOWhwjjoCiCppO7MRlixdjecMRWgry5NgIoUABaI14v
DE4dGl70qOoJJ0vWNUX97vbCNMyaxOMsnJkPiDgOsNbvzNQN4IWwDTQUgwqB4n6gUN2xJACgtVoT
Naxib5KrillR59ePXTaEc2dJc0y7UYoznHHHA8WKkNWS+azAItjj01pkfwtX8r9TXxJP6605eFJg
PgyZKpWSrt3pGQjPBReZiXcE4AWv3A3vI8oZ0k2sI31sttHycTsjHY10Rn4LUVwEx0Z56Xd66ek7
Ur/5lVLp24CSVG1n/dREQRjOOo1pTgbGiTym29k3nyPcdC5bmYub7jHp/AkRJonNtuykNoJuf1+L
u2VeHpX06FgzUKdP/pfLQTydYV24om0Wy/PFDqLyQLDcsxr/+DJw7SQfdTOHUtP+fMByyDqqT9Gl
baNgc6iVSUUT0YD4TY3lDwzxy2o2DXOk0vfxk4c3fU4H5Qx1gRKO2vR6AzssYSPtTjsrA2iOrHc0
qzseiq4pguj2vccpTVZTGUOvya8ysJs+szT1Y32DK00VmSLZ5EYDLXSRUvSEuR5wkhPQfk8MW9hK
F7wVeQMv4vC1p7aywu5/aoV2eNfhSuAo5SvJdhwPXLuLx1smIwoX01OptZTcXskygnVcbwf4obRc
38kIkFLixB4nq4xv+LbYfcZKXZ3z4lZkVD9Yv2oU0E/7Lcf3MCFCV8dsdBRcqXqUYEHNji6jR2Q4
QXZoGuMwMDcy5DZd5rXK7962pIxk/o+sApda7/8i9xjSIHtYNarFHsKRowdPyOV1Wztk2i5EjeQQ
HX40ROX55bGpPk6Ca76e7V36KFNbRyveShykbzTE4N5A2i2qvhTvNaA6bc0bgrG+1d2mefT/DVxK
waz6H157OjFNLgQXER6KEzqLY5Ogd4l+FsO6s2tEeX/LlMJUrUlXwp9FLSP6bDNwTEYImzgv0Grk
qDySdDXMGs9iMtoKdFve4sWVuos0hcjlb7SzpkGFbcnRZO6HcAXPDc/E8TmhVAqsrs9kBJljfyS1
9ZyiZx+ftel/CS7Tpb8+lT0OwjKDtC6m2DqlJy2wC8jz0+HoGEhOa+3DSigmcx0Iq8nn2ytF7rFB
Ck/SrAOoi5vaHTbFLka84uLNF3jCTBXsnsuNVZqRvGuIxxC352bkWlQDoZl/+DXl1SWz1K/qQitU
F+O06YT/KeiwXXAxYQYBWiWI9ny1eT7kuUhU2aDa5aXEtzy/lC7KjeGFIDcLV+N4qPG8JBq16POd
Lz80vtNgqyh+GQxmPUExmrfJgSXql1IqSa3MgxVn+vzX/0vZ3/l5R5RI8s1kt1Gf8SvHUp7bz2qE
AZhWU+IwCrWZRAjU95WopndZJQg4GCaD6xXVBGvEnRldi9xk4FZJzYX3WFSDKKPO//Qa1Ea9Kx4D
K5yiKT2J7C41krqeKnHg1pXKaxI/wtUkjqBqdBT8BbImVGZ1tZ3yTpePC3oCuQ1SCF9hmD7JI+kL
SYt3g43e86mEQbsZmrjzDlzsl0SHC90P51k6SZ7ir8aIhCNNMTdgSOb79mY+cx79AckfbU1+0npt
8MJ6rUWNFbVtq214O6wR1ruG+uOeEjL934eOz6AHalLS+0Z4o9l4d5y8pT3eMpddJw85i2P+s444
0hEIIdIRTk2fYY2CprYxM1vV+u0V/Jslp4beCclGha9h7+zMLJ1Hpi2oTUAgBls8gWfeubIGTsv1
WKa1yhNr6hlwnQtSpWpFDbH2K1VaVqp5Z17Bbl5G3b4D90OdWRdg88UQiHiSyOaC+uvg3jGxmOHf
EVOIYssin2M0TWebebnDDVxednxmqwY/EW/wYdLgG6gzBKOjMt1FJxzM0etG8cthGvGYZ1jmLCfa
J/MppIzS2JVPlJ2xrkRohadAcG9gmr/ppI/+Zju1GQ3LXM0Z3BhI/6xisMlOvv+36fsoYjg9mfOF
O3AWHSHFrXifH2wB/co5OLgFAFwOeow7k9CtRlZ+1QqK/2dh1OUBFSqGb6i599OcIwKcJfdGEyM1
fZiQPV6MMklDLfjOX4YEbMv1zU+QiyK8mdEzjDb54wdD39EtOy9bMokoXBfBzrLOs2Gt0bEM/90p
ZB0mjo/O8F4Qf4v7/31aCvFylvte8NUXg5gIvHdrVPYhWPVf62XgiEZRenX76YTBtViI7QkF/6nQ
XiKvA7MQbMJzm1nvQjI9AJRgcOE/vSPyvGL8Lv6ZYDJgk/SnKtZzp1xGvBvxMSJU4OSJnJ8FAgrF
iS31cxx+aKg7e86KmgRB6phbunJJKUmCo/ulx/viz6JAmuGBw7mTWhKSYuk/8nsmI+RJmFOj0PFR
7kdI9VY1TGcEZaQP/qiLS2JHSzvkMsD0xEqQtdcZXfqjpY1CXaucqdUphoirZxzfNDu048NHPGtU
1ItvUmSDelQTOc2XtvpooUyDNKKNGFieBSf5elke95nT6A8vRA2NKwracrt+rNeAii1pWqCVOIZn
3+eu92taen/UczDyYoNDQ9i7WsGnEBFV6H/yCnWS8NeYWgzxSdlxcTqzXv7ta8//WPhMlLtvPM+e
jsBYj6FoBMaTJLD2bn81664amr4kAnr+nqpMOEeOyC1xarsvluxCdW3ZfwaAlVzBf6j6gxZ1yh2Q
VRobxzPdiU8BrYYDJACR9rvW8CfyF4OFa1uKfN+y+VCJl2LPONDYWGhuH/mXvcHIn56uBsrrw0Ot
oyKM6+lAT7Qe8M+umaLMSk3y2RgP0Bcgljo0fjVUhlOfFLq07N2cp5XqQnR9O0oMC8ShfZC5rKXi
CGBOnNqXSvE+uJl2eauycq3eiSGVlr5v/isiIUkU8aKuO/kno745hevWQ9I0GT77N+b4CwsJdYbF
fMqpx0Ro90FoMk25csgaKXH8mgXj0vLAezH21e0Lujc3/C9RUUueaUem0828EOJ0m268u6T2UxzQ
B1IQp7XCXwqgAyoLOLCayykYBzzlRcmad/JxXeDj1sAUOSJ3E2asxi8hv08VWAUO+z5rHo/2eEoq
a73DO8fDyNFFZlpGNtoBwAIbSP6w4mzuzI2jmysDYfDpLx8BfmvDkeYDjC1ON5FZDyIbzqOouLuL
FdDE5dCWHGmP1aW7fOJXYFKUWc7igyKwWW/qP6qOkr8+gofq1TQ2NxOKUB1+AEGRsRU2TiHpPKTy
KvoHd7IH2z0PooR0Ha4vVpFfWZAda+DLDmBSpK64cZEu0mD/AhNphWXTojJoyuo5zPoOmZahtPkJ
FsOAtxfnmxsWhSijUGaX96YeojP6FmsBp0eloi63SgNPGgnWGX3crmtxvYKiMFodUW4z14ZRS2/Z
2/EqxUtCwD/eaJw2fgCwwGdv8MrSB5mRF+qcC7VIpwMcrWIfghANLPMQUNK/1ejYeiL/+IOLoyMB
3wiKLBCSoBLSZNt2htuI2LzoKF/itkNxswspGcgkXsk5+xUpQKtTNCvmTx0D0fTpOtrhdSMCchDW
VdOc8Z6Wu+Psw53DD0STsU6Egtbxr8SUkV11pM9YBozsKS1icHk2vMrovs6PFIYOanPsr1bdIvVo
2wVPiqF5VDmjyONBT+BHB4vXOHYzNeSPI8SH2xCQNnXTfBN5bzpDtKqjUL6LilIycydcvkMrHdw+
+cFdTZaOEV+QvQb0oUvGLj1iM/jO+myZQaTC2IPF52eqEnCbMrXg+mFteQjxxwsrZOZSnzTSY+Qt
zMl6eKyxUdK1jwaKUttMsDbuR9P6hV83ErKC1urvpgFqPKfQTAp7MIeTtEdPyn27VD/6HAYLmNeX
1Kfgjx9DzRvu4b7oTqY0+vQ7eif525I7BcKLa5vRkM1XH2yc/ELtpILG25kUasysB2X9ovzBOmiJ
b8gMfOA0gZUIzfeRlXJDPV6GeTWRcZrrWB7kPUP9xybbK/QBPxWrVJeeSzHXFFQYpyj/O3sE+Yaj
skzf/HplzWXOg5wCFUkizdXP+OLGMufeAAvssutWedwFjKrtbWxZ4L6gc7qwNyUVKV1mH52Dw93o
2apfl2dDlxmLmCGcLPrYiwAOd0z9+tUasTGAmmdbgfLlqUl6cogXTGhsV06ULVxYhUHf1AAwpexE
2qiBtPFqJbZyvlT86+KesnEQTUR4+jpSmSg3crJ82V1pOyDDlFhp3av1TaT+VHaW2TyGQMfgltyS
u1xHoo32u7//mzeoZJu2AZoaWTwh1Jo4IUHibosv5KajSFXCpOXmD3w1x0+9F6LztI/0WLNJHTYe
m+dJpbfyPDvv70yXkU04QNM+MAi8WaEO471oUyG7VgmkpHPgtE6eZGRnXCldBuiSA2ij6F1zY7GQ
zN+aKZJGDhl7TqNB8n7fN5y7mCm2hozfbhr5VgJXQ/s7kORuGDUUeAvDoQcrig+1r/xp8Bo3r6DW
9c3o+MMYOK2uPaDNFfgR/zYoPcOz6p03op4MlX2mAIOXEUShZljbKydbnDZXbAg2FDQXybkj1LCr
XsqxrxBJvvf0EUvTaNxmiuRXAr14663BZyAywLDfokzUGPs3gCl7gmWL96dtQIVwqzClYWSseav8
belLthsIEVCwOitnVJua1oJy323KK28TetfW0v11P34ZVSGxUgiW+syJl/HE9z4JrKVyg88wtc56
vEemtNa4o2AwMmvlz/62M2J4DMWhWU0QGMQt6BJtzoFqsrfi3PnNiFDW8uANink5nsFiC+XYw+Jx
KATNB9dIilS16j46lJj9V4cEqOX+0NVnHZrdYqIFG79ym2r2H2H0J6fv5BAOFQGGruLUZgMLckWV
4G9l1NMrEMrZUyDMN+U+wjNctzirZ4Y9LQ1zKZ9/DjZbwx2QtPGbxZbQe7sSaAVD2bG1SfotNHBj
qSkXtdzNQjYLm6Z/QKUQKRQOXIubueF9Y9WPygCc5B8LzSAXv/O5GIj69dB+ypWbLcJavADNmMbC
AhwiiIn+BCMSSiwKCaw8+webEdQqAb3fP/7piiEW/FRe2Ux+pt3iVHF28LIYXfErLikSNbEqn5j7
vYaithoIwvqxRi+3eMU9CnAUxuT3ZaStH6geJpeOUN9w5vO5EkFkt0wM7mOnalfAIHIM3H1Cv237
UpjZsYjtPH1pDMukmweP2CLzG11q3VysCF6aj0odkw8FZZhERghTT1ZAPwXrqr6i/lxevIaU0ymO
Buwac9DusuGNEWdPsaGVAdA2S1QZKMP9jK+DPsv+TPvJPFWGTjqfSZ4tISWXT6K7vfeMWkZPscsI
UopbrNuFMdivhaQGJGYUDxGWpx7pE83sd7RKXr5+/gKobB2sPIyg0IwwIcpqMq9s5R8JoGhwwBTf
fcZF+JkglyJYYcorvGOtFyD6hIrPreBym9/qHZ1e76EmWS5HXjFlZYZvnOpyYaymspspHmXXATNU
4W0Pew6zWafQvwMr/h72l1xetDwTp6/Pu6QheFXMiPnvhNEwFqIfuJiARXRSwW2cENWWxuFEloK6
Z5zyC27M9IT87uXGU9RQ2B37kQ50L3FT6OBjLl6OePJH9IK2jf4IZ0vESCCXA/K8p/+YcmqVu58/
6FkitCDxoo6QBKtLgRIu+uEaVziCKUQZzGTo0rgWBBE8PGjkLQczO0d675k28U9GsXmHobqeVr8a
/mj2YhdReH9uF2kIDVwV/qi+d5jSm4sDDaNA7C2QQdRbGi96SbLfcGl8gvKTTKR7IecDcFO8Bzkj
AE1jNAsjww9g070CR2HmW3eZUthIV2derWQdNopqVSBcf2iZ2e16euRgovvqx101U28lHIhO/8/6
G4xLRpfUXbIowJWceNWfoc6TqFZnh7wYDmez4AUUEujqzzVSxqQyR4cOS2rosgHC5XkGEro4tLe9
Qno0j5Ie7MAPypA6Z+m7oj3S34l8IKXnGRWIFgZ7cYlU+TJ+fpGTc/ONcZrcLIwy0kLZJQM1gCzP
sxDVGP6FjKY2KgtOSH5rVvhGV3VE18d+D72M3LMzhlbdCgoqT3iuH38bOePtUE8ESYc+0Jb5Q4Yv
E/HsPtJl2LAt1xcEKGfkdl5o6bJV1Xn2L9d0Vxfin5JXFzNlIRnqupCPsIvGltfwfJAOQO5aIKzN
JGyxPWwdbJhD2g8Wulabrb0SQ+qzcpkwOSfE0rkGkXxTGi+Udv6QgjDLmBkPY020VfqDvuYGOHq+
99KJEcUH/E0OqA5MGxE13A9AbXjDvF+tv0G7GW8ePknj67kPGZ/gm1Qe5q4DGdSK6lZQ4tCg+DTE
dkHIHY03HfINdRSDrozTss4Z10asUpwzZ4AoYfdMBx5nEg5DsvYVSWS0MzdCwNkp+Mu6aOEWV3QZ
YSowcNgz7d/ECE37IHdwFOFI8g+qjRegb5hYPB1iUMoTYlkVB5RwM/GooKUPn/Cubj3qAG86nrxY
oDsBmwWm+uCHd3l9JumtpHgTTDydbr8wBS6v4+ABwnOpyf59eTZAVdN0PYkD6t5fz90E6KdDWpg3
P58rXEBYq+3jOnivlla2gPTwDIgkcfX1LhL/V4q0ISCtHGspMYfXlAD6oxq77BC9HEzk5OmUR/s5
z3OO7Th8QHsp1K2OYc25tQXjHE4dyX52BWswvU8mB9jEbwa6Rye6XT1lgvB6+ZYFbruqFlKi9LGo
eqT4Vqp4PYJ3WBB7EwbiKAv9RTd7YRxbekGrO5Oei7s5icunNEdJb5a3VE+2bBCbtKQ/grCxUW1V
KlYqnnkNtIDPLxgkoD+/JTxtAEF2Y9Ew03YJnb5mdzspvAEZh286U1N9I2b/rAP/qswNWtxB8VuY
EQISe7oB755hGHPy3RGINBgAfvmLBxXuHgPDA3SICW1+6OmAyQ/6Shr20BSVXG9sspW0FV2ycIJV
1XBJviuyvgGeHqX4Cginz6+sl8r5WFAszKtLmT+dQVaRGNhCtb/vx1hod7aw22WgFuNaLpAF4itv
1xzp5toRhp1ZdidgqZeOqgl6qC83UZL0Ooc4Ze4xbNVJyZ1C4y0Mkc5Ut85m4SoZNuljxGaK0SBj
F2/5Ej4nkNoVzbKF6GW4iZcTKLOYXomF0wVXrRp1oCue2ksU1T+XVS75PInHs8cQYFO6UvkrnNc3
xYmbUTE004vnVK+bdP+zjki9WQYphIhg6KwXLzh9YHquiejgTZW9p+sUx/NOORlCcefC5sJm8teZ
0CFCeDR2DA2IfAvlAR53pd1iXqm3v7COFdNfn+e9Ws3dOGbm9lXosADKvdUfLq/SvMjVOGWGkTlm
+2wZzduUZ+LlvjgiwJCYRYR2k88hwSgvbBSVVGnXgBLcg4+9Ui3C/fc3sD8bAuqb8aIWG7+6NtOb
auNsUWsa/fy2ZrOKD2hwX/v8AJvBxsJKh1Yf3YYLfyG8lZJry5PqsYq1Vs5gzxeHE/zZzt+hwDI6
Scojl3Dvm7pMBQ4FyW2LNESv+Ae8dNcJeYTxCYBrzLKGic5OBPwEScIIz3YO/orPe5bNnMc6vu4I
o5MvmD8//Zrskw4m5SdASS3Pteu5hj/Ro1JSOz4DKsRXnSsjBToeKRE/ppF2Z4O62luDv5DkqH7I
J++dCXXfx3MmuJqYEP+ywcNeWJnm5kXFiGlYyhVwKY51M4HSNFJjq1CtuswpVIqCAr2ZV7Xe7P0w
qRA2oQ6V8qEVJbs+kZR1eYwWWG07dtpnKkJe31ZSyR3l7IOSDpqCj/jMwYm0IFgKEa/Gh4Q3AA7K
eiQx9PgPn8FIWbd4NAZKvbKjjEATd4bL+wdb5V3pnuM6Y3BEwAVwhu88iseVgpoERCxVrKEUnwLV
OE2TFwWtVqGnlfCe16pt9h2a4+Cy/4ylkuPqHsThzup0hjkl6FYLxjLv7ElA/TB0hxu3zDmeZFvs
ChDdzrVQmaZm/jUjamE02Q9cO8Ud/o1BS0WN/nlFR8JoHvfcGp4gQDRG4YNHld8feDvYlf8AxLUr
Nvvpc2RmT1tVSZFDba9K0jUSc2JprvOL+AFsLrLTpPxR9VnRSlOl/v3fK1J/Nr8szZZXHGYs/AcD
34NUQHrcpqzUQZmR0lD/cFqDRvsxZKaWcKb2NbDPke9MLTRjllK+5zNuEqaEKUMgCG18LPciEm65
ZI7Ky+wY2txoTASHe4GS5o5byG5pVhSuGnR0oQCIf8xK18CPbMs7fbGiQtVUdSBCJyNPQrfemar4
T1CZTGkXC9i1e+7jmAkLlkM4TTPFdF0Qzy7vNyKf7XX5SWl2ZZ3eRvmDuGLwjFb+QMbhPyFe3YKA
b7Mh60g5EZS/FCeGMXuqNuAieHXNsk2Ct06fHD9w1cYE4W+YIgxa6h+jYy10MOyUeRIpo4sY8sVt
01ZLOyOSSAAIGXS7EFg4FaRZUJceCHa87yOJItFIxltGleFc813CGTgfiO/8ZzpQsAcVCVR/KAC0
bCFruxuss8sxjaTPCgv3CRPzr2oN79ABQYidbwkqCMruubsGn9QXmqcsaANO15NN6l+6CWUMnerk
rT2X9T/nVZxLNnrc7r/rC/7geXpHCuQgiJ3nt6BpiOFlkZnVCrfE819MBkjkfCSL4g8QQ4l1Xn1i
wp0vsLqwkCuc177s83HoNqOOQAoekx8XqOuU47K1IVqTuJkTtSwQmqvx5XvJbPq914Xj6ipmWl9w
WIEDFE7K1/Sm67oJQMCymgFhn8ev/kn0yxhep/cjLompIdOqBzG0B9Cm+wHnhwllelt0M9/6shMG
XWRqkU79OG6sKx2qZbAsFtV9ZGh/E7bKixRAxxWkEe45H64bmuR+7T5wmJIN67EgmIzC1FYtjf9q
hUyF2w4lHiyCaisG2jwxRSK7jO3veHkbJPFA8ZHUmpLtR8oL1vPnQVPlWFRHm44tihmEQBqVPdQI
nb57fz6hLJM8+B35Niv4z6wWqmEFb956J/zj9Fh53XFkoTyaRSr56qO9J/gwnhGUZaFXRpgJbw3B
QRX16clo9/IenCHo3FWzY/MVUjiS5Ll1BciufpDi9YBv7vu0q9WFor37J7uYKU3ZU12jVAd5SAwb
CR/bt8uqSR5LxffnBTTd0dOwxzSTTBhjeR9Han0t7hA2MebToYkG+xTDynlbDdfOYo/GNAW3O5zO
1t84QcSTqS6W4Mz+A3ZepVVUXx5JcKz72pkQQY4vjw+NeHlPETrHi+Q9B+d3vSt0YYWuWdh0AGCW
fgRtfkjXwrNX54bRD98A9QXM0Jf8tau3jRnjs5Wg2PRe4sT4ByuTLlGJUJlfkU+QVtp7iNBsJNm4
r1vztk9NXcb2a6tG3AighhPmmTM9HSDoBAkrY/YGlH+JANmcxDMU1JAygJh04sgO5Nc6if28tu8y
C1PWeF1LIZT4H4QHrFXoslxVHG/OgxBg4MwZE4C7V9IWxzhFX3TjpBSFm4+rRbATIyyKnArfvWAr
RRdvsCdST4bCN3GngS3zE1Fg2Dvr5TVFFs872BpDL0cLRFpwjCMjDXhlOfFdGIqdcbMmxMtu5mFV
iAoqX34UleK/BsIqbe0YPkKf/zQALPdWgj/bG2LI1z2jPtvSIYbhIhWhM8GpjOtqu5nrqO+EoKFV
SPvUL3p9558YzorKyAMA9xHPDE3DiVb5AZEZtbLyb4t7cbcqS4eK/FBqFJo4cHhM/tqB1jf12OmC
ZZNOsgApSQVmFt3jAftQo/09kLklCFNySCSWLCK3U6sn6kTjmsaOUincmctVrjAgU9x3deNELz1k
5mlZdSuDEgSUwyGxjihyJqML8i7CX5m7kC+UYt3ahdb4TXX5L9n8hMU81kWaSChhzrpTM5eiyjO+
n9MsaVBtrwiU11zLamGwpnqfr0GP8dVlYPhmyr8lo40I8fy/FhqqOOqJx6fUTB39ZSZXAAdSdgHn
h8C1YaMflqBlxY9A2a2H6+RJSFSxoQ1KNYFJJR3N7MK56Vu+OZlsS72n4AI7KbNpPTdS2lCFd4xw
X1GFFLq5JGDSW43qXDtbPYZll5IhVHmArzM1MGPFaqXIuDTL1LtYYbNGXxgsqPGfvAdH+5sRsbQU
m2bc6rdkSahd5VtVcCVb4DCfKA6QwlaAoK43XYMMfy9Bt52+bJgRVJjnyNFzhtkwROlMcnE+/uRW
usrgEKOEQhJBtHxBsnTR2el9R+Wr81cbX9lJi2PrWQWPmJl9tOLsdG6bbcVX1+18uGK7jNrYchpD
x01VAItKGpdW63+kYrW70NEgKChQy3Yk2gVtIm85recWd1hw+nzIFqoDyUUGXgRLyvaNHUoj748H
hLZKOhxpUM5cvU2fanZLga/h7VILlifMk6WV5lKvE6KrudbuU7uiOh9mJTsVZamYGTX68T7XDG3n
YITERuftu9aayb4mi5TPRj0zTvOaBWi2qSUj3gx10LYyGMVZZUara+lZfs4ICWLA0fWRbcpzXhHJ
c6LmCbABDIOhtNfuEkmLCsBrZAKX8Ykh46XTFTbRXvautaL0VHQj5LV7eXI6Zvf320R4ZQBnlysl
0deLMR30g762KEuSEvST9UdXqUk7wg8AJm70oVmVOvazk5PGURQw+VY+I+GYYDK7r3d/JW9kzBLa
oidopBBmNdC2VhP2g0oXThG7WYVqdlxpFaR2ynRNTab8MPY0Kn8REFo0DWAQkizFdUadKl6gKPqE
RxnILcjLL89rX3cNcPbFL4dym3/+1ehfN4RVnzB0YwVWA/fE9qaEC+aG2gLRpVb+NG+3XLgQT/EV
BPkhMaqYb/LiOTxXY+s4xMj+IQ+NS41DQf6bNlMrBMJ92h+4rS3o8vyAz8vVPkrsEbrRlrnqExVL
hd+xRX0ISNd/jJ8iLQFXaHRKoiBVdoUv0EvHcm86JmpS+mL0sWKoTqzyxZfpqMOUXPxitXXR7f2a
AUeh7hgLAMiCXCyYAr+PQxeOJV25iwAwxrt2XBPjtDyMqGF0fRZnLYZAHFF3bgxxT1x+p+t3kGWe
xMiqAQG6xc9b16WYmUweVVtTWj6GxBpqDgZSbJKNiwFzC2RVjbJHU7ce2+g0FuiGEZiVghYbf7mt
Aqu1iDEi/aKtVcQ9a/LN+KR9Ph+1RCe37XgGpVYkrNzJxkB9GDA1Xwz+CI9D6hBDaES+iGSuLRaT
3cJ6XukJigTvaPkr/pk6hw8Mk49A3ioPBAk1W9olHtuqUrcW1jb3etHER4lJ1WDCc/9W1BZ6egbV
Wi2HbHAhXGwtYQgEUG5pYG3DBQyotwGCadafhCB1kKk+eiyCjHj3aSOgQFdevSt1STXhqbO44CCE
Myj+NrlyOEn00Hi1IQv6MtDfsietTMSieqkh7el2+BhRhV6T60Qsxp+wfj4jwuEFvLEAlpw/Ubco
0eseEOTlQPtf9m912LqFj1trnptvIlhHxVnAAfeePQwVqIQ6yM+YWzwucPNMNv2UEsdvyPzlCG8L
jOfeNd6o+gwtqr3Dc8m3ttEgDQCTFDj9mvz/eq/I9SWbmxdsrHS181YZ/C10wc0TQtzDWlDXE6Jj
73RGCHLAxNDZKuS3vgukSZ7KyTWFhc7HJr3J0+Oku8ZpozteYQO2NsiXgz063HhiDl5CQJe8wCh7
cGvPCJJIt9PDKKOSBhj/3+Mgg2qxXNAMvqGFLrOD542udVi1enQ6OcgmIlwyptQfhop/XfXXGKKF
Dh6HbtQaWIn00b90xPLklwe3e08NX0jYW8mQR5SuS4zcf0uq3GUabFE8g4UboslPeuqGTwB64oCY
kxDISunr0CfZtv9AQLmqyXInV2SXIW6FjM7hFTnA4rhnQWJpiTpbK4APKoZT+PzgfN9hz89BUJYC
kXn/UHaUVE8gDw1fTlfSWPhUwkXvajygsE/YYoujvNWDu4CZzxvznmflpbokev1vv4A8rREQtNjP
96mXeOyTORvyzNOKKtfyf8c+05DR01lEHceK0Q/CMMzUG2NVKBf0ygsJnCqoRwHMUiURV7a4YMCM
laALMtsP2KdYap7KmKit4A50PjYM/1gVhQkbalOkwro0vNalGt/N5pMlvp2XKjsc+TNLLeLoxeOW
g6ZnaXypPhCxJi0IAv+EaswNiXevvxkHlq38dSsQ6tF7OI0gnADjaCJFHXK+Am3Rvzh5vryR5KsC
AnZDeuBbP7+JoZknF21w3wJ7a1m6Q5T7Rf4oRFjHqjyV6mByEFvhPdwVQzKRmc1QVJyb5oRklK7Y
g+Nz2wwxpHmcW4QRCXkhMDrj9jZn2Z/iq/Whpi2lEDdDO8lzp1eOk0YSO1vESOwt0EUCist0mdJD
o0S4NngLsO422442v+b6448R6dlCyVGql+YfIHyXn7mdOr1KnffBV7SVi9Hm8yLNTL32eVOHwMsb
bydhDm/zvRHJkfJ6iQAodjWpMj0kb9S2MCfyPZKbYkRXV5/e+hLYI1soBaP0tEpLECWiDKII3B/0
8gaXjRnCx3zgUJhHFGMUg9RpIu7iHAwZ8P0nGpkjyc10R+IRaXQzijyEx3PietJVNcqb23gwHOBT
oPlJFTSOynjhjw6tCnNBHyi092B65LY60ne3rpJ7nAXZTFSPChr4k6/sEwdGUfEj+8Z1qZpjvNxX
ZGOSiB+krhKuqDDTgX9SMsAyMeRkuQeBeGPVopi5JIo77hfH2NSTK1SZb9ArAlp5jCdKrZ9HK4zW
06IEuXlNnrbKqs1YnaSpg+TdwxIHuqzMOpvrc4KYCuMp77RDb1EIC/XQ2xQ0Q40qrWMRFe9uwt4v
F0wC2L9Shz7TzVLq0vaqxsI/nUDU2DXZLSSY8dOdAgZeNYWI1TcNfIZl+hz7MKSfl7AoAvRraJsJ
YNVYYKAhjpVCdf9UYiayww2MA5WZCz1zbl0ej8+MqKEulM8UcZGilKb9A76+Q5wmA41TJP62gZ5G
I0X2KZmuKDPnDsQqBUF/QoC2ImiOaasykzO6z41L5ztugZQccj5TTLoAPH8gDRApNX1FImp1Muhy
h7xv6vKFUus8X1C98nYm2/GJ1HGo3U85M4yjhFLU6cONnMkIvltixNwF2oGk6OE1sU+dXX9uTVk4
SoIZhYCnzWAmKX8h9/S6UKnqqY0AvOWXbXD3yoikNkBYq9EdHHjzUJZN1vh/3/R84aC8e+k8Yza7
twfZPxcke3tKf9+maB+OmyHvr0PIzKX5jeGu8RyXw84JaE/dgniU8za0GndLqrespOekZjXWtZ7N
AQ3ywJZNfJOyY/TrQFrSHRIg0pQO+DTY013oSYpnKwjd9RuU4hL5hChiGHHnnqESyEslFoi/2Z0w
+N8XrXI/X33UFgt6DSFCItJct2vrEOLCYWbhgCm5T6uP2v9Mu1bmbvBmSIRSGM6HdJVcKyLRzhyq
PlyRV/QOJagWoZQJ+trV6a69j7xt+YqvbR4zODP+GOQXYwM7nXrNn4RRkt/JfXXAyLkbkxiDhIJU
nMRCBhIa7oNujoPt7Bo+v7WuLKhN+u+3BYzuucj39hovUIvJgJT1xHwe3pwxmQsDf8QpTvZw4l7e
xoTTWZtITdGdSYvQa7iu2EJIgTijFe5Fh+ZMklDODR5A80yxi5UvzdqgALUoq53jQ4BLv3wn44L0
N98BMxnPJr3tBF0rd5wpZuaR5XmxCoAxo4ba2KGNE6gFS7P7YSy+NwWtKv9d1IqsW3JEcDhbcshy
Dmswc6Sxr6v6OifXN9+H8J2Xm7Y/1FroCkLW++Z/xbVH1o8W5HcvhVzLwCEgEfcP391ssHfNYD7R
VweXObdF2fUZ8x9T4jrULZ+74VRW10oq6vXFAeYevScM4uPjeWa9RJ7ylEsHwq6QGo+rtY8cWFes
v+qEh0w/5ncaTM1VJSqF9FVzcMb9ydhH9VLDTwsEV3K9XB7MeY+fmbU9ADEZmZ8XTOcrY7QQMAXN
PBWvLegnzkjDjqPkFZu2a6PHVAUXeOoZV9mrnEHPVr0BLsbFZfaFVciqU8EiFmQ6D/i1nnrnuNXt
2ffM3QdPVwCUvtf9Pz29VDNiIsigJuoo0/uYypYXpuwdmNNLDw2X8OwmnWyv1YrIHyKf6AXD0blk
Ox5yQwNxzT9Th87fOA+rx3HES4GyJNFz7/PqF7puRqzOrur15bLlAqJLVKKLLWy4aVl+4/44YvWS
haGJIrHh+zQPU65CFuqRvoOgyuoA/P4AQSBUrEMQjbjmT+TRNMWS210gp5G79S8GgHgj0tKs9DGM
O3TVfJ8rLKB5Xf9yrglITXrbKtpGerM1ZKoJx7NBpp2O5MbliP7HMSLhV6X2b4XuKi3mT+NpNq4P
VKNsWs9mv/Qma3cEqqwyzUIvle0RiEeNoedzfeuezP3KN6Td6eZ6HncMs2oJOnJZMefudNhgxZQN
QuADqvMQnrJGTx6XL52/PGnjqhdq3S6BwCzwhiWc+aIjzNuo/gASB8kGO6mMYz5xQPg+WQ6D3yNY
QhdThCXNzkAqKODVbaDE0b5r0subJ4gC/0thaISqUrFMxwW6EZjxCk+fCoDpuiRO+nD+UHyB7Mxm
DS6NirbwT4Pf4g6dSIg+gGTYrCske8oJqBOFPsqwL2SVEReK7Wd2eHzMARKErqKynMmOD3KQRxdA
6Oxjw9uBw+fcQKmRzzm9+4NvRvysadC8h+1Osym+PPFieke2HOsZXVPerCDONE9f4YK6M4ELDi8v
ISrVZChcY6zZFIOB47WegcMMlAXr7PYrrNdkRk7IMOOIkGU8gjawn4/Q8HiqkoxFwaKVWx1XQBFo
Q+doILjjQRT8c+QFUM4tElYIGETmu2GlwqcL7t/Rzw/KoPKaudn/2M5NEmwYruQ3DoPieVsnGujN
8xBC1G6IFYRmmOZLHVGb1NHj1pipO3oO8j8wenshukEqoRkaI5KRVd1T1Mq/stQFCdSc9mFvp/jI
MGaW4LGPO3p0zzfkW97SFA79O9RodJ1cr8EHBxXCVY6adcCiI+l8I5JcgOkn/kgRdTkARoercgW6
RYxI7JQlJ+p0Y4B38Zsx3JZkbXehDGBdvUYkSyN82Kfm/a29Xx2MT42iuJ8Q+dSkioU1LnssCYbz
Zoj8dm4rRL0OQWmpFDTTYq90jrd9PcnkYeQ/WYYRojw9sO5tsRCEwzl2EL8YzDJc+06L+NfV+ep1
T/amFqCJLLV+ga+Q3O+xxKF3IZMPVGWK0sal+X44b3/2owDMMcM7cOe0Czyz+ntOwaoqbso+5Qs8
+NPj99FvNXfsMt6a9PxrSJsX/zYcQX2W1DCNyQRhuEkExMw1DS93mLptnSqdsMJzene7pX8Kvh3J
Hq5yXwqGoV1SaZ3KWbp8GQaZxrR4DPwYS2PKbw52fU1EPsOMHnLGoCWm4Q3g8ZoJEw+kO0lI3Xo4
2QdkBu8E5OutaXbjSZ3bS6YH44xbQL7Bo9IA3lxdq+1HZUuP3Dq2dHm7lxEgyLulysJMuzfWFVtm
fAxV7BrPuxKGwDbs2LXNuy4VQA/M8AoRuC5lQ/MYIyaBMZ+K4h7ZXW1G48+y2Irgpghs73KGcXGz
AQ2CQWe5n6Tu4DZoy3pRoHnASYAZPfcYviHdGpJtslOhBYrUkyROgD6G7DyDGmaqvrNJFfMh6vvt
Rijnc14Q88FIBjMPQzqJXi+FVI6EZ1um0CIcQZnOeYB3j4cbhqT98TEaCBd+b7hrumn9ysqnNpZJ
uZO345mRltPga3KfgtnSylquJ1i2SeawSZIVcHKzuAoXhliHVD3UOGLSnWEU3Y54uJ/B175RrMue
KzObl5eGwyjaasoklLzn/NNlWYIToAeSYtIEar5l0CAI8Hh+IbZH8fGkUz+DQjh44kRNtuGFHBIA
N8gSFGMFsJOw9Tu5YqJ4Px7oyQfElNNtewfGKC87d2lWpfRTWqG0HJbcSlfTFjwKe90SDI/VMX2J
ehbKDp4/Ze5JW42gWVHwEjbaAX/TxKDOGy5y9dERsIXHD2SlW9S8Rs09osUUw8aT9cMrq9qOM0ox
cVayqiG/uwPYMNrErvz1SGiYXOGS4QIXM3ipEb+uS9wUdsDfUPkoGI5Uld9t+HBnGgj04JmgXTVC
8gToknLhgrfhSW7CRfckTpJ3+b4TKkANF6SPXDCCdGTD/y/NLhvan70s2MdTWN78w2xgt1Qhl9IO
5Hh6RRIU/DBOjigkzTpLmgQ5Za7GiR2AjM/wQGjQduCjhqxpelTgnXtslOyQziJWl2Pfd76+x2Pg
hPjhO82n0qwuMrRd6ngTfyIPzP4XqPli/kMKz8gpi8ippO85T+43f6p1h6UOyajPJNRRajsSuthS
EQqtj6kQK7SXhdsmV4fhZYUkOlX8wiUoDceo9i6AyTnEdnD5Y5FkQd88IfgjZd6svGouXr70B1Xi
QOHh95d/n7QZmN7f+aM4Yo4OvvmiB4bfvcW45Qi45VG7GE0DQ9wq10ORv4KqMlhiKnp2tDwg1kaB
FgihA0BxB7BcfGiYZV1wTJmmUf8GkTpYy/F+hxPqPJq4mjUYy51B8fBB1tgYfFnUIQuLKHMCtYyU
i90kWRUFMPCu/obKQVG8ceqQKRCGtBT02HTnWhDc09sPXv/dU9M/KJIhHI5QjBwmpdTG2IAylwp7
PQwGDV0iQPXk293HgXyyN4i2W/wat7ICfsOYm8to5JoJhPFbRa1Y3hmfVcLwOsSgJrhbpBGa36wc
+GETgPCbzraZj2kDyy9muoSq2XdPx8lIb5IwRLWX67g3b75HIeGBzLPVar6jsnARHXWov0Sx8bOk
xWzgcoEjB/0bbKghQKkCt+3NSm3SoQfKigIB7dAA8ag9+1VcqgZ6hDmDAfcBWRn99tjz0SFQiQsh
n4AaqIVMoIp9Hn7s5ohSKRfN5yBrMcro30wEYqf8yAHB7dW8IP+EnWG07mRnrQMgHQhEY5cocxum
5kYuRlIbMh0VJEvCCJP7pjYhytHAW0QpTcUvhzUubMbz0Dg465bjyesm7nZgcZVeZp3WYrjsRmI3
h+oaOX7QfexJei9zkl2C8rs86a15RHzH3rrCrO4nBLV9Ntzfrisl0WyFTCvJ2z9wjAjp/29sWlI1
8hHsy+iiYEsrTXIavgTxpxap1mhpm0h4JgbYWV9x/0WS09s/oanUxKIx8cUNg+8AAUeP5jNF3uJW
CNfyLigpqBDW6EipDBHjI97qLgDgZ1m+bQJeftTwAWJucWwcQm9TcF7S2TB6tMNguta0rp8lnt02
ro87J8Q7uRoEZt3niw+bKljV2EyN5J55S3rCyUHXdvy4CAiM/ZMeLvnUcIagA2lQ1QkwF6/jKIMp
8+om+YdgNlqhp0AurQNIPuWkiE8wPGpFWLawrgTVatAWvsExt04vKHLYA9n8f9kW7a147WCS+I/8
U+nRj+RLjvmqbJs1SJRfZq18tTcpE118E1kM6KFT3sphYyfxZNosYbf/A8N8kqM8cZ7YJJqiXvX8
WeQyqoEc2S3qVGvQqe2lJF0H6/bt3W5/2aKx6DjYakPNmcEvv/W5YlXCnhudmj6RqAl/P19BhAv+
/GZjJHADwObRSYkRfB9EeOOlHs7ZgJQRPnEsygnB+urT6f8tNnSJjde48e4G2pWmaYi6SCfp7+S9
iM0HNnW1lK4o6CQmBAX5m7Lb25Q88moWeaXE2dvaZj/Y6zvhUmDplLsSxNXxbnAD5EQ0YJO/lCVT
0Gs1fQTEIqfEXS8xPGabd+Qkqdkd0vPvQ4QboW5+yuwbLWyUY6Tx5OrBc6jQ1QgXPP8ua8Qm5xov
flzcrcDdPinNxfcEFDSO56z0ji80wlaiij/6g1dvKZgMZwpD3ZO65oi1hl+ZulfuPWrXVxf16fUN
SC56d1z4weuygiiP/SiEA0RqCT5bj06pdj9jEiHi0EbDVTUVenLmZHmtllyVc9a4Qq1PUbCKpIZz
4H7bdZLhXnELS8oLvpfhi5EzeMZ4+sZKH2shp6ulB50xg5rzYaB5kBoldjBQVvWBceP9Q1d7UTMa
OXwOXND48OIlpNFnlZ6HJsBjuIU8cg3glJ9CRHdBQKXGUI56HVeLsS6lwWcV7bok7XFoqSJhY995
hL7wpDSOnKqoFDWKNut3rCsVl70X9TtGJZss86+FpRa58M7r7HIdAVsa4yeRkO4hD/JmwHY70Bt1
5iYws889xecfiK2Ln7SkEbDlf24suDHzFeq/NEwEGsxFTL510aFZg1b25w5uv1YU6Qkir2kcd+Ca
OZBY4yejkt8UNt5t7bsZEfQkL1Juv8YrLT/YhRgI3jcSgPVYVLQGTPCVgTgZDNt2xzinHvc9dAZo
exCu7rWrY/ZCJBIkcCWKxG8jVdQVoXuTZsHk7akIn3DSpf1YMChIlaSfirExWvMG1oSqfiIpiZgJ
b3zEmLMGzA6vGnhn/sZ1J7OHoi7AVE4ZZOGCa6AUKunQYigqEYBc+uDsrq+1ZLr2wQoI7/MxxPTb
+srHxbWmGMceuhnrXAA2Bn7gph4T/PI8CWtCoSb+4i8cml9uYJl6hg24whkNRohNHoz4X/ZzaVL4
E/9nbsZpzLnzxC4wZts6vEsjfzhvgvVQAJS0unoa4KwWyWuFi/1X8QHrzzDnZ8NbqSoIh9zDaWT9
15wl5M0l8+3XL1+BDaMo7fJx92LRisjA0h7tLslY3MpGempouSVzDnhtc8fBXQqRCbiZgXgvQz4R
9MwSZRFD9s+DZBTNYLP5EeQmXJRJpTXiGP0BeR1+PMA49z3r5jlDER+TC2p8ewsoCqHAr2FAbQXX
dFg7pP9df4NyqGm0lYGTpXyEiLZWh8KW5v1oIDqs4wjJiIvNCDLu5CwB0Jwgp5YH54Ow+04/g+rG
2zq35rLKHfQ2AnzZ1SZPZEyd3KStRD5CGv0RQGn/GvybNRtdFjMVXyMkTxZaQbvzR+REjZkCQTKY
1h6XlHm6Q3mjvyTF21+JglrHQRfZ4U0VY1X164+G3jCtIDDxRTnX0D7TQo0FSyfaTmbTX0I3dgU+
vmYROYcnbIhFOt+YcH2aE6gecG8FspLH73JPRNQcO0BYFsOmlhXk3UD9B/YYnriE5TaKDtbivI7h
n1uyjrzeE8pHGuAhikyp0IQmJcyoGsTNOWf0RJf4DCx5LYEzw0f2SynHZxd/gi43js601MnDXdax
JxVTvP8XbTGJHpMClNbto3euivdIkrg74q1gwkG+qwZmsAzmSiDQtofCy0EtMLu2xhdGro0aCvB8
5o7SX4kC3g8Jaa4QLYyiBwiP6yB4YLBipAv+rsg7k9t9MOZkxlVdWEBWKmMTzPlMI/izMpwdyNLq
7uOYzjWmhh+v/pU4kf1ZmIk8lsRXnVr/vlwpUS3kkeWYA055p9w9z183ieDR98FkNa5BUkJ57Pj4
Hm7cdrQ9RXW9XDaWGFK3S95+GWR+cqr6b4Imf1gf8g8GXrlf1ywe/eRylxksM4mhC4UVe+6urP7V
0iG4uukUDOqqWhSsJKCxYxDws02FMQb9DC/EauVlhdyS6V8B9raW8iYQWSVuhmlWR0rSvlrGanBS
y/WO/X+zdY1ZkVLK1y2U16HP8qQJxSNsTqRaHbOFo7HtqQwlB4PRZ4EmTg+g0cegp2Da0DpbN85O
B7MS/cqKZYRaZqBJp2wFyaph42SVYu0nCW+dJFKdfMGtm8sn6YMccQBXCoJuSnNBSP7E5pooTFPs
F9jZUmFwRDtRebxK8myEybhOUC7xZYpEnQtKm4aJjDL27DPvRzBHlECTtoBZL31gs4/wv29yw5fW
zW7c3BeOTNiMQQJSGDTolYoTD5uJ79QpaJDnmhX1wbdmLtH9dPp5FfyZdAfr/28Ol9lCkgSi4BuU
EEFQKbOystU6TmTuqjXjNfWNwmJzmiJU1hmeBLxtj5dl9qnpTIbgFA5PImuh61Tf8ZJ7Jomdvrsh
BusRvW0GzEumi3E3Vlgo5YMXlj+fcsxgLRd5JA9Rnpm4YGS+4o+cLNfykpt+MINR0vKIKNqUd/wb
pdPEFzVatLtjzzKLXC17jYEka/SfNeyYI9avgU8mf9m2IkIQG4i6cZ61AsI+v9F8gCCgxuHUQmHv
sThhq0sZZsXOWrF5bBtDjDITNL0yShGDdRIQ2MFXj5gKKF9XrGJ0rnCxEflTAhcVM5TXUz8ELhb0
8VZifugqOPiCBWtTKechePH37/PhlJOMJRIMfb615j9wTInOzeWoMhiNSXckrMaa+oR6g0wb1PyM
6bDQ3AVeXPbwXE7TKyGmefDtS9kVqeUFGOI0y4soeBIziiFO8fstUG+pQrnV9JHMA7bV4+ImbBpo
BAsYh5xaEx9BYPpHhV+Bt2bWq4jaD+3T4nfGAHuXXkXB7rIA5TXAl9pHUFzCM1xkZ1zsPJ8TSwOx
5OGllx32EBkTdQbaIl5f/A2ccTEU+/eGc/b4iJP7KCLB2FXxUagQfESpuAqyPnAc3z/5vx+C7X0C
YoMF06LPMRKRzKCgwDAbS+qKCll0slPotINBtYEcyqBXi2c3w/tSHs6stlQ77NbbksMmCEjuFGHd
aF+tm6x7Mg6RUmd40mL23eawLK3CH+hyGKv9i+IUiwsNWOHjdEiWFiRud0DHCyoqIEaeL52cvRd4
m0PV9jIeq9SgDxGgxdcRQyxSRxo1r3xkzs8quGdKHrINJ0VJutyVgssrNsdhc6ZDOlszPDIJ2vdu
fbw+WcsN4/GtMj/kVvjbB5fYgCiPUaiseA+zxxpyUWkiSPepW3xrQ4LOgZcWepGaaQem+AUly0MP
Z6QPMDuW+Al+4YHUCUFIL3OJ+WoljsJLP/K32R2Cwi3tDH9/yEUSOe4e5PCRlVMKtPqx/8KIRuij
Rep5BXrW2I77kr67E1bJDvLZCD0lylbb557HrdouSkpPN6Ts0x0+4BaCRzizkmerTqdVBTOKGM9i
8gNh0UR0o6anZyYqBwdt5cmD8O3Jc5vrsBLFLrlkd+VXzZv1U5rBcPskkk6RNEI4V+cDb9tsreXN
GZ1cwbknJps+JkLlvi8zPoARgm9azgUl+w3GERvPpF6ZqUiFzZyzHSNIYUpYrYPOxUC2ah/EYC8K
4eKA1YsC/enjJ8nnJlfs4ZA5F3KEQFMYZECdqFuyaDmEEB4r7mtVqNC1StRbPvLE4SzMBBXWmoBl
Zs1vxFQgmY5A8/5ORExQnNYd9XIQiM4EUadW4ROyay8MlgD49Q+20Cx5Vym7cqSXPsoJOkhpQic7
Cml+SghwyieWWGPu8m5chZyliT+hoNTPqDKRS3TojZbUvEoT0gcz/9kwphoNZP/FyKDoLFClU7/2
b+vynO9qhYDakMIOYOCIZRGSyAU7GIvfeYgt9X6zH/V9TRzA0TE7aWlCUoCk9FpqnI/m0bXZgXPC
YTYcji1uYJXkk3r0ubER34dCeCf2dEzrWSZOjhvKCayD3pBm242CuNcOkGuB1hr5Y7Jd2QZeTfim
QI71ZEAEFAqHBxG14IXocBuFplTWrO/hn91q+IVXfhDMDlkk1XjI2l760w+1X37qkoCHbIasW8hP
dIDR3tw2uIgqwdY+L3I/dOCgiy8rm3kEUEJuOWd/FX9QLyDWOf0obs5gWHNqTL3mBLOngCQXCncs
eiPy51Ug8shk344UXT/q5RCLs+KCvSSOpIlFKaWaAO6PrH8uRi4l5H/RUfcijMzP4vuB8LIGUrWo
zyfBnk25vctzDTymiOjZgne+4l8J73XE8doS0vSZKK5TZgI/E51+IA5OpMsRx7DOOAx9oo8pBCeG
TzRS2dd/6UV+Mbv53e9EPrbgPZjnO7wGFnaWA+CCE9kAkVlQyCZed7eZYHkk5TQuH6s8J76KlBPb
xutyNccm8JyroYMR1buKKTJ2p2PZ9cnbnjpBw6qh6m3YWa4s2kGwRo647kRRTDMsDBUBd0kDIulf
HPdb0EYjnMj6UI33J8PVr332alIHmBdNjQlIPO379rZBCuXtJMdud/vxtoj7tzcFBE43fFhlcBn2
MA8bmFNR1t8P0dAzC0jh31cRyrpBhDezactjIRQL+stArvd3qCX8e2Z9fiFuHipRQcMz8cg9J2Pw
KHL2IKT9Rsd4rME8JVs8cP+O0gHZpv/wDOIuSsGvbfLZdHvJ2BU/kJ9+cmC1CSTvfwwzAcod2XMM
Ip/RTbmcip5JULVBe5qwcKTeoeS4YIO6J3LsGgzROMWgpGybLHjaQ3pmYdtVvR7t4w8ixm0LFGox
YRRz+rDHsJWJtgW23rky9IzSjpOhUXTzD4a18KaZv4wxIpANvxd9b+itqT3aqUvSXsk3QoXawS0I
5hnFlp39+bnDplSdbxtiHe2cwjUHCv/Gzx5S5yF3qdOBEQdE5LfMnlVOVRgP36jfuH9m0PDYei1y
O/uDnsEW2gcWHFeU0CuRAreTChPjJ3p/CYcvzf5ENtXaFGcWv2/rvlqtedRruj5eYlEOrZ31MUln
0I0ySgSvFpM+1j7Fl0e0OG6CBNdxP+2pDF3SwiKbr8Ng191hSyFyDQRxo2KY28VFjGN0jesvz2TL
avriaikTl0WcjwciRScP6ad8oSpdDmCo/sDC0E29E73b3RWm0i+ywwsCUIIcKESE8rDM/tLgxi1J
CdIOa8Kw+p6MtZHQNp7T2+fXnklAq8ju7xCn0XrlcV6YmRFcwckcOFfyp60DyIAJ3HXbF0H3SkYH
1EN2QzUOloUnKkxE82dQXGMu8qSmn8af+8IyUzOiQZOycg0GWj2n78ZezMJpMJCGYuzVXbTmZf7j
5stecG8sUSG2lZ3jxlcTSzrnL1mtzyZ8q7QfKZcFhZvwFPqzjFPeM/nmZGf1m8ZWdWzalbcD8/f5
qlFQMSOJPvvPFvUlgtQ6iIIm+J2l7FlpYumB96hR8sunIQLACI+eF44aR+MTdOeM+G+oZfpqkStv
oYuw+FnL3hXRpxDn1/x4DUkT8IG2Q/lZohOwpgcQ0DItMsi/0txek5ZXDbLn49035KplA5ecWfxU
xTG/WpgMyl8GXMnhY6RFvJmqgjsGo3luBCgesmcEfdciIbKmk448mE+S3t2gmWuoeYNi02lJC0Vr
XDfECfu6fFjhP1QQIijBkzwJR0JFsGmNDWKftkBNsh0nCY6Cw/zMFcGp30NQYSCUIISx3VZTYlOh
ZKmNjBzE2sR3xxd5+U+kQ8AVV9uWuwgjurkGopxDWZ6rAMq5AFFlNG4v6v3hqhyMGi2MyUasU4EV
qoMZEk9TTsFnscLVfXC+7E7O91li0oXbuMeQRNRTYg7Ggj8KQP9QeHtIwZqIF92G+bz7XoqfPYLn
h98p0FGGKfZ886VGBK844lsSu4fw/KHMP0mFF4CTd/p9FHX//rq74+YW8f/sJWwf+eWiewoYhBOp
rEI8YqrKuNao2GNKq5nwIi2rCQ7nFS00uNlApDzavcHWUIMuOn6KBjXhAIF9UdNi06Ubv4g3Ywa5
UdYGorVml0JwAdA2YVry05y2phKe55xCFi6nbQ6MtJ5/LbjK7m1d6BmrCMl0go4UB6ghevQAzbZQ
fzfUNA1WKhp1v4DEywt/noK/iW+IG81Q4Ky/UcW8W1O5qDbAC2fm7Hy2+rWdz79sfZIvaQ54kyns
KLKIyU4rBsxdly+UsX5TiPHs33XgZCpEU0BHuwu5y9Dg+mRitneY0HoA2l71Yo5yxHXhhJW4Nvw9
NDMCgl/hCAqIFJjzSdYpUFFpWaasN0J35nTCrVHbJsK+Tw7nNTj/60zAZuAxkQal+werrd/fUfeo
Mza7tKZqM3Dg2gHLqz8nZW0Rmiu+Y70MLlmsfkIn0a6pkqT/RaZoIDOxmYIxHezZr3mFYrEGf/ec
a0JY06OvnballqYs2GT3h6vEh8zvYsScnHH5Jt/IRVCpQQHedA9SCSW0dht9gtmXn+rD/TUrc77q
ZPLdhyJjnV6rZJ77CqAc1c3E7hYs8OdN84Ru/VR0DBKibUu/N2eQWmnOA0IoyK+O7wdFh/1LVW5O
etithfgaMIfXvzRo9SLMzBajZm8jkrkRlMiZddMUaThNifapDddpL5hXW1YyVA0uIUu7KfE2uucx
/8UTnH5jLo+Gr2vpscGEMexmpjxecKWaBkzVBwEx6v9xmvWGxBe+CaF+4wxshRe0Qg7OgadbZ77Q
6ripdOMvNJLop7kHHMS2PGWUEYfcPJjdvVzId3sd1aJmvD8ptg6O1Oor7KQV2qLVCmqk0mqkowRh
sayL3atCp/URy5OenB8C7oHLVc7xpwvnkceDHTgaSo1OT+vZoZyTcXlrX+aAsRsrZv1J0PNzXT66
KgHo4s9myj7LVgNPYLaaxoNpxj01nWBa4pzVhPlNV2T2WZAxi/khw3p93KtwFFWxgMvOntg73XmN
N+4qivh43F3zJaMiCBPS4EUxgCzgsS6yzH6zSdsiZmXOiqgNAKfTRQDEtAkOWpzhkdY+dkMNlJsn
sZk8fH/CH3kqe98HYYKxaSCQmfrbF26d6VSToc5hCtUeQTtiLFnXWClWC18kKnZ30xZ3NUqC1E0F
KB3ZhEO2YHb8Fuj+e11m5e21cCZFc7zvv0lfivsmLqVYb+6AUBfGtjmz9p92JffFISd3onDRVFB9
bw+0/Y7v7BVl+NgX0YnHP3xO1ExhdGnxdWLBT04VGrW7iATVLXSolwQgrJ2Jmi80jhzm72Z3egj8
r09RRwCWC1GO7xufm8q03Bx7ZoMm8HUG40ptDWVH8rJgFPn25LscR88hqG+DiJkkyv9eYgSY8Y0T
xzz+D4jddoQ23bJprFbj9S2JKxbNR6SynqjTWxoE+iAnTkKhIzLCkXGvekbebXMy+7Na9FGICqLd
5Zj5TzCnRVWh3A/FBfcSar3L/4nylckkpRUe9M4X6PmwKcN6pp30xLOBly+6y3fXM5UKteXw0hbJ
CFL94sh0z8wyzx9I9YNW4OPyusozI4kvJ+KVlUCaEEz4wUj8NT0iPoiwgosg+7Ixsuq/Vi7VJ/gE
w0xqOaM1+1nJkLuRAo4V717b2B2kF1zWNVJ0y+OosUhuvXaDzmTYnrrpaGZQ4HM3m9cgvCZL5XQu
mhHKzU9AziEzIJDRu31xFcmV9ytY2/UT7qtpotKqeKjBX3WZiPvQrB+GEJiiHg2amOAlB4dxC9m0
pp7tGmIcNZwKpLpyTQPiYqBqrvWIeALdQKNPTSriqTFCNyIY0iqXfhrPXYjGLnt+FUlqvIoA76FU
z9Aa4pFP1r2UuRS/16J3G4O4mUoPeQCt1MagcVmkBKS5qan7yK8fMcukOPdZY4mbx3fsn8l44WwU
40a88VJZnAjWqlczDtlqoTQ6NcjFC2FoxyBBcc+AQmMoYhdv1VkRA/Ry+mAgSOzeAij4vFs+bQW/
4avwTtmU/eh2WSlxzIzO2vShiaVj8t6b4PUGjjAzt/9sozUcgxnUNXXzpb0IYKojsyQQWgCA3ylT
y9iSRw7N0kw8xLaVgL+jArDP0aQCP0VEUEJeHCh/SkApr2DoTI3b6bBHSEOR48pq3uHcgjlkz2Hp
maTnhwnmo850YaIH4lZ4KyZOVCDQr5Bd1H3zMdDbb3JS1tQ7lbgkIoG10OcgsUedX/eLaxvjkRf0
KyCFGKtbytVLm7OoacdM3+2d9MhLlWRr5VY8x7B6sfi9nBnGnjvT/ivMy/Buq2SGqmU4Ti4Mbb9j
aXDmrXhZJ8zA9rOXgZ9+ZefrU0LysNdoWb1rXJH9IY1VbNlSYLP4wpjP34xrLL2G4KIqq3/Z5f7g
3sYD6W5XpsQlDGbvc5PCPakYNqbxda4+uMZ8xR/m22SpRcRt5PWqgS6tME4dEpK+p3C1n618XwSk
d73EXLWAxHKdoH3sNifmx6r4Nymr8eHW097fXO718g8p7xvdEnSn45LuLiscd7lQcsWXNm2qWUaK
mPzSRBe8/he61Cinu0loG/u3/s9e7FMMvXv2yEw+coKQ+80kEepUHnS8/ZJkhVIQqPcyBQ9SDvsJ
dvb9qdDhDTLBU1MLZtw8oQ88s+JAjzSfd9oxlTF6upvwz/TLfa4XAIFUn255stQQcanBNHoTEFJg
m0S9olahIdWVzPmdidcGZRHE30df269Einr8ON9TzxAVow9e26HfprPa2yK8tUy1lIuoD/O0uLel
SlcLSukYeI5giteD2vVgvTLt3jtSpgHcR+D89+RiqQ7YRNwoIt8Vka0iRUKvZ5XYM1urpNbsM2mC
r44Csv0/MyVlO7Oxbq2MTHik3SUwlwpKsTC6XzKpKyxs273QiNrqVZp1ujsdUdIQbuxm+Hy3q+GW
alp9mMHfvhmQg9r/kGp1JQt82nwDyYRqNgw9ix94NE6EBmUHSmDIKC1Fl4b94qxXAjNwJwR1xQQH
wzf2Yq9ry62fUckTPUfOmi6R3AL1NPJu3ntxvxemlHZF4sStkSdHxrfiXIeWjsCSgx06yJkasAVG
QstSRReOpL07HXICdFe1V979M0WV3lU0vaTpcmaEu24U8RJNpgWvwixgagdkBfqyT4F3gjkg4d97
ekjlRW3BEVbgvr/p/2wH6GG5MRc4RjP7/jaS22Fud3nk8rSqU5l64qkBFBX5Iw/ibvM9NEEyXAcQ
/DpuSrKyxV+ilZamGe1NqtbefeC6HLn7q8B1yBCi687vpHlhroPa0GfwVeGh41P74JNoYeUXx9cM
8W99G0Ri2DxVtl86CkdqQpia7UUQlEE5L+QPXqMunk3629h0pZnzIYqfKGtTlZvU899T+TojCp0j
LOD2lHfR097urEfVD6WZH4curBnL7/p8n26pQpmVT/pvfLDuhtR8iIK2TjakV0ATfIf/1Tw4Mmzk
CURyfKS43ZLSHH6fly09k3CZbt+BbwTYybMRQENzyyh6Hpv+yB+eq2kVCdWX0TQReMqcyjwqB1fX
RnPOzbHO/DiKdsUusdna9nd6452QlGnqnRAh8t5BMrybR7MyUN5+X/caoJQgu5doN0a7ch62f/Nv
1xac8ZhxFG5ev8mBNx3kcYbUYfsPxjvAMfn+luTvHR73/HPKgh2eke58IdNp9KUMnDri0tHHXEbq
zx3MMgAw24eKXMjwxODMYeylg30Kfjk/GZauXwAGlz29YxZ1It+5IKhtQ7YEebghQYNOxwyWKyyv
9UwdBAfBkbFA32vWmITJa1HDQDWuWMF5iISIdol9qZdyyAoLEsroLC3+oDnLTgOSe6DFA8mfGKdk
DJenKHoSfvlGJjhwcNPaoFbZSeggIs7k6jQR
`pragma protect end_protected


endmodule


   
