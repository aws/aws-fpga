`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2024.1"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2023_11", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
DFbDCxfDNaPu+qRK7QCZEyRz4q5R1Ckv3KnrNCFCMzVcaC2mC0wemx/2K6iGNXDz1RcWFQKkJrax
GP/QYLEMnu0tbjNU4nHcoHr6lSLXnW90ZeYpmOuznxEqH4nE5TRYyWRFUFRqTtdVedn306h4fTvz
Z3+yEokoN+oBJmYfzQ+rD898N5oiqc6dz43Bx1xtlXkRGsc4yb4/YnX2JgsGETi6HDPP85zrg6Rd
eXbjUEzwv//h+X33IB5i9yYewX/CjcFtEordRlPJcHiitiXnsSv4wSHyMEArhwPF7BM3WR7jA8rv
Wk6T3CCQG//3qsMjxy2RNSt1SFh6pWaS32/IXA==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
qrnjYUM/58hBbQ+CdMXfLkrAwyGUqLf7oA1SIrwuz1M0nAu7YCyFqnhGX9WzfPdO2hLskQMmBJeG
QV3B33NEfQexPfWp0CTZYZ+hyhaVML/OymT53Vcrn1mJUh8gjUQvpMWT2RowA+c9PDPv7rbFTemz
d+3KU87Skwsv95TmcaE=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
XhDbqNzKQvPIQ0QhlBUARnjul7hoo2mEJQgKjv3pshgmnjvV8hfHQcivW4PpAqki4E4v/H/mETdl
YKAskZ9hGn5VRPmWzPHWO+4YAt85J35O+uMGNSbG5mI6j0aHKy6Xx25O/oM9b0mwHg0pt3CRNWIE
vizA2WFxXuGcyXTeUxg=

`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
cr6oTGfvZyFvwk1d5AqKASZhSMeYtMp8o7CY9E39JbEXwAOvrCSX6wJLhqiV84Be8SZbSxSXQjnw
SXg2AQyZcw==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6304)
`pragma protect data_block
fSDXRUw4tLJwUgDStnaezJmdfsrsukLbnRosnvQqDABD817/HzU3XEb3q/GBb2E7Ok2B5Y6fscR8
AHWkVGX9ZP+LNIfXtSFr8W1q0im1IM0KeFEW2qBspV381c1hAQ3O964955uHqSNJPvq623gkf0j+
w6ehcMZm9Wen8npOxLaxEsajEfuBwUjn1g2C3KnCAgtnSzvbJcw6zDGiW3jnUQjjYBQi0XNjqcKh
iOqr29WwC7c6gqKBU3IXWlwF3kt0x8CRfSLaIzmDKpYtIU+6vVhZrqA8DYKU7dTtV+dSd3e8aC1l
IIQjUPAI9Mdaq39/4OYxCpEs27ueaLIRDqVVzPAo9cIcKC1pfFmlcrGSwjhZMZLoVKoA2fGJ8rnp
3iz1ERam1uwZormFATUS/kN/zmNCF5mrTm3hxn+rdAauERW67LegCGlJ7gw6Yb1Lq3CClcQUUKM5
mlOXM+btT4zNQ6Dp0qyoi2tuzk1llq6Q4JLnlGfE51lifeczXirlHPeCxFMn5+djuTPshbIVTu4e
RQRullTaOFl0FX+eDtYKYpb0DEPLqXBq70gFRJetGoK/SjCNFzmjZFTD2HYCFGQDe7+OknWbzinY
FNg/2TDjCErUhYr/Qdhu44MNZYdw5eQtl21j0filAIp5nhtbCoDwTfJm/o2JCs/He1URWtOJRRvC
lCdY4a+GCF4NVDfF7W0iEjzzk6YHqNXgUFK+ATb+tQiM6OVxtXFQaXQDRMU3JmRKWl8d8UfRGXAm
K8vgrn7sDUPUqh4lUPUJNLHOYYYoDglKIJfYc0SXtORad7F91Ou4ecSp1TEVyCg0u3olrCFhTo79
FGO54l14YE2vFEPScAO9poWPhtaHm2oYTy0DzeUg3a7xasbJIWw8ACcyYmCpPFcRtl3mFzrDG8OM
PqsvQUuhDuBiE/uk7b8m3VXpBS2EYIVx4XoqXS3GKcwQ7V4Ml3lO+9KhMgBHoDPUPFnpvhEEQf4M
RhGXADBbOIitJ8Cj9Rgyq9lle4EqHLAeBSHBK7ccs3fhoZHLkbPlDWiU5N8zxIb59tGNGC0PSmX7
RF6QjYtg2Oar6IJsfurgzSQnEOGr80PgR7+fB9vRXAFJ7ROe7EHVKQ8uFapVnrmkRihY93OLeCRp
7YoR032rioPJ4xT8XiCDI+kQqOPit0Ay8w+0iDvwJNLKpUTtqDivO2JSZR5MBXO30abqs9YHRI/j
q+kMI4jp+zDB55HCno5kKnW3p6FfiH8nQhUFyGhFHCs4GqWksAaQ02+WzOG4k7XM5xZvM07tgzdv
EcaiNr4Y+FNO7ctKN2xQemq2ydSQiaiHxnybJ2ljGmk2R1cDyhYWioBn3qJ5OjKY1l/OqAC+GVVA
1DkknV3h61FtnSltNKU/DWD+Q5ywvlou3Tdb/MNTWx8TU1ORmBEH+JIBN1ltHzgC9XlsLpCY21bI
EV7oHuFa3EcEYGxX/S93JEb5jdHn6Kb0xahDze6Ol3AKiz0k0P/cqGcBa6AQmU4vjKpx9PpQGOqA
+eEMTtM4Bu2gn5MbPajVO57jMIc8fJ/y0rMADIzu7HYBFfq1jHzp21REfe+nM1+WaF2OewlM4KAh
77yKTZslB9a9JJyM09i0yKP7tZzh/mJ8k3Xg8Sy35hgQRVKzjgzKTKhTJo7jPZ86X+hVT37i6Z9J
pDjI5aAM+o4L59Qh6xR76fapDk1J049bEge8ZsqroH/KLP0Msmv8M/ImScvmkVo7aRLo4c6yx+Lk
tJHYcaCcgrp3J3hwomM1iBDggSgqFjYhjPxbhwc1QMYUfa1tft82HxGtHONWnnjWzyISzvJ9gvjO
GoK/XAPUQxlyEb6fXVhRgxK6oriehBCg2PwwuZlwxVd55rNd2E6VjcjYZT2Tquj+ZU+F/PEKwCfG
xO3zzyYpYLJ4k9ycIz5xfyYu2Onw0VfJvq89Jg/Cba0hAzvvduvIIhkdDzD5mdiFghGCYj5/rwMt
2RAEAeKLuNFhrO9H0fhQfxtJqEY3IvA/HRrpjm7kgdmuSSrYwjTq2pMXKsGMwdn5LumBiQrnprDl
JNvU4IfQqJMtO2ZK/xcJoc3ZEaIOSV/GG7r/zIrxycHu4JRHt0D8AZY/6Cgz1ewmmYoYGipBtKbI
cFA1SZDnZHKD5ou+MjI7e11ZrZfGy4i5od3ANQwbrv6XcIyw0/4mV+KY+Pm+LfPNhljx+0+C1Bh1
BQlRU6yA9Q0lvtJEYfLGYFKkCW8G8BX46UGqq6wX/tOIKBMe6oHBx2sEp12UcgyPkPAQMoOBbx8T
rRIdLM+cCNa0JeQDJH9yuapOj2kCFAzmHEtFDQYz2b0tZYru+lEgDAsURqXnOsJ2Kkh8/W2dYi0v
Ydwk8lWgQF2sPFBEGK4kc3pfvhOTMXhvECustFhR/to+KBWzsm2Cuq/E4OvVM/VH9Ckc68K5Y3ij
Bb4LTcfblXUjuPe/mE7Iey2lKTDcNwEIDqMj69bgEFg5IrbIotOFqXXsEUgEmUwENKpha4alegHp
bYIMRMVUEwhBDEW4P03UA85ZM8O2VWULy0nFKzhzWhuIh4E587lYfge9phRo4itO5Yl7TURsBWf7
mBbdkxOJW4VO8ONgFcwh3OS0Q6+No4TxBkFnd6JuhcPnumcOS+OXZLlu7q2tDcp02NlXyteMJvFn
lHRRvgr8s4ZxI3xKytIw6EnH486lHExP4tJaZo0EyJqkq7pyAEuuuuS1FOqGatprQjnQ+kRuECa+
0PQ/IfaP/wmSm8uv5rpWeQkpiX97gbCdf7GeAXg+71yxN+QxMO0MLq4IRLx/qU0JQntuGozjWgJS
xXtdlA3+tfYA3eVsXsnVLKKxYEr62Hjv7fZScrg4BYAxfrabANuGzkqD7IAfsC7oPdpS/GRMqkJe
w4umxe8l6pxBAvs4S4mOCDjOEeGpBmGXSOWd9jZFptr6CLtR8mdHxmk97tBnxfZMKXkx79bxl2c0
9hvPjkupMun5LL4fwgn8mayhJpzXzxHp9PsUIqo99fDcqfsdjv1k5+0WWIe2Jh3AdJJY75L6+egz
N7V6DaImQmsyK6BvKOkPzevGX4PlN3nD9+6cUZWDSaHnArd59SJfLna6EemrCtNqpHnp+7qJjUQf
TJz6huQ9/pkYR/48E/5JnO2l2/nO29kbjQxsRiHFQLv60x573pFkrK07LBWLiHGePvcgnXHOteTP
2XwazHLGExv17hFCWcZePJkVZAhiiRJgjJ0fTfJL5tDe19octV13J/ESD6JM8JCjMhpZ871ddtfv
94zyKQC0B31qg8AZ5nRT1epzdPxGA0qEEhZG8N5qE2mT0bnFOhllcc4kRSpomOfCvOX0z3yJUB8G
4SzMoo65FgP8lIL40KxPuQK21oNT4FYBXfJl388cYdUW0K5h3v64aWx3mPtk2sjYKuDPjjX7DSnz
lTC5cYEOdoRu3jwHCfflF9z9/m2rMmzy0Ppq9V7AGxo45Q6frCCWWhNaZa3c9uIRBWhRdBQOkJAr
y83F9ZyOi52Kg/a4+TlMV85OauAD/35rVgIS2cFSo/hCtAET76L3sbqt9xdWNLp9M72TNNvMueQU
ttQo50i2YKuf6HZhaPUZWknhRRKIi6z+RDgdpoPHY3YNiMg7DkIR+SNHUCuHAWFkdi/TPqUGN75x
MB11X0KnapcYVV/w3aKCEfCp0mZRzjLVp3IplkVhI/SjLbinQGSvO9q5ELD907sCTHNto/zP9DHa
OzC5eyTe59OO+ogvbVkY/4M5pfDnVJgS9gWVTQMi87N2UMx95DzH7ZIlJfNIWs8A3uTKzF89Q1nm
4D3gShflUrSYO3o+yeh7iNDGb13ced2uW72VjhbPID2koeJ7/WJQnVt3ppChT2NvCVMg5mRFFJ8D
A9cP1qjD4bfxII64lbjHmtPE4czYhxr8MqDNpELBbvRDBKRFCKgTIIMNFCnwLFk7vj9XTb5RUak6
3+Z88tYyTlJ0amNXjFLwwCx43cXNAW3OFSdPFP8ujQUfQ2hQDm9/KB8km3p0Y+KvOKlaoRXj6kgL
GFubc1moHU1m7omD5UxDbk8KPAYMr5TeZx8qOCmBVlF1+aHE5KdgpSo0qGVCdgXJ9aIeBgXpUGmg
gBg7WkBI3iE3lftNknqcgkcYCM8UAlpwmFF2g33u6odIOIxvaoOqoAo1ZMH3c0M+MUMKLszwfemK
HugUT07kwK5E7FSUW0TakI2hc2wu4MWiiH/mx+l35Lijqnmpmhsal3qHtksaw0PcPnnN+FQHSSBq
7yNKXTVz7gbOmmXsJQ0MNkOwLAIwTBP405XSxcSp92ZQ01KzxZ04b5o6wbBHR20T/hv9z7mp2J/p
7q0SVgMCpM7AEbQI/ndAFhMW9w24GB8wCbOU012ks6ZEEINMwJ8JAQTisI5oudDVINRd/WMmoF9o
S8iA6PQOBWaN/fCYVjqhDMi1HECtfMUtVGHRSUxTXM17X/9JhkzUvpButKNG+V97IjJLvc0L/cFk
YyAhs3OMHJP3w7dFItHI8+iZ0iOV+wkcqNzNU/KfY0VvGlZJRpxlgSCKyupygTguj7hDcsQzgeRV
eFtSBJul//JjnH+QHuamE+PRyB07m+wwSfzcrT/CNkvbnRpt1qgfBHuAhsdeOLxv/fdNuuu/FFI+
1iWLWor2ZjcKor99yKw9mZXOct5+lzwxCQo5korCpA+CdEu8UPoV5E0HUisBcBTzA5hhZE6wl4DI
8CzD7XnbgKZccJjAzPFnrPsuCW/byiVXngB1Y+v3kFwpFB8BUGC6FaaZtkzdEmYI5WxwtTcoXw6K
YAeSml3pXMROn4RVwSas6SeAKAhyxB+IbCSDHkpsJDXyM8FIyd0svB4uAWYzBirK/g465fg2EP5k
rSmDEnaKe9RoJ68EX2Y0OrU+3/XpTJGSWjECLi8NoqAtPe8i4TiUJCRCnOpNtBXa1AvFuN1L8a48
cfCUZp3TtjaSeh3ptiGKJSUJQyZCpB+YOE3162X4IPtsx7Jn0nTkWTbUo19B4eVbdR1zp1CYE+xp
Eu4ZsS7ATDrNPFJ9+YbYGdHx0NsvW2+SKE5KKEbqsrGUIFOLqdKdTxWAYvn37jA+9IkeTyKH51V7
E/xo0e7JRCWlEyFOZc959TnfF8qzdEdgh1EDqJg3q/YhOha0A3IJO1ClBSCy8CmnSW9a7AaBza/r
5tZ+vBVard7U6ffscsRYg17aAEcbfhhSsVb5QWU5x4cauQbVgR0IkIkEE/WstB7SK827fXyNn8fV
MP1hIWhTTvLccgFOMaDLre8n9W542D9LTPpG1D3Zi0EugSJOqE8ufL2l1/Z2XBgoBXJEuJJiqW9W
uZ2dQWJE/k5+bwU9WRlWO99JC8zU+T6hnNy+b1L3oY5fv1MaS4OMtgkDH9NwH3efZxEwqQDPohMm
o3a8GFo1CMFNN/LezcNeoaZKJHSySm+D2Id+l6mNpIBbSCt8SKiS7lagqnlysYqc/PMPMbhy6U/B
/g0UDyYgh5VjfYEl3/qKjTACz4qgL+PcRra3sHSvOPkBr+f8DDd6/2y6/mMFXF3HntS04a3PfsVu
b7gFlPJPDIWm2l0MDUDqeSOlv9YqFDgMXdckq2IppcDYhMyNjm5NsKKlfJxQqaIEDVM/kn8zjcZ9
+Adr4Bn3+KAwZo2TMZpkyPne6m559ZxKqeqJW4eGnbI2CSU0ik3DIBNJBc00l/YFsMklubw2jWe1
QdubGLFDFoEoFNz2pN/y2X7LpotqS2HDOgFNf73awkza7AmkGwiXrh39dtrBXUh7mu1RRNHxLyxn
U1ZleNoHrsWZCKJFnNJ/4KND/47zM7FHzLds0kr5Z7/eFsu+deIfF73RWymlwulFGMx8ggX3ozuG
CkMz/1Pm2ePRYBrKdM8km7AeUAwufMgci2HNWyEuQdWKSX+bMNBrPT/u637h/n/SBAnrGDXtk7t5
9t1q6g9H9V9lm+vP9MqGBG6L92KpHtpi4f4bY2vc1jMcg+CVhC/Wcxrr+/TD+9eaUjSjatSPrxOY
gRbQWOZ0CFs76y/duTLoWvhWlzXzuY44CWRVbBXiMBtLjtmMbBl10/UgFSz3ZMP1XKTekgGvOmC2
962KOydkp2GKqmTHRPVtRvUIjj7IEO3kIntO91WbDa8PVMr1pjXozS014aUdEJW5Cft8lYDua29z
HxGv4XW3yC5lt3eN0w21S+wKFUXs0p2nW2RRcWuiAWLOPDkm7qTbrwYbTEgf73Y45PLtp3fWdgBx
BDKabVmNcHLMj6An0B12tsaciOhQYt5W/+JgiH8Kpir2kwD3q5V70DNyxCgwimF1RBQXyVxSTXH0
tuVqPkJbikuNXD4PCqaRc54m2kZT7ST3v9wGZid/k74oNok8Nj1E0qRG5U+ssWisZc9ntYH8CnA7
wRfniu5yfYAZEja4LfRjBnid/GYtWASgMRJZ+b/ZmCfc5bDOD6qjgTGUw3QYyZL6MUztQRN24HS5
29eNNlmAGAkHvfDU+AnB6ByUrnBTrJD9BxaRaN+klY0u595/bi5cl8fBgTypv52zwZ1onWVAKOvv
RG/kump3xfvpD8IZj4v54ZJo8EBJTV3+V9wxBKnKhJdaar6CGzeQbhiK/cav2ltxW4VUTGfzBlvk
swHfn73CyAQ3pV7bURSGY1Ba1AWY4AOUHFYS//AGairw/jgS4mmRf3fr5imK2nAYqb9JKpAK+/4w
uk68l47F8lkzVQW3hVGLtcFkbe/v5GTiLiCI13MYU5pJiVHikjrMJCEXQ+1SXCXQlwrk0SO1NfZX
sSMBW7n4ttigsni+zHwSGGAvWvQjH9auZbezF+l3SjjV4u2abd6f/LEvQsFL/2X5dKrRqVsyXVw3
y/C4fakxud5gXzmVTnKdrHmv/Mu4EAMj8e9jEpH+gtCBAiqvynHXyLJDttEfd4Zct9iXVr2zho6J
BDG60OFwRCtvnsZY6LZN6UxkVSJDsScjVZuGqCo/4OgCU+aubvWQaeI1XC+6IzOPzSRZGRHwl5Qa
AgDBDCrxE7Rdfh8hIftYci1msppahGgMUu8o9lH6EvdjwD1ceKcgwSEW0S84dP70HIhy96ekBvl+
LJ4gl9CcA5eixy7Ih0evH9Zf4nkspAFUIHM3kfJkgDbvaomZuX8meTtA9DzHFqeEM8Ms3OqFPYAd
JQR0fRt9V2BEGarlZtX9DFuXa2Oops6W1uiAEqqPZY8gW4mFzpZVQv3SSWAxEf8ncYS/yx7KNw1T
/k6i2J9vhVXsum6rcnjc1dl0um9MyzfW0L/Zxy3kBSQTVO6y6M/iF4MmzWPayPbG0ijWZZd2IhmM
2wBMklEKx+8Z6D7v8fQf1Wu1RlTnUuP5+9e/elIZUh5zU/g9nEygS/uze1yd+jIpANrE+YDLWLEv
3fNEnRnU/MAD0JduTvha6fWE8KRAYyTUoZYJwrqECIaMJg7IGppaHmriiTHiT3Z6MTmGTrP9ctbN
SLCNkjyZaXD0LnXB9Cicr+ESnbwoTx8Vm/G30xWYzBx3Nw9xnZbVWdLN7s/2a9T9kERVeObvh7d+
xGglUvaoDO++QHBG9upb7MFgUdPY9iyUTpgsuA/S37tIS3nq42bweG5slfKumYVoG8h76BGoqzvC
yWLYFfWQsn6Q8oMXcDvr34/kilqAENP1lnB24uubnuUoVJ1C8t0mJOvmCkQyus6X9pr8yFs0E4y7
QwjtRCJ1cFXNLYM6zPto5bWOt0bWtR/knWpFWRsfpUdryRrLugsYJmV82S4dBQo9gPDQpdZGZ+9x
8Uh+lIcZwXe/1hJK5YEF1dV6kA22KOQ1BB/0sqi2/DJVQcBwOIvA/pLwiD1igFDhIa6RXZwc5ShS
mZmIxEnFePvK9jiU5slitdGxPF5h7Y+pFrxc/nHmXqe3yDIjBjsx/s+CH+64QufCz1LDQWMea4mt
PG24hTwvQZLp78kapEDuCRiIp1uybwSxBtJMcY+51gVfQM5AFYUVrUxcSL5GHlCqk90YgScmYogd
04yv8zXp91913A/yT0okqJsag+9/0Dg8/oiyCwmKPdUDOqG1F4Kph2Usk6Q2DNXx+/xbZoF9IIHY
krstO+tMy0LskclpLaOnaajVd4GDehvfbRFSSk5yW4ZvLdJA0W0KmnD0PvbGN4HU2Do/GAYVjReO
C/RamUtuTz69gLykR0NL0k+aK/BHuT4eUCewcW2TH2mI/Bn3MNNxuq0eLexs1jCEul9/6X6znKr1
ScYnDYPTevyZXRZxXj0ssmToRVvg7fQ/BDw9p0cadX1ABE0wcscqxcfe26NEwEyU4uQP6k0HJdy0
9LepzjowL9QvU4+8Jb6pcDJeg2LilcFMfDTZq9CBTRVP5dEET6ybotDOmZVgXUpwYIxgcGYTicKq
0uxwnmEJ/Mfx7ajG+mF0KUDWdUIryK46yqmKrKtVaQAfkA==
`pragma protect end_protected
