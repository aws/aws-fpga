`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2024.1"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2023_11", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
AqabqDQIRfbU9cV8k7KKMpKHGzJRRsQcWGyFDVUtzYLUNvq0pEscsry4SrsVmHuJcFDbr1PZdaq0
8Rav4erIUVcIM+9dDr838E++mmOA8FxQUGy1iuWA7ZXm0d46mcI0+Y/Z47ca793bflz+hn0Rpxmf
TCanVwykJwbaL+ppMfHmeOrGvWlze/SMKWhxCnk/Cwf67fDS9vWniREq+rnhU4pSutZ91CyHjVi3
m04kTQ68Op9bPbEg+DbmN3ZBUB1yRJMr02OIC4/PaIoRZpUlde34P5mfiZ37nz5UQak7EWzdPkei
DuvEEHDdCB0ecBTH316tHq7Qp8bF7CGJJFF4Gg==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
g5BWwR90GTVv2amvMFTb8oS4p4LtlNvnq9HivRrD12Jiw54dpITRG/8p/alYWAgHscdAEWAbLwq+
bZuwdo57qzsf4iM4QQ5N5zUqWsaXmkt3F9ekxF+3E8kjjOJQeqqMs5F67NG4YXbwjFT0JKyY+Lsz
QcyfdoBUtd812MsWKWw=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
AcAD3AhtRsXAsCXlRemBCC4YS6N4/ImGhFYGz+4YGmNFRlJrBGwUAcoAw6gyL4aYipTVzs5ldMFr
Lja0raKIlKfOgUWX6ShLEutZZ5MEaRxbhM+mWnXs3AN16M0pHIm5pVzmF12D0BpZ9XCAgVsqqQGm
DtmCfhtZyimW0NCnShM=

`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
Ncm0wIzBR4rRAGfWky8UPv+QRedF0wcosXTVY10OcjjOp98FLbPEX0nYR1Eyy/uIip1n9d1sa0m7
Ux0HhtYIUw==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3584)
`pragma protect data_block
SogxMtZqwlEks7iIcPnavog51I0LUTbXgylwBsa/YNaV8aZR/qp/KveBz3EHso5re3B7UeimpYNf
GH8VUi8tRumqtmdsotKlnwgscuNw05k0rcBRlFsEKi8L+4vRCLv/iNMGCI0Nau9T3CksGlS79q1y
8AYYnkPvCbXSO4G/M36ayWYTKANnRhwh2FJng2NLiL2rqUALS22tj65EMm2dP3uTEW07IcysQ88g
wuMhmoV0KYnnWmYRqhbrDkB1v4cTcC/G3u1VMAaEbmqVZR2DmuWU/vmduPENV3GeA5kX0fwhjNwo
CDtbCiljsw+yhnADrf78fkB6aaELXsfHu85Vk6HJDDmnzUh/lyoiVNsXfxHdpamVcV/bgVNqHuc0
1dgD80Z1tXrYc02DPWCADsHSVrCsW/lzRziSUGh1ROBfmz3lqrpjjLPg4h/dXZ0i8NKWSAKU8CUl
9z0fNFEnhYNSD7fotou7JeVm60o2CZ3YTs3H2SzbKUE2Sht4bx1Ob78o/tpP1hqMEPfY8bPjfhYN
yqieG+Vt+iXVJUetmczNzMTqXUKKScqvpr2B0iJL9dU8jSq0PtL1AGFyew991fcvvJcwkaw9Y0bF
VMtyZm9EO2u9OaJYjZUhzY2L3yB8EKtz/lR+gBG2n1U7f28JmsepZKDsb3031QzjinXHUvgFkmZd
wE8WoW+Xs3EmkzMV0M3k5UtAlfqSzdWK0LMkSJXuTVHmOykTOcDQ0JZrnjdxkYUL729xuxmlEPyt
RmD0N/li6H+AMnnPRfxqxCkug0L5yOfrXMpT06xd2KWFqJ9RQOduw/IbWNGCjCAT2+mNVZLzOG/K
xA5USiUtIzA0L1Q6G1LnO3n86sbJ2Wp6KqWcN0jYY13xUnl6Vk8MBGeSkScw6J20MxN5CnnYRmqw
T8fpD4+/LikhDrVxTEAmaDclRh9aEI7+kjICdycai40NHyGkMSCaCEcOKII+bXc9wl5+5NHcc6Z+
Og8EfWOsoUMculXweXtEFntRQkU0BlxKvHXNyYg/nukTJuZmw+8GAf+eCouBrLneFiUlEOfQLTiH
KzrpJyty9anVc/TK+3T6MByWuZglI+0vRdhyn09i/0zSLC9nA/ldvML5pmAftZO/AHCqsb6wPuCf
iV6xT4l1s37f/tfUwp5RNFSvy+GmDyoXHaiNvd9y1RMONvJA1TqyDwdxDuJCSfRR5/qCziLeFEa3
RlT9auPxQFRtFP9aGa7MvLRgD1erGPPW4rtpEhVwVAhmcgdxPg3VGVfliDzQqJnUAvFNmwei7VMd
h7vom6fL9/WW0aiDdRP+EqpHj0rMiCxr/6VKhSjheIlTZzwSXig4ZriBMeXKjKdCto3B+dI3BPy9
fNGsE8svxZruce3N5z00M/ne0N/X1vKkQIOx8lUsHjK+aGzKSgR2O1ldpo9y8d4rU97llOod7S5Z
8ym9UI1FZoekxTbbG/mHMGjEh6pkKqxGrcj5zZg9CLhGIhGCS31klkGCKNiJwPIqiSgiZLcGVSJX
qHgtox8ajFV2Fa20aWMqbwv6ZT0hGxy5A7x72OVdLY7nnDe+Z5NcmqBgYO5Je3l25Sun2i4ZTMLp
ihSSVIIJvXtUN2Kc/bWboT3YVhhd9i9iYWNNH2UvSDRqyO+jnFbAUTBHizO0rW3NF+KwZos4hSek
kXcvkW6D7RZ5aMAXwgb5/UVG/kJgsIlU6by3bxK9GUUqjZb0X8yyptHkP3nwGhpaGGWf/KkUVjh+
IMtD0lJ2wmqE6+WaRXC8HruaCM5HaKKGnzf0Tsr+m0mCJw4Fcwj/xA5IM5WrgMr7Tp5XYw/7REOq
0eb5ICNoFOHd4aLT4DBECwEIyhWm1f9pdYHzbsIRYJERMUfy//ZJFld7F5iHLFFfV03vd0cVTa5i
fHYLLtv5QH5YYpFTicQ1xNxjkHgSIIP4V/UuBuH4nlvIt99VjAgNAxf/bY8ceUBlEFb0X2sZc4YP
+v4Vj0utwoS0mg7NNPi5SJQcURmV+KbzwYhnh0+DB17G9RIZoJeSlD+avZrs6gml9p/xEeaXOj4w
hnUlpuBDWx+foGw+W0HvmKtMoa0RFx6B4eIpWeHuo0kn/v+KeH4hbNyRwouIE2EYOrelmCuQJ+dg
sWJivqBC+LhXOXucOUZhTWur8p6dL1SpeE2fzpfUg4rGmJgyFRES6CsSUTJVjl848WQcgEDYeXhp
6U6gNP63Drc4aXph7KV2KcEnWcxDRuDtCmW3BkMuFIB0JnhbIhZBDLFCRdBXxKxk/SNXuQbn7DFr
aum6Ct7Q150vIzeejIXk5+ZqxadapDfZI//UYLkCH69z/1nTj/iO73CXjCozIPDpi3ZRooL+N/e9
ZuuiHy7AeTRfOReVplsqS827mGOxOH78Oq5G6k/14ffGPewtWNnsuXPHzQf4T/7HEvMsrjQlzkde
/V3afYB26yc3GI8HkD6UsRXI4E7679jFCpaI/LLFA9AFpAclLdQkSmUqIbHjP1w9CkVx9ES+kcmr
s32rwW/WLiQV+t918hUMr75kWHxZKAEDtyz4JYB+VbeKlrg8XZ7089O800nZMPWGsRhx9w2TxZCO
roSesc5OsSvyDDM5yHxxM7Cl4dSCSekC9PZww1TG9cgOvqlI01MDfLYcTQi8Ci7rLOTLJ6aqbigE
8xgOR748jD6Y0ufOmycVdPu+kwy/CntFNWmYyjJ+C24hrKVqS7zkbaLN6Ltq6ZfGGGooRKcM8OFV
fQ6CADITONGtUib/i8EGJVlbCPvPEzeivvHaZZ7rjZn4X3Egs2N0cWoYP4zmTNonA6mz0YTCK0AG
CactynVqfjrwbRMbiYOPYlC36Z16tZijWHTjOGwJo7ORVTt/cSxNC6/zADG6EH5rOxqwkH6r2Ovv
rvCQJQleoIWr71jqkx0zKCzPMLdNLv5rylc8OjmtgmfQ3f3JZgfxNBtyMyKE3XPuLtqneQ1A+Qx4
Oog8XChwYxp/43Z7U0d9Ww3TfFgWMZb7j12m0bYSwxG+2nW0Q0LNWJYJtQ94V8yfTivaIIbkD7Tt
JaGsp6QSsCYQFZ6bFB1Lk7M9TJ/RKHlt0U5dCMOwTRyBf1C6aIogb+1t+ilgv4Pc+4BRZ87bYvcI
hU0JTLSDPdi4Xrat5RKG+4+W2Yh4dfeK8HJSPlmonzaFfPBTdlfAuUCwHti2O2yjSdXwDwxEj3C6
dNQkZ4nZ3g9k25IjK4cvSz6P50y0QTV7zC+nK97qLgzpQAjEl1l2ZHkTmcP3o1L3sp+Wx2TVI2iI
HeNZArbkJGbZVwIRym/zLzrb7a62KdkEkSlz8nHwwKFwdod1G6g66pJSgIprL5n+Um1wrRmkbAwW
56hpVYi0x1B9ApyFJUVrk90+lEQUmiAhyMBTdrJ1WLI3lkITSKMfqTVg2VFnlp4AvkWBIUu8ELck
IS6u+nPq/egixcmpSpqZ6LIHfz2paMjSbzpeclmadKK2pnnUBGR0oKmJXZS7syBO/EGFd3e53itD
1i3sOPgYMv0Cv+KQcZTNaHq2J9UbcLloDnv6FGrk/6FxvdYgNzLvqSXDOdGvCbzEgZE8NtEb83f8
igxp9T7CDPknRcPqBmAs+FLQqcrMxPTxl0U6lXeLddDkZZ3cCVPFx6FBaEmtiRYu8oDGtAZ5+qBl
X3XEu4jLJEP3x+9dvDy7BGpC7eABVJYRxKHX/YUcnDTipg9P1aoBTaqrmtx8WUpj9w0xotFHd+Zh
S+KzUsJiofZ6IKUQVUKtIvfmFaE3/7N4wjofpQSb+CsNhwVlP7OS3o+f8KoM/3q6mmDr9iXN/eoT
xVLWtobQiDeQr5+S6TSJzyWSKWVhPlz4ZScva97fLHJTE27AsCyLWgBQv88LVNiCMgXyabcIxi2h
77jvRevLijYa1EVQyRxucHIXW6YqYEGm3K741t6KWhR3MqPiB5I6bf5sQOum/3QxTZgcLsaqERg4
WY/mx+iTAwgO7JCAiOF6o0EaxKrpfpLqMy58qF7/1IlIzShrsdogBqW5kXPslefJrc5j+F/a+/TV
cvhS9AHYfOiH7lVcmTbVzUxbZPod4YdBLWaclGewAicY5ZSM5uqCQYwkWVflf3A90sqOjpoEgv7H
6HthDmJxC3J4wUG9KsIu1LMujy4nnrJLmRYLk9lagLjd/xefr8KxfbC0vfgMZ4o3Cvtd4ZV+KpJB
PpJ8gNfGj0z564MoxF6gryyLb3VEcRqBGIx/DHebQfDOeHnWp5DpfADtMtVpy49KOLpxYVCx6DVd
VkPj8lxUoLIlzxHWIbrQYp+SUyEWMv5F5gST/uFn5pEYFtIwozfkKq5r7EEZMdIJvbvs06matoRN
KN9fOqRcvkWWyC7oS57XCpOvlqmmpSb7hFyXHKsMT5sNqCwwx6JL0JQe9ydhMibhY3+goOhheCVv
f7yh8BezqGcgC/3it19w+1+TRa8ErQtYKpQBSw7Qf57qgueG8m4Ihn8jHplAoAAyl1cftetpcBds
RkLpB+iu9xSi+pTijOrsDVWv4FFs/Ouf8s3YDza2ci696ZIMVKDdsU+PzYVVgaPbHQW7pr8WA7Kl
IrFBYsZx/sVwAy//siEG1ETwlbBFSPEHpn751Z4MeHbrHDmyjQEN+dagzfBCOJJICRjFOCphToDv
Av8wiNtLfFueBGgpd5Lv/UUU5bBMyXI6S4B5oyzUoNr4TU5/RM32cxlef3eUy22+/DrYwBsxog06
IgTy80e6zYbcOSKZoTo00lZ23Oa0ZtW5pR0CK+fHgWi3FMNLvxo3qsPUjtBAS8lA1lc=
`pragma protect end_protected
