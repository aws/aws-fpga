`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
FLXKCKlQ2DH7e+OaYz6vCHJq9N4+AuDRc8UfF2zDWnuiW3/eL9Txkr22DEmJOWucQGA63+hqK6ED
X6oodKcuKVZ8we3OBUtN4wb2DkSL5MEnVWnPuYvU3R7sSMecS4Do4ntSLIupVJMsmDXmYSH3bZfv
bWzlRI4iWBE4/S8EnsdbWpNlvr+B5LS8WMnzMoVn1PSiLd9NGhciDxChLq0VJrNZC3cjJH7rBQjU
Iqr+XSIDmMMcbbS/a8NbOWtt4tQeQXS/+jIr2IgjCicVzkyWwuLw/XQqmpPO2ObkGrGGb5i2vm1C
hBk+LkhfCaxPR0zijyCHapzD227t9vpEZERwMQ==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
QGkvBx4ajSdIlJEuqUzTvJb3B8cs8JYix2lQ3jcJKhK/NOrypYWO4PqIt8QSdl60dreb5hoT/rof
JNIPnx6ecSRLu5+1zXuYZ1AiAi9RpKci7533bE0Q2vmOO2eNYOhAizdS+whRBr/O+IZV56EBgN0g
Ixn3Xfnosw117aLH5MA=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
a8ydM3+5uDMAiT3f/Xk6trOkIyKZ4lYbJEY0Ekl+hpqjJITOPu4+SNEH+mjt45JrN9C7Tf+MY6kh
e8QoUKgFaFXDR+cV/RZuIfi3TOQleUc6LExSz0OFUkfmI2T3f8F8n9zfudjcLHiOesQmrIk8lQdm
NwC28qHuC0ZsZYVjq+E=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11968)
`pragma protect data_block
IWOBRgNSetM0QK+QtSTUbbJImF9fQcR5vXM9Mgq8Zwxs3ygRaKEAzeNbo11g7QVPdg1FrC4gjlRs
SwEBSytKsP8gmkZ+ukqPtQLEAQY9QyH83OTBt5AJ3b6fDzzKx3tErfHuZrTL1neJTmzVoG1s0a8N
2+LT/S6NVMYa8Xf8L7OgXQ8Y9H24T5KOO/d4tuqs4OB86AtteQ1hpDm3nh6/pKjjSds9qRbvjHA9
D3rcdwI7V1+YdgkDAxX1eX8mSQ7nt4WtADI7YrqMKPFF5rpwcuVUs470KDaqn1qGN1TT03g4QNoi
eVraArD5izE4KWJIBxjq0kkevxfdBImTBc9v8/DeFWZXaNY5pLKS/RZ1u8AlYwNaS4QwX2etja0B
rYhyTnx2oUi1eY+SLN8rw5FKfVg8OF9iEZ/McTxzTf47ScjDdaxgjlE5zoTlFbt9n2RyIPAK4Pya
xxlJ7NpqA9CN52Z9rghBgDZSUp2p0tFFRNLHYQsCcpyLa58zVGWe0JZsZZfPTx6Aciw7iJBzWfEE
32wTWOvYLUxJrYMKYlsjb4UYxTmWnxFDSoocsWd/GgG9H65gmgPPZuTdItHbMvEt2xKGfKaCW0Eq
jjIk/TjFiYFH56XzqLYNnEzKgAJnYt7d3CBkw6Aaxqm+3fXqRJtMfMR3IrdW4Gs1hNTyt1Ndj7jm
aOBCs0QQID+SMYPbPEc7noZKKFQZf0/Ndwv1qsFSSeqofHndWajA09CfJPJRqSIlDjVHc03K84sF
iCmUcXnMfU7xSyfwBPofdVYlJbJbeq4Ne4MrnW/ZphDpQohJ82bwxPtECeJjzYYAlNZ5rpJOBYcY
h5ksZ38PIpcSs00DtflhROoFAfncJBUoQba3bRHQiJKd0YHaXKim7nmVyOmdIn8330HwLOSS+b8t
+VcKSXIVdLAwV5dVqeUxHHplvz78fJn8iqAC+1ESuefj1T1HND89zxycRiJB5dYA3M0xyFVMxbgh
6xAcRFCQ9eYaqeSoHXFHe6pbT+UqF+yYQa8rFKnR4G0YSo2Kx5R3pvnXmwOMNx+ZBcEFXm1GVK/2
J6zT/w+NJE73pGgAAW8hBHTiiTeJlc7qdlpGRc9I9o1ClsMe75ALSwoPeo9ecHuIso5Xg1H6XiuT
skiYOn9ire4CvKNpP865UbTj7yWyLT4ftWwroV6vYjmq2hthRfHGxa6m+yZgNvhumwBadLTwi6kS
sG5HmY3r13Co3H4tnuiDhOnQccRIfPgOW/upNuDhJkHTAftm5Rr45YzgTkvF80pE1GffwBJGNDTf
Da+uiWhMFKpcmp4HjGFA/zRl5BNxQn01QI5gYl+9o0hmO/EAXmzlcyGzG+7yN6l8fd8bZYHuO1q+
Rf3inu0eIFCvHc5+iYKzV9+m5S25AG1LkwRTXCibVBWxqpP1pIqSsESjleBbEiimhII8Hhnbsk5z
rO2sbVPrNWGNZClyGxZCU9skIev4SB4v92uTRQIams6KmM8NFggbTAGuXhtsYL6qgeDPZbLqS+EJ
mZOUEy89Gnqoh5qPaFiWZS2/F2n/0MdvWw9Cx2oCL8cvzKzqnetJ7t2yOfZFS7Won7tkFTz+WMTI
iJWM2eTQOm24osh/Lr4mrF+nVYkslsfP9lkjgH3tsB5rT09p/B/ghxmhqmp1p1WsONaR/gu3IiYm
4AI5Am1IrLdfIhLskaaCrD4EthtYjbLrmAWgEzn21TvJYPiEgfly99AKRHK3PCOtV91Vl8mWXubo
oCk6Fjfsu1/yqHE7GIiQDKSKLsSg7JIPpe0LcJirtx+mKePFhW8yNJd+4eMb34kJFb/RXVO2kvj1
ONakPxNU17P8+0dhfFJg9TLwyammS/EE+eLDTfuuwlxUF5r7zzEQCHr0qn2VHavoApuwvYVyZFq9
SA/iit4SLIpL/mfIg/0zxGgI3GcrXNG1NUm4U59bhoNpV2vhS2Lf/nQjLNaiUoclCMBzpafGRaCa
DuzXprKpX1aAlDY27z1eqU0dpbWFUaPduBoKH/quifZWdkgjA05mpCVX7e7eRUgfuQTxFCoIi1SX
LQG0n5O2WrHsTjcjgbGekEOlnnXIDu9IsfpcB8TFAJw/pdCp0GguwDX6seJ00JQ8DZJR5R6Xcsu6
1S6mmYvPT7s+h1Jl3Qf+nQz5h1veB2sBoOcRT1AQcZxSK4QUC/ZPdBUsuQnWha34RDYpeiTrf3YX
MlnyvJOkbuMbLsQMpOSrX0FcjVnXImByJUEpaRVIsqUEKqbGAVJa2QJyjhE9jvFA0yUoatdoRGbc
I2PMffu5f6gd/+FV6I8P/HgEH5MKXgMuLepCpNfgnssLAJZodAvqmgItGBZzVepajri037kgSXIN
XLKmWppW0DfkrcxThWcQ4avFBooug1BrUjoy0fvzgtoDRfCrOZEapkD5iRk/shHDgzfG6w8m9NJp
vwszecFf29tWZ8kKP6LrSkkBBJcdXwmx85uFR9qDIzbZanA3MzvCEv+wvU5sB2OASX1b6vAyOe/m
XUMCbCh4odbxZ8wIB6UoiBgAdWx/dOeMy+3FLanaoRZdPEK6f37HmIftnImZHvLPSReQ7ILrfNr9
m941k7vk5NENp510CpYEcgZKuUBVHA9LdCNiVBNrCWllCjBbVPbqrobnKZWC2u+byv0ID7Z2oLHD
PXfUo6Alg27D2g+UXukXNOSiaS45ki/dT97unLvbSnks/NnUPVsR2c0luJWEuqvDzwjRPFYGI9Xy
F8zjbymfaHbGJZXBiKrmUWDSsUWm2gaACfLzaNINd3k6sl2ztAsZSbfhMf7K8ODBuUfdcqsZHNaC
Jx/qiBNuNIDHADETC3DDno/XTLbRQSLHwinMgdciZaTPQMPWag0fvQYpWYSzhP4cmYk2Ubj2GMBo
X7aqjpatCdZrwfX78jkkgFffPQR54SyKMG56tBBZ8pM/9guKY14r2vlUfatdFCAsGl6ptYJs+Q+z
xKebhsepLJySa1NMV7H6o9DtQyfqVaFGA4T3Lop+GcFNtUaSyz8vF+PI7sC2xeI5ALuz/9aWFkc2
EC8RmVZovMd5RWXFiLUTTkhwXh0bXiDhsFQupS/qSGQP3JlcEmsNZ+6UGhmnN+L7+fB10Ze2CyJz
k9ze7NWT148ZTv5rH7GzYIskMM8T+EqofAInrt9tkdCETcNzjbMUkNMbm86vy9c0hlTG+uZCGjmv
T4G973dTMUeozIDoV3B3niJqC6dVN8jgCzxGWkRclTKSEpcd5tPja/xCjGfwuRMmCrvne1gAECyu
uKg7x0p61PdlZuhd1Nw4A6nv3/5aA6cm67LUqSB4f7Is2eAlDVLZJWEoApOJI2xnnPphw7escH85
v4vPCFdLM5yPWwtBzUYEGm/RoQGkXoT1gCF38kkzRcbLdjgHheTUs1lSwm9deubVG4bsqP2+ZEUo
bLkA0+sOxbrRQEX3jPcRaGbnjpz2OQCVeRWf07mH3SnItqk1aczB5CiSr79pPCiNZ56x74cwWw0z
099B7OWC8aEubhCEzgobo2+GwpzQb4+hqQyks16+IV7tgRP/sgTWdcYTItlqND4NBXO9EzpQR+f1
7RQB8gu7nRJOVP7F8bQLVWtLtIZKSMAmDsZI5Ca9XY2HXw/phZupzJW2nSOT/CyfsUU5STVbieGx
8SjWRV/tgd7j+zaw9Aw3Mx2cj5Za7SMFqYDd6Vwx25Q93iq2nA41c1PC0xXx5PhQnYknNVDJLf8o
EibbogNqhOIF+6iNOuE1HKcZw05XLxYQEgafDsgn2IouHaQAZ9upwv9nu7v6ZJd5LeTKJka/3xFN
GJbyt3dSzJZXUkec/PwEhau/bfp0XiudlMLWq6Ker7pLrwI8gKckJSh8xmEFN6y9gze3gZHk2rkq
VMYclmubWgdJJNsefHvXD+Wld/voqxIVq/6fJJLZRUzDzek5GlstHnQKU1JKXRqCxs3GRab5lhv0
K1SoJEeDFfR/yRBXx+OE29cVgXCol/TT+XuDEGguUIQnh49PB3SY56zLzjQwff8JRMBkSaNLzTyZ
+oZDRG+WVQ4i4OvlaAVfmSxWxyOVBvFi/DSxRwxoyc3VQGqr1XZvc68xlIlTk1IxIG9lhz2XS/tZ
r/CPf1j2KtpGBsl2DrkYDTdat3kkAuqF/LIzVoYEfmIjoyyl2yTYbEQJik60s3KXmGIUQoFQL8Ln
nBV0Lo67Z/w21LfdeJpP4vVQPK+jq+W9invq7gO3uy0it3Y5u+THP8PwD8SOFLSvwMj2ukWd25ZX
X8DPtIWSMtpvseihcU4ahJL07NKpp6UHRDNo01xgByleUfGUVveIUTlhF9QLtqePInjroXO1WXi0
92Q+i/updZBqblCnnE1/aTP4mOAbwvUJaK/N3uxxHvWK8XN+vfqvgoLf5Dv7L7t4KsQj/r7NXNwg
vaqYtJ9mgFkg164x2OC96ZAkKLtx2L/M9aWe+JjauwxNzkJAGudwbeN6FKh2k+CiZJzYFWCQ6RIL
cpG2x+Nf7CzyOWahHVEsHdzLD+qWAVIFouGmmBp3jg/dRUUGk0f46Rs9cPiHVDH55QY6IC66/fo2
4T0xQPqAqTQ9MkEq5+iweb/KLqGTYldr0N1OezBASwmLBtqNapDeyxkg4AEG1TLzVUa45TTwywJu
ajw/C4ZmK4VUs+l+H6GikFwAK544h3gps05aMmvPxlb7OIicB8vD+ui8mCehETlNJSJXVVi+d1R2
ve6Ts5DQwbh6w9iBYP24tSy8uaBYwrTOSmoLrJqw/ZsLxKNqWJOoZkGEC5iMURcqh7f6uhCMh1dl
E3YCYx9/IV3s5mHfQa5HEGPLYfFkhDOi4Xa93CmBNPYLKYibioaZaP3V8FmZvmnehzPXz7O9lYmK
D+I33gIViqPh2IL96mVD0VdAsALhh8HIwmKHrJ8889qqxftqzOifNSdD10WfrBe9aKJOAiZyfx9C
BeGGqmgYU4QN6b/wBlPTLUY/sEcB+6mJ0WZ++lrSScom2QfSeP0TUc/a66TdqcW2WOiHOfS6pjFu
pVoQcI64576INUh2YX5RNC08Z6vD92EqwzuHXBqaOVtCB7sSd9WDqVoJnKlMaUcJE2xDGtxSj2ef
/w6dtAV3TweM3BNNZ8Z0za5JbH6t5PzhoqPqVrPQ5cN+wF9kBynlkG1dfgqa5gDbrFacOzR0XcSJ
bmhsWrzmr/g+RrtOda7AcfPGsl+Cs/jzYj8diIP7UgaRhyYbnszdxWjN+bKHjRVBOgTkkQQPObaG
fwUrbuqSqBwcPlt9Eu7IF3PqZBe5dJEOiP13xHBwriavO758L9bXY7JpU2xc/QNiK7DiQLxgAUuh
Bn5UaK1t8JiJxFFj3uClLmnguPqHu0YfxnKans9+4Q+qwBb902X2o1XLuQIm67biRgJS4wiws7JU
FRG1wOlUleUweJfNklAUKCrWoY48UQgHXZ28QM3HNn8PQ0QiQiO69t2V97xXHNbpR6KB+UNjhNIJ
kmfet9QGofm2eJmrClM3D9PH/8Yowho9B3CVbe3U/cg0kgEQxfHTGWVC7yuk39oHk59l+4nwlF9T
AXBHynNwzCFiLvlT87GNeXkrB3r1DHn+7og3sjNDytO0DTRDZr712gqA69ZjbuJ3Ssqb3Khr+PI+
y/Pqnsw1FrU6tlUvQv892/lx4lufJ6YWjPrG7e1tC0R/4qi6mLVPpn1lrwySAXZT5sEgo6Lw62XW
+iG01QDDRw2G7sTYNV3uObyhkhmHqeuQTJM+GT5fgN2xfROyVqjDJrw9W4IrJh7FBwUHzMr1j6EA
d85a+M+iSUCRaXWz24kslFQJv+fRWzjtgA5aS4tNXBSElry/+mhq6kECce1cKDpRKKK71bxpoKEh
F8mKVQJeI+hj2jxv4+PXIWI5VPxsSAieMgJqkf9ppYwLxEVlHrujIIpB7vb7/ZXCwDMawuFrznC6
goRpx69VqPq0VWsHIU18OdCF+dmUfPeQOOvUHB6Y2dxtiyKbQXkyL/BhLp1ZWvJ3Cm4sUrlcNlch
skj+enJtgdgQfzbfu1y7uiQS4Q6CF9Tcnk1DKktDo03n7sSu0e9Sz8Eu61BDoCMlsfpDWxgueajf
tnrXNaL+ZQ+7RqoBhB0dQgLYwakUWIWBm3NkyslQ//gGeAPRXx1k8zUXTbOg/WH3S2OwFsP9ZrT3
KpNDvwREwOCWEL040ZjUqIGHMk6AgmPU47fJdb02RYjJ2U+bhX8I+KKm8Qn0qDek8FJKuReJ/6j3
eGSPiThfbyecIsMq3/I4tp752cu3h6cfqRgKSwho6qlp51LqE3zXvQNc64RcuW7g0QA297xtIYVu
+ARHti1LM4Q703t3ilvR8MKrStAJwYfqhmHPWGdMNpebhMtrYfU0Do1DPDGrGoxNR2YbdsvMj0yU
uI8e3O8f0C2rgvsXbvvkON/FbTX/RaGULvAzx/IfFoDw1bsPwsWXrwi8AE9tgw/iIyMTYx23Dw80
xvRUTLKC4br84l/hlbRd+dY7aGbvswWsvTRYvq6JIc9OR+PkkrbY769wBBowSHayPvzo9VnTHScu
dLVws2sJaEzEJb72XIXBTCCCKPnBJKYukc4IJPbkym8X+3umoyJAIWkUj+YrT8l+tE3rfuy8vt97
KkryJ8VTczlYtUQDk8ksLyVmEyVILUPwXhV9nb7djZL9m2nvxVyF348ZZjpr4Dg4gxT6dXo1+NuD
a2cf00PPy6/2Ip5t9DKGws0Rk9AjsDvyZe4F/2AlBV1ckLZ75gRga7+HwYs0Wwa8xry5gS8oFm35
zkJymWvUwdrTeIPkp5F1QKriRI6wUrKQ5+AQ4PfI9N0W+5YjZvhXVvf29wwsAD/EsB3ZSm+FcJS2
/JANHPeCFNi7Nm0sCGwj+gAMOpw2CrOG3lRgjBou76pC9xDltIzWvQ1BELhDueUC5GtFW9X7qpYB
km6nC3nUJOZPIs4MYrvdQnp9NO/NH/xKIE/8GHe/mJrHtD3RlfyGG/mULoXP5kiebfs2FB4gFZL6
2b0yEaKXcP+jmpnRtGtAWOZqaJrj4Qr0f9TNiFOEG6dXPb1WicPy3bnChFyR/Vh6IMrPIddzVa+D
cFQaMJiOT5Vjiu5mguaPtCLn41i7P3T2Li/tZ9nv7yutVUE+dFx84Nurr3M+cMtrLu0T39egsI9M
TLML+LS0E/UIKstiPy6Gw6/BMoRWW3482420s267B+2fQzqAFhpowSaQeriwfe9UBL+xzVCIbN8C
BsU1jyz65x6EN2gqR2NnMm3EIP3lCk7EtZ3Krjq40adbSU2Mgn0E6gkwficB79UA/DHcaENkhibp
EpAnMspQ7JQ9rMG8CKHDw+GrmB4KUN8XWbwYCXPqzKNwpVMUtMYCrqgEPeJjiQ/KBpmfsLMwHrwS
sbmoviDkGjXQTU56PcjedUR4onlZHOR1ZRtCmKUFCbYEsLkh9ZRm06HttwoZqU65qxSRnAfmAFJJ
B413K7vEBZu8dr6sDNc88JZlTDil/p3iYHxb3w1k0JdrbHwLMyKXfhUToyU8D3DZ4tKE6k8B8sh5
LS5c6Bo8GhYjlAzxbJZu4mcIpppkbtTPgv8gdFZeMCdXw0cDoirTANXgmtgCjeK0kbS2O+aHdVK4
dFPu8qENum99ZN+/woYjX4X5SjauVPvGbAzIStrSFClohoYlcablE3ro+K7J5dpvAaHwVBp/bkqO
3sCUi37SL04kwwGfXckmIA8uuZHdjgm2rbNfoZGt+O/qhvjWzX7y19ZxLTpo1gQHB42vP7cijmEl
Z9fZvHHyAqUrcf0s9uXG9xcFSKEo+XDggWY03FotC3jaWgNBFlNJjhDZKNZjcQpW2VhqoekyWsRN
sTgqc6SmkI9DqGAYshadiDSH4MmprjbaPlwRzu489GiieXTkCzk2fXSzgUOf8/elxzcu0+wnTLeu
Oa6cZUfYepiPXb2yGxY29HWJr92gJm47A82wiIGI4de1nSccnjR+DL7kly5AEB/DceEkBzuD8/Yk
qYtrAbIP4Z04bO4+HaoNIaG0xoA6vEG23Db3LQWwaiCvD049m5QO556y9UdP9Dss6LHssUm+qzLk
V5f+Dt0zJQ8F1cUyd6t22CEibDW/oLSA+/KZxtFC9RtPE6Gck+Wa1UkBWhCvDuizEKenienNscMo
p1WzXSA577af8V8gWqFHfAOTldxF1VypIkBaEyjHf9DHNJgukd6u3/R8HYISaN0xigmyi+u6KjX0
Wj3zE108eMFLEPtYAxPfrAO1p5CJvagMcIEONFPtxV5BSIiSL068htGb2GtKzAH7N4Zy/AsoAjCC
qELFqbqlbfmzH0d7hI6fNV5VsVSGMtrAziShYwE7dEPKVTL5PPi2wvBiUb5F7WNitkv8bXjiDPLe
zQv/WsAsh/buSgkvTU/4GKOT2+h0xnXZDy+L+iY9yi7xv7Q+FKZt7t7Q04fgHOy2XKry5nvMO+Y6
6m7PidgTNWvhYNMXJWL9tMxttfX8M7pYSHgRickQIrVp3fvxc+W/Mp75fSNWyy+dfHgu3IecPB5t
n8xM67Gvgl+eB2p5uWsOLYmnwhVZ6MzrMw6ogpyGegroeyMCNxTT3Ybr41deC1vQugnDdOSM97kQ
erOjFSvmjEIurp1gVNXpZcsv3CDZDzy/fLeEbO4iu+GXEhnw1sY5ZZuJBpvYHHNN+fL+Rplu3l1a
aMx9QKQpxzPR/9P3BLfv7GkIWGNSfRO5daP60XyIOeSmJvfVxwnj1i+gcB5SUZk/ZG3sRIJoc/kR
ZO0rRiXkIwUTQf0o2hqLEc6cemDIS7bIZjT1raemJYbBy1YslnU3qt0/Nicb3D2NJzR1Q92fU+bh
AF2CzPuBfSpsTZ6uEZ+ecLRHf6Hofrg8EG4a2c/7fBxtH3Co75RUXe1WsP0Kv/3YjaihsC6bxcSS
pvC5bsIOso4khg2/eZuzFHkwuUfpZu7yH7Vt2rvpUoKf1liiATXxL7zeGtItcSDAAqj7hvuV/ZKO
RImgHV4xUTLGco3/uvqC0zK7FkGDhkQQ9HHo/cJcm6Scrt0fETl3M4k/4j40XsuUg4/y+kGpaatZ
nAQZLOJqFe8WIE/Xei412Tx4QKhsRMYc74BH1S6tdsagEaFCnnyx/dTLF60b71878EzZS2eIGE7B
YQ7Cfsl56WrzSx/3n/IgwpnsWUasbo9kc7rZPzqQIDEQaGDOP5ChdarkypGYcXkRnJTWlSkHh7Gu
HkWt69e8Rj6rmWpA2lCjwZ5m7KzGwK3y1sOWSVgIBteg6/yZfKXaKePntJ00U4mfwmCK3mRhmtFv
mXRYCUmLiulR11ZcXZlx30w0FvIG9aKJOTBHtVxFjxcibeUPeGNOU1g7Z2SNCkUFj33R3cEqaotf
r01EwHDG0Smi6eXlty8+RM/DcVUqHdKKHoV5eIWaxvVNN0hOeo4MIaA8wDQDmLbhjO3VrBicRROB
+kAM27qoxe9It0WhlBfFFovLYFEhaSxJMkWj7EglqK2xRk5ke9RFxcUb9MwOoIPO96Q4+IxsxGcr
KrbPrRNFJfnw/57zVGmR38bTnC1eNjKkLsDNRG5T8vUfVmC2jE7ud4wC5ojIAjH8V9UgTKOF8BIC
KWR32tqXd42OOlmy9b6Wiu4jNctymmv4yoRJiDwhvt5SfIXfJ2bEfCYdZx4ycaJfxyjH2TDJYLXc
S9xQ2wI9f0CYBECvoZS1u9BBD2Abx0Z6k9OeEnv2WSZ6naSyXZTUX1aLyf7bRiOQ0s7TAKuy7eom
yw3OpyCeZs8BPnUczQ3wsadEOplUERNZH/LNhNuAJMS//1N17+tcaskvW8lUBZ6x1ny/GlBLbsuA
N6j6iHTOzUAsk6cUpSL1WUqxF4ETgDfHpUEKditAet7mDsy/yK30vt1s+irJNtmnNdtQgc85RPcX
DpaUjSLhQ2m2jXn6eLhk+tIPd56qvYxdHuCrhH01Eb4TyRmC+2rdWJJNop+3ynvhP8n5Z9VTfArn
S02J0p1m/TKDguGOGaT3CabQ5UCF+fmiL+E9QQwj1GoZvH1vueY7OfM19PFVT5YoC3nsqM0LKYdo
QeGx3CkqCV0+xLMrVQTFdSgghz+3tFC2yX5GNimr3zcH6reyCSNg3xDZWuKHVBr1tnz4ZkFQawx+
VebugTfXvMsPxcUnn1KS1JpmItcFhLY5dfoEZ58daIVQqrVDSDz9XMLd3um9CVpJJsOrrEGoNtSA
3YK2MKHotXaaQnu7PK3RLo8DTInAQZnvufy8cGgS8b18wktEOTZAPToEBkol8empFjHzqMa+COyJ
1BFVRz8w2i3/9qSF2VBOg7ALDh6hbSp8D6SBU1a9LOeV5MLpiHci4/qtSp5UzuKdtOQsf+KyqiSM
VEilCDAHiNhy0kh8RV555Nuxe1wRxWIAqo/Gc/8peEB0ps9OK3VcTPGB8slKhwvSDjxQv6ncShLU
pxBo6yE++SMHH+Gj7GRg0I5OdEPn7ZrWteiRiXBaejmoyab+nj8pQmlLWN/nCCycyW9vxr6165sx
O5nTGYgd0NRKUfPOc/+dav+sx2JkWbf7HnD4hMiNjpk5EfIHITPauLYr5kHIjZPM0Va/iu3l5plo
5wj2hPJlrNpl8vJRTzG42YJvpDyODPFZ9M7D1kc/TdtSxSawJboHMuw52HuA5jX0sjJduJlT6ey0
tz0wBrX1evXDjNjmephbSrpLGYH6bmbpRA/GWv+FDKG5xPHL9fMeehnirQrSp22P6za/+SVIr0Qy
zky1fHoPxNH9nRXXEI3SJXwjZvI0wSy8n1anfp4cG0S4fXxE94k5v5AUscaRj5OmYta5fMc9R3ED
egMbLVrQ7jrf0dddktZNGTCS8f5jpGZaecEY80exniRSOAnRn47KjiADSxxkVCNq1N0aJx3VQDyo
SSVqihrGsgikbkl+JevkPnrNXbR5YU2W9NLW1JkXRA4llpe8QHMC6dbUg4PZAnvtOkSJ+zvbK95x
Ym49V/OEjjvIpH4q6uU8+X0CvB1OFvrtpWH+XxwfeNQz4uOYkXM7ZZG3ICxuWWNX9pvvw2e8TMVw
BrEZHyVI7yAWXElRwvV2B8vxmj8Ivln1WGwHS1dbogm2TmzJJJZehXTYxPB8BxyGH32f5G9BUqxP
MGRMHn7W0uds0nOkCGYqs2b6fE4R9hm0WMGBoeFnFJX7u7OcdkXKqnZf1h6NeL0PUehYmmN2375N
0ECG6Xw/AU987NPrHfXf3mYlLZBlsuzNd85S/H8A0g0LJZ2yQS/WUXQp7IE6rYAlX8Us3919UJdx
Sw3WwdkwjJFbDPc2ftiqdS0CoC6mVP7VoYb0RYmfPgtXaA8eP4JGbSCVFSkTJiXJkaFHDbcGwqdN
/76++u34qOJfU/JRiA1gKiTw+rNigVWG3Z/UOizsE9p7c05ejq2J8rJKwFRnpuBdkYIxM1zBJGtX
DCVjkS47DqrRg8wkAMji+oRURC9gsLRMy2AcLmFtnFSypOJIdZMVP3x0CHOsoxiad/+iS7pdF2sA
QF8pu2hA12nQcn3SJZymbRq2kaJm28JTuzgCH1zqlPGd7lpuSEyXHCCKdWgGrUa3QKuwHZ1qBXsH
vpjkAT3J79vbIJMwpGeT/UqSGg3pkWa5QVLliibZhSCNo4ihHCE+Vl1NPdYTdjVxEXeV1+AMct9Y
eaaXMWeC3qaUR8bCDVK4Y+3WjB4DD0BsB3EHFl/lGE86uNrpzpTR/suizeTEDGMra4utLoGJERik
HmMl8t+Pwngibn0obMSX+rFj0NLTectd7wb4FK2tNhdqAIcViNor1qPg3JSY1w7pxEdXkReDf/DC
H7Dtoe/ZRnBBPDaSGGpOo5iGkLGstw76JS0zgosMwc5WZsDKhB+wSpMDPV2TSYSwlVTISPUImC3J
awGorbnmNFZtKgbNb/Dxgo4a51SuC+ZvYl/tI8HQPA9lufcg+MTLYGNvThZY7JcUywn0gZ0Qobxu
c1xxwYe5Ip7yHLchwU2p/k2oTzIbpLtPIUfxhOXfm+RTjgKyqkMuuqi1LwU6tFc5dbcEtxSmY6jE
lzo9Jse1WFywM+nppi9CSDPg8Jsms44g9RQCHvZtCiy/TFOB0rm/fWA0L5z2f0vvaT2h0zJfGoZn
1iB2TkyruOZn3UWMx6fT5NM2d3ROSUvEfHNUDL+emikD9yfYW3Y/LT5ZVnVVgHeg7OPdejiuuvM4
Ed6xUFA80X5ayWz21utB4AfrP7ZIQyTzl44clabOkzO7E/u1wnXmkM7MIDz0tm8WXAzKiZ5gHGAp
tyYF3B6ZgHo8ekrXDyWLb6fQBsGaoUUSKwl9nA2O9MuM71l+CLq8SWUbxgLIXXwjiroZMhGZAJPc
uW0OMzg6sn5gean8yX1XtY7TdyFWPhOp296w+UumY1R2pnESOXNY2b1KXorhtyGYk64yTnLU0gAg
aIIcbhW6F9p8KwUF7cGpmzlrE2na0Q/sDMTGLw5jxwiPpE83D9U2yK4FwTNy5qrQ0oE9t3EpK8NK
Vo/8s2cZZuSIelNO3UkY91qs7o+zjpvvWDx6Kq+yvAvrGWfjX2eVgzewOCA/sbVivjRM344ARPKn
4G7G3rydL9xeZlq9VM6l7sgxDnRg9/vGuZkEIw56ztaoUps3pE0u3U0gFQsC2iDBZ3pAs4OGS/sh
9z5BCC3BWLyFP5IQHZ0qJ/EBDwaXD3vPBHviHm3wzxYDe4OOv0lx0I/PxDJLbqpHMHeC+D6z3OzA
DfHy7SMqFIEB9MDL2JPwUIA73w/ugwhH/o8hhewq2xJMkASwlllfMWqXlBmCkPIqvb03Woq8HAs2
ziBLS0+rSUGJiGuWEH8jQ6YIBcZo6ouzFwHFwbK+i/pjGCPg4xzEe8q6LRsQlC458yPg7H/ZsBYu
GSiHy+O98OklA8EaEq1/2YmzQTjxVnbf3NHRRIxKN9pyWgdxB2sT/PMzYr9IM9gqjoTlpaUeeqrP
2GjJV7ZD83qeh55GgPQigQQ5Aun3sGc5EY/1blAakfbHj5o9BZfRV/Fs1lM5xjbgf7bf0ofrZT2j
DYCHAZMyicFV7hTDDr0eQKXv/WpGrRUxb0gPNRPbBEChk7CJPrqBp8j4RjchqKH/zRaSnSzuOYIy
iAKQEnbis28Gqi+rywBj2T1xYiLfCju6FKLmwDPr0FPhkhMY0u42+NOJr3hSAjMaS7bQEaSoszwI
euGeuLXYGqK+MGG/e6VDsbj1zFXtYU7xZjorQwS0rGhQTSw8nDI7ypr767AdhPX933CKRaM8AzN2
iaNa6PBsvdyuzQhtiMHDMrv4aJd7ivrqbdoeODF8XL70zhcN+ZHkz7cUql0LSadRC2irvm3RgdD4
ySozK6hZTydmgapqTDpoAYEZGXF2avlqq3MPVPuOb6tXWgoDh2pVeW2SzY/J3jc2onqCArPbaaJU
n1nejiUDckNP3jWbwffM5M4nEmEgBdBeFPRRmwR2FVHwTbGsagxCoEL131E8WLqXJ03wGkLoUOli
ob4HBSlQfvWWv9NBZiKyrX9AVFLy8kNEx0flmPruyUQV14AiqK1htztWPq1uA3F8m427ORwNE2yT
Am1dofIrZ3ckjQ+AP5GFMCDWX7T94Lc1L6Q5uau74JQNjdDhFaZS7WpPsp5iHqacdLSEqV/maw8Z
HedZmmw8+g6p4PvvnH1Y1fU9/cNm4KicksHnUcFO5cmNcNmWrVla4JTwc8/GR0hbw0gIhpH+iEbU
kuiQtsvycYsiZguZQyb005sBjARPi6d9MeE9+NO6SDXtUl+56SgoWocR1oDRrC3WUkEYhDIv41cU
97yZYYghuPnqR9Hl/KfmmTIwTdTL9E3q+HXFSTHYojjfZtxUWm43t/v6saBQWUo46/ZJvqR6iLrs
m0nqSUixoOYNmsJzDGinEWrD6ob+4foGYyBDAbzqfNSyELoopqOOIaB9hgIrcb0RBY8tHURQQ40S
10Vj93elHT96lNR8xiyJeRTm/eVafY0lzZaXF1QcwMDdGDR9iJh94/jEOgEvNclpaD5ff8IvLT2T
fO/Y8ZZP7WqdpRZLNVLnyU3cmFW2z/72rFgawsuXizxFdTtyzSpEYPCq27TOqq902sKzj2IL5GhT
Ry0QUmEtCnX1zmoW9Y/bj4ajdJDr8jLKBDZ59M9lvakDw62AvYOcwBThsmSGFHV6LL941fpv5+HP
Da9y32pPjRmzqg1mwZ87zszCgPEbkfIsTeqE+0tVkREx6Vly7XKa3/dPPJmoyBEph1EH/wiXEz8P
xcb+eGEfGUhbVAPGuA8ocikd1ZklvuMmyxOluuFvV77PR6pNYwra0WxOoRCgC1wJelQhzd4rL3+F
CZQyGdJ/859i/FaWnhJB1XUAs8imqdzpBo91xlFA0vkAm3FSs/f4vr+Wire9ZefWKd6B2Lwjun5r
GTZ5668ku5t3Lgs+YaYDdE2jKGEXvawWx086ize0qtFNDlpAZOByg+YOWawp23a9JcTTD1HbY2QG
G3Gt0TBkNDPUP2FQ6IFeI3ZXr/cI14DZfUJl7g89AdYeFugdrnjKlUR4GyG7aUutOI91GjgIBWWg
JyG4zrBvusWCyE6N/amE4Lbtr7d7mLg+cSD/92x8AyDUxB3Tdr94A8RFxwRBHDBoulJF9501prI6
9+QB+makL1AykHJfMFVFHjv2khA5sQPw76ZcVZ+kJNFg86NIm7YdGTD4okrWLSpYkG5sI/643l6G
SM/SoAQR9NBmOPSgzKkN9mHN233Yb58rr8K/jhN2VMm+Jp6LiqVDbINBB8Zz66BWD0IZI+xhDBey
K3hM66QxW3H/ag1yFYUQOPIN1YWZzAT0kEg9S9am1pdYB4j6S8X5J7bBNuEuL34pXtRcYtDd37Vs
MHnUE3/cX/7uZv8c+hF3NsWatAy1ZyOrwAcPq0XD14Q9j8kP2CddaOka7EF21UGlgpCLljhdHvRC
1FL2rYXVVbUOBPqhmTFoNdF+zx8r/WjyVQWfkeh18/FSoCE5F+5+uKTb8RIxnfMF2gVtqY1rxz9Z
k5fzg+UsAOuknWaVNiUdI5e/dIdXurgajNuC9W6e3JX9WcXDxYde1WHOgiQafnw5uF1fMFMafDA2
jfKs7BYQrXMLNOx1jG0TbVqBFZuJuGbT65CnmlrxOD9vAdYZnTB0WxbHTXoIQ3C0Dn+Io81gdu+O
yqt4kVAtVsam46wNoThFF4TggZ8ziNV7+vvlHvgrpBgNRrbh9T3cXpy0DfaKgKRQ1AW5kXpnR0qd
NjlfQb1me3u/Konh1OekNGNVqv0u5Zng/8+dv0X9GX3NAwAcDut0k+R2hNNB0OfKoFvBtF0WY+2Q
ZxNgY/O1BsjtaQ85IowKD66Ef03TAXWqcm79yUnbBODM+7w9gwY0WWLRNe76fyEkAhSjWDsjKNAm
DVRSgPql6r0YmxBkNKXwWiTBxqLaKN+bTCSrV259PZ55RVsX8YxtNrdDdpAoGGBP1yqGjXqnQjlh
/Bvs4N6gy1b7JF248TfKRLmMW3mzxWBqsI9plF61jiV4IWkJkvovEUibR8428tFIKQ3C41Xuauhw
ifS0wBqvb4T2UhpvKpgUijsdSesvLgq6QqDABeMkYWh24TlDEv5e61gCQsck5LZpu7Q3VVN/S09N
ros7CHP/qw44+zFA1jngG+SL5XT/TOojgemJjpZ18mBwpMlamqXuWJRo3PAskoGQa4ONGWLF8OSP
wW6MtDXY4FtdGitIJd/NeoVIVR6Z6s0gDEcPqLVxErDAiinjGbAkZst2gBsCOpGQLHRgUSX+uMaj
F0xWZ5b/VHbWG7B3O5jrfcFnIO4I8jRji8QRS1IvhhfN2g4vcIFI/+yz56LJIWnzjR3E/V6KCMLn
4R4UcWc8Xg8CiAEGuKVwcnDtdi4xxPoLN7TIWv5D2Lg4E9oOI0hJMhEmgMTywjZ+PT5tD1dw/Dv5
JwkBcyQ094qJhFlR4rCEsKpYiupPRZd9op+I4Jpa1UvZBJPrMGnOhmc62TUdICSmOhX6fmZrZA==
`pragma protect end_protected
