// Amazon FPGA Hardware Development Kit
//
// Copyright 2016 Amazon.com, Inc. or its affiliates. All Rights Reserved.
//
// Licensed under the Amazon Software License (the "License"). You may not use
// this file except in compliance with the License. A copy of the License is
// located at
//
// http://aws.amazon.com/asl/
//
// or in the "license" file accompanying this file. This file is distributed on
// an "AS IS" BASIS, WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, express or
// implied. See the License for the specific language governing permissions and
// limitations under the License.

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
dqAQ0vauFZeaDsj53Rbs6p/DZ/JTW4ruygPimSmUvO7EqWX1gfEOacCSKTREiDt9fTnj4YIDhLyb
rl20oSdslc7vQDHIFq6NdbEUmfwh5QWKclwA1UcR42xBmtVwuL7ZkEITrtvLK2xe1PNUYrMM6q3F
5cQe+eO3iOiGC4rw32x9ATyL7kbnTxvfxQlsoMWVzy4u5og8dW14zBIw/Wxx0dk/fxpxbYTX5hyy
kynkYlOmlbcRFESplKzYXfBTMUm8CVaQkSuwi9t146xwHX3NBSisHi4bNqbXwlQx20ykxIG++n0q
UsvpSczxuvHa5n+BL/8BgTCpWodp1sfTg5Mlfg==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
TGpIxw3a7zS4TAGG8l4qer9m9Gi54oT9vttHhgr2Qe7ZYy5vkq2r4A5mJ6Gc/dZ4lVSlDiLbU5Mv
C43Dncen/YFluWA3d2kKbYdZ49t/mbxPXTue+g/vtAmvpVb4vB1sekWfKNWYGla7pai0RxTI8Rv3
SDbIeNsljJfC7K5Pho4=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
JmNMTw0qB5GOcERo9W/iS7pE0XRmyJmKQYWFsejncIaRcRaeRjbWZFkJQRFrgw7kPoPhGho01vaJ
SEWxeDWDoiUNJwarz6aLXYv+lvuF65ZO5pa/2MWQdYIwBRE58Wl9AheBsEyWjdqaLST5vKg2e9kl
wxFFOtcu5WuCHwDK1RY=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3920)
`pragma protect data_block
GU/1HPwDdmfkGUdApvCKFGT7nIpD8xdFBzCjeuQPcSrAWKWeneXkjQXTvQw915KNA3WcBNyZsu9c
8LBFSp+b9RPoOTLqrmbjprx1nzh1rbTCYQrsy6sM9+25RferJMVR5i77vqdWObAbrOwDMHB9mIMM
jA/KJ9TZ7F7NJXXBF6cffsfLpNFOYv/9S5fStRThYy+EvB5iiWCjdBFz2e3w5h1hKBzFhVstdoSX
APNnZAFjNovoMV0AQO2JArbFGLKPGXDMqSB6ldPoK3bbIGEeS/9mcbUOWsz2x/e/Ha5uaVGMdArY
SrWsRdtrdgzzP4oD9eKO/W+ofQ+CD/Brd+WmUmdDX2pltzzg9IuaQcjWOiiz0PN9Uj3vgvyf9JjV
a6IqCvapohZvd98ZnEzqrBpfqLvYRV4MfnmrXtCwRg+0VsuIoRNHhA3x00GRM/JYXWgS0akQZPw/
+dJ0+8SCLIb44sWWL9k2motydCxc/HBqeqRUGN4/FMVpkJH6/p3IOWJ/em5cX+Z+tBG1C5vuhBtD
2h9abo7OPwFG2hEjIM7gSG/9jrGgdI5uu4x1ATVIDI7uQZgasTTnP2QOsmfQqBJSbH7z9NodJ0NJ
qemgXYyJaqKNKql0IhdW9Ac8G5rZlMj/uwj0lx+bEkK6vWRYiliSWzClHTPmD8tvrAKfd87QWink
DcFGg59vIKlOFh3FFhF/r3xltU72jHoB7HcivmDup1wdaeuYPLzQBH22SImattY9s8s5yDv23rNg
FJmzjZEzB2EmYVj7de6QAGjFSHS5nYvMOcY8wfbnoUeCVllLwEXCaDD//CbeQTHv79mo+SzSyw8q
7R2pVSZb1PErE1WfPipvCSU/YfU/oaUnAKETu8FO1vdQvcWx3ewnYGNpwooXZWkCJZDEfh3MFQH7
mHREYoJDvbVDOUyudBNDEAXYRMhD5bvLzKeZQQ3wghrDhFr0L5jqKmjfvZqRYISpVLLu58ZD0SHR
ylrQiwzLvfBDJcQAmhIGd4Q4/P2gUaoH5NQeBIiTpmhxos9GHlYomQV9b0cucGLqGrF/Satdiqgd
+zNRRfZlO+7ToWDiAlQhUUW2BiQ7mRyLrWZfOuQhCCc3KUkGhfuvHzuqEKac9lG+Ib+bYO703HEP
bBZaeyBQHSzMJIKtidXz4p6HlEFJk7+W3uBKpRJMzIskLJdj38e40RDgFttQEZwvikZilIi/WKfE
uoQZTqAlhrd8S8Y/vS8O3JSGDo3RI2etrcpdnIMxbTUdQLZd5tuPheknXG19w3zhXEE2vy+JPlmq
YlZQNrHP2GJYennNKj6l3aQUX7JjE94BfLjjmL/170Z8DmoTQjlwB6LCMqbVUfzbLgwzrTqh7Ps0
+f646b29/nW2xxyEBKJ7raTtIVGiXgp/hiMH+Y5UHkcqBPGZfFyPOmteYe/y5B9elECGZ85a8lV1
CWWfH7tYkG6HXP0XMAzZgH5AI8u5pH30hwuJ9j2f3aBpJX1z4irR3Co2fN0XHI/ZSAoZzQWURZlv
3x1alhpqL0IaN91wUFk9aenhV2lqeWpIRf2CZnqZObGSjt60CICuR7ygIPUbVg2iWhH6Ucp4IJQ9
5+bHkOmLcSUB43PsFlDMGZqu0KQyaXmPQvOxqGuPiSZqOBK+sbawwHHosoMGdQdUK0FyQI+dBeWt
KKyr9AKS3uHa2E5IpyuqenfEdf8C4OBfKkpQ52O2d6CYEGIRvk61VGNQZ3dBNlBIgxzQ0W0dTuh0
/yLH+cL1MjbzfmRy4CWArWf8yu1Nk5Rfk6gtmUms/imj3lVoMd0wObKMA+1Ey6WKrDky2bFmzM+S
W49kpDFztwgCEzMf6KNqMlcLg9m8vYm2h+zB0zZDdDiMbp46Ev/gLsJ3hGh6BtpHFTvH9vqXMoLg
pY67hY9qlomwGIXSRwl1fGnTznUNrvxMZFF7CPt9vSnvyiO2FmBtMUzoEvqICPbUQVkG0zGesWme
816AGYCWAxV0x5PpYrUhRdvTjDyuLk+SJ0S8IDYUJEuQajGLHR7O8Eur3XkYQzgdaMkvUQPgczBI
AVAbZbUJwVIoI8GcWEOFZu3uPvY8wJvXMrmuKIRgSM4KZTa2vtAEOUULw5NBqXejcrD63gijwmt1
gbcI/5T/sd9mmzUxuge7JsM2SD4kJyFfwI7wzh149egi/MHR94Eszt5DnnaRJ8YCWfb+wL78jA4M
tQBbrwcxrBRB1/Anw3tD6QphQFhRcevQryhXFadNHpDGk6tChDarhmlBcA3mxOZ3xW/h9hr2iCIv
32N/Ij1u8b7sNkkFkPxofxNgrOXQ1k6+LwuXFRGPA0xjuCdY1d5MJ1DDHszYR941p40xyTQCF6a5
pa5QQvu6DSXANSnX/CmdtWDj0f7rqtNZiAYrTSLxhLncKNqyZSVqsk1HX3geD4gWRActd4X0iV1E
XH52ZS8sb76FA+cNdMEhqUT1KQThmBXPEGqxA2LbmMl774/J00CHk+DRWhUJEEV37MCj73WvKBK3
+VkqiFtIKtXdwTFpc2iPZi4lVDPRx8mkdZUNWuogLwDtncXQyR1OqDRZT73nYhctH0GshWGRr9An
zYBDXKtPBgySPGFiX5elVjD+5Y2qvANMTUXBGN4lMOMx5UAjkhFt8TG39yjlde70GbWE+bhPnfKD
lXSsRFWgU7TIzc0B4HiQdLyVesxLlFSpsCWgRB1NES5n0ME1vCUBf0AECKRkOqI4EzR5rvTuadhx
i7WhGG+YlUGpB8fYDL3SzONz7nMzstCwVktYj67qcCyoyD56jAYaBOjnTV7chBcQwIxfadMup6ke
uen+IcIwnQjf1X03dnWaXyVysgsXcDY4xtqefWJNsELL1Xaix2NZwLmQZKNcyPa32i//SpbSiRwH
hn6eH1SsTVPGDCqehf6PwvnZHMHwKhT7fiY836YL414zIxUs+SEHb/s2XmLe7EkBjKd94eG82joj
ziYNIn1O+fRpwOS1Vz0CUsaOwTA4XFPZMej+oNACC59y4KYXT+ZTbsabyn32fSQxN6jpc2uT7QBe
T4b8I/biGoGy1ZMKMIf7YfMQKVc2E7dqk9huH+mWCGKI1L2Pl5Csppt0xTpZ0K46Z2/HJKnYYNsP
TzxepJ0p3Cy9qWMQwAq01f/yOaGudb1KrUvUw8g7RNTgzOeXP3LegjNNf8rLr6jFx3j8bajNFRGb
qsmLkazzuEjuVwYLTyKw93GMacdDLfUzpOqFSEkwhEeJQn85fXYpVdF56nzRMvawHIyGTU4iQukX
XlC5iYIyikuw43mqnNlybb4MgLxkYw1z62la0v966OiRmuLTyzPCX791yCsmtJONttpA/NF+IeEz
MamuzeoR80TzDsP/89WzPebTBvxKK3dlNnqkNA5ycjdlvSjQC1JPxEpwsa34Dakxn5xH0NHwzFUT
BfWM7edSvY7xOMGlM16Um8Ux90prS/WzMNpuvmnBBoFuplYWnylVnSDip71LZZYkeQAXq9wW51hM
ZUWPQhzn0l6lUNhDXAxTIy/Kah0p0cRDAfDxx98W3wKFrs4StxF6APF9RGQ9PfijCEfZceu+Tg6O
Gy+JIxcF7q8hU50ihXCNqRiNBp94jI3Enywgxfpq14kuKNC77cjYD/PMLkXmd/ixg/BTDgaSrj4/
KIQ60v2KuYYPk8y88oBLdX5X8sBMwJ35vYNCRHT28hvdf6ecsqALWLzbtuzVbQDY82hb6pttzo6r
YYQIx+4hQ0pJu9ot4WTZ5+WTMbiPL8Q0fiQAgtBrQiPyquLPNc+emK5deS++ziqJCteACu+TwYiE
LD8rS7dgrl5oERbMwstB3k5FpSHe6tikD1yykXzP1FAsklRvZPgCkoHafMOnBEH4TOWfJhjv7tVg
Ia1lb1qrvmP4kbcXkHQce0A4eCqO0f7sIlNle3ZZe6myNyvh/SLQrRsSH0XKO3iUyoJ/mZDCgXdB
JpRFuGzLD3GreoBrByaPGTgFesgGv8zM+cbQxC1f1TPEbfmqKlFiLWsP10IyJgMaS26lnjzY+cFc
yeM7AD1Z/p0vu51f0AIN0UeiF5WqS6I4O4HJCZ3NT+DZ77hFnDuH/8FPcXsn4kV5hBJujaD2SXOP
psU5digRT4253K/3sRWE6MoHLhoX6Ut/C1AbBolAsAP5mE7ZEz+blFcTH6B+KO/P+TeiL64qzVN3
/CmlQqSnexjNjECsdghN3jzoigUOkR/xSVDV8ZxhE3S2WKQo65Rdb7DMz1egLcyPfOF/7JnurUW6
tgz+32uys/4VRO81hnxRA8bf1Kq7aPMshz4eSCs9NyN5Emi3TvPK6yekltWt9K1fmLdj/j6tnNqL
6Yf7XRerdgVxBPZjLHsGetF50HI6flwoSqH3flhgnWZQ3F8UGB9uVATxP4zadJLvH6JJT5FLtKFO
Dz8psPKwKv02Rj+MSuIwo/IOotTH4plPEhSlsATMkOjuPbBuM8vmmz4FHru2eY65/LpUHG0A1TSW
rBVP1STJrw/q99t83lzz+8sT2Ru1LX6yaqPnjVjnOkZwLiqv7+nRR/cuVjNxvmrki9/V4BQ/imln
3v4rels/pmBpmSj0HCdK7zYii/6lDFLa3VgFGbTg7ZI4E4Ruf/zw9MUwkmPTA1HxeTwJAEa1h1N1
HX4NsKVeTrhLyIqfxkHLwAnJGInyFwktIfVRaTc+9YDSz/0zi1DRcZbR4VdIDdIJpghvtXJ75el/
PNbuIJAR6ohoaq8lxtzvvvJJujaTNmsvDTRK4Lx4uuE6PVEl1XzbVMQMnqV3cZnkCsHj7jtP8B4a
DwO/DnQz0qqSzF/5nO5Nn3do9t2eCmaH3caJh4ZhBTUMiCP1UUtI/zGF1RUvM6ndkyUnIr05WhS0
uCzmrydesKO1PrsGsIRZq/JfZS2fuH0B9k8dTNEjp5DA1RSeQRckVP0CJVcFnt5xY1+iEZYwGxKG
xKs53N0luRjj5vAmzaqj1c3Vanl5ZTomzfEJJEqJ+vUf3cZGVDH9ZjhNYwLaZccWgWnb642WqG1V
J2H3jKhFTH3rvnRgWN9Jens+aHrAExgZf/oa+v1EWz5zIaiSPJ63tU7+iSur+8gfSfXZmX/pjXQf
R5i4s17PXQCX9BZ+j22wzH5exeuUer7bXdTNjnLRGOB8utt4LKR1Iak7Q+74RBcoOBplaN8DKFQO
9wMN5ZSrb8sGK3gjptS2i6UqL3s50CDnC5JUx2fc6Naez5tsJ6Qo1LUlONM=
`pragma protect end_protected
