`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
T5WV3Oo+jqhyGp26BMbmUPJ4LktdsrCWXdn6TYhZStoo7g/3GVO8NswF9uqEGjaRNCXYFPxRwpbx
qxQlZfPr32z8B1CyMMmJU/4j4lrXC/AG0bNi6ZpUVu53C7mGALI/nZdbyR0PjaX/p/ssSiQP1aPt
XnPhThknLDs/VTrRP24ob3/2iBvwwsSmvcF7R1SzV67FsfYAB1BLc+ddmiUU94ploYKoQBtEJt5C
MC4/n7lrKVPErLKV8EAF65+79VN+/mvZOkXm14UfubQu+Bh5pVLG4c8GitEHwMFVd2R3LPFCX5aN
Pj7nKsRvVmmAvR4YcvmqQZRh0Jq/rOpVxdsiBA==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
dKI98HgZQ7vLlFRHkgnKTOa8uVJwKy3IDXpcZby359vhfrZlKe65T2yMX7NJFHQoUvkghdSlVGwz
MY066NbNfKMIzMXfR9Kh3PsH98e5ooi/C7dY76hiIKtzgJjsqrG4h2nMpj5FMNkIlTIf7IfH+7eg
CmLpbnLBF6s8tZ5L2AI=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
XgtJtWaDHULPCtqFvZvxWwkXd74+OVMoQSsg5Y7zoN+sCn2zbSavdBW2njuxCIPS3zuAEQbqvohK
QePfPtTMRddyLr6GfbJI6+DKhyEhpE8uyrNZSi+vZy1YQh/795tMI6Ai1n7z26n7xazgYymy+ANL
qO+snsnsrKnHWzasTsU=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4208)
`pragma protect data_block
hJ15R/8ygDBcM4WDJHNA0Q1enCKjWITlu+oUIdkDw4MqQ94eJ1ba+88iCmpGMIXKaGvwPY1GuxF3
X/yOd+DOTXvGmqdDMLryMVBcpHkf8PSSIP8fmqTxQ8SBRcQIYRr7lpwqJx7P9GARxGhuxBMRDVxs
HZl2V5ouCTrnuayNtyb0f8NmVAEmx+RkAWGWAV20TX2rBjuXBtPpVFwHmWaY7LmCE9oDuQvM4JBd
k0gHMy0xh91UvsXVeQTDPSgagXzcjk1KOJvxi+7J4SkspW+REsRN/mlk2r8e3rjccjT4rHO9Z2qT
8b66ua7GdoEZ89ViZuW/rlFGON3dY6QQzomBM4qZICR0SyOG5Li+hLtXl1kHxYvaK5cRQVH8vlDJ
lP8C8/wo+L6ftnnn/HWTB87Ag8dExblUkyjBNgj3kdY8JNu6kyu1LHbQtzdGUsi2Nhfdy3cYWIPe
9QWZSSfmF+ETQolY5Hbie1x5pWv88gRpsLJyYjGyxbUqWN/jylkVmb2Tko99NPZrqFM5DAEii5G6
3X+dK+Ylj7Pr0dZYlw3b79UK0Lpsq5K5cRpgX0KcowfXZ2WJFnfVvw22rYMQMXHVT887f26SPq0i
RAvYSV4VYWSIz4eLUfP0FFW4xfRTAP/KNMJ7vghXzhKlIBTljQNRwyKxbfEbfTx8s5LhJ/rY5//4
hxGL3ADzKUiCbvQk93M8ICvLF99Yq/8HjXgGYLTwbFBKrAYTEYCHB0zRl1q5NtNoooPtgl+0r1Nf
UjzP8qxbm/A/4+yoS1fNSNvUIWVCTQsL26GoCy5kKicxOMmmE+I/756NkCmYupW/qmR7nq87HzLZ
1v3AchOEEHcW5MWiaIzlGwCTPdPOAVBTIvxLwj4oEJZAVabdjresrOPh+qV6RysY/eZjMIrrH+SV
3USx8EVsGUS7tShIiqathKtyszhEto2x3t78OVtHWxiEY9CKwSHkAc9O0fAnONFc66rHA/MBnKYZ
UJ7CpzgtpMQD/LyyRlvjj1s3MYlSAGAijN1vTQWzavGhL39bMiEF+c5R7ySWeuznuX323Xzo7bOy
1nUfzf/SKBm0HOF46JFCZplLa/tiXDku23f1thi45XU7lVG7lwCp7r7YQUoJpZfFKKRuI6MDbB6e
6uDDT0552UivXpKf+VcJzUSoxP0FiDq//LwqknsOpyuqU0i1r51IlZ/lHoSyHgKMKorithJC7F4b
CuBYM68ZXozQcM4xZE+hTJ5xYwCpyfyRKZ9vEIveVIIvGTbrAgN56lB++m7atbR1P5QOxvzPj9J6
8xGEMN+tJaoa1xYq/LUb8R1h38L/Jfwqd8WyZt1NEUT+ob9XUrBwGhKhHrQLzLVdaIndTFGPSabK
tmjaNaH+0myOSWoiQZRBghXZQglGwxynNlMPdurNjEzfh4HnBOiKLMQI/UhbZ77eSDHyoJdqH3jU
KWLXsv7o1Hv7dKxy7OgmNun/zIuXYs73vE7+8qx16m3+Toy6hkvJ3YNP9FY7z9GoZHPOyxyaJsRd
P37FE74zeDT9nRvVDz3s8XqhRFhRttn5JmK3zZkcxQjiW/t3gsCfMQTrdwpIEdRRm3iEua9Lj5YE
kydhD2Xnqr3gLGK8nW8oDfVpHtFizLI0bgdsSuBkflzWI7k2it5vSrjbAqf2EpaC/H2aF1mDtm1a
gwmMNz5w9lkFEf0l3ZomL0ERSDIdmKAV9jt985D6L8c11A0eDH7CJmkqMIrnsUfTzUMWuuSKhHKT
G0kkRExcd6AQ2eG3vs3K3WcWFFTMRcOYPtcv5W3MMb+wcekSQz6F2p7pAOSxXfTLQi9A4SbMMQhu
LeryOIee1ChmnykwZH6bbNzaPzlnWHmzn94tV833PdVbiAtXEVvZGqIbjCjyH3mKOK+Pv72s2Lks
9fEtJafPJ3RSFu/tiomY/Lm494cbDz3AjAPlxZhxB4JnyX/vWZqF5UdPxgOl9Hd1Guf47IfiBfEV
L41VMLIxBB87U0R+h1BkTxMQfwCcuG6eWwu4VySD4QiB/lZ/Qi9ASOL6MjXK+wDMWg+OBC6Euf7E
P7qdJypSibSRCWuhzU3f/hSFzr7U4iOITsXATwF1vbGRq0ej5LleVMRw7tOEOzykCEwiLujACxGR
SyryszPE205WveQd3MtTeNopmr79nNoyLAO132jhiaklzMCIpftM41QdPGYzTEuI+HVplH4H7sky
UMBwttJ5g5GKZiRBOzOcCPVFPDoStvkCRN6sCPq+fKvummE4S0kJYJ6QifZ12MQ90RrNJDtPK1g3
JiOzJ8fBni8PgtYJS/q5v8XIWdXRhTn5hE+Ej/MqizQkj67iy+/Me5mFSrjdw0K5eqMs+4yOV77R
efEr7GCZXt9xMaZbiTUr8KTTHExyPrIyi2zTQgg2G4AvDXzLYlfJE2b43M2r5GJHuhgmjeHrDv59
T0ZRjgT103eYeiqRvlVi7X44Z9na3Y8lSE/bmAHaqfvnbkR579iX3k6ORSPTc/zXBqFJj0D+KABK
KpD9x21XFvgQ2x77FP6atc+32+xWwF3BZcm+3tAzd3i861c2mq1RWE1CgwIcOCaST8gX4b9P2DNo
tyHhym6D5tJk4SLB2FXemnPc4YiJx7t87zV63UcU2fk2vtXirOTSV7EzsySGwF8+QiFfV+4pzcFg
KmYUArcjARHw9kHVp1OEZHYIdMVkgU+iJkKdXSgyPQI4tcGzGeoHTO6dKdoLGdlq7V/Ggiu8u6/H
D/Ax/tJb7VhWdQsA6Vmp6uUf6uqu/9UvQdw3/QooofLrAaF1ipTRJ8K1iQN/pIXqqljcio0BeLUZ
oGCVGYgN9JB8gZrsfSef3tYmH//TXfO6u+74dUvqbZjCYFXy2qaGNsP0WQhmmX94sy9+NGecsrV/
jHozCdrePAJQaZfAQuLZMgU347L5GpLxwSjsKBVToPIpyoXoyqLJzh+uWmxMY82+rrQPjKNhCrAg
Ork/RTLK3zvydsL3o/one3x212YrjjCPEjh7pskRRviI6j69TJJW79WkeZqjxRXmkWLSXDU1xs50
NPrsif3CA7JkzLeC5wJmbDzW414Xelshtry5d/86TvsXxslmmB49kbgCPujmpK41PObmJukHwrPd
vLwDMgczZ6HSKdcaLO+MuTZRVNuIPzfOV3mPT3qn2Sw9X2DPlhmHiTWxTbLJ+G+9o2+/e6DaECh+
J8NwS8f62W7Dt7pqWKU2U4HpdQNrtEysoskzMhVFBAKPEDrW5bOu3qXBMebfy65Yy3UXWYE7KODo
u2G2MsL8H92CUKNXQ7tCi2iXW0YDnTNdZRwUgboCrgSiy0rdlE8OGCZ8dO57DMfDY/B+490WZD7E
WAVRnznottFS/SYYcDetNweQK84XaLJt0ov4WAZyTuOCUJijFhmM9yG3kic6fCNaRAohg0G2VnmZ
nu9sGg6dPLHYwk4RWHWcY0oQGAs43MtbKpaSZnH6HFdJ1Py2j6YeFczmSW38tLcGaRa72O9yMqTi
dgrKb7GKbRqCcXyam2wnNhsUxGbSubGlN+tYio+7btJHArFyxICO9KXzqoqpLY3w3w2KMUjtsw/Q
QI8U6U2bxv5LTn/YrIfxL23u0jjVajRw72EWF/e6H33Y2uaBilTGrMAlReDLM89zzYdjs21DJTV/
3MMll2RrUae4gxZPa9xe//Uj2NxPPgkJekn/Ls61AknR7/Vaz/PS9HM5QtfSWHgoXPV2muVhouLF
Ttk2EEf6aYIc/A/FKEQnrkbbN0+TUUYGqmASKlf8YiCCncaIW1tYrZ3hrZQyjVlu1RRZebxxxm7S
eibHDvWo/BqBT1E7DpwIVnc+UMz96bs/Vq6xjmWGElf81vF7th9X7PmZwKAKfSDMk7tIHv67sFpx
PXWVNgVSl1CmfOXpyR/Rj+GwodsUBnrzgNtsojHYIsC9tSKVYLcjAtlTagpmwaiHXavYu6pdjGuW
wo1unCpI/21VWuwcd4nyzzLNQiglYVzKgWB9oohpnHqACnwjKAkR3U49goD9cE18WXaCl95cZADm
sIuArh+kMfcqg7XlqztwY64gvVLG76jh8Vp5L8cPn5jJ76AfZCmLtIeEBfOuMT+UY8DTI96Mukde
QGTouSQNrxddhq2pKnkDHjTGOTQWIPmFae+578bk3kmRjbOY6ipOy8Sgr2/YLvPutYLADFV84JQ0
QiauSI4R9GN3t9fvsxpS58cyMDnWLWUPodlqwWV2Q66LLR6TvFtISxH4kk43zN/hqTRwUqt8Y0RW
entcpNXM27geDQfDTnAAcWI1Z6bpHdKYtT9YpaKIFnos7fI9MoSw9gk5pfryR7QtcpgMxm83dOK0
hGdZb0IFmUl/GsizS/Bi95fiYlM4LDiBNM1i+5mX934cPbl6wD/mKOU41xgYSkGaAX9TfqQYnTVR
8rm3UIVEMGtHemb1A81pdrrpIpaDiQp6eUw36tJPtgE++TJWuWhfocg/FeymDZDmtDv86J0hsL6M
xb6xZLPUaNGMn70eNvapub0kdFqYOP/2p9Erk6Uwnjm22SYCeeFTUpLUYFNKuzNQ21u2HJ7tb+fc
RcgRRMI53cufqQ9JuaMSqRi2a141DmpHf9bM52VIlSr3WxNFfgEXrJu/4Vv91lUJGeddUh4fvSOm
GsX1KmYA4TPKv1MSnxq/fH6OXwL+4vgZWGZbcVG4rJEKNjYlDzqnzyVDi93lkg1bDsO65bcY5ERm
cUDmOlVV2iNHASmEsStFn/OAOPLb6biJD8Ij8vaaX8zeb3YUiG52YO4ya8uch+J4BbNpzGdAcdWf
3gr8cYcu/kos/8KwIrx3xNAoz0DBsa9iNtRAE/4nzbRVlKVVVvp9by1Rw4F4AIDGazvId/xpvS4G
k4uXccFM92YMsejAI6z7hrMDL7R8D2zBGdTMBF2qYAKMJIJhdbnRkZXzi3TyeH/P5aAw5wYE42TG
psk7U9PEXFEZnEoPz7LPsvgGav40h2giYdWBpMj+5lQQkY9ev0v7Bc15duYhjWKwWR4oi5XIEccl
+W3FwNQ966HMVc0GmHfJ2IdqsVaLQbyqBjylxrQgDIzMmcumr/TGFuWwdr8tcpXhtyGnXxYHLw03
lTyEzcwYNB7D/STcTrLZqcLRHqQOzD2eVuwhPuG+jr92RuJOaQOldezC23M8+WB9Ifs0z0aiMxc3
Ing6bBeefGmfZ5xqrhd1aMFtwX6jA8aCieCFnNKIhOdKHlogl9vwDQzQ/lZmUuMOzENXTt4rkY8e
JJ/5EhwellEk+7PkzdosNbFJgzmxsp3SRNow0MVS/5KNikylVINeO1nTDPH7tpnArObGbAbickxx
c+5WnEDGtCUlvdiQ9MzJaaoPikk+LSuyNVban2y606pCs9bu17AHFqhwFOQGDk0wqvf3yBhZb6gJ
wDZawDxrsmSrPdoIhcA2/0Hhjf0LIE83GhfHoC2YFgpd5gXf+X+T0JvfY5QpiDqNkly6cOv9QBku
xzxvFv8XDZH0HBZm9ibJeWKyiztZEDlsynuzxGFS1cpx6WEvDrKKRFCW7qYxkdgOm06rJ8Kkg55E
+gyLWu0Sd3V6kng71KvanZKQjOjF5s2jbMgksjcDRPrxxQLqncH4cBxH188s5p0=
`pragma protect end_protected
