`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
X7Ap/lcDCt9P4Y3yMp9tdozJADghKxUr0U8MG7RkfxjrrHbIPEW9HtE6OYrFUVtsNvq6ITpS0t+v
vFeB+9wCN82bredOkzoHqSEdFijaLObUNPyRfSHKT1ODlXU96y+peSt2S/pI5OgXSuoP0+10BdVu
3yfQSCibrkHZHnEvUGCD3LJWxubC+l9WcqomQbd369MUL7GSkrXMdj/Kgt/zFhnZAlBT1RJrV/9W
4RVj1y0TJoBtECYZtwQWtJhMLDL70oCq23vYUVt1c3xnLzzESPkRJx4+Jmf5f16Yol1DfnXl9++i
FFFQDAkth2VgsV5j6DFlsQt/fW86hpMf/7dFxw==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
KLp2ZP0OyMs4w0hL3IKSR6L/6m3KemRegwkbxv6gBouNw/n1F3X/KPvT6c7BZb5FQ62l6h4WNPmX
tqZNzXmekfbJ+8f0QuIOhwSChes7997xu8V58EDVZObuYMUvEzc6JtnFRL/UsYiMPAQ2VoV/sKZe
Tfolc3Hj2D2EIljm7Cw=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
YggJi7VL7yilmca/WxYUwMY52aVEwuKDT4cSf0fBabbVSI5Yoc/ne1H9qSiTiDdCKK4Frdn3lV+c
872OMiSApL7sWsYZ9XMjFD7sxKN17iKY79ADkcDspDTtr4m7tDGbcpPcuKfzAH6wqB6LW1/ftPPV
+RzkjvwXtMC799LHrbA=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1120)
`pragma protect data_block
6Nw1mr5bdFdum9PEh2xUPz+T+jT6WGAhJbEMuYvOnXKwL0ONYXDPn+nkzFQiM0PsjYFXoQvYzOH0
bKw66KL+zsD6HvZHNCYMLtbZYFyGP1Qx7ZeHwyZ+w2npvMxfO3/erTP/cbeQQa/XpD6l2oSuKw7G
NL3m/PlVXwhjrzUivL0ARil71DAjJgxgCsKxXKcvvweRAqIA9AwrGuj/uOtdVmhdSwqOo2UW7rMD
cjOXVFuJ383N93q7nM23yMnXrhEyPYoVeO7nEqn5bUZovxXwsH78h50eLQ06PULPTC6cFipTRtT6
w4v8YK/BTJbKs99xayHKf8BgFL884Vkdn6fXyy8VNNYFqPoFer3UTlOsvXyQ/7bJWb4rJnbpY6sd
6TRPZRJTsi7F7EgM/oRP2ueP4fauJBsQTGmi/zhHNvsRCudUuUZ4/iA1Hr+JrV/hvTYsPWOuL/v+
BsLjklo5xeg13qAgZ7G4+EXgNADrMCa52JFDKZz0QoA45MAv5JXc2sCGfqdJ9Oxg1ksFo8jV24/K
q/twZOQygi8B2ypXPmJRc8WLJ6qBawy5E7sfduE6Q9Akt+W+Num4SUklTj4nX1f6dItHLi6gue41
Kb8o8njask1ex+ZYg1uOvI3Zu1+eFO6rrloq9Xag+DcfFWin7FzOp8IixfTXa8P1T1xdd+PIwXGq
eX7KyA7iqpvjq0dd/cALNzlREkBOH3schgxYkjICUnrbPsBOhOmCooKBBNl2e8ZbF82XvmFXewgm
mZ4T+lWWJTgydtI1mqsb7picmyfBdgOZPDUH1/vVEhEOGCfHQzUzk4mQ/r4I2uvPlJTLaxPWW3ap
8YfeqIl4sIG9xlDZrFyHfg2gywuKdy/jXbe+NCnVdh/8ypEBl09Zmpc3dn7Q2XGPXyIDoM7/MDyN
1Bc0ZVxiFQJHpERLYAvNIYdr7XGNdRYC0bK1CXqR733EVGcCDoPVSBoAC2h8hMMF9QNcducQQog0
wEH4o4C64LmVrKGkZW7m2eFMOgePu7VwxwAK0PPEzxvx98GeguUYwS4+FbWVgFhr8H8z1mlwg9Iw
RWmcn5qynXggG5CKShq2B9O3MMzive49+8tNebekGCTBicjYMHLTr+fjODIOkU7CxWDTemTEg2Kt
wT0Wv1+wRSV6QZ3FI3fL5H9BmQ2O9q7gQjN/l+Mj5Zx9YQ3h0sBdck6z3WNjT9sbJCVsauqTeWed
S/3CeowLvEhp+fR2d1+B2+igzZ7TGCBdzHsbZdN+YIbFGLDrfLm4HteajCSFYhUVPnZkooYtd7fT
DCK1kouGkZ+pQs8ldQbq1BWqwD2JfuAuV8N50G9s1vsZ8paFhZhFFNlhtwUxjmOlBi/gCypcallL
DamWj2E3Y/CfHh9ezPrrQELdSsRZcQGwxDJHuYce5eWETKSrUDlE65ON/EEDWDCUCcF15/pX4vFV
8sYza1BXqnYyIgU9QmZqvpVVFuOHQi+XQpht2OB4XebbUxRV8Q==
`pragma protect end_protected
