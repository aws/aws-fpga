// =============================================================================
// Copyright 2016 Amazon.com, Inc. or its affiliates.
// All Rights Reserved Worldwide.
// Amazon Confidential information
// Restricted NDA Material
// =============================================================================

module top #(
                     parameter NUM_DDR = 4,
                     parameter NUM_HMC = 4,
                     parameter NUM_PCIE = 1,
                     parameter NUM_GTY = 4,
                     parameter NUM_I2C = 2,
                     parameter NUM_POWER = 4
                  )

   (

   //-------------------------------   
   // Free running 125MHz clock   
   //-------------------------------   
   input               CLK_125MHZ_P,
   input               CLK_125MHZ_N,

`ifdef SYS_MGT
   inout               SYSMON_SCL,
   inout               SYSMON_SDA,
`endif

    
   //------------------------
   // PCI Express
   //------------------------
`ifndef VU190
   output [15 : 0]     P3E_TXC_P,
   output [15 : 0]     P3E_TXC_N,
   input [15 : 0]      P3E_RXC_P,
   input [15 : 0]      P3E_RXC_N,
`else
   output [7 : 0]      P3E_TXC_P,
   output [7 : 0]      P3E_TXC_N,
   input [7 : 0]       P3E_RXC_P,
   input [7 : 0]       P3E_RXC_N,
`endif // !`ifdef VU190
    
   input               CLK_100M_PCIE0_DP,
   input               CLK_100M_PCIE0_DN,
    //input              CLK_100M_PCIE1_DP,
    //input              CLK_100M_PCIE1_DN,
   input               RST_FPGA_LS_N
                       
`ifndef NO_CL_DDR
    ,
   //----------------------
   // DDR
   //----------------------
// ------------------- DDR4 x72 RDIMM 2100 Interface A ----------------------------------
   input               CLK_300M_DIMM0_DP,
   input               CLK_300M_DIMM0_DN,
   output              M_A_ACT_N,
   output [16:0]       M_A_MA,
   output [1:0]        M_A_BA,
   output [1:0]        M_A_BG,
   output [0:0]        M_A_CKE,
   output [0:0]        M_A_ODT,
   output [0:0]        M_A_CS_N,
   output [0:0]        M_A_CLK_DN,
   output [0:0]        M_A_CLK_DP,
   output              RST_DIMM_A_N,
   output              M_A_PAR,
   inout [63:0]        M_A_DQ,
   inout [7:0]         M_A_ECC,
   inout [17:0]        M_A_DQS_DP,
   inout [17:0]        M_A_DQS_DN,

// ------------------- DDR4 x72 RDIMM 2100 Interface B ----------------------------------
   input               CLK_300M_DIMM1_DP,
   input               CLK_300M_DIMM1_DN,
   output              M_B_ACT_N,
   output [16:0]       M_B_MA,
   output [1:0]        M_B_BA,
   output [1:0]        M_B_BG,
   output [0:0]        M_B_CKE,
   output [0:0]        M_B_ODT,
   output [0:0]        M_B_CS_N,
   output [0:0]        M_B_CLK_DN,
   output [0:0]        M_B_CLK_DP,
   output              RST_DIMM_B_N,
   output              M_B_PAR,
   inout [63:0]        M_B_DQ,
   inout [7:0]         M_B_ECC,
   inout [17:0]        M_B_DQS_DP,
   inout [17:0]        M_B_DQS_DN
`endif

   ,
// ------------------- DDR4 x72 RDIMM 2100 Interface C ----------------------------------
   input               CLK_300M_DIMM2_DP,
   input               CLK_300M_DIMM2_DN,
   output              M_C_ACT_N,
   output [16:0]       M_C_MA,
   output [1:0]        M_C_BA,
   output [1:0]        M_C_BG,
   output [0:0]        M_C_CKE,
   output [0:0]        M_C_ODT,
   output [0:0]        M_C_CS_N,
   output [0:0]        M_C_CLK_DN,
   output [0:0]        M_C_CLK_DP,
   output              RST_DIMM_C_N,
   output              M_C_PAR,
   inout [63:0]        M_C_DQ,
   inout [7:0]         M_C_ECC,
   inout [17:0]        M_C_DQS_DP,
   inout [17:0]        M_C_DQS_DN

`ifndef NO_CL_DDR

   ,
// ------------------- DDR4 x72 RDIMM 2100 Interface D ----------------------------------
   input               CLK_300M_DIMM3_DP,
   input               CLK_300M_DIMM3_DN,
   output              M_D_ACT_N,
   output [16:0]       M_D_MA,
   output [1:0]        M_D_BA,
   output [1:0]        M_D_BG,
   output [0:0]        M_D_CKE,
   output [0:0]        M_D_ODT,
   output [0:0]        M_D_CS_N,
   output [0:0]        M_D_CLK_DN,
   output [0:0]        M_D_CLK_DP,
   output              RST_DIMM_D_N,
   output              M_D_PAR,
   inout [63:0]        M_D_DQ,
   inout [7:0]         M_D_ECC,
   inout [17:0]        M_D_DQS_DP,
   inout [17:0]        M_D_DQS_DN

  `ifndef VU190
   ,
   output   sh_RST_DIMM_A_N,
   output   sh_RST_DIMM_B_N,
   output   sh_RST_DIMM_D_N
  `endif
    
`endif //  `ifndef NO_CL_DDR
    
                       
    //-------------------------------   
    // HMC
    //-------------------------------   
    
`ifdef HMC_PRESENT
   ,
   input               dev01_refclk_p ,
   input               dev01_refclk_n ,
   input               dev23_refclk_p ,
   input               dev23_refclk_n ,
                               
   /* HMC0 interface */ 
   output wire         hmc0_dev_p_rst_n ,
   input wire          hmc0_rxps ,
   output wire         hmc0_txps ,
   output wire [7 : 0] hmc0_txp ,
   output wire [7 : 0] hmc0_txn ,
   input wire [7 : 0]  hmc0_rxp ,
   input wire [7 : 0]  hmc0_rxn ,

   /* HMC1 interface */ 
   output wire         hmc1_dev_p_rst_n ,
   input wire          hmc1_rxps ,
   output wire         hmc1_txps ,
   output wire [7 : 0] hmc1_txp ,
   output wire [7 : 0] hmc1_txn ,
   input wire [7 : 0]  hmc1_rxp ,
   input wire [7 : 0]  hmc1_rxn ,

   /* HMC2 interface */ 
   output wire         hmc2_dev_p_rst_n ,
   input wire          hmc2_rxps ,
   output wire         hmc2_txps ,
   output wire [7 : 0] hmc2_txp ,
   output wire [7 : 0] hmc2_txn ,
   input wire [7 : 0]  hmc2_rxp ,
   input wire [7 : 0]  hmc2_rxn ,

   /* HMC3 interface */ 
   output wire         hmc3_dev_p_rst_n ,
   input wire          hmc3_rxps ,
   output wire         hmc3_txps ,
   output wire [7 : 0] hmc3_txp ,
   output wire [7 : 0] hmc3_txn ,
   input wire [7 : 0]  hmc3_rxp ,
   input wire [7 : 0]  hmc3_rxn
                       
`endif //  `ifdef HMC_PRESENT
                       
//-------------------------------
// GTY
//-------------------------------

`ifdef AURORA
   ,
// ------------------- QSP28  Interface F -----------------------------------------
   input               CLK_QSFP28_P3_P,
   input               CLK_QSFP28_P3_N,
   input [3:0]         QSFP28_3_RXP,
   input [3:0]         QSFP28_3_RXN,
   output [3:0]        QSFP28_3_TXP,
   output [3:0]        QSFP28_3_TXN,
// ------------------- QSP28  Interface G -----------------------------------------
   input               CLK_QSFP28_P2_P,
   input               CLK_QSFP28_P2_N,
   input [3:0]         QSFP28_2_RXP,
   input [3:0]         QSFP28_2_RXN,
   output [3:0]        QSFP28_2_TXP,
   output [3:0]        QSFP28_2_TXN,
// ------------------- QSP28  Interface H -----------------------------------------
   input               CLK_QSFP28_P1_P,
   input               CLK_QSFP28_P1_N,
   input [3:0]         QSFP28_1_RXP,
   input [3:0]         QSFP28_1_RXN,
   output [3:0]        QSFP28_1_TXP,
   output [3:0]        QSFP28_1_TXN,
// ------------------- QSP28  Interface I -----------------------------------------
   input               CLK_QSFP28_P0_P,
   input               CLK_QSFP28_P0_N,
   input [3:0]         QSFP28_0_RXP,
   input [3:0]         QSFP28_0_RXN,
   output [3:0]        QSFP28_0_TXP,
   output [3:0]        QSFP28_0_TXN
                       
`endif //  `ifdef AURORA
                       
`ifdef I2C_SPI
    ,
   inout               I2C_FPGA_QSFP28_R_SCL, //FIXME need to hook up I2C
   inout               I2C_FPGA_QSFP28_R_SDA,
   inout               I2C_FPGA_MEM_R_SCL,
   inout               I2C_FPGA_MEM_R_SDA,
   input               SPI_UCTRL_SCK,
   output              SPI_UCTRL_MISO,
   input               SPI_UCTRL_MOSI,
   input               SPI_UCTRL_CS_N,
   output              FPGA_UCTRL_GPIO0
                       
`endif //  `ifdef I2C_SPI
    

   );


`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Wd+2kFjzXcoXxV7AjArBufrtM6IaZnr7RRnPpPPqPKOuMyuLAa7Nfw2cMgn+M9zETUHBaT1hT0Lh
HLcgs8mHELP/0MKCF9M/yFRVQjl2W1mSRMxXsbz+pUxu6END/aGNjRTo6UyK4OtzoBXW8Kjzc7jA
ZAzEZT+7QcgA4WoJuWseAkDNNKmtAtExOoqCJiOpK2O/LbZFLyLi00bGKZBNc9kydqlN6YyLH+gt
SmVedqoUjgcgqdpZw6lF0vbWbO/GS7+ozQOoVIkmvKaqS6ymwc/MZ3Hqi5IuWKxJ5X+ONDA556gL
brVMJHXjMDaaUW56ZuvRbS/XqBCX8gbvixrhyQ==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
o8rKZPIDht0nAxe4GSL9guH2gTnKET9ksWci1h0Q+1yJeP0gj+XXsoDjHHrLTUUtrdIGALbUK8+s
AiFCpyJKNEmcxIHB63lxJhpIK+Q7Gp11ZtiOL99JUlYWJMkQMDU2VDA91trJLuXmWSiRdd0rnyXk
9WZVi2xnFMctfWXMECo=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
aUo5qevXaKfnlN8wCdo9xoCE3co3Ir8KyjcFTIHgo1QkfYD6tVDOTvqX/VuvPS7VfiDa/1SmVBu/
XPS+n/3lGqw4XMJNPMmeKDD0Q9BmqQpt4pev+T+gQY1Dn5opDeoztPGWm+nklIOBUxdaOk2c1cMM
SMFV3eLbWJRRZZSexFI=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 39168)
`pragma protect data_block
pN4baJ+xHlF2CnyvI8kTTr+dMoGAvv5jTgNjhshvatOjkX1gu9sf/wL161ufcPLp7cdqM9zbN+M9
13YdWL5jXITKtpEKY1uAS6MKkcpO/V6BVHEG6r9s0MmoTQelpR+z0eIyaa1NCREvrF3tjidv1+bT
C3pGaa4pPIqZsJ8MIuaFsCQAUA0kqBegdESamSzEWAkxht+pr/ckZ2dnz+aZEGLUUx4liLA2hqDG
95ZtFmC0trVnH4y4gTp+AbfxUuRjjA1E66Y990xR2AcB3Pz05IJ/Ok2TZNHig9r2Tv0P6PaNV7Ux
jlDGCVCYBqLZY8RjTSc6Ho1FxEAzhgCtHBRwvA9+iamG33iAYd31e3HQisThOynorN6UMcWyfvFs
FyMyQ/vWLPrAe9Tvo/NqfCQDP1F3ysZOnqallU4akQKpDLxfM2tqJznZ+uc+CtZoXzAXjvs4XYMe
LDzE7vkmV1VL0TK0n+3bvjsQ+MAIzLiXjRtYr/VRMy4ewu2BNTjmF3huLTVksvxnsh1UfP2K0lrf
Eb54TJ1BDxI5WmvzerjRDCNvT3TZPEplnvK5O6Hc2dQZuR0y1pYVNZxins4BTogrWh6jXxuzYXLN
eAfHt+hYlitZkXqPRlONfKaCABAQDgF8czJP7TtSoyl8WGWZmtKZYDgIDEU9xoEol2KaOcfurN5R
3IbsJWUeSDDdugXYWCSt0TCM3+cvo682Z8Ig1xdeOYZtK0T6LctiPTO352sFKlrSHWELTIexUzOs
Pjeto2VQ8fnqMvDxr7kTUAyci95oO7NbQUIoZnX/wAhGgZQNot5mOtnWNLsstEjCokcSDcx2TY74
/2aVONGFZLxkjq4/uyQ1NRY8q8buvRkkh9mSDFxThphaCyW/iJ6wbKXSLcyvmyfRmGTJLt6M50rk
1BEPmlb2dZroZaWuS08ZVhImTNKGpfpkrEo0vtJUA35t+t8DFllDhi7bFze/KKe2xH6vUgE5O+tI
aa0q9uhoHj/h4R/LXbf/bSVzw7zofioGlHMXfY78sVgRuCAH3LwqDmi329kWlCe5kJuQtE2o0JYB
ItK62Duh5D93Zotx7gmxx3zBDkfPphSmPUteP8KVLSL0J339PgFy7pDIWqEgGy6U7vmHQ1C4vPCB
9T55H9cLPXgHJi8pZNrx0JxtDlQVv8FgdlUWylBaDWsCRoQ/G9RFF58vJyB7mQXYi+xGf+w+5Dsj
iZUMVrTCqyLr/g6CWrE47nWp8Z5ppGZv0JIozL6Xr49VtbsPhfk9LhkXvyaj/3ng6oYJgaVbDOkW
VNZCzMBkNqhFUTdyXu21QDCloSIeBmlzGMdrxPwoXp0oXqApaIzKqvmXWxNfmM4REtS6w3PFuMe7
mOQfmc9ElgSYJK9pmWkBgENjRLfbLUGXL/c/lMt3MrNk+6oASI4gyHcOlOKUNFbXOdF9HH+uBM3S
k1vPhlm+N8iOANlzo5tHMXqN0dkvahDNBHfOMp0AByi3ENg6RxUAD7mmcaQvsu49ykiHchCJSOsP
XIzV7J+a/vULh6x+zY8KzXSGs6HUXLu3kuZCCHL6j0SJSa5B1jCbKnx3xrZ/hCIQ6FZxqSrz2bN5
E+sWzy83NW7sLe4/r6cE4IvWEeIxRfrX782UflcnMSu9ld++4VMcTxJnm/MEd0VpLdqKDsyHL+FI
N8FDaUcE2BaaLChvjq9TDneqSmsLrgNYdsEddEVazaNFD/FoMC7KEvqnlMZ+ihvzXeYwRdJGGMY0
dtEpa0zh+J8k0n+6r5qdyvlb8oopLXTbkIBM8QBdgKmlL6K3JBodjAhxcnm7nSmNLYdcqizYVGOi
4MI4RI17jWaRC0K70vGS0ifbh2JE4fMJK0bgwKDp5vE74fmdcwoapKs8yPwjE6J4JMTMpytQXZKP
S5QGqGHaz50thdQcd+YvALph9T0RBhenxNRUu7vtmgFQGhLUwA26lY2QFhQlXLR8SAp74OkQJwiz
6WrQkaN1TsKpga9pFJc6KbVYRA4XRgC4gKmdBGzGXjlV46eVf0GjEqKNrMCH6oxvMhQiA138otUY
WGArUdKfipyplbbXshc9u4j5qBFrcASX0hsOzdQaXcvrjFJFyvT/eihMsOUb68mnLzdDHdImNe9C
Iu07GoVPN0zdxNR2/n4PAOU5oZLjWcJKJS8HC872fAgpNYBhnIbU911/pysLiN+Wu1OdbSz9u7Yi
T3+2GZYlRlZvB2puo/STYqHrgyOeA6OB3JLtcndgD9hMPsjxL4X6iRYar/ZA0sKRImY6ZHM7ypDV
I1C2B1wa9z6zYkuaXCJpFsc+/k1gQ3P0188G/5G+4HE1Qm/vLVbHsBX/8/TD4BwMXVuajAmNc1dU
XQr1yUiWO3SG81iz5GrjVVhD2OO752PX9QahFInWO3jn52IyqrBh4HbiS0mtnIJCNDpam16hddiF
6VSNc1O/TcCpIo5/7tX3CAsDO5ie32Fmto5u1Jd2Om4m36F2LG+A/Qr6z8VaeLFzlmzkAsLTKoLw
lc5cdohMdjETEeR9spYMcxPFcauWI6BLS2047huWELT7y7ucIG7PMdm5yVV2+hPUV5Zigl5GNWjI
McX48zX4X7GVrCuzTdfZxf6lGrcDI2424NbqxCXtSidkRrKHzF4CjlxeS7e6IsnfQOjMEOarACSl
5m+FQPx1yuUG6/7x1Q9XUeeS7UcIAgNm290ckDmOsEqDuyS9RJviBcC+1DbY/YqSoHP+bx9D/6ze
/I0qBus8tXsherFY78V/etlxzT+Vwkk6x7cyvce6UZB+ke2Qinz/037kb6FSDlVgKiHBd7GAgnrY
wlC+Yj72GexBWj7D8XDeEQuzJUTzuKJA2+KLB/G2zWq0/V0RIn20+Lgda6ljqfbc5zKd4wIZs0hd
aqcxjp6QAlUIRhxFdjIMzyBWd8uiy1ZwX6wF2JzaQcF2O5gN/L4mWEGFcpuCxzCrpPLQvlC/SCsV
PCbMc6fhLbi2mL9EHPEoMlDr7NSE7fni+MUg0fzAbOlgWNSC+yoKU5qluZzf2SDNKjMEain8JL1Q
EjPFfdHjhlXXtt26R88qxlI429aL2rdGZrIt4iBbk4mfDBjmLjBi2l2rcHQOJe7zp7cfDb1oWmx0
8txkAMC8Z6+u0Vfq4yUO3IXMCb6NiWFwBmlgtpZKxA1Kxj5qgHCgqPR9havWJx+jKKM1Pppdq2mR
xG4YT4CYREYfVGNWw7hsVu+DF1t+Ck299NAE9dre4t311jErCuxfrzzcAANfV4kKTDfa0XKz3Yny
0Q9FZhW8bK74SpeOGYPtcd4/lu97GwIeKP9SIVh1a73/5/uhjddapzldWIkAq7G025HZf8AwfFzr
i6PamWUjWDYqyd5Z0qNWow33rYOzUIDDjXf2kpXRAPdE+medUAGfgOV5nt8K8qT/ysRpbZG6LbLB
TRGXLA6Y93X8AODN4lrbjsZ7u6KeXec5LRk7JLprs7gLfw4oCP0tIQVF9AUW/McoqBEqqeGELFOQ
IpOVq4u5xN4fRmvJLmoizYnusyZRsom75vl/BMH8Ig2J4h13N5/6LHlNv0y1W/HcglkfTpaqdDpo
SKLL4NqL/lxmfQJ0GzNY0YqEKFW84FExvpLOlJg4tl2XAOsnxEXjLRcnuyIWmzohk9YFt3DgpwIw
usQ4DPAXqtl0osbfdnSk12uoLpn9JllGLojXEYNJtLmTIlFjqMQvTxE41lXaedcGR/S3UtOqDwzB
t1IDd1l50Z7cWyNpOnbV5XkUuGzRsP4iG7pGRiHy23g+VZ+rmLzKO+/Vd5EiarFfqK/GtdYEmSUk
05OX9yioUYkJRSVCUW4wdsw7xFewKiA7DOe1nvQ3VU6x8WCjDwjiSyytN9C1/6vvGWm9TxmjUOu/
adb99pdNeksH0gMU+d9oN4lNSRJpnjbqCsil9hMF4WxE64PgGvH7LYd+aE82dO8JPfcpxPY93dVA
m2P85movbO+qQzV24wQRgwEzxRgkqSg3NuwkMOANXV87RisSyaMoE7AyAT9jTaGwYDBSWpIH3S61
/eMqvSK92/GFsFTQDAZ0iSD+NNzjoZ2HI4rUDg4P1hMGLDPLuUvW0ZT9iTZMIg7O+afXFONudKj7
JnLl0jcLvgmeM1sRqwZyBf9b8uwZkkOj+ogufA/MnlpsUuSQ/C9kptoCGNMg2d6XOUtxZB21kGzZ
vDHoj+Cdmmhmocczvn7E8+szCPvawjwXlRUEbioxX+O6pTJlzPs6f0GdoOFyTMCNzHmrNuXVzaDW
l7pcbfZCpAWcToULhQe6MgU1lHTyOKNSNXcK4uIbtjlYUsSirHhkjkI+3kZS2qA2lT62xV4P3PI4
TnWjOjkB1n0E0eQ2jDD+NSnuviHE8zkwh8MSUL1UKgHpX9+vOqzxrXjJ/4sKlzZy5mbwR5+P4QKo
/yXZCaETlY0qq0OJNhTYRjacByVAd6kmJ9n6AUdqTCkcTaa9rOyhzrCF7JGLOL65oGj6N+3pDwgo
xaR1P4fUNGzthpefqPSAsD5qC7Kpqfjo/mf7SvZZ74suwe9im/hSW+f/6ktZvt+n7ECSTA6IJlhn
ADlL2tp8dmNUD5RE7YNIgMf+uaxXrxPWuajCskrqBHZ8XlDUAsMiJey5pLxDY4XHKF5el7Z2Uauh
gcCUVKsoKR9ougKbOFlvU0r4NLan2uEZfTV8b5Jr6yQMna1Y3hKhkvP63dA8Zuc0PeDFk7Ad78FF
pu2jnyrdA04P3l2OnCKbzOZlkwbdoslF8JqPMqeer/lrNq6pQKaMpID73NwW+hMdmD8avlOAd22R
Ezc29rJGEdbG5zM7eXq6w98SZMIoloATcqAcrj9qnobqGhnA0EbPRP6X68qqITpVAXETQek/wNzf
dm08znFWvSFdArfqpAXvi1Qt7O/fdUIIcfkaBwOZj30cBfk4SQsz69+KVspDW20dg1jdBiCVtB9G
x8CL2XqHtTHvEDvGXmT1E13H5RFyC6bfrvuABTYt28BRfjuJx+dk6gIGBtw2ziNawZKqyjP32DPn
vCgdE5AcJQKCmc4xiroDRm+NO4xiYg298WKR5IG+FyX4W620qMYZHO1NPxL5+n5ybQvqdxHM855J
Pel2WtKS0xX07OemRL4UGwpHOccg5vE4wSJKaXwXN4F6lEJCo5OHP/9f458Nms2DKx73lSCeuKc9
TGz/tT2hK8CH81ckUqaJ3POa0N/kI/asGYrZT8CcQouqf+WO7YXPt1b3TIN2d7CdmGmAg8mwx7/x
vazDR5H3MyvkBfIoc3bBCyoOQG7IWTZ9vv/9zNFUVCp7oC36UM5Cwl3uyQAnNE7QrmUfpoAuQyA4
BFvPhMSNNd48ilKsDdbMuSV0W+0v0mh3i+5GJnFsBQ7rMNQC0E2FXdQGAu75do2Vfe/CpGXW/Kcn
N0A/P544J/drxuUxXsFeOJl9jkfIweIdZLzZ4ScpCPobMNPPguVLvt9KLL4FGaxGxwhAueKMGnp1
scmSN1yFTxhn5lGduj+rhY8ZfIFeXe7cahru4Cv6emzcLl99VMESnMNpxSGRuHGlEwATriX08BZH
ygoS9fxK92+wU4L+gLEBuOl5ZUb9eAOASbPoObu+2p0Z37KiOg55i65TeSk/wdF6uYb5GT5CRkJM
LoLbiIIuLcEAfELm0U1W3gMj3aISEI4sH9Pwa682itQ/MxS8bvbpc8MF5D51/+8Aj62zEddc/H9/
sxhUrTx1aukwaqjHvRVId0lsGZhrtqBcAB+VCiRP3UCW02Rdt2/h2xvVtTFc0wWTsuqSjFNgt1Ls
m9ifRoMafYsr73liduqjIIP04Iatt40Na1ZLE31f6BqLFx7LxsxoJzhkKr6pWjL8l0MVnDwgaqXg
kM/dWqCC6xpoeYpIgTwgirVhDjQRu/UatEAIlcovjES4SU/LCrIMiQRqlz8H0B9okqLLLl23Kb9b
Oped82t2RaygGXEckpOCbJzBEMFx+5HZQWk0Gj+OrQJcA/sO5ROli/Uv0Bo9lQgTZ8445nFi2kux
zsU6kHMtJxLfJovG1CyCc2L88pnA1nk3af/oXOqdDA07p80GcaSW5C/B6WDfkwpib8Y/iKx+ElWk
vb874l9cGdb/PVwh9oF1bYM4LgCi7WO9mf1KFW9HyPIC+VYSDM89+icI9F0JToQXCjXx5bAD2M9l
hskzui9B6QGJkbvYbk7EIbdU2/b07A+a6wlZQLVrWNaPr1WEBKZl2GZBcVnD2A+b+BOnnIRLEhky
zTvjMpcxjze3WH+NFDfoAzQ04SFvncTbzyGFnvSclpCTjcBpXdGnmR+WRco9bkossQ6LoR83T5sZ
jb6qgyYTxIAIxMJp1dJHxWSHdtJlVi8hSBBYCnPGvOoLfYEoSPNX/Ibaanmy2bG82y0OqGJQhGCu
H7xY0oW9/h/HhSUkFJCpqKi9uA78usxEbOt8Nm24dzpJeDmXAmizhNrYcWQvo6eH1nIsV+WMLk4d
EZqpm34SJwa5att5dWfeLf77wQCQ/JMmlOucO/Or3guRpNR/o/oCPc3hFOLdsiB0c41qPRePxEE0
Phqa0A+mRdRXLp3Y+rhxp6rYBwktFjEJZ1nIEOXnatqwhMOLNxpV0itPDxnQRruLIYymWvNV5otH
m0LFCTM1+hlvMyw/X3Q12l9CwWXjlvoAd/+muOka1lryqABMMNNv0L60U+f/hi/CgP6Sa5mlIsz9
0/5VMa7/2QWtHAUWuEgfvxEjDtzIoCP4SHG8QpxflxYELGCBLdFajw9Kp0dVptifVyQxK6LFay3z
bFi0ZaPPUBZJnNXYT6XDQERBAYr1FFIK1SuOaNd1llMjf1Ig11/fF6+aa1bR1vQ0b8c3XAoUQXQ0
DXsWG0H9Xp2VI3C6oDqMKZo3ZDeQMdwCW1FcrX2VZVLMDnT3HWg7LiPA6eIgNeU/6RqMLMSuhNhb
R5rlO07eFARJYSpuBad9L0pbnYe+2+yKgJknkpUVZzrQH+P4NrN5kkl42hNpnBwhsJPNejWoZFL9
9K4BYTccVzUn+aPNU2soelcAGV2rV2sYe8UmNjwmp5moghdvPoBkNKgsPtw71K8CFC2xdn4dI8DO
zY+MGu+uj6jhMSiLlwFGtnY3JYXBVNktUbXR/IdUjAW5zmaTr3d0XPWQaBeBTm3KbuxugDAs13vQ
sTR9+omnhnkLnHRFzAooLPNIWv4c5I35IMoIOESFsG6eMNkIyEwBs0StgHffa70FqQSwqkzrnKZ/
A7vAKZXIrhz32XCZ9Sk0pXx2QIuHmaCJKwjSWqtx/Wv9c0pcY2EwzEjfVGzafgN58DXS4gWkdby7
Yhla2PLweVzWHRLnmitSnrXu9to05DmdXlAjQfw/5LaBNt7hF26FQLQ0MRL3NEsARlz72fsjNF7Y
8TFZuIP/ydaZsOleqzMArVYm1+nGSgGI4m+5VhRIA8E1f16AxysZXVv6LUHF3qayodsTnHqaWkfk
iHJy2El6iyCPHWLTq9qS3rLFZ5HWsGBC5JqLckmWqsd24EbpmOS6zxOPt3r8jLMtajutMmzBp/8n
pT9JOkUKHzkKWqJyUqtPrHJidAAZAhrm9UvlGyl7SsMjzbmu77wKqBY7Buv2uT8xk1CAt0Bgixw4
QTLdPw4z7AoS2fwE6QdA2v1E9sdYTjDBkGnDY1+Jk7jLWscGldowmkM5waR8vbzt/pJQvQNOwN5p
v3rZulzzTc2ggb/dU6HMIjG79LmP/qVxgpxtHOWu6CE+2y/Q8qHIeCcoZF2tngFcKNd7dRHxc0Cm
WPTDunb8JglTp1T7yPtnmEGQROfQSqSzo79zm4ED86i+XxB8b8j7fSdy4xgims0MaCPy4cYuRhuJ
0CdWAJEEQX0vFKMaz+M4hHI2fhYPIqlSmmqa3N26uB64oAYOTzJd0tutA4v9HA8LoUcJHB8lIjya
aTyVaDO7Q43nrUlGWNzZaKM9ETazD9O0D73oojwIbrf729zmqbRnmnBdn6pBpsxtaV23e5wN2VXp
Lh60LihEzswwnkFydea7nigfdNUF6LQs3BEtWFLIFViwnJalSvE0BFjsosf7CCrcj6m7vRICgWdR
DWvSTdWC2xO0ze2AJuAE9k8SjJC6zbF93mdKrPUQ0re2gZ0luTwBJ/sYHEdBdE2QxU7uqASRFRDK
If5vTOgnFFaGYIa4DqLFbdeu6zNQctuIPYurHW8p+RzS3x3t7RVHRuPB2MHn/RaXFDdewwcW2eMD
DfKYm1nwZ0Rf+sq7ZxxJH/6RJJEC5hYtFa5QCl8/zszYGtWnkp+fsqWsiLu3KSP7qt5tYQWtM3sS
ZWx22J2z4YIjAZPcjGi3OwSZpaisYbDYZ5pob7kf/1UZ6/G7t2cYHB4CkH/vXzCjQkM46yfaAFJy
jKo1kiYvKtlfTNAbezKLATHOnAo+caIfVXTpbpzBySq870ShzCj/PjSeyhJzSs7QVTvH7KZd+7p5
jCz4c/roJ9uQcUaAPOIOxfF8JH5259bkrUO7LI9SBRgMOIN9CvJXULg7D5LRCL1lS4T3QHPrtqf0
ue0WLLb6YTRdDvfoVR5JYTfY/XV98Vt2oovpEjfKRjUrVDPREpmkQVrI6tkBa4mWPLaNa+BUDUUR
Vj5ihnYTwmvVYG1wWSWIsfe9Y5y3QNmV/lLeLrIpODnpZRHWBc3UZdlaZGkiIus9HK9rcj/k6z1z
DGGXD1kqBfORwrm1/uM22WnoOMmhKWJlzFslgcdUJwGSJScjRDRax//XmCez0Jmw2DcHxfOdzA0O
z10pSeyxnZvRvgds0Gj8RJnXTH8FbIIznSqv5BGqQ/2vMvNtAXXF6MOubAv3xhCw3+bVxEMECSVU
JTLa8JqjSZFHbf0kyUvtBhwHeRs7tmEGyvnN2bZGYvghQwM3JR67aC4ouSNfmlHom2JhoFm+q9/v
qrF25CF1eKWLsSid8JfW4N1gLAsfeBsSDco5ORsq+H/0UYJFDhiyDzAXMujZ0cYFvkUNJh7aieeO
R/69TIBqwiAShRdsCifckU3NMEqmVFmZFC9xaKSxhDlH5OFwq1SzjUi/o7kh0ojIvTuEbZnA09zu
yfhdxPSrLa2tJUA3H7SO3vco32RL/Jp2SOtlabATRKCcBJf58+1nSEpkE6vTAQkb/Qg0ZRskXquB
wPqRI6N4sSpFhmNkU+TOcUFoaO5tX/R3bWUd5QtwNLanlP0wWWyWzWGOSWqHVzT+v/TLxJhSVc30
UM7kVFS6TUyytSxqiNkayiwTrYZJhmV4I3JaNWJS049l1yVzqoHZMDkWKQ0qA4FE/7tp1OiXoz6l
2b3Y/9EaCkMWJvJ5krzwfPEz3d3kPuV2D2hSNhb7XmSW96ghrZkTsItQgH/d18wi16ABdVOWd+jF
R3yOqkLVHjYRUl1xV7jri07iOQHlFGYuSPoX+JGI4S/LZThgFZSSGHCiRvDtRw6aSYd1FflVMAgK
6tdD/bP5hJwCq+1l88Z3NBY2Ws8Uec/2ho1o45/kt8e688RwdOPj+aPLQLFscVtwPqeRbnyiC5Yz
30k88O/y6RzUaDNug0ym8OTx13Vz391k1QHpth0XKFDB6RXnGIDSkIesqKrpJNWUOKkFNSbSC9IF
14M1SwOBTdgvz7u4Xh2OCIdMFw8NmW2QRcRa8k5EQAL2svH42Dw7GTKoExoAw1wFXJrTGLIiPds9
bzaO8qWLgPtsFYuKnFvMe2adx4oY8eOhpj8uiQeYNPUlfpo4dqILgVOB5WV3W+ls3L0nqcyjebJK
MUAMzNbX3J7KufP3xkzutcFNHZluu/hpBTYJ0bAUHmu4RxylCGP+PBzcOS6ICT6lqLBvcq392Oxa
cMnkgNywHPahEHWqM7NWiUPwbtuG+4xHGoaYoG7eR5Ipd4ZdNoyF4y9oN8QR5Sm+iXK4kYdu+7+l
Pq9TJIGgOzFkN3d97bfUrr8LLhlu8iJjRcObTm3556Ok799b7MxQEDm1cZkxMWTkHsjz+E0r9A5S
lhBv7knq8r/a2WfMtbUIii1XpPAasCz8auh+tXwsdT0VwHlD3QCvlL3mHckwwtjwoPGlNVvQZSYp
bjBDf2EgGsU0/fssJtkCmnHsWu/gRtF/h1NiVtuo/53VIUTXwLmvgmhhuNVYHVPMCFx4ORcnCU1D
JFgdRnjuExqo+qzwq1VLLZd/3f2JyG+JQReS7kIhmYtJyzK++dRx5NMuT3VKRpzreCFhyEkOgjvK
Nselty2LO/cZ8ucbfJAYgN8xrdIblkj6pDbRuMf2vfE9Qx7lHAC+VOgx4omXeUGNELK3LZxzcIqx
6URSvBXAEr2n03oChiziFzYZvS3GMJXYLReLVKo0a5jfiYrS/zwDZ4vGqlocKYQ4rultb1bypOrh
Be3WKTpUzANbgea4SE1qQz0SeRveON8ezyCLy2cc/RR5PtJ6Q3J2cn3Xf9gEqth1LkDMxMS0tbMP
3Wp1DSRm0qKpPb7gMYD33Txt/RKBIb+rP5lQn7yLMm09U+Zx/0Qv1pXZ/I9OxoheLefCnxdkB2ux
LWnMhPJ2SfZGC4Y8I7cgWk7gVT9e8+ifTCTkEfqEEVghHcloFzakA15JNb+1Devo1cqTviZdHQCS
aJAKyvBEZuDd1gqolZEZVPMHDEpeb9OfvFUHU7ynTyn4ovWI7hu16febtrEH/roDMlEfCYquWRXn
5Gua618iDDL7sWd2TZrnTrWZNlgIXyv6zR591P7NBH/ckYhJwjwvsdeq7sO4n6gMUk5rl7MXRKcy
3mFEqxIacaYOAFgWpvmv6N4PToN6bIHuuueCvPtvW/QlB3a31g+/iAiXCesF40hibMui8zeDivL7
xBzPNPrauWX8I44W8cljndZdDfpJUy1XtuwEh7wPAjPzoHwlnbNHR2LQuLMhJZxAg1brP9O9vGGS
IxPD6Tt7Gn4xGh8jpy1OxiqtY9W2R6AKkR9r8DiZ+rsSyKUGYJPfrbaDGr3H8PhDZ8Q1jCNLPw23
PgrSsZ7lxOKMMhddSQ/Lrdf0KngCywT356Z+cffFg10NnvZOQAEKgIYEQAawRoKt1IUrCnAOkuTp
X/bVXVaw/bYxABtjNVzyGdiRwsNAXacmQLMDlA0zcv10ZX6PGpsxawjaSk/MCY3+Y5783aVOAVG9
ei1eGeGiOIKGX1y8SQqq3brTTqVIbnXgqesGOBu/Oe9Hq4G/ZmFO7Ey+BQ36yY3KJV+yQcW4xB9D
2FByRXWO97IX9VZ8ucj3YaHhw7ZNsCxrbJgtVTy61D5+nIaVpJAVjleYBvggX6TwsMT6r2FN1WHK
hXg5wXEflyG0S7h0336ZXHEJdVJ0AF+eoOLDACl68Wns6poq+4xCRi0uEbLBvTpvmWYiEcWVho0s
RH6OaUmXgwneCfECCvcRiAA63zQbqoJI5R60mwiG4qlU4sB+NzXbUY5CtmnruvJy3Rrbbe6evaDi
21d67xVb+Q5j3dMl8LF+GoCIQSIZI+yI5As/ATyTZ+6CyAntM8VuFqj9YwzeoM7aUsIilg/0g99f
Bemn1tUrXwx7qPBnmC9YyySswd82fGe5x8hts9Kr8v5dMLJHflvq2cclYz/NbopIHpTSEQ0lXQJH
QyszdyrajGF8wATvgz64xCDWu5N0AfpJyfmrl8dNb972znhZabdh5etWbN9QTRCnSNlYxMJUD7Hk
1P9k9ftGBgMx1GWBJXWwkSVr3K8NWexveo5x0lj/ZQcKjrYXmTjJ8F+IDSNsqvcQ2fU22D6CGYWf
jmKQmTQ1AJcQJGLsoS9K5PSGlNqJJwt7juM0FQ2gzYvZucghdFgnByY6Vkwr59Mf181H0ob4xMPC
p/7O06FxvV+lljCBh9GEDfl2hKWqZuBbXfo6VC5fKtL/q7cKsWMKd4hJ9hBEq028/2fuK+G+EzIb
pr7HqJVGh8JAofHKb0TUgTm6L/yHLTUkES6Biru+yR+A41uDGy/QQ/b23MToWwQowSHLDlTD5VNQ
y72KnLnZ3mdIMx00lLsrs2jwWG28o8hJYoY3bYXjbdbTdo59a55KAEzHdIIjDrN4zzSo9G5vuv6G
dDyQ4SOoDXLOebeKZ7vJON5NlTFWQOabW885M2Z5F/zLqiKW1Q54AWp885xIGU+mhN0YXrQUvXnB
kmnUX4/boCdVgGPqfPX7V/jn9qWfvUL7787iGHlazaaBgykhP3VuOFQekoGaaKzWPZwr5b3XTINY
5GBoWsrOqnwcks+7JfNKPyTGcFV88vZftDzcCFyRNb0Y15Q+MrG2ZGjXa6CksK80UfFk/oIJfpQ5
/6YEtYRd/eEXTslgNxhfeFp7j8/C+VI420Xy6fK095ekGsvjduNeWLc0KyTL++LaOlLVTf0K8lfq
pP9vdlSZifGnZqZN9j+wYaufrP45Va+Key46HnmDtLW4fp8xJu9t6bG02LuamOYuJKRMMcALJBBl
jg1d5tHLjuI3uEsJtI+mzYIo/PpEHa+EqTddjoGiKOOuhQOOlI18Ro2FBgFivMYxDQo1aCKKv+32
/Vc7J7K4tF8zgzBWuiM6sUEojAk9ClVy6vMbKSogX9K4YwGOZub/ecniIVndD3CmQ3nHIR2llxot
DngSaWDkine5CHravgM8CECrshFKgd0RSWjYPijoKBRigpPkZqmvrRFvCPbesycHMBPaNqqqb2Mv
Q/0vzT+2A5V+m/926VYeu77ih1ppitNfBq410NiMDb7wE/UEfwSf3377hj2bsiBU16Ti3KHl4WcO
yF7W/5oR8qXv+auK9l1p/pi5fsZsoLe7gkhTq1iX/alyy5OPd1Wev/4VRzqa2nYNmZBKO33YHhtw
g1ydYYoZ787eWDFPqyuDJtNbGzT+OjJfA2laabK/MsjWhMK52BIm/vEKbQKTmnkoSXwHHXQBuRnN
W9PE7A5APls/kUZhlRW/gJ04VUgK76kdVpArDD0FEh6alCzSVmUHuEJYDGQv4fjQJ0wKZFtnvU50
5wpLUJtzx+uTualZAxlMkm1ZT6MfOH+5OFPuz73E7lUGikl8e8YA1W6aXoULp10G7npemn9gJbDX
6Om60s37qCI9MtWAKSEZxENKVIvsdQqLM6UDiF8wDFccvA3WgvA7D8f+QbYkDOrAvinMldzXUO75
Jhg1X7Sz8wT05jV/9071KXKUCQBgdtAYvqoA233YUb34y+RlBa3WZ9OQlegfJPNQ9i4a1bDKMR3b
X3LvSgj9XhIJr5g53AMqpAV/vJ5nOEvAfl+Krj5giwUW9NM+s6IyFwLEtBtumDKGey/prbo5XzmO
7kWigyesu+TzxJ3SlEo3oP5uqjRx6NH0gwKw8ldI4WXCa+LN539mPulx6fcaqvdYLZrGnagr2v+c
JM/0/9wwnKoxYqTnyhf+cIWesxWEvRa/VrGNV+U4FeEH2BsrTSo8dZ4ilE4PxhxQ/m+3p18tYLl7
v8Cfye+FKjIRwc+e2t8hbh0JFVKQNgqBFN9YjtryQJy2ybDN9xS1GfKkwJBcY95eXIDi6JYBiQ8N
RreSok/pXZF362M1GsG+5GYZNYvdWtdtzibB5AsvpEqvclY8krF33E+wKKXGQwrlUwrGfSQvRoxi
YVPf3cCsbpPpLsX870verBWOqZF1WsyqCzAz4doY6sSJntEB9PdmrnYgVRgWg3uwmTzCkgATFS1x
Yc2/KvhvXPkhPM9FzLxb3CbH+DMQOGz34D/DctMNLP2Fjpps98Yz15PxFTneR2XkUV+ACjuFKeaH
pUYaQeSaHwOU2Wxm9nMQASCmKGCRVHmApY8jS+p+ssAY1Llz5GrINSqDN1Qp8Gu63cr58Q5lwdnV
RDJNZx7xkvzduTLJ7kZz+oYerdwLQD7+UVKFvLOHlYgFyM1G9kkWdqekG4bPJ1SEyUZ/j7abGYLw
hsRbAThbK4gXlfWc2QnuoflaRht62vdEFTt/oCTZ2PLUyFIdBiOYdJWyPS/wI33eDQPShNyYZzj5
kHPIdoh4fdPDyBrS14eIPbS8hDfgzzyRYztPI8CPRxX2UK/6ZIKYGR+nVzO+3kn6gkh3OVj9lRYB
NvsF92v+t63/7dHDZGiH/NrtCD5fOyedg2Llc6OHJQWh3VCvrheNkQ33Nk3HNzFX/uw9rQiX2wkm
Opfwj0hX91OKrQdPndjGP+2A19XpvYaV/mtdU92BZayKazS1btNfaUh+RkqA2y7HlXhH2fdFBSfU
gJwS2u6fZsuN/TBzqh4tVbI/tbwYJzxVHhYM03JDaL2OAVYytHD7G0vNI4/+M2VaSEXeoMfgvYqM
rg7gyrYunu9LNbCbkjn/AsnkWDJ+Mq6SoZxzK1jEvK08VXakPA0wG62M3vWemDXVdxliIqFX5eAm
7CP1ZakKTCX/qJN+JH2H1by5lGPWCP+5oxlpJFuVdQYyunBlJ6nXCYIEFU5Rpve0BNUXYLmvX+LP
u9nSQOvOs7lAMKHnNDuaJuOX/bHNKplX58IPzkJOPxlvpV36z/jwECpIJ7uKDkn9a1tCiKZCwVNd
DYM+FGgS8PtA6epYTWoNjLa7NvY2w3ZY1UHYmrTxMBufWUbRPSCeav16WSD3coyI9YtZq2riexZa
ArVwfu2wkI/A5fe8gBkRz6w6b0t86JrIMYS8TaCKEAvw6V9jOlnGIml6szmf+zy2ZOLr6Q8WQ/zc
bmmOIL0t5Vgf4k8EOHdBlaDVtJHB2ufxT3BiEPKaR8pFxCqHzUWCDle+4gCBE9kPzKlmX5aisk3d
kIZRE1IOunUOiaFrAYwz8bLrxF2nDUwhZKsm9xjoUBqE+Hda7W5Zyr1/rdziITxjXK1UJKFKX2k9
9o7ynyEn55QRy2/6eoGqJjSmqQPYlShz+u65tYC/XyJKmrHP3+CrNGHj9/I0gqdLUx0P4ler2ICy
SaQkxFVgO7ycnS4Uj4cAWUDD8btytJdWfuzAkcBQnT26CBlMXTYuTHnhwRc0WTPUN9+L/b6VJtCm
1aPafYR35gZxr51a9DLYvGGTnsZgm1OsRo+gsZ3GG1kh1DSYGeeqyOq1lQ+9UgjakPCO6m7e6oSM
qZ4IX3/tpTC09sly3jX3YLeE+e6QFaFbEiMOrQViDkD2KHU4+9kwy202siDYGnj0UOnoCO25bdsO
Zy3TzyCECtnBs2yddk26hIEgep2qBsjFHUUjvlXm7KDd3vwM6GjOQY4U0LHtBlOqvQeOpcbMPCpp
qgDz+uNavNnt4x4hP/Rgb2uRrbp9IMW0ZkCiZ36PzsZ+lL2MXdfK76IohRJPBOxDcnZabvzEESqW
lTIFkdCSJuIcic6bAIcsyuOTYBgcDsjVQlEQjOAdjfF+cwd55xD4UrlerxRx2J+bCrD/JT5K7eAC
6khB4jqZ4bfQ+yKOAHrS6qYIisQsMj3aNrociq9W5zLBamGRXpy0ukOhwXbxS+dmpnwLW/9Xf1Es
TZt1GiQvJvUL89iPRUiAod9UErMtk0+ccc8pohuV+2f+e5GXl39WVV5Jrp/UIMHrQ8/au8eoYcGP
W4343evIxjR7wV+pidLsHVaIpZt1xgJBTmAa7MMudeSVDgJbiCqD+ps7rrCgX3SJj8+KgOeMiVCA
eD+WF/nzDOmPNe8ROy486BgEcF5ENjbHk3+MTmTMwCPAFxyZKYAQ9bOo5NV8ohL4C/Y2Hsgjsv7Y
3iM1tKaH8IMa3efEQCkVObSyDQoSlq4RVAyeinotuvO9BDee5sBlqI1XAYQPn9Hs2aadQAECvXAz
i9ge8OOcI2Ua9kLK6F9sNKX86V0HSaARPSdOn/iAXQYozMUCmM2Qaiby0BWeT5X6YV6EsM93fKwG
GVG7LYitxGdEuEijOPUYHJsPgeLZXY9urKxvZN6djqoQtBy9UilzfkOYQxZGtNAsg1wJtyF342eW
KtAlW7AvMTMP7vnzU2hYLcPvA6U1rJDuUHcUfWYl1tWR+9qx/ldu1QY3QSikzpd04bMKRTC8IPMG
aFbTayVWGsH5I78jhElZSMdRyD28pv4qRcyCgjojbFhMUIv7WCvK1VgyJrSq2JjIj7a40IsbgaVu
jaycc307gthl0RukoC2PVAHI8KDDLwC5guCpTFC7EUY8DGmTgz+xckARkSSxv4N6DlIr1aymLquO
wGJYIZMuyiqYICETgluL0H57fyWe+AIiaEI2imAzoQleB1LFY9T7EuNrV2ahKUAWKRA9cGlsMcxv
qiOtzdq1118CyQSJ737tB0BM65d9Of2P/jH+eOX3Y2Y7Ua7i5hw1G29c/pGa7lXdJMLKux+JqXBH
K3ADqxaZwQSDS+ZLHTk4tt9aV8alr9e+NnC8zh3ztlrR/zL0VmFQLOh5JpUspNzZlDz6ALaV+V+J
dp1Zq3gPtYEyVd8ERA/uWj2cNm3FfAWAdOLjZYYBquKNJsw7N3MRI5602Mw44N1K7BqZh+++AKn4
muivBA64oqb9GZEWEjee1T++p77cexxqJasBtYnTl74xp8IhDDNhjQetB8QOA6unLtOzcQoG1Hno
MtL86r6ZIIsc7K4oGkDBHJOqK5BNGj+VBWOfobRXfAXCqSS52Hx6I42qoSFO/F5npp6RQIHNBpnY
VAfDZO9etHWyCT2UWb8tUI/lZdUk0pbyT9fH6mYCEz1Xewa7w3jOkywELIPyZELdAVqPATDOBlW4
y1xGfvOpo0Y/x//IujY+ebLFvz7Z4o1NB97i26YAFlXt3cwpUwW5VEs1/rFM05A7LdeqBPIYJDFJ
QkuB6ftprw0PwJ20bHDdbpvvc9OVyodPRsDhb6pe6vL3A4vjwwuo/g+f7qSgd/1kQIjuHTK41r9J
3MbDu1O+g4dahTqyUbP714QhKNMn64ksfIFZLU/cyGNOiW/PbSehRPfXpcUmgNa+PeMiVVwVjs6y
03UUEEt/lLRnTgcqa7lO9qpanwXSrI8JB1WLu6yMhq+5hr/0wV/HN3PJefLURTDIH5ylrYMBuSk+
CGY0jg4g0YUOpHZBbp1cUqLiPgJu2zT3w8Kj0k6XtgUSQzRF7V0q0EzHexPUJPBidMMNCZftZJN4
8joA6v5RzJWlIyck7382mRyYeaLXFGQht/Lty8IwgazDuMsAUi9Ugc+CFXmMe608dPVna1XE1Oor
/fBayALI9chXgO6CnvmuQ/lq2znxH1bGJlVvX3b8cEP2nyhTtDK/PdAN4rBW5q2nZPVz76lC4ZSK
QTxeO9V2A5lqQsxaFWLyM6fpwK2kzDkKqqLVOkMkznDr5G5yM+6+u3nAZnXHgoNLqos1x8HUxFzl
mdBBUSNbcNvyoaH0OYgqDiDuHubHnKw781JAwCVak7LFzJWJLyJ1q86rRJvtrnK6aTvdJY/AcfRg
GfvyGVicwiwslK2pVC1GSKTX9yGwEOBWUeLvvODlgaefhUEq8RJzmyILPDSwoA2O9/c3DmllvrP/
44X25FMcEG3uAsFQHzQdG2SoT/E3RoLabPMncnpk4lDenEIAuYJQPKEmvlDadiu90zQlpbd0YNl9
wj7nJcNMlt5+BBWtWUHdnW9Rdc+LfwIkk1ugBIb9HoTh3bz7s2rfg2446zJR34A3NG18aTrlb28g
L7GSMK2HE0Wi+CUcVosbRoEGrRJKRVgR4bAjMbqARFxFJGWktes+/WF0nKBJYjc+gLfJ8FRKLU4u
VkZP/KB4F15t7H1QNy8HSgIicOnVEzazePt3IoVkZReL+kHVZ/EA2oixzW8aao+VyoUNKE330iWw
9NI+QyzFBD1ktcG0jSpThR1ZDUsmgCpLXirLayDojxccT1ytyQ52sqlQC66StCgAhmYdRgN+Bh9S
b7ZLBDGJA3XmuSWYplMhlRt36+AY3LNyNnhNbO+JMJMoEm1nmGV/IQvbU+hjyU0SLCGmIMtALMKD
S8O7DHR7rf+QeXCenCDPk3rZ0BVIUZ7qyElANpqaB2ca0v8wGbyv3JcAnHUinVqWvW+Nk1ZC5T7L
Uyfe7TkHA2yiOmglTXjVcM2mlf4ILmqMDSXPp8QTxjLI6oOhmERr/+MrVencGDcgOZArSdjtWazQ
AICmC7eDnMchpwA/eI6AJEJvgnScqeQ13wLgXD2hcOm5kJvC4IWnQQBKCCDFTJAgF7u3iMWHdB5/
z7XSbYiVAOcOgYzwWdVROl6LT69BHB4+UXZSxhmE6MZ6gSV8qwhAYl+muyWced+v6uLmNPq2T6io
dflc8x6VpiEzn8McrmkZFx/ZOluwd3zbzOsQ+aXwttH9WwujnE5E37liyHNAJuruUe6yJFvItpFe
tN9NiXfD/mF6jD3Bnu/y1PQlFPG3pQD0G55cB9Cn8TtDo0RGPDupcV1XD5bI40k/N46GulidG7SU
50kvinw7+hYyemvRI5PSyJ2oaOw50d2TogN3G+/vYSpzwQO830AvRy/3bvOumQGky4VYkUzdnMSL
7Ouvqi9rTG2C1slTGexkfc64HiEdBUyPcdMuvEkRMF0UZ1poJ3Gu5cvaQwEt/AREYMRvARDFI7kt
R9m45/32f6IqoHjHlUOYgkloPMTGYTrbgcl0LdRrugFhRGv9wVMRTVCGgq80mPCYjEtAlLPB6bPC
AobHN5QgIF2wjzLhN0uEkD4T92vXB8zx9hnJQdR8g13kGwOh7GtPJMU5z/T/lA5g1E6aZGyeuwJp
7mTzRgbLaTWTYR7p904a8FOGJuIjb7165Zt2dj2mJ9t83DxWDUvRKHkiearzqGPlQWNs4Xi9ZceZ
P1rWHnElZnLzq8ZtPkGNdN6fmyVJTMqzUI9QrNT8wdVUb0IA+syT5l3mQHyGCHmF2sPbzNi2+QPh
6CTEemxsivUzL993oz6YVD/j0CszCgbGCeWhUlAUcZgfU66kB2+1x/zz5dYChDaEhauTh3bILikZ
LkEs8kzHwPal0ZDeG8jwFJag/Uf0Lb9u6EtWxZZYmU7Utqz7P2cHY0vRnOqtUiskYg4iwJZ6qRZU
MiSge4nPVt9DBD8U/oKTF56scIdpFd27Opkva5INpAmxwMqOdbIeCwAnH981cMAHB/GEMRSPqnS/
pu5j3TiQOKr3PUF2MJWUsNKqzz7HET4wPrUxKbZUB6QJZufERA+lW4gh/1dDGDWOfpgwaEfQErm+
KtIG5Q1gReVG+UsKBpBWuNWo1ysLykhtOdiIa1RcwuILhv8RgH4Dw3EKWfsfaUeDTJGHmDK1U2ej
I/AlLu9np86BN0nfWe2bqP3P2U91RwvvmGPZ6wNb3VfIeSaAGO9NZAT3YlUJAVtYv740JJTwp5OA
4ir7+TcX+LFPpSpm9uxYXmAXnT0X20EwDOWpSyShNW/N2ZjvCFq/5P/HIUjvW+7C8Tm3wpMbvGYp
aJZc7NpPd2CFoSSnq0VdO28jx2yc6o5gsByYHR0I2ruMcgpp34rwCo+KQQo6PFzQGM5wSkFkxy+Q
YDI/q33CsndjxtVJXzpCMNMCAKbppqa8nXLBPv+PHUxdoLD41hA5pAdaPn5x8xpErD7z9mLM6o04
2DAq8/BHS3e+mW1dxTGFzEoAGmlZMrjhA5MFhTErAC35xhwjgfFMwQZVp7DjkQBi2MMt91krrdP8
vsTYIE2iQdk4Fg678ualXuE6I6CzV6JsIgDl+zjleIWzOhDqkP+/ZKmvp6uwgIhH0psnzCZu3PXM
4Nm8pv5cp/RDE7DYsNONL4hmjOy669GKCrN/aSkXv6vXJkjnUHFyx1r6HaOxTw1mZxDF/oFwr1Wg
80lJkF4aMktzdXry8JfupGEDHthzSobZbEgKO0dWMrr5mxngWtKwj5uovHUQ4flNvjJPqKyRaY5V
OLXd6pEasfQexQoRtma3O9WmqBoX3YQOhW2DBvzyFwhPgrkTWczTg1JbPXOJ1rcjSeM5aHDgai49
yR6vkzMElI8GoXbyzTOdt9jdw1KmF/w7oUe3fiFtq1RBIofkSMvF3V1nKBVtRbwl986ET2niUzya
BXSODeCm7xNtc05vjjWuh2yjZEIOxCPfBJEe6Z67ckt86hVP5D5GwvVdHUIn1IuxilDIjqoW3Qlu
BTvcnX5w/eZFgiCvFURmzyYoFKxjalyAzAmPd0joJvgEqZRdZOHAR4gPdpL6hUagoROja1xDRqn4
yCSys+93O7wRWoKiUcsnKRxzTenVQNCLVCaZPzpXJygAA6BXOJiuI+zHg8+8cwy8+vVi1976VW1H
FJTOuwhVc+hRPyl4p1b7F3sxyNjRfPlQnqH0RPxWIQYMgL3kLFNPA+ts7S4mCmOBigG/aDg3mHmX
g30OJyHEQRaXXQ3YcFqGjqE2JFVI3PqZWz9VE9O5T6xCAKKlmAxHdxnsaFaRfugTbJR9T5JLp/8+
OHwff3ln9fbPJq/3OL6jZIBfO1+aSFLQy4/1f2EmyDuqS8hJ19BAZd7kNQ7JgWLn5CFAV/cSCxdI
oJBSXm+nb59lM4EPY/W06eAPZNhsAEOVjjzB/Z0GZRQKEw4FtxkfrmhoAaL+vBn7PW1v1O7yjWcT
LihpjIwpW92a3jUn9iM+4dUI+tykZqAJ2m7nPoK98h70S4d5K+SGjemATCy+jfXamIK+IuhTJhPm
LEyW/cKGE68gJAzmzoLYMapBV0voEoMAD1d3SarQU6HYMiLQWPHiTxPUh7ZV1CWiWdV+PzpY9/lF
pVM2yD4ws2MfgIXYalslovEvA2DHjvCQPmRXM5ij6cjjLZCZxNhpdR7iYoedzeeG1kcp50HoqUUE
MtHQ/BNn4K4AwSn0l2YpxeCmlF3xEo3LiOmQgHZiWcw+MlPFfAjLn9fG3Kx5+bnnZHipAN3E1280
Zgn6tJwMUEYYIOLt0qRn7e5SzbK9ZrjErWQNDwG8Gbe62nrJLR/kj8yKxvQAle9Eti7HSBXdW9+s
3VUzjlwH/SEXjamVIU4cAw/Y6H2UObWIyNlfj+qWgSD1JlMaeHlv4J7TT/OMwZayyEki84xtjrWH
qk0UgvbY6nAxtqB60MkIVuiNovjM2ON302TfQgAhaOrBCDRc5H/QckwFs4Kp1r+rNa8xNgHV+wwC
7IhXkhhJ3ot3MWoEojT4ZmWuIXfAiMNVLzSsPOUNycJhiv39Lb+XsplpQjnZhi37T2v29CkQbBpA
8npjXbggqai1v3+YcbgKvvxlPxYKSzLKKmvcsZevpF0kbtAao29KmS63bNetnhR5+u16ZapeyhW1
502h4E6iXOGOPQRaI0IR6Ptyx2ZCvrvh7Log7VeLKvsPW0ITysqZL4UVlsp8RqEk2nBxMgsvtP5G
GhPR4VjpLeWAJ1ecSblJJfYaBVT8MrxJz2YRCqlIjn4CwlTNA0wIR3IC7wjVLHqdaccSH6is+wpJ
HlQP5+fJsIRHb3Ijv73Oy9kmFWfGA7o1a9SFeFMeU7Md8hEPL5VjLD6fucpvSVoxRRqPIBDPD4QL
rOrqFRPXaT1LFv7VwyvY+VyY8yBnUM/0A8utQchbpBXjCYfIGH68WcAjxY48Zs7afEesdBoFtAl0
JazM1c04UMNLOtIanAy1BIkXlaaJ9nq/E9U2QLEeAU24xoj79C57mT4gWhbOpneqeTpQJKTkQuea
p/2+tAkMLbMUOP7EWtCBd9EC327nrvOwU6GdYBfGs3/o5AIHGQ4gkCH4amuk2QE4b8HSs4jHTG4n
iz+g0rCxmSMajYM4f+5o2dlMQPOLcFxzfbS53jq6euBX/D2FT+KRLz4lYUIGGyv/lCNNzHerCC7f
2D/ZUcVE+r7tDVWDVlsgPi5Ui0cg4OAlSKwaO4vgMvN5cNyG1i/NVNcse4lEV5KjtLmRZR736MF0
ga9xYYyNUGzmf10xOOw9WGGBQWWPQ5l4mTE0Vq5Wq3w6bbWWLhVE9XTRd/w7bg8sdrHJYyo9DS0l
Q3yclISaaW/HIt6gmYB4OGdmD1N8rvFg+8cFZ5DM1V1p+AjcrqNzCAcLeUf1dS1H0NTDTaomYISQ
SQd2WgHUMDlsbgGIwXY/zl6oIn8dYswqKlkIA8CImaBmqcOJVzUFEXt01n/dApn4Eu8JDvlCF77R
os1lJShewqWOPNhyaN8Bat5L6rAe9ky7xQPw8bo450tfHuG4B5bnFe3qf60HS6PMcaGaJwwpvZYs
OXnXfvVAT5GSq2Tzi0U/FZNRzXvXKNBgRauuDPNV3zVnmkvQNPB0qGNPBnp39iL9L0tN5ZAmCs2w
fJ9/UA698uRIe2Q12CF26aX1Q5zzM09B87BL2MKzoZJ4g1wbo6vf4K9Yrq+wbKLHrXKWQ+mqQ1xC
wyZu6WA/L8Ccfuxihwt1cEmCZsBOV3GCoQ3p22z+lUr+JL54zfoEOXWRFyz8EdinyAE4JXQfQGN5
BiyuA8OxlAoeetOCscSL5VApYcsJQZro7mXUB9s2tEkdbDgnN6PEaxiTq7zlUtCGZ/KlGIcm1mE0
lI/DcUl6JAjXnvqYJR28FbBOqKwByTdsABS2ioHBh5MqO8whQQ635u4yvdXuYzoJ0FmxFkipfKYI
4GuC0BaFAkM+R2eLQA1K5KO88y3R/CkuAQifJdHeRSF88rBqMoIgJW/yxrKZP05i8Lwlb2dLQZ5k
f5u8LPY0igpf0AJOmh6AjaZYqudoe0zkc1+wuLQXoHtVZ3YXy8igZ4D4DFQvLHlLq+0xayKn8cal
baKijHhTU2GliRBLjaHVxZ0orbqzbCHa0RSxSAbH+zVAis0ym5q5CAyFNtjjDWzs5i9NIkzcvEP5
ZAe2UJRn3AGI/V0Hb622vrT1U9zRz2LVMM9qDIkD+lloIXc7dEgIneI5yKwtSkWvh3P/5mfmUjKG
HFFI2dagaJ1F6q0inJcPcGkhFFtlsLJARAsgvRPTWm8gIH69OwmoMYqWX+iIJ4JWtzuz5MBvpEDT
1Q8T/ftU0bUgG1ta8jJ7F7lXdpddHwqlW2Cb5P/EI9iXlNB8KDtsY7YkO+eGcgFvPCUMxk+JeOOu
ua+wbYg5Tf99ZDFxqobz18ApOSQB+z8st225O/mLUEH1wyOUvyIXFvFgTOMBNTwUvtaqAv6qIdqe
ALhl52wjUAdO2YWNPrd3Jf8f6rSVxWV6VU7WWHEAOpcptybqqfISy9GkgxiW5g88wjFXEwWgkRSY
urP0yrnKWe5ojWVY6OfiI/Ne7cGiYAEi5TCVga+6Q1MzhrK2P5rK6MlN1S4CgLPCO/dVmgx+otSk
EnOyyzEmXSUAIf1s2t5x6EmSEFsvg1w///H7NBgC2xz7TQM1jvOCPdAgclGSZWsT3afLsXVmxAoe
vSPysbtY2JK7B8I5cY3FzwvPSOQfgu9PeOXOiKF+9OxkBicvQILbUwjsjVkVkGBWrtDx2KTsrV6O
jPzpMOHFfJ2/TdhuVbvMouY1FJt6xqbSD+uRIG24KG9ivXdHEkfEXo3LqTw9yE8FYM6FCHSjB0pv
fOV8BizTNax9Fh9s6qkJjLZ/tsgbWZpCKGWcr1YqGl0pxwGws/sfyrTjjt4GPgHTFZG8z2a0JZmh
csG9ZreKvmKINKAN7WOBUCdjbUBYMcTcE0SPPzrW5K5ik0BKNHwjMs7JoouBKFgnBk42O7Ra/w9H
ans0GCrP+k7BFN7iCkfLrSa8NJNbXCpvElRQFLvLmBfBHQM84b9BnSFouGAdGcm2ZBu2kiAF2We5
o8OPAM9dxVfCercMW4dzmGpXXVKwkbq/gRv+dTJGt8Vdqc5Tke+i4014fvafmrt2+yrzOQVAMyKn
qR0QcBwarZvUNLO28MVfuh746bJ8voxBqA4Umbwzmm2kV105yJghgrzmSJ9b/pjZi7PqX9a27UI4
/jPqwQiQz6ttI0j0D3aBmkOs3xM6ekUO/tmv0SXdRuDCx8dVs5x29bvBiYbUnkHP8+mRVCdw7eRm
BYFlETpy4JGJMyf3kj1DYaSQvqFQAyADg9XxInD2MLNofZbtle4WDYgkBf/FM+XzLYlxHOVlW8gu
bd00JIzk1qhFzELDsJ0GVkGX4XTk1pKmawmgmF9IVXr+gb/YDUSZ64w8SrDtr3vZgQVqCYrxrUSG
/1xymSIhxOiFkMU98VNtNVo1D2tsxIM5kUUP1LOD+FbhQZQi1YHgKEwk+wI894bmz+dVRBl0t2Iw
UTHENIiuqAke3Gyg4MmHRH4GAuJq3duvGeRbsb9VY4resX+4mwWXZx209t/SzVYp+ccDK8VF42KF
FfYbV4U7n0sWYuSb9nMNQqNFt+dU4BaUTtmF4vtr4reR5VM50nWwhLCxfx2SarCFXtzz4hKqzLCu
EOwSbUP+a91i8Cez4MVEcDx2iSxKMa9/5rl9i2wHlbi+T0wXrxKCedJElANppJ0OFxc0i2Y/HyeI
lTaJhaQhg9NOrUCxYFO6oiYXe94alf7sJFNLnLo8zecwEik5IEFBQFaqBvmE+aVjv+D3mrXjVqkP
EIRZsrplM37S984FCxx86D3ehg0qcO6fZOZ6vYntjoG6tnSrnbcxIthYsxs4pDgkx/QX6OWCSGvr
RwRnGF2O+gvPf/1SyaDoV9gD/dhC7Rt7VL7SGKClJjgOL1nbvSRr74sWIm3lmsaUQnlsScbGEktl
6iKZuMLL3PaGNdNmEwtx2pLHKcMnSGhQUI2VgFCVQT/mGEs8I40fLxRu86a99siG6zjTvuAlKLg/
aZ8klmEfWiEblrbkLslcYt+bfz+mvh+zGX54sMX1N/dfsfJRIGFeLNrm4rKj58NYnzhDO1GS9zyZ
0DFAGOOj/AlgtrVyQNmtxjoniOdnaelPrI4RXvAsHSeFpREUKTEs6IW3wepSUy0Cte5p8EjJRrJd
4LNh6k3n8z/H0ay0ogxy6o+R0fIEh/1/Ru3n5/hCxhVrtgmoKBLiKxgedHWcCrfm251NFhAyTA7n
FpgThqm7q8JvV/jgqbqMEqhnOYd/zVhx71ikD5u4AxRjoyOPs+RHWXyrMzGJO+5quzdcZgF7ngdM
TKd4d9hulBnh8/P14E6BddhQQwB8tvw9/W2SslCFXwrS55eS5B8NbDmAIsmK2ISfXdsr9YQoZJSK
y0GGKWHm9UrcYl8SAYrtjObyQ6eSCy1O8/6vHW08LByelLP8Ickmr0Oz0pFxznOhJJ6QJ9GwiJl+
vuZJzgJqqtnPbv2/owg6Z5NUOOl4l3kN75mP//2EjY/OhoJxVG87C+RBCJXllvPSgE3BskP4dPlD
FfAP5sxTeHz3c4LuH31gtMrvHsiRNCp36/qa8U6G7Un3dE3LsSvNwvyB8N0LclOO8keN2NrxK+qM
5jFtUAytzrxe7AQ4FWQeHL+Rd3ErtfoObzm9zzQqY818+U2k1+wk3qAc/lxS5tphRyaTHJZYiynL
mNonImwJSCy5Hqe/AKb53F5nAtNz+UokjZdBQ8N6dGPx8JEO/vLCtdPVGiIqKXT3a2H5yIrM86D7
dcyXzJMZY8gBR5sxpGfztL7zvU3s7bDbYMa9U9+8is9LxxAkp8G0AC0Nw+9xTpofIuYbEJtzBzo9
SdjqEOzQACCGSKtGRMfgE/6lhsTaV2FTHy+dovKDYsIKEPEjPJrwlo5yL2bi/v+gWwSMzX2oRS/q
d+MLXu98XZGkesHcugQn2TQO9XVaEF6OiiUQBR3tGT87L3RKP8bgWjz5NLXzKlHVlpMGk+Ee+tEt
RL+c1c515QI6QQzy5pN3VeevDLayTNZwd5r1rHwk1Srxnn3p4NQhmQijf46ghVE/BCLOUOXg2yuY
EU+94Ebwp5c7U7UIJWt3Eu6HfX0m/jZ//Z8JYth2TXMPgC0D4EadZwcm/XTi4vf7NhUdNV7IPNBX
BsaYYNPId3/N5gMIrvZOE8HCzpNhrzXqB4k7643DVts4V2iVJcwpGy07v9RMw9yc/QKwdpNiPc9O
Sgu0AlAS3GzmLdbinsLdeDCBK5vw/SkiRRp/uP0sst3/Taj5tv2Sy2ioARwYL1sTVShPrBYq6NoL
0qLJ1swZojiKPgFNgiPQIkrwjaXN6YE0DnIX+iZ9ThB6vj0R3tgIEZC7/9fJN+6D/J6J4Z7FrWKw
oH9pGcIygmZfFMa+Ja/m6dey4r/bHVj6GFfiYWtQg6F7+v+vZ+tIF9ODUm8pFxNjtAOD2jAUjZHY
swLhEqxALqfQL8roBUxMtugWo01eCJ4CSbnkDc5wzmnzLv1U//XjJ4sprEA0KXQ8TRztTs5QPd87
gIYUFmIKo8TVX/m6xhah2BzBXOk+xfmQFLAAVudU+/J6w9ZyotZoO46dQScLWTgoCvJtAimU6+w/
yZCdWlAJHidm+zVS+iNccMAuYd7sPBRAtbLO/zMz1Z92KcbwlFFuZRHRYVJj7subvGE1r54LxQpL
TYQfmKuE1+p3KmxRLjf05BvbvrNDcPcDt9vzQyRitN0V2PSWwW0yJNDOBuxL3sAHDm/D6STlwun2
SEEtPIerxzBHZj82Z42oLxBeKKpbUQR6aDMOxq8VgG2qpdr5p9244HuAOBX3YtbMM1kP7H/B5IKj
X00N3zf/eI1vSVtlJVaR8y3QWt3WM0v8P58XaKkz0twWHUQmPTY7eecGZy+KfoH/k7KJA2mT3ZvD
XWqGv0zaDiL6OyjNC72MjMh0BYLVayG6i2uBLoUQZN3O/Ubi4uP+BOmeQXKZMHmlqCdPBMDrSotW
c4NwkIQW/gHKpu+tnQUlaEELuLxOJTyvKFXlcvt99+XHxR6ggP9fqXDQePm4g1O/Vl7LAZ7XP7UK
kU956qGvGvrbK/xWWck7oOapyPG0Pm1ayW1+beMRbhL20AVG03JdQshAOiR7lQ32/xx1NvVc0huz
mxr0KeYscjeAy2lMdlfX/OwN86S9hhfHv1QR7/TrKlymCeBv9oh8IfdULLNU+pceFz6eT1uJS7qP
I1UMDyG7lUctxaqh5u+3QDrqbRuQHzt/iixn41ZySAfiluEvrZ5t2NFV//uK4RYIyowfzkV8g2NW
FXm8s7kRLXeb5y06Jy105mhZucZPBH4gu5vYH6CQN3AgtnCOtL0xFhPd6MdPDB7QjR+rBQGocMSe
Qp8zdWxubLGKI/aCdLHmfQjFF+qiOEkrh4ame76HPp9/jUwgp98hXD7DeZZokbuEsvUgzePuyPC8
YwbRkO2c6Xl9zm8+6MeMBTfimH2KO94OMEvHwbg2nJJDMn3qJjsnEOfEz1/RzE9+Hp3yUBDoKfG5
prwIf+CqdPus90X1wdHzFj6iA6qnaFlbt8NoinDgvo7VK0aXjHlbSz/M5p+TNywGeW5ze48bDAlV
vE4fSE4E+ALGLLCDiJbOEuPoIiVm7YyvZsJ+bd40DSGagbu2b7YU+VTKMUHaS8wFRSprpiQsT8j+
wlYIZ8g4yFt6bWM9ow1xaPmhLadBXzZG9LsZf5J6vV7x2Tn1exywVggWU7GAA0fx4maSBD+Kt8CJ
FwcLGOC+a4v85//u2ZumDY6byzGTRIgEdF9RRj2+h3S6ufZNpGhDHjyXNY3nwhvIK3u7PM9/W7Cl
TrdLpPB74vCBdFQbJMzdj9XzFMi4hgulPom3oEh62XKnOVYtmNyi9U5xlKj3EzWtguxj3APSNgKd
bGsTM1ccvqt2S8eF4QXKtpy/aX72euL0+DOFVhuOVKjfh+QGsAjI7m1A2n6Ej13XyXP119mV7eiL
jaIDyxhN0uoh9MfuPO15YQ7qNOfTwZdDoTxX08qSDq98SZuTSq8SnnSc+vhCIi+M5PZ9F5c2XeJY
C8asqNYRjhHoSFdXplgCsSDHGWAw4b+BLPOy3VISSMAZzNYzrwfSM1/5z5XztLw7Goi8tjoH9ID+
0wO5ledE3FmO5spSZfL8WVvbs7jUXfw1t9qOjd58bHkvU/9l7ScTnalMUchih0gNQJ1Onl8L7/+B
k6IEa/1ZEJx33+H1+gkcHU5XKmodgzi3i3MG4wzk8EvrxUgxikp07N6fbgZeoW+fBLWI9N1Np71D
1vFhY+K5AFUz5MQc/jbI6wagCFnUrWJepQsfk4m8TF0VeifBqBlCw0z6VB3+PNlkYybd2Ahi7NGA
Lf0cUZmosQzkz3DSTfwXjk2hrlSLTdVJE38XG8UNHdkF/mMPcMiPNgL+IrVJNfuFH2cvxD5J3dFq
2tGiQjCY3fFTPiwkSjfqPlUtt/wsLTa47KhkwD/bwLC5byf6XuwCT0hjAi/gGOONdV+JWzQht9xL
5pp3pYHfPAiyIAu3ViLKkno/S4n9wo5BPCwURFCtUvAUkh4+nyqWUfgoDUq9kvzb0dvauyXZab4M
V7uhFHbP8eQMnXDYJa/a+EBkMs+RL2EZV3/jtGd2h5pUlmo8iKHF/WnYpj4JvtOBUBIuhOpcEEXu
O41m2aHq6uMj3Mos8XSOIHJ1loTn4oRvn5Zs8Ut9QRha630PLUaaoAW7hp7riVs8CTcSA2dUpjIS
dLNcWE3uQSHsYexTnRF26xKoi4Mt9EC6CcsM3CCnHuPHxJaaVB/zE9CU2qPttwXHL/1lAdxSuDUK
wotxyH+/2+PDnshZM0lKQZQ6Geiy3RnWFgzzup/jvAyIWnBTYKufvqZHNn69pd50I9nQ0vxRevhh
qhSAY77L5YyrnZKLU4cqHjxDO3z8YkFhmUZirA1fS36nFq9NMQ7v6cXz7Pn5wi5VWLDSUdPdSfaF
03+HjeM3obLGpjHaLm+IsAIfT1dUrth8kqqH2PIB0vA9nvJYG6CxHs5pEygYwc+tnKs59udq15qK
0jc5U6bGceqKKRlJo620SEE9pB3qhx1kc3qVqecUqb4oh6ElOBNVF05lsn+QCpsHatNNuNwjHOSK
CGyRBUEI23+FH4J/nqkYoAUKXCaEjGemZxNpHbgw46qO4ZFlfhv1DxrQGA3V3Zf7dMKuJZMHLbZ8
BxbrgiTpxFfpetuFGqt3lyLuW8xnEthLxZudmA4ex3ug8lpq4FY8Vd8bTYeE76g8Z4ZFpEsCYURO
JpU0rrqxVYPIOVCqKdK/ApWbONMRLfDgcoryGxZzwxDYhSExwGtM378Q54w3m7DAlaKBQOKKJd4X
OSFW/XzuEASGfP1Gk6hAy2WPhUBNVG/mH7u+MsHRMl2NeRdwVTS+TDtOAuaToQ0w02ImRtqIVYyI
DmZ/4nmRHFjjDPTf/jxVKevW65sNEnURVjY52G22ZFxvdVPKuwNSY2+5Qs4ZvQ3RM4Mm5lcnaLbg
WPtwoFxEr8zJiOYgnmgbrDay4js+IrLd+vTc8WOYYbAUd3RJRrJ32JL+vhc0qdoff1EJe9wcYT9v
p+PRmkRHt3t4Zi4K3QE2BHmI2x7VMM/ynbqF1ONDz2ZcfG1YOu72YG4nxRLtp3ZVIYQv2SuDy1EB
Gc5kTFq2Zg+m6W2yVKGcL9mzJ1dszIgBkbKrY86p2nydRxouKalqxPOJs9WZQQiVFygc3htc6M8p
UB070kis0HBDpEvYZgcboQtchlWv+Z4qo+EFt75RFCWAytwh36DQl/3wm7DWG8sqrFeCUOhSGZgd
e36FoQYPDpecdPADBa07zc/Cu1Z4FDrWa/U/vJ1EQki6Ty4FztmB5rnmYgHVHWEaEWAxMolChld6
Qa1xq7wGyk6VKFAmbSANeSs3qadTVHF23wddEQkzII2Jh5sEb52OIDx7E1+ThoLGAxll/1yIEpZ2
aPDjBlnCVsxF3OBSgrv/i873745R9gcw/A3gQz/4js7EGliI0FUZD/fsROrW7tWyUAtcL/Zp9+Bn
Rme4CyKb8Jmt5G3ercQgM6hMaUCaAkZ+4fLF+g0d9Omo9zVO8i3mUJx+TRc0lK2k5KiU/wJexWjc
N5hEAk8PWUEenXGlk482KL+ZeuV3LmEyfxnYk1jSHO4pXpQHwS/6h5J7pdZPj0n3AF2j/CvPrgbs
QPyI1WxLReBFW7Q59wPIw3in/k2AZA0QKXJ1sL7AtN2LBQ6dOTOYrevQDnzElAcbD216jHpLAJra
AbRnSUh6LA66EQ5DUEbkfYnnoRta4aOe6IJm0+oP2k69hGJvCgZqSi7qnl1usaMCZrfinzkMErJa
kjahBulkKra9eDO3e+dzMe5Sf7e0RfO9b4s5wcb7e6r0D4m1fE7wOLh4nCbV+UG3kqSukGdOk4o4
HzdkG2dOU3Qy0RY+PBTEt5Vpo45fOoDGFE7sJsFYc54Kmkq0sUxGpRdVR/UM73pEQm5ddNUBXEut
q1FWDltSgAKzkU7ZwGRD8FX9jz3K/foxOf8DjeZr7zudefswWq8+PAxMF6+L2CKgt/bOisF4H/Xc
ct5oaDR0Upyc54mB1WxpFqcmMg0rOVQFAie5+npH5deI0/mK9MddDQAFqGRs1vrKTTHkKDOsVpmO
huaqCSCirRLwv3/4RnxWM2wMjBkLDkGYdFayrt33oHjerS1TrYtlkSAIQTbfLNSRlMksyolceXIC
SbQHTACQHwJoXjtCom4YwJ5kxGz+yOV3gnK6V1tH2bV/8p7zixU9RAeVB5CDK+de7FNPdjlGbEBc
n5g1lwnukXtTU1zQq1k/4NRUB0TvPA+IgAXpNfml4/29fEPQaYzSFPDMKjqoIKbWb4c/Lm+QbD17
L7MVx3jrsuUo1hW3dn5E0+ANbmkEkU8cH+uHM/yFanKW2jHf71fBhwCKLbcKdKaJibBZUvrcEMZk
mQgx2bsMYLlnBeSfdsw4BA5iX66N3viiFeeI2pneQdYIxgzUGmpFqmBAZRRnx7MMHZsckhvVhQoY
h8znOiUpmHF85TVJ0H++TFatlEhLRRpVRzQfGPmMKtBEqRJlS8r8H/a1kUiUyPIUhLy58nXCOIO8
Q7Aoaav5hNYQxnHhZXtjLiF+eFqlrhoj+dkoP+T1VN8AWWVpQRqpGex8Xg/+AG+m4enpst3aRnj6
6WbMIyZQb00rYRacAXNf8g+XnmgWp6iBpO29VZPFKxhOwykD7hWd8sSr16rxM4DVRsi3Ap9uBmH9
1p9nETuHrzISnkS+Tebn9IwqNqmA1ad1/adCOoBus0dzRJc5upmtSa3DwQ1wggMy75Uj6QTi3Jas
B5TCUh1m9Mc3C1p/LzVvsr1nJg0Epd2gDpbIsZUI7rh3NcrhK/b//j32M/T38mdRU+jMjoWffECH
4h5TEXpDMvKNy9HjKVdjC/0zvrB9iqmi2tMHQgVcgG6Tm69tVyu+YenvFCOujkFAmQDkK6ZlUj0k
Dji6nkl2MMzxnBbvIVQt77voxlaFhNB56LuWpp/64RKtnGIjTkoIfnPIKN0Z8fOb30EdavEcvpSH
d6gkuWmOb1I1LRhGDULYtS/N7tA86tYuBxH52pMWxdXbnZwNQTL10r0J5FP5PJF+ZrHylZ3kuIAt
1JQHXo52VO9R/JTZInit0mvtwPYHv8r96yXV0GmeQ27yg+CtLDLW/bqzWShJnitxKkICSUe8Y2QT
x5vXGuz1Il7p5/0JEmtncXbajVY88y2g7/yq2bxCVQBw60NoqN89AaPVIEKm+v1CtyD63jHI8Hxd
EjADfqE5YhcHWEFWhDXqahNLawRFoKSt0LPKCyKFMFpOVLn1cili3BzUdh8p3D65oBDbGOetugBI
VOIqIXF8mKBUCWlDLPjAjidL6U3spqH5yKzujLQjcbfS/NRkyUnSDbbOnxSvnmZ3c62pXP3QrwsA
5jRqccE1kO2HXTXDu3j6DfGu20JlDmys8aRzwpEb2mLnCLNmWcrcjFaCjvrHec14SS0Bn+0d9WmI
LRLypVjJ8EyuxDN9jDtT6XmCcGlNN/9KnMy7OkiA0wixvw2feFNBPlfaHH5tB+aOp9hHLsXjILAT
zMilXCurUpwbxg8l7V3jKtNRMAW4wsziwvzIVHuIhlx5o2eTy/xBGjnu0j59MrjpVZWTtxFJDjqt
gIQQqiXzh6wlUsxvEIQSuBv52TWf22IUKpPjhKilSdddhMqd5f+qU3Gl3hblWeMQqwcLsz+WpKiI
CxWN4da0wAhrnmnLc3flAiqkvKarcuTyuK4xKjw1c+M1X6W3v4/sHoU8VlWrzkpF9NszTVMTGqgk
efJ9zCyLz3OktmYtynhiIWKQwJ4pQDNLriVuZ3PFxUuqcWe/tS955iYzDhmmeGDKhVIrOcLeG2Mh
UJwMTc8DKfenPnX1d95zorvg1Lesvle0vTi9k5ExsiCvpRQACtL0/4yZYW+oV5zqw/UK5S2Qe/Wm
8m8vFxcQ6NJ0/BZNS5tPVLDtoEbQW4vTALq7kJVS47LQ18FR0NWFb3OlX8LHNVZUVIRQXOWJ2+8S
fufqeseft9hAcYjmLdeCANOwl4STpqAjHlGHd0D/++htVY5eY/2ncsNu1iYVWgZGkL7f7ugQLtg/
3xHB92q6Y0mRCa8t5ROJMN2pVO2v2wNNERM+JyjwyOdei6P04mt/ToNg2gyMGQQ/nykRtyGcM0VW
oFgeOjBDDqSl8oam8Vt80Sf1OmmDrQVnYckpTwC4aI89VuTKYIXG2NkWvhmilJ6YYmor4UCxbCrY
dnXL3Mg5XJdQE4joTw5IBC1pDil14WeNXPEIcgs9gHfK9QPFelZvWUa2z1DRgtnHFNJ2/9SlGR7H
WkXS0+T4luf91gB4CmviEMd9OCKsGL6Ct0PpLHEhlFd9zNUz2Y7lQBZxhWGDwHWoTCZOEj5BoAVe
lDS7BFbzzIMYUrj9QBrGkzJwUmAAA/peunCCr02UiJYzSBNxKZ9ps+Wd59EzG4pWvFN/l0ngrFrW
93FypKsOHSeC6zd2qHD+twCYzcU3TnLtzlsrz7twdlgqV680lYfuEGRnMuUMpwNHzZNkyorInxV6
8gknq9bNK6rRrAwHTLGAPUsrvtlv6yJmTlp88puyYtnptxQNf8VC3Klu2ysdSbb16Id3OHJddH3i
7iBp2KPmfglKV9NtfTjU6qaISuj0XoYebUrP4F7KYqqvUND1lTYIXr3tb2NrImm1lziQgrPJb81P
RQKlg5DY68yfJnT02rLPAv5eiSXOHl08cJDsy74n65wtFeoU69pxcAJEGwHjrIG6b0F1tLFIJPcg
/0gjDFoVMone4Ap0n2yr/MwxLhH5XWYzbogwHLThTqZf/NuX2z705RGTg3P7adMXliJ119WFhnCM
L4cccZO+LK+UKLdyakLgwBfRVy2arjQpZxkYRU2PPVvp0jNh6CnD+TRtDVPI9Y6Y4LB4sprxZ5Vw
Q76V55iAmoWQ2RV8KMS02wfd+z/WeSfEf7Lvc6v+m6oJGuIX7lm5nJIxyB+oe73IUh7Ttc5QU8Jl
o6Kb6S1/63hs9GdiD5NB9+MjBU5GIBoM/uyoEc3ZAVe1KsdCYfS2kQrbLPybwGnI7LLV2T+wbQzI
I1mI4HmYL4eDIXsW9aVxC+DiUphJnoq7dmPud0JDlWD+HQAF0pfasb1sDS1sYv26hhVbNE5eNlNX
hG2Sq+VjjRiGiKum2ZLDodB8INAOKLH5XOX8TELZFJPVKW5qTKUbs3tTpdXrc55aECgpEVkeqZP8
nucxh1m62TPEW2jGMxpldmPM49OxoVNsob2x4BSsjBdxJOUiGCOG5k8CXXz4sw7ksaNlMHEdW0os
Xt1G6MZToYXZmGclP84gy049Ud2XYCSTIxUbunWnQV4U0WNNHT0qONDdEac4rteP8yqsstU+82vS
LwlrT5uZjeh2v3qbdyABYCiABwJ3x5bazEqOqJFfNkcR11kKcKrX31tkcMat2vzUd3m0E/vntHle
i00J3QPbKKcOAS/+75f+hN5/oKqyY1EfHOSuOGa58lMkrgmBrVO0P7swsC+GxLlekWtpitorxqH7
z1oku26yPi2+xjLIcqbUmdQFzAUmSs47elMt1qv8Qtbq97nXszaTmzc7if1M2EegGGYZieVJc43h
/R8KUeZ7pm+Vw0PaAo1ORtChPjo1fDq1lfXyLRHDtbkvgCgC9khhXivf3sl7uD6zF7oZ95TZUVIN
ewqYMv7Lcgmogn+GRz0REimJZBWJdpNWGnt+AhprxgNG/tMRfIdqOUZd46dbcYkWNgLwmSsWlaM8
HRfnMBtDZcNEIpDsMFk0k6AYLcZO2D6rJ7YhT3lmF0VPIYDRNiXTPctl+q2SNoEqVISZEWkjmRjk
KNbL9hZxIwHTRyzVg2jyQB8+wj6OnaPhC1K2bsxJoKtmrSrjh/2btrJ16zapqw6w+wGnn89KHGvk
ny6Fg8IYazbq8Rh5xRjOnoeouf0kA0PHimAcxw1ZC1fhMw+q0+8Z0j1t7Q3C7TDKyLUYSORuPY2G
FdWArhHIsg1N+8txwuztzRjA4Zj12tux3QJOUR99U/eLwGw58Q5PSvhgRNFw8yv+wvTmvBBlQT5p
tDcHYIYX8bTn5GccUQhtjZHCocvJMGp3lMioc51hQuxV18kvvxyI/OzHjsF2i1GlCVQlz8x4AdXF
+2ZKd2imnXm6Rcf5aexHXNCqhwWYRG74urOLdqeLmdhF3Hfrs9UUCj3YxOn2qffLUb9YUHUgBZNI
q3XdT8tsB9UW9wGxKmPQK06HT2oqPYEuu1lwr+sbYW0ogdau8zQXta/HJcPbROWGN1Ff6NZqC5m2
MMtIfKkY7Dq+d9UjaIw5OlpBA6rnwjHjUS/o3Eb821LbAKgxAxj1en+nrw9AGT+KAjDMTFXn3xrK
TfBUAlIVksU6bvIuFacwelZmloQ71lT3ALghK4ZQzc1ocpjk3APQXXw8kk+qKsXw9A+7NTC+AnEv
x42c8LZnqOT4t19VdcZCqVG+3bkCq4nnCfFNtrzeTz0lHLXEfzIyZlPN0td2S9QaFYqCaBNruwYS
9uQJiTfa6kfdgxXhOSjr4+02vhT/2eNYQPqRrJB4zuXUl2K+nNV3A1Oc0J1ae2argP1t6GyQLrI9
EA++Qrz11tMFplo3brxFMHBsybW/UZ9EriSehb16MqloPf+u+QDNz7BeQNmQPsCDRr7nqNbMfSKo
VGgIfGVEV6Moh/C8i9toW5TixfgUveOf+xCKE39LVMrqUimKM9mKjpAMOp1exncCUqe13sH07g85
QV12W9bsY9mpS1+VHop63Mb599FcaIjKIzO4j7q+g3Lr40AsTb6nJ012T1ITyPzaBlJ4A9cIZC3a
rU0vOsGuIQcUBkJCGdaOuAYZEwXYshotsOGGi6Bvo/oDzSCEoYVvGQze/k+YCNSDqkH/HGPBGRNr
Vg6WY6Fq9R8YO4SQjp6gh+Hq26Bo10sKnsXayQqQv5kfp3POvpBH9E3QUopv9Ju+TZl6jLpokEHK
OkG5Qhrk4hMQsatWfjv3OIGHvwpOU/svdlGft5CHo3rMkmG2fgYmdIdgJZcOPcRufywkzQ4GvzNw
zQHpay0ZZoxZE2Tw28hTduDOLU9cYwKnMUKA2bEVKTlZuJ4qqWXSy/bvqn/xvMClAdW2JEd/sEpf
z1D8CZYHkzL+3xzximke+ABeuSYu+ThTqteiJurm3M20Ccf21xBIm+TBQRHvjamuRDrBMDN637tr
6beCmkXhWmQsX5SuYUJBWjY9aSjghrOsnzA/pGTGTuca1Gq3Ds1a75Z3iX8oIwwy5xV4uet5Mv2U
rP01Wb9+Lw+seOEZeEx5I3k5hbzWF0zAo3SSqFzMzQWb7+DwjQLxhV1P9PUFlisjnauVn08Wyid/
WfX4Tz9Ckb03OeugvcqroOTWG1R4ZefPrkSQz4Me3eRoxAEd2u+c7+8fEpvmnx83fDvsIIbu2fvb
U9ZTrPzkZ0Beo7NvCOETlAvXtdC/7F+sHyRsUoBVDCWvSlQ/dBCmqRTvuE6VstbO/2feez4N1Svf
CQMgqyFn9eVqf2Bpjbc5/u0RleWW/DNcRWElyl6ecYlaI2rww58gEdLoOxOPdOOPcDqbEwVXgZd+
4bLy5zZAPHZPXwdqjh/JfowtF4Asfgcv4nJkgUOWANJwmkHWufhS+oVzVKYYeWik1/5uT+DenInP
WurObej5UdYJjqolrEIJO9S61UJ0WbEVwBFb4HknwQO6fjFa1urSiD3LmhTk6L/WKSUSWk9F36CS
AyiCgVISMgiDFK0VWF/2DMecttsRQ7s7/sfjQ3X1hagsRlbwwjA9RvUPPjs/XwWcbcpEE3uGOJEo
8uMiopwv5fjxb3TML7+SicxHfD4wpF7b9K5HaCBfWKiHPsk+m++pC6aU/RfJZEu98M0u+ZT+D38B
wJdVupMk4Pw9gFwXIz3XsUeIfH7GG71r8oo6lhoRsIukHGVGR5OOaQC+yhEmeHFT0XYcBF2ih7ZW
b655lhmxYpPO1IKIquoZJwR7hdt9yNJfuJADL8dVhiGobvvULpkN0oR9Ti8xkL9G8xnQWqW1GTWe
7cNySqC8ptRzyOtQH9V+xTrjerIunYBo+PWmRxd2IHemE913VjyNjEbI84aV9bWOuT1gbSMKQFpT
oSFZkh3TwYvvKFOQyt6yXNAKRV5exLBzQKA+l/UKY3Dg/RbRzcUod1jqUhqfw27GLle5CUD6Xcww
QBc6KoeleNuR4nd/BV11SAc3PD4G1f1BPqYeZRzraseTXvuSppl1CIKAGtaOr+oQuJNEzMEIWmr5
Dt/ku1S6iKZW4g3mIm8Ka3QNSI1tsTwy4yDVgIhftxP6cd8J9metB3nNhOgjYuLWowA2dObXF3gm
MQFIsbXcwc8wFgfNwQF2240YGsUUTB8Mq2szbEUv7xUP6zPE8SbCCJsIk+ASK7lgA/bq2r/v7kBJ
2PYI2tTwkWvFcz3yH1DlWGnhhMqVGPVdPL6IwEJDMd1DN6dtB0zDdPRydFMVMpvh36UkXrAkziQS
xc2OSBzpI4E78V4WUB/MhJr9AX+QgD6F5d4SE4fE/mX4YcRCZCljhrnQTLzCtH1ouEDjvXaUSfEv
xwkvbuO3jACmkaAxmfb87sRXr0T6+zPRWrxZzd+L/j6vuXYx4TfPGbcp/xgAFs5TWE4zBFMlzGuO
l2hmSd8l6iBC+Wx2GFaCTKV3s1s3zsDfc9E20eHlUQNnnEWqCt8j4ycvFzyYg8M5/TKIXTW7+W5O
cDZZu8M8Uat42Q8a9EsyOGWtI4i+y+gdobz+qaqHo6wxtRsZ1S8UpH0QNhbjOwT4VqURZdGr2gYg
sfnbGNvaYNWMKPTESpdqr82FI66lYHF8xg7q3ys6/eh9dpuQ6kB9kSY1WrNO/z2koHZ6H5BYsV6B
/AlhPsk4a828OpN7ygu/vXtsc4f8Xi+lmJ1rh2IWDDZcWt/v7e1BYckcBttyvR8eeZTwV4lpmvln
HdfyPflgYJiI6PN3gXXJjYFw+z4vpfC+cHyqSAcpvJ/vD17Mwvtlp0zHfH48RZolfmePRZGbam+w
sp1ZzTQ61h0hoNOsC4RMrOVcnD45T6fzN2fOvt14ABaPPtkW0qgci/UNS5xZ7+Wu9sQY1U1QzQ2L
s2RsNq1L2hZUhcGY5khjODB7rmxf0d3e9C589vXJz3UhhqPu2gyZSSRQEXL4WQIryrc0czUz185s
c8I9x9ka+9BW7qyzHvJjafqhXduUUdVQGeLNQta0ibsxCsHzuogc5uCwbMuYUFDY89R8opX32Y3s
GTlsiLpf8DCz0Z5NDIwWNXQD02MuTXzMbx9gSkZya9KXYXTDMzrizwFLP+qvgEHby1LHa2Ug0Vzs
/p9qe8OMhPnH7/oyIVF9UiU8cXqb3tkLOThLh+4/tQb883u1quQuwzlcyoHL6df+P+KUTeYTPt+Y
5UinD40sG/SZpgiOKDuR2hI1vfVVTn75MVUs2kH7RYXQOMNpaLIfvqtkVsWFHoyG4P35JgbEeKva
mWlq7q+/4q6yR7O594ease4Ke96rIBkwV4qoCLBI1INMtD+gbky0h5CD7GUcq8Uc+WkyzaQjgsbw
8F5NkZa3jOxv0vqfaCLmgX3+sJ3JnxXYM3DQiB5QSZpRuqG65jdjFJP7j9HAejQl0n4Lpm7TwzVX
3C6/3emZk9O1Ld0+90dZLKiL1yTdfk5Mdx0L2Qg9EBmQc80BmuVIlsivTB8rdvxFEXwAGKZxk80G
QOavNpX1vTOKxmLHYQ5ZpqqjLDfrC5FP+Z+WV8KeLSJNgf/zT7s3rPL/BLmeUniU8uSoDb/ohK2H
TjxIY6nPZbHJQxRpeewMa4EbTBjOIqQXQuP0YJBWWm9bxoTJgtj+dOg57QZb99ZSuwn+dx+WrwT3
tMC6MKdQxbJ5RgTi5h0VbIGWVy3sM6yZzI6yxtjELlOXMwC0+dIrG8E3j14uqCOhr4+O52u1f7ZU
VVj8h+02OS5QVQdnPtTbmMHu1I+3BnV2D4EVktbU92wrqNXYmFX/mghxhbkzdYESaYJL0SVSFLP0
Y/YaUlQxPpn+/caPzzibfcokr6CerdmXku2aqgaFkZQx0A/YJm1uE9PH0J8rvPfcZXSTuiZAVH5T
UCmoE6LalsmEMSRGOVD0C/oaFHnsSL9UTsDw5b1Rz34OBmGeikxkjHOG9F7PSNnP/cSmfsy9fhwW
8BA6XhoPrbj5ecHGBiRsrY8EP2Lr39J5Qf/XrqPJvk7LTm9zrOkvoeZzInC6ACM+CTGh/EOoIgW2
zFjV2qTl/lV1zsNhtP2UB4yitMIfFjNToVelZXi2DT1Ow55/CkmiokaUhrPMmjBml6zlTg38OR6c
64rSbvvgz65vuLnB8EvjNEJD9JxwbD80cDECobZ8fetI4ton8gqc3A8RzGsT0W2OdlvFlBji4dY5
D+U/p3I5YfoBXby8z19q74kfUWYwra6I+P5w3lJQcyuPo8JJxCQkn6e6eC+d+Vo/KwL1xZuADYlx
GZawZsYu6EOrzRq0sp3Oyne7Rjj5bj0kSrBWci+UbTteA7XEmgtZeoTOq+lbTPGOEpwHfPqK8T4n
vuMRFV6yycRsql7WSdnNcT4V04D7RzM0Az0lgxJkP90OGbRbl/XUAAyXhoBXfa6hNH0mD8mjUFLe
oAYNk/5SWjlCNTgb97RrfoOZtPqbFYEU+VvlNYPy2f+8YdBrniIYvqnMPneFfjr/RfhhoP4MitN1
lXyEyHzLO66HZHCHdVebS5durjPCPbaP6P2qNMARQdKCzY1wEBBJU9xaSRugHvX/Xs9QFSIovwCY
h+sMSVJqEPOlwkaUtrUYpweuYvRJ6+zLtUYOguGREIyRTn/dJLX4fhqYTk9VWS3kaifPso/brK7L
edk3pzLQcylQN7GLZAYHVkrku0ppTjRwKKjegKRlfZcTftltHjE4aEfgvLTNM1eGSbjaONJvlEQD
HItLwjgpDecAgpSsbzMd5SX3R71FtI3kNbeIZjMd61oF2asvQTuABJdwAbWZBxGiJWkWMXc/EVbK
TGWgO+uBDKqak9Xe4IP6aGMSaS74FWQoPByn7d7aiPH6N5JujKuBARdnuvz/5I74SbkYku+5lHl0
vp6sdpOEW6byIxIR29hlXdwZfN5uaK7xXO7LRYcRI1XhJ5DVzNTKgLgFaRCEwWnsjrbjdq8LS66Z
3TXtX/LSCAgISMX3BF6HNCqde7YJy0MaGlMBs33BQd8hWGwPiifZRaiOGOEoo6IPN4HMXXapIkC2
50sQTFDTy82xeIGfyUmRI1oVHi63SxUgZ4lOTam+QIKGPkNDUKprPBkVD6y+YyO+gc8Mzok2SK2t
Im60mUikpcwgDKJFoo0QV80PGPtBdQFWPu+7OCaCnfG+ExumU/B+N6au2osMza3ltV/ISzpFAR+X
2aUBrg5V4VKO7ecm1BEofDu7FIyVD47NvMGsVtSd3HkBOyKv+C1+zG9Sm1FwubP0iID64WEuVDYM
EOd4eJH+KBm97VxdqkQ5N4lDgHqTpTcG4S7coaS+8Ud+28lT9sSzVId9fzNbUmW2KA/Lhmz26q/0
vizeEuOzkuGFsk5KeZnBKp4KC5mMnjOJ2YY4xeYzc8erWFO4mL0m9/z5HwmaT8VH2oFt3radkkvW
SCIeTvQL4id+QGGH2ubL1i0FgedMwJLsRD/xuhYwiY8mcWV93yLlfQlyaPj0TmnzsA++1moqjiMB
bNFrNm9nyKcLjmIPTpO90oWWfaK2E688ktAsOdcZ7kfHNXH243Dnzkpr5xdMOzPTUXJ15Gq1XnCW
kaG9L2O0UU/E8VMY/hwGWJNLxTaxN2GoPdmQ5tgW4G0pQ5TaVgcgND7UF1ufPar+1nnTFKZoPpe+
6DHzWQDAKX63FAIogfYsrVhuVt12aB6JuzmHR5R6aVqWImAU9EfrDPvIuxGAGrWewFboLjOkveBJ
LtYiCwEvMpnmocoVtMuSrHwhRFTlm/ZNcb0KKbilZts3RJDHf2WlQjmsyNmFQlEh5chjQghghctl
DHyPDBoy4lJu/7Xn3EHrG6d/9i3fhZGeK0y1BM8Ie2QdhskEGtWZCCFEClOBxtmmB/wk7VeHNxBi
Z0+xhBN9CSUrm+/7vfzEBlKrGZD3g5zeRzWKdvlkJuNNM5zVGS8dDYXPxPCjr52OnJ6r9wXgDj2+
5ZbIC2OmHGpEy9YDaDwQhanOrjOUGwQvquQr/hULsCl/E76/t5OO67t8EcIRDXr7TuFhpAknpSL7
LJf9O61WkQMese93VkNjBCuY7txIMY9J8mhUswDv5ORWGfzW5fc13g3xaLTFSwrgmxRPzDbpY0XV
MhxA0C1MtNG/3W2KK1oJS2J73mfJsQ8AqEk63aTADmdtPBhs2tNxcJ5c2DYwnZrOIIYEmZJLapTz
yzRPZFYJ6lCyXGe/JGuSCvJH4kb0VY93OKtYRcso89J227eMsNiysviUm0laO3739U0CJBDzPqJ7
JnJF0nUrHzpDjcbYoFsP/4CaQMRtVFrp9174OCAxtSw4S9190Qna0pVcpZdSaElkvOVd5bGHA3SN
iVCwkBRbUFOZ9v2iUHJYEhEsnD2WbDpuSfy5YGIUfRqmkBy1TgVW+i9Pt4JBtq1TQV1Jkh0sGG32
P1RHxJxP0PooGdM/qzXeYNpMhyBqsu/NVq8KlFX2BCgKam1E8g+YQBKlA9/qdppVeVkeZa51SYf0
Wk7tGI7rwdRmCJIbR/nwCT9Hnt3DHhPun9pVUd8YKGsV03OBGD0pVTU4wfYLvh+oAg2r41TF02kb
9YIWpIkAHE5FqoGEEl19uA1IrFU5de5iZIYJd2B9qVU7mTzJQ2Hy/rj1ClX9issYMEKs/FIa9N8W
ED1O4pAekPJxKTY0A2OdIxPr3o6ZvV4SKn51pvjJxGQu99mvK3FskyTQM9Z+OqDCEvL1aBBXhYNS
i/KpFpwbAtGQ3DCTOWk1VtGffEjsKBGIzd4w0eu6tf4C4W4fSAPZ/dhqojTnk+wDd6QuPCu9hkWb
O6dosUSxv9jmi2B018pqtHLTGk0M1h2PRHqcywuqoq5YEcNejiagXuZLr3wBeW7iCDzNKTBlwqV+
RtZ2MPTqmi/zG0A9NePdzZ3hfWUmoJzzYzqaO9qydmUfsj0mO4PivB+/Fp6WNFPK7CDF3otxiiok
W/Qv7UNuNpwJHjwqdYIjfaaKky1b80hlkxdUzfrnCycww5iladFlNW4rJuWWNY9NeKaFzFc9mUhf
Z/+0VzTXrYIgpbnTKxNBr/Qveq/rTLm4Lco5hywasI3jE+yGj5kqS9kSdjep4/r+wG0ut6O29Psc
ND/ggj6PLtB2pSNLxnxFn9xau+aFpPIWH3M8ysP+EIDXKUNDY8bKxE4ayMdVRfONgi/VRo0MOQkU
VWLj0G0ddYVT7N/5+gcM/VR/eJrBBrP+oxgwjXYHO9k/wTdGy+K7cFMveRe/TPQP5T6uCcy/ai7P
Z5c0fD0K3t4mgE9K/Z5BCl6sMcpWr1RgHzHqa2QvVVK03VfMHAYUFhkeGuuDGUUIYBZWDQ8WjwrF
cugMwL0jKn355f+AaZIhml53pjzByzrLomuhgOoGl5wq+7gz2Vxo7YuApFGJjAl2KzaHzXL3XSzr
AHqduljzci9++jFUCRn0m6NwpnwJZdCtJ83RzmvpnuSilUlar8hiHPUChz5kwjAyxxXdWIPKQN1c
XnWu3gvhYj7c0F6wwWrm6fcDb9pDAsbiU7LoDld79otSBZuXNBsmSj6jWV1PjRtoUOoJavfsRp/5
fgXb9jmHdrPIiIgQwiajpNk24r/FYXnAOXL1m0PyZr5mmMhL5HzoOHB3hs6ZZFJ1H3AFlE+odYi+
8m9JBwQOYHgfwoBuX5M/vJrUPDzfoz/8mocv/l481bGUhHxZ1QlX9bSmZCEX5HC6/rm3BRFT2Aa9
x9n8xPDY1CTsX8v/O+JjdQDVq9CyAIxqoQRarZQ1ZbUeMauJGbLZP7ctY1zBj3kVLpxdjaWWONOg
5vA5y104U7IGXr5FyVnd0y3biILOZY8DVFioKS7xi6tUoLJqkl4GfLLtEyh7Omxs0f6c5lk5xlWD
gYptfOnc7b78NJdevhYEOpLO9ROXjvl4AS2A8b/XjuC5wbonGk1q0RuK8e1su7uNzGzbRRp+oEVY
daW93sldO4xB6YDUwXNoYebn8LMdGZoW9h76jtGbIqVZv+fZx+ECio17Bgm5EMaLvLVX+hqKj1XZ
Ra8fQnfuDBVFr8uqce1S017eQj9kWqvrPwbin7nXXA3nZ26IbTSq+ub2THdy0QCHTBinusRKIgeV
nzOFBj/FRbfTPxY+Eh5JpDdJmuPtoR4LKhSdeS/YxY70ZlLlsqchDF1pKDG2S/b5VUoN7CHWSMa1
X+BBNUZDCLrkRwjpaXU+oiML3Nki9Vd9vrBvODvzE3BlBTxSxI0Bx7nG8YBxntFkInXsBhiJ/MYf
icd9UZw+3hr5wf0ark3T0ke/R+5Ni8Ub/moQZ+r21dC0JWkys6tNmqHdyXHdE2TpUsGo6t3MoXP/
ujLlKHlaWHMyrxErzn1p3hLUMEu1r6p0d/EvZFN8zEJSYiW92Q/JWGg+hctU1JeCXrmhy1nkGSJT
m215HjsEfzhM51LQkuwhqNYLK8EzOuMi+/lD5WTkAOP95XCnwbvpa2uOv8Y+IIAKYlqmMZoZxDQa
VNDUzHrLs42RYaeMF9d27eVYYTKibvRtpc+a2Y/ZevK9RIQcJlvBxj280ymPrbLpWfZaQqxO4dq8
0CJrj/pur8Gw4AAKMw1+4lACReJjN7jC4zKLTaKmrd4jq4df8QVxspqYkOAWwZ/hg+m9ZHVvPclX
xuZiBdEAix+2DQ29pdeqnNi/zYc9A/eQ+ooI12t1HJy1kU2jC+D4VVW/Q4yUzP3xHMBdPbJMomhF
lSTRLtybJhqKdTw45eR76bAlNbJh4mrbsjpw4CAaadyc4gZ5FYuasSFi60sM6jTeF+WxDGsYhUEj
EdgK/f2iNU8efnr5fh+nIF96UeV0Z8aVv91fuHfdavydqLt5X48aSkoqn8AC+cUcs+2n/zqsN0Cw
0k9HRDo8o8a1I2wpKaosZ35KTGNvV/EFuWri8olYSIj/QXtYz5pC2KGVC+n69NIRN5Im4g6+Dtde
MqavzzWRQdhdq3aRWbnKe5DmM4qGraUn7S+a5Gi4bPty1GLYRqcfGu2p6NhQIQ7W5s24RMa5o5F1
//MmOG/8l/7rjXrkJnmTtI3Cd1XH3RHXH6ALbfglXUtRAI7e6Mn7R6MU/s9QtFLKMY6GOXAnURyd
mIk9QDj8fP49RuOLPwzYk3FwfXti8etGSP2SHLzpb6IzxPGvDt4KqMvFs35AedFbY+vJFoqp6jK7
rl9Gqfwd1Qyi/r7sm4e4KYxi+e7lN/IhJ6/OtDfSA8VOByo/IAsl+JJLEviugWRbenMl1RdjO4VA
kPOq6mLfDNC97sIAv5TqTFztqrTZjW2ySY6eU8J0PHHzlo4tiJU1QhyP1ksUVRTWS042PpKtFA4c
w5XB0Idn9IF75eEbsgtYiSm/TT3kq8LWolpf1wWvPB4mjj5LN7cJXCA7PiAT7K/OtD/XWPjG/38I
jWm0VtkFKXTg0fMl5LxCyX0Hb6Aq1uDio64/wJrlLNiuOt16GxY/O24Fj8wvnKh4bXBbDmHABSfU
bARYI/J4GRC0rVXrHqAsnKU03RIxhh+IR/HiBec+4itovlDyfUNntmYtM4hX2Pyu8Kvar/4dNb9q
QQoInSgMykJFHnNiJF5gz33P+LlpZcj6QNMDrk/KkXBluym2c07h4Ta+4aGCPwR0qzOZ8dw4tjJ4
7MLKptrYwpAFdRPbEAWOQsb1VqyOcV7zx3MbZIUWpTSvFPu4oEGoApDgcaBcuxmCm7V8SN+k38Qh
2rMXUlgp3CbmX61M3koKTodRWaMPXzihjTBFJja8w8zBl9HewZJxRjAln9T33QKJUF3epzQcgc9P
ocSLFWL85Kxfkzpg3fvmzCFyUbhEl10R6g2t1vrsiVCa8BIDeAqAvtP8mdseZWQSKZYTh+IrnzH0
WQFppBExuJjvQzha3jmiuIU9IIHXRdD/cWhwHmihfS/kYv9MCjiSX9j/C90bHN7OMsyHSei7OMtq
8/nclKmeoBJ4l/oYwZBYXjxPreuzh2HXvl45GXRy/ga1bJjbqbmddWgiHOaSg6Hxq/D8AE7bussC
rbuwNNO0WihvH2aqOCjLisavB/+TqGOyUvqcBPafdKYi+R71g3hZC36OEB5uDqa+52EVgZmj1zHZ
LGNofoRzTH29s8ITfh4UO+H+KAzE7crhpJBgTfWira9xE/JHWNGSaq2StmUMe93oTMyPFy/t6rpu
nbD6rYybkvucrOpSxVwGJf9/+LGpEeMCwXyaR5vduCucLv+wKj/Ss/2aAZqxgt6TeT9pZci2RcEO
0jIy7Clpn+Y0X/13mtllRs00cI34d9bbc90tRRHZiIEDH1PGzvabF0vmp9DGo7BzQTUaHHknpaST
6ZDZbNsz0FTH+jkCE8yMTNjmbTbLIK3ALOITrvQ8lbpzU2rLUuOaPsq0GOrRbvcp3J3a5Fulw85L
Da5+gATq3Vehrukn0M9ZD5fHYIVuVZKIv9M3oZEh6RzU/BQ0SKU4paV9tReGeuFzxHWUpxLLlOfG
DYsms02ILY4p8A3DuG314EEGs3/yp8DO0wbTtf3yUalPSRvBpNWxgGPSwszdAXZVD6hTB6Pt+4D0
FRkwYHYlpC11j6ocMD92tOdCvWaAFJR2NLmgVr7xTGfIIWjXM4UnanwP3luGtjUUy3cAQLCupJUO
P/3OxiL5P1Tx7tffNnEhVBmFNQFhz58JujVIu27R12VWyUcqJYPVsKqcIK5j8ktW7Qxma5p5KgQp
hj6/sWQ01sH6y6hxeHY9svtaNw+eFQFPdZSwPhX7uiqsLfKZdYy/xCatR9Iq0QHYQC1n0tKjO2FG
1g6L8162qBTKaSDxKj/yFAHHUxBSn393rnXC+HwG1VHlH91GWHSbRqYffsJeqlz0RPlNjgIXd9lQ
u4DombKNkpSmEhwFQgWmRD+Oy7GtEoxp/7yhg83iFPqxAqvO3N3PVCOc4imdnF6jOrVfDQvqk7Dy
IjU/NWy6YQf6thtBl9FBCyxU/OK9ofm9FQIcdtk+kIpnDpgUEC+BRl9d34u5IXvpVH/70nziWFM1
A1VcmMnDCgTPDY8OSiPd7UtmMQICDBndAz94fS1pxX24oN8jEm0OwKObnOP/KFbHbEYnhXUvXfs0
cmozPRYx8Rya9Dsq01EJiAfDF8Mu+PuNsRTp2brWRMW0SBF8gErwjJ7WPdwX83KlePqNhGLLeiCF
QuekF2EyIP2U2PvW8lhOF+0puZePOHpS7HXdmNHO/YEvJIlIDDdAuMKJLofPWUCrkS4mZucE5KU0
rL0nHO7txKbNp5mvvSVGIgi2FhOj6upUfviNtGGDi7JONAXhEhUX/dz6M8u0hGSWsUqhJXOtRaoQ
0sZsbmEoqIh3zwfWhqQB/A/z3HJuyBxvAHLyjrXe1XI05uklkKFojGX3sv5i437QrdpnX3e2DbBV
LznLYI96doUtgUHv3hY5SN/P48ivUhh6WBFw8GRVOmc1hAMipNW8WiggxWsmFudVVRWfahN9dxtU
hPX8uLkFx/Mlw9AnEWjYd8IoBDQ+GQaxthqCZbOOn42kjnfz2Z5yrfL7Op2zmedXQHlLIpSzJTqe
TvyWW6bmtXxdWhvjkddSvgc/79DK4FquzdNkpBKHDomoML9sXm6/GKP7OixrBfysvxPWw0V1SP8x
DAsKPLaneOPhI6+XeAFHTQUIR/xmEyVeFhjeVAtETSfoHoZu6mlAfj0hMdT7Kf/yZeEVSfEetsR1
Xvaqqa311VnUKeNhcDQjYHAeQaxsbaG1pgIdAjIe7NTIxSE/H8bC+kLtiXDBM68+hWhY+GW2Jp4m
X3rWJzYdACrwmQ6EC84XUvfzlE6xo8/c0ZUkfoP96K/HPhNLA3NtZVW/8e1OeMZX7wnBrs3SwkIJ
xKOFA5UhROJUze/FSpGXfkkii0y8tsS7uE2Ua4CSVKPbvn9cC+xuck1cGGosaPeSioZhwUXwCT9d
ENcMj7cLoQzEnmyCWdbn2Lonns+totEBv1Tf1JnMC8M4gm1J9a229Mr+3/JWNn4Qc8LhhbHGLrqp
1Bb3L4lmiPm/M9jrRH9jmyHdMcHLxII/bYGTdCcPjzlRKPcy9lqdrknO6GPH326afCXQaALIhPhy
96BOK/jqPyiB3PwOqwEnS2wqPzX6zkRVTG0Sxou+XXm080EIEkUncyKbht6Sef3xEHrVUSFHE3Cr
wQi5ikGSb0i6cLrALdgVHBTAUgucnCBr84Wz7e7xqzWSC+mIIOQWr9VK1xpRu5y7qMNldpbsy7fB
jrVCV3s6tlWSUIF6tibAdKTH6ze7JcSYlRS++enkU6lnD9FDpePXDD9ZHo5J7oU2VWvAuIjwUOHJ
P5vZJiHL96YMOcdVY8+ny/jXXROih9I8a3b7N8wtuf2PJ158QtqYThN2zVi1H4dRYmavO/bN4Hqz
WUWVG1IhYxW/kvPao+3RUAxetG4oRL+nP/qACMZKQk7ePEL/+9uL3RGMNNE0G0jIdzEel7/BZcxo
BIourUS+D/6DDnww4yCkibR2XP3lc7FkWM87q4J4c/KvHBOcnlJiNGPTDh+h07t/hXimEYjBQtNq
mn/ZH0P+P+pGo2xP3MwJ2Y2DBNkkyqbD9chW+UuW/j+pqFjFmE4XY4wwyG7QDQTqVdRs0YJHrOUd
Y5umLvomlWHKp4uy2naBgQtF++8VxbcnfqJKFkTqRbRn3l/sjEK8X9N2Ux1khXxEuF95RoxmLVO5
6qf/5juExXFXGSiSutuaY4VEJwwU/fqRAkfuIEqlIrtIJJm1N34Zj53DdYwJXPyXrxY6zcaL3DB6
3uvXO4sfpvDzk/qc5ebZ7vR5p6IZpxuJvbAR5XLQfVYKTpzXYXhuW6QYRTkvi+zUSykbVS9+v0Ah
jHOWRK6ViTr9W44bl7BcfzSyTWR6CYLLfpLj1gYUBcKTi+/bNrFhTzQ7SgSmuC8URwOY6IP5rucf
VAInJvbjBXtWjvZ4h1LWnz+slrzleyR8BsDJ55nf40yltyxkdZsr+2RdvtQJlES+SIG6bXFvlaYn
Qdi515N7VaUn6jLnlzPdcliBBcBQnxgeLb8RV7YyL3Kq56/5tduhRVb7k98lbgoYKoifXD0bq/LO
VXPEX8Yu09MbZ+B4UxaZ7wpKVMiQtkqxDRIGaSGD3XIUDD8/zmYHz5Fk400nxtx9hLiEaH/epVPG
YsK7/R83tF5RSyCIhnFo8we0lq6BtKHjwdtuo0sd1E3WBXkyRX4mh8ZOwBmrWFh5h2wLP7cjI8Qc
dnr5lBpAd/qY6N50aO1AJpu1/llYU5iUNgxEGmjgqLzVQvjDwQRonFGxKFmiZM6dV7+JyuOCKC6C
UaqMWpjN8qz6MOicoBLS3raEe3MqZW1Z/rD/R1TrObfeLd/EQsme5joqXiI8+2zIKVsYIEKeXn8D
3TxwW/3RTIOqxy8hu1DgZMJgwCXyq6ANAxAIENpBa2dnIRAj6yZw/j2wJV2NbHh9PdkOYt73YnVE
fgXf6Fr52lsHyoh1hwUHJQQXuheM2QGIb9DbubquxCsc4TMp+wQ8yTR/5hK9rQSpsuTU7VAeHVSJ
B0f5QUaxN/ufI3cVvnbGlfGo2Pk9mMDWc0NyIGGOlyIJErvs5qXWwygrx6LEnEzxyZ08oP0F1wDG
1cXf4SSsJ1rFcCuojPdkM2zKsDOoLfwy+0tETOqxOONyAggUnVhln4etsy62i7OTCVINbxczgeXq
M6lNqgsxCChh4SCLbK7D+/nBRTc83rWZSuRXILf3RtTEXfbTqZi+pae3hDiojbleEBC9rC3qyiT2
Wymy/w4F8W7bsvMUS26LjGE4I2/9ZFm72dtLX3l9r46kTyOLW37yjFL3mjzNxl0tAzaA8YIPy8xI
aei2augvVrk9DUX3yz0aW9B7OY6PwbnimDRPTa5GiiO+weIGYxAAd4lonjwuzXd22mf2kAidZEBg
d/Y9NZ01/KRqtQg1v7aklc+AOCJDwcpQobvJt3XUw8J4YTrZEPw783HTkZRZiGBKhHSHFj1+IsQn
KyL/yJhuVBjYNQXTqcUgK3mZmkfntK6gXBhJJGgE6DlPusx7opPBQXTcDvfYu9t09ePTsgAzEYaS
tX4ubXy7Zw9sCgUC7FVND1tkDrnBiouXgdxSuaB6l99gkdZKq8V9PPWLSTVH1sjv57ERl9CTgs++
/Wl+3r27kscRf6OsFflvBtU481fIAeGupRiUYrOLoYiEyHnCxkkegCC/i36jZC1EvL/wm9qfzIEn
UngzxaJr1f+cMbJF8J5hJCcvhby7bzLUs8jitnsqsMd64gf50IXh8W/tZ2MiWTZzG2qRFjCBsKQB
Vzdkitrg3XHsD5TWJkQtt4uyU9GTj3jI5jpvstG4CkHr0DPxC6otiG8KyOYv45bdSg8LkLr1OikO
6cN0ps8ROz+R12FsRwM2dBcxDpkv7sFf01drzR5DeVD1dwNld9N4QKZZp+tZjQStVR+CiHNErLtf
0d5BtUiyU8XKfqd9QUzynM4wFIryax0LMJ/RgcphuVIQcBfLjM3Lwd3IvCCC+RjPczClnimmQYAg
00MrSCwiistGwd1S06L8r2+y42hqE/lDABfys/W6g25fg4HqlTvdcccEobMuC9jO9z8HGLQuyqVE
m7paujKtms6NnHoPRMfSWGHKylXenPyTTiPUqV4a8olq6XLvmCvuFie8JebHoyynCgj1PfWvi/yJ
mdKBqgR8xFgYlRVuIOmwH2oI7iRvKUExv0X3Kfv3tARveyCjrXHa+BgUlkAovs0PI6AzPZMy/mIO
CSWEPoJkMBTIXCdgQAPS/57dx+fRuH9x9lpPbSYvUn6da4QpPHmic/Ym8LAhO77uHZteG915E6zA
luFl3dVS6sqocCY7hIJyajrZQaR5fCBUssFUlMgZc6PAq6Rf5/+HYCeUEvCSL+6qC5YvX9UHKykx
XUe6gIM/WI+/x5YIYYoEZPkw+vv1fL3zb+iDQnQkMi6suSGNbYy7laRCEie1xW4rEBzuAut56UNN
JPAoVLOpw6TFsbiZY2i0laJbfN7HAQubuJmNPhKYnZoShNEjvOGfVwhrws5gccW3i1w+lk7i6XKN
tYqk68gFc2XaU0PJ8Mg7IkJ0og27nINx+M/jXZFdVOKmsCizIdqctXoM+WOTCRz2itl7SP+qeyvj
c85YbaZyqdYJSHiCZSSe87LUjrRFjaS24H6EzZ1hppefpAACw1H8wATvLquBfK3Zqto0w81E8cct
4sthfZIsxpAJXLIrOdAxgoAMRd+Z6i10BoZCIPumcRp/4SIPqFGGghlrnQqXiv5XhYFq/tBRb2bk
+3ATZfUOc6RUe8Ea4uBeHrllFuq+PUKhL+//HZemfGY2SUGNmBW43y+Mf+BWgeyP1Eb8LNZ4pz3A
Xm2E9qWdTlW5HqVRafEx0dH+pVtLSS+cDpBb12dkDIHRz3Iw6K2dkAe4eT6AEDsJFbhu5ptIkls9
oXZjAd4XVucf+XL3ySXz29u8ba+rYTT/x6qO5xDv9th6/igSBLTORFgZeD6SHJBPYBTG0KfPvWh6
s5QjsXZwHOyyZepPlA+WG3/ZAMuowzQI1NFsYEgLw2rUTtLhI4SguJW2FmD0UE2wgDwOCozJ6S2V
nTMMRuTfGOwG+zv01svnq/yf+TjUF1oobMqxN1MfPMjBPPeA6hm5TVHzkai8kS3xbBMzsukxjR9G
yHYyNRhWt47ZthAhZGdeEucQoLyoi49r38brn8Ew7+cTDOeb86SvOYjjhgobfiu/Zp+qSiM76ND0
2SB5OEQj9ddqfE2SELa3J0kRuYwv1j0D9zPunAY0fG6ADSFmOALURF8b5tBGIILR0vPhTMCcklwB
lrGa1EYfHBp3vgFMz+oR/b49qOG0EIUGG3D9EOIw3phbGDR0LYmP5PyWe2goMfjc6CxLuL/J96Sg
vKsZf2MNeQRFqTkh9fEOCztElhXlj31l/JuFewMbkvWUZ2wH3eDqG4WhNUk4+UElQrZcAYTsc5gC
EDU5xIyyT07Xof+BTCsTPVDTyF8/7/KREJCR5lYSjg1X60o8s3eEvQJZTvtd5UA8O4ANE92sHPk8
JDUAczOVFziN50kZJoLiPsbNJOkxjGvGu4Z88qgUW4Y2CzK7T6q0xBdrC5L2nW5tnC6dzD65PDak
eZqzwWZtp2W4Bx5AquQwMQ9ONyzb6wGlR/c/ZgBG9nmL5ct7V5aK/VbAaCM0ifsThVkX/7MJR5Wk
HmotQWela2Twx7I4l01heFa4rqsptevhDRpXQCQy6T+SBiMplzp1S/JTuVymUH7mqrh20TNnyh6U
iPf7LERLihSU4bZxYCMwOa/L+bV77FAbhq9iwfBei1MgaJ/n0bW3IoI3dKiAN3u48Tkdo3AOw2E8
Bicwg8y+iIxp0Q2zQh16aP8FECuSERQWA4v1C6Dfcw0CV9yuOVQrlIlqskqiSRCgP/kFKu2aEXIS
j2QJbV0SNrv7xCUGN4TiUysGWVTU78UIayRq2X1G1cRdZfRbP4poEePvR55gBD1N2fZnH2OE90iD
nwJifxTvS3aWBMfwkcUQ+KTb6zYyc5TUn6SUQzMRWC0FQ6sKQqnLNBZNb1aS27FbF9P/Q4hLT/Em
/pILTvwc8FQ1q93IKz08c8R7SVGELOgbaiTN+OK/RbcfW6YoFpGKM72MTAFgxwgUJFZ02A9+g2px
BJ0QLQ/bCzbaYJKq1zYjxFHJ+XsQt6un1+9MdS5I4HNM1TVdCLWxjtc1zkJBsdAklNwaonOtzPSW
8L1L7PTmVrzWIJ2chlPQ3x96rUtg8y5Xk2+KpXPNKKwclPVEqWVWtTfKJq7+pjMoyAlP/J3zzQiR
iLwPf6CIzjDkWufzwJR8WFhE6zZZN2pYOyuBx4knquicQuyxJvBh/GBEEYq92r27c+PCivKxLEHA
N1M6h87XRHKdoG9ceGnqnpamRKMceBhbXi106+roaOFwet0UDAFW3vPOq1FwQ3IuR9aSgJpSEmP6
OjgLHaFcXxd3UjESEOnTMKiUqz+VXSUa3S9q96IrBV7usUbbBoN2zEJEYY1skO4trImxfkFTkvvT
GwuG5VAgaZLp8lF61xbt12ifbj87kCN/dN7EHAqzx71fH+siLbjRZCPFSmiye3ieJ48DOIoDeskY
AHMmyNaVGyGlk0oBpR6IzM2VJz4SsKl6CzyGi8Q5Ln1fU8ijvudWXvSG4kzKkNbHPESbqM2Y9s4p
jvRLGyRuq+OEeC6Ojz7UPnyZc77J2G/qw+sRAxFq2Vpv48yefcvd3opxI7AWEJ1blgbZsRqTI86O
CU2xCKV3Bjsmb5sws2a1xYcQDdUlyl6BJRdFVssHucfBazKpj9xLhrrQLVSOMJd2b84tg3r0aG3L
HuODxOFbTZJDShhWMKrGhoOHzqPy44AgPrYISfsch/vAUYZvqovQMZs56UxLugXH5xQrwkte4Afo
12YqvkfXNmTmz2z/GMJ56/WnTDyZAeQG4gEznxH6FDEuy64FYfZb5uJgkAJFx6QefWgXo3bEZu+Y
06pQdvl5FbhG113mikf0gziNCMKXdVIqq6Gx9Zyo0vtz9k7cnllscEutS1ecpDJQCEQORy7X/JGV
Zl/6+6XuLBJfKVJnxBHNIa/1rsljudRpp1tiPRbvvoNE1pdX6wvE5eMtsGr/5yEoLAgRCQF8v8/T
0M2h1SMRtaIhjmvsLq/NsADlJw2+TgoMahURZL0wsdW9BzfFIWdPFqvwgwvdIQw5Jhuk4tPuUAgw
dBebSX6nKauO5Nzz+97/1/xrVR7u84QXKVTHssz/tAOtWetvJM4hbuGvsxpmBoO1OOVSIvLHSbcA
YxbbqqMtgxLBnCQzfhabzyIswgwNRPQs5EFkkp5Zh1x9JVxTkNPGYtP/YjMXzphC5E0xQDDGZPwf
ViXYD7OZSI0NDAJldnDekxWDQgSuXCYvbRvyGsyFyuP/E6G4y0uFvHOzIInhucQcegQzZBAty35V
HpvYQVw6CPDETsMXEW9vsVj+Z9saJ4s9ZKjaIOnLRenQ09o3FRFzQiBmL/Ts8H7rZQ1C1a5gmpcx
QxVF3ysFzVGxGy+wa1zGRSlC70hOXl50YdURNoMgOgoA5f/96vNJ1XCVxlnjLBL0I0/N+LqWz0OP
uA8MJ20AHRRG
`pragma protect end_protected


endmodule


   
