`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
msjbjZZv50JwJc/jSAZFgHjwLuzGlmmvPd7YlgtBloDVfyj9pajPbehofJBf5YhKGs9srLlCVW12
vA+syZnNXkKUu3NH8toOWofvb/eIOOVBEfOWZ3ucMjZXuTJATdn3RqCTZn8H29vJBdK68TGPRvEc
N+UJfhpH8s7FoEf8va1jh11DTU9bWLxXD1B3KFLFR4xquovDQBpiEZKJx/cfb7OhNiOW9gehqWp+
cuA5KugO9yXXuEZNVxmaDqg+kmN5cY4iSFujXfv4YcHLgl46bCPu6+nWj31MrNOE+4Ooot3FaH11
xfaTtUTTjrEGSFQX/BZ3FsHlfwqQoaah3//khQ==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
E3lpVoLNkpaySRn42M8E+cCL92lSO0H6HvjUB5X1vjgVvQHyO2W4K/XOSCLq2/c9vhC2JCFSNF68
j/pWe3juIaN4YVxd5amufuUvOaqmFUZuQFv8NiMjde3/bav4eVIQWbTwSWzYtrIDvicF97DZOUs+
azlp+P5dFWFNV2AphU8=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
KhlLXUIR1c+L9PiSjHzVec0VZR2e2QdgQK7T3o9d1mKhTO6IQ/WB+pCNmjQTecS/zduS6DrPhnKe
9VglvEuuUuzk6R+EX1JhFlpXPzn6aLK+EB1bt07zQySl6Y+6aYDRh5Q7V2tHf3iEjeww3WAPUfmv
Ipy765ZQoB1XjmSMLYk=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5568)
`pragma protect data_block
ck/k2gHjsRDT+qQWZttqkEMjSz2ogyhA1A5bay9wgi7zr0Dd4oXCTZe9+TWJ2D3bg+ddieppP40E
DmCm+cvHOcBTweeRTGg+ksF4Jqf7zC8pTy9E9dLm/5/Mfy2gLFHUnUyIxK52qFxZyq6tX1m4mBRq
ABfx7wFtw33cHzmSggG4V/duZrCV3kdhkbf9GWkOKyHrQbR7vmEvqrZ+Rk3RrDvPySVZTNGPebR1
X6dgX+YbOqikVmVFed/4rmVhXsAv+3QKsludGGPBfxLQ+zkqAWZZvc4iiMQD9PMBzDwMpZaJHmB6
Lw/A7/VeSNEQmEYTXS+Ri81xIjo750hp103L7AKP1kfRXrO7m/xMeJ0PwLXsQLRD7VZdNnHO7nlM
HqEZd+RpXYHaCywQMEPz88hj+XboXjCBpT4sP0G3qy9AigTKddWUPXrNRwSs4pL4Dn6bvKrChKQO
/qHX+IGWYp/LLpF7mcS/O5rtJBzoyJPKdiGxJCIwASIE9Chz6u7b52nQEarnfkSSOzbFXouwFtIb
nGSf/18IKxuVCxB2OVvgaauF5wpOPSo5OFbdGaX4RRDW2mnRaTPxi2FW9s8oSiAu9GCQWDwOyUhd
S+VfAn0pwWG6nWi3MKSvv9qK5aB2c6IJXoV+FHqADA9Oi3Tg11737njuXT3cul0vvde9J62tvSL/
XsYLO5zuoLQPjpASN7hQkIKFZtwL9zRDuRDg7S+8u7w5//G2WbzjW5BEN+MYYdD7beUUvEOZuxP0
673bTaq/4EJaWbh6KLcUmL2aTfBIe34EF9pQdv9NF058m8+couQX56K3b1FTigVQqyh+hkPRfH3P
qYoJjBOB8Ce9P7eR6ukI7J+e312KyTEO04OFls7pJ58gHDe5Vq9ABJkAgOz1ZOsHqYFwCiR/5tWF
AaqYXw0wIM+bkBtuxDWTNyJkg7D/yN17PTIRu2rulb5/xm7aXhNbIWZWLf0eA+GpmScIbC1A5fHe
wArKbs0SWIqMU4moEAR1MLT6yXl4a22u3OmP8QZZi+aV4K0spjzG3Id9sfMXFNmeSm6mc+r4/J0o
MJZ+S0aRdx/aZJXa10orLhGRzGKLXOHYslV0vV1MVXALUzRAjxjOE79rtbKpQmUpH5x8my9ijGwL
jONm+q3qlvO9/5viWsvpbiGKUCk7tUNEqEQ2H4zV9dSu/wOreQtVYE8++agZRTPWzqeKbPJPb4ZD
A4TZcl2+XwE6kXLGx/zvkkTDrj2HpapWgovSy+3i1ebn3RgK2fE1XAZdCz4CpvO7Vk5OKpdyWmhj
o8tFLYTg6sWAc7qxv7PQ6dx/RbDdggTfr5FHxQ1zlALeQe0SoNoFXDkt8evODcy5wSN111RoUv/f
KdueYI5uRGZ12VGLyvJHRtYmtkc8BAQJ6V/w7raxFzBIaX7mhKOYTZOmB7MfkJo62SI5VPkOJzTC
rnoyjbve8MuZYz3yMCviNCt7CJOGw8pPmjF7RnjfBNf6u11tujayJU3LpQWTyfS2K1dG+2hiklvg
EQ6U2tPrGQFBgHmrH4GNGzwgTuNuDmsvLbOBeppUTrIJjC9KwqCiUEklBAG19FTFwXWTZ1XlIuke
7eeAmp5f6RIGlL+0fsnlSLh1V+hwIiToU5u97S2jGbA0cabNP1CaiGaZuWi6m82wA6e9mutldrJg
hS2ZqcwbJoJ1lQf9tbywq2h8rhmWYMpHPo75k262CwbZl0UKxE5Cb2OgsIVSgBeRwuXAdNXoNRif
6DN+ESZyhxU1/ZLei/fqtcm/v40p7cSmSdFBmOernalHr00X8+V96J9UTHrMHTQBxl68a3qT/W/r
1vwoDqqbZ6zRiT5YKm8VSbdQ3DJgszvNy25hVY7+eTmwppLkWCXYiNGmrIzWA4aZoLtvXi5odxPL
3FyTTYLVkNO58svdkRdDgROUCElV9oWQm0u6MZTpMzDBaxGgS+J/kSNall+VRF/KZRef0oP3/l9u
kKwmu9c4TbzpO889iy58vHqsrytgMqEvx+wwTqWJo+5uDTwTpgne1ZsA78+Y+DFp64kSzZ4Gr6v9
Dm7mjVTcDVD32S2v8xK4vofqEB4zIqXpMNTykwQOc8u+0+Y9zqcd4YeJKy6Ow49EKBHx6muxSxDl
9NiprgrDLeAB30olVLZO8AaZ/8KK1Zyj/RLS6qOPYi3Skgvby8m+HETjFT0RWBUgeSm8JzyqLC2c
er+tG7Jo/Q00dpYuNBP9EmadINrlra0adSdrdoES8J4XMSh5izfOuOeAg87oESgwhkvpVswdzEj0
ps/8CVizyiY/HVIPfVjmZrKfDA9zmCNms+bk3NLOPUW5AQU426sBL4vQ/mZahJhuR+rNQLXTBKHn
9h1QLGvz7ZJagCpQUshMswbMwnt30H4tsWafAYqxwM/WQf/aDHGx4xx1IBO00naez6lhvA5tCYUR
PtPcMqAWKAgW5aOxvwWgkLqPCr5pWq8tv+17/tcw0Ghcl6eIrHf8n5urUTE2EgtljGTj/D62JUkM
21oK5TjbtWDSS0yWZxipl0PPuvmVBdXzpceabxnvHWTnEtz+nR00V7sH3pIhS9nle+KSkrAu+YqZ
4LhajG6obz/zDcTGG1C1GAOpPT+TkOFNZ0yjIycq0TKMbspYKBM9O48hvs1T7NXFN8PEOePqS6jF
Qox2pSa5PH6Untj5myWKsrn7CvkAbve9hkNE3ORN3OQoMHWiYL2fLmEhtRlMWUvaaub/tG7bL9hp
FNMS0MyvIeKcgUK8mdoF8mW7sl9IseApHDcT7O6e0ZjjffZMEpJfzjIYaQjkugAKv/oGxrET51FU
43PKEjgGktsVLF8dMHPkBjLsnqNO/uXX6osssrBsrtz8bRq1X4mOksK/DjyclfTg8N/5TFrl7Wft
SpyDkKBFGjd+IBKdjb1cYkdzVrdyiMAk2I3A9e9rP+Gz7FQ0ogykyw8bK1oB1ATqs+qlCUvE2027
/IbNU28JguZ6qWeLB0qN12gVXWoaptrLKqyV0rSeo5N23U2VYcQNxzrx4sUKjliWPG6OqYlZZQO4
ipSxjpKNU2QneFt9Ke+ySLOTFqU0ZbbM8+mfVjFgrbc1/TWSmaa3UAry03sxQuj16oYyh/1GywqC
CXnujmJL0ClSq1Bd3lHVozVypXR6u10VNQfeIKoUT0z/bfj3+IJib3VJm4EICfQUx0UBhPxCJyQD
5p/nxUReUQhVu+MVCmMTtFGQ2+33qmmOmRgKto5+xSYwOg4cxCgYNanoUrSE66ailLI5wQMMl5ay
uirfQU4KQC/r9r8C7uHevH0elsTmMzIQfe48JDHntkIT+6+M8G3l1tXlfoVzpgZQnJfdlJ++Lw8k
1wW6S64qUOQtkUuGbuZ7fLTf24y8oCtP52QbwpcKIgH/nXcSYiAMkCfYZM6iiDD1eFPksjOXRiO0
MyB1uNIdJp+79G5SD/9Fvw8PCwtAZjmVm2tOVg6JuOaBKVO3ndVPvQGnGw3WCs3wMjDYMB+0u8gb
KO4fl+g6sD025Nst/cr1ri36kn+gyl10b3Zqqes6L1ffy96Dz0jphQTJlcU6L8TCfuulEm2bB0O7
VeWwRVAz2nxB4Ybt6NwRoiZlByPzBQaxRCWkLhmdx+00WYEGRmZdv/wenr7/3p/XDMWB5UPpGQZf
jk844CSZmD+widPGcPJr6TpT8ggGzEcRb4aX/b3ea6z+48hKFnAnRUjSvWnQdXiVAOJXRrZacpnS
69wobsLMxNYG4odoeIQPDI7AvnLBXG1lVy59YLoFnd0Vc1gDd1FdwO3TcNv8784N/30+Nt489lsY
ggX1LrvO7L0r56BQ9T/kHfUhv85lsc/VrbZqmkR+O7yZKI0bVhxYjrTsXIm+WR/SAOB45kee06WU
CofkamajbIi5dYbtUJd3ms+R1fi15pg9xNB9u1aGCXC9Yhowc1aurr0ZJPrGYWwUJtUb4Gi0ba49
dhCwCMSucVdvqgcsj8aBZQP1WP6lznPXmmgsCXfjMbuvj1nr35eAqMqiA4LqY0/efIeGkl2qLmZA
1a4XgGr+RWE5agXj69UWHMRF9Ft6XuNYRNxIP8Mms1UA9UGAYjpLoq25Im08QkV1rTfVm3chqY5T
wZERouvgDgjEdCj4i6L/y7QG2k/rA7ycWbjpm+wlTrjnJ0A5slND6ETqy4WI4QaBziUrYQtrB5q1
fn/njl728gNkofBnaLxyX8B5ERpQwau/IPlhUwTPRhpBIFQtcgJ7iCK50TtzA5YpbBMxrc9FRmyA
hkV5Sj3iiC9DUa9EK9LxMF4vhJexChy6d0UKtBC56DM0hu2wJP8rugscSgUfnooUJLK9+KLwPHay
EbByBJ6rBJMhh2s53KX/x9iWKhcnI6a2DtP8p8JRdOHgk03vqbf/1ad1g/EIAuSHCs9tPYPYE697
RlGCUxV8vJzXgvR0uqwE51z9TDzkRD83f/tyro/jRnm/YnAtkEoKiNmYx01wQ4m4vCSVem/JGhAG
2PFjCF/qPXpaImXaKGtKX2Sx8k4+J9h+7jeeBQ0vO3ubj0Yh0Re/iAIL95/x0nPfjYNcw4cGawWm
ipjeEmvXQuwuiMHRCNUf51r8vxQivfn45MrZQmEb2MGHs1KVOVSAxdfDmdMaG31eEqJ5xWd6lARE
z6TtuIAgopvfWYOfzLGEb438iykHIsRmSgD2PUVD/In4Nuw7UDJuDPK2aVHyL1IC0P5q2gNRPf3I
5r9qPvLsmtigga9NtUU1RUC7sgoZXrCXoMDPiSFmhAoPs9gDcA1Oh3iWX5ZuHMtWTpH6v/UYrLJt
AY4fkreJmNeW5iMPfJ3jhuhz/rQDBs+IierqZcC1zfv7CcFa2Czbn3tbE13GLJuAFbHLAIMdH8Vz
obm2RaAWpNRB81VvmPzIeCdMcpsjEkejWg+Dw1/3EkD38xAc90tyUV4Nq+7OKfmb7rFVWuEyC9y9
r9jwcPIV6f+LWBlbcDSt9xJsmdNbVyGiY88E42sUbjRcfV/XvAL0nuTqoSu80tbAniwHHTjYTuXh
31n8eTDZTDAaYvmn+3Fqi84EeRCJLyxuwAeS3dcuhY8IYJIpjOMLY8/TnIuflquMI8eGG9bVUDYN
y3hZwuXhwO6lkwvx7EfKs5m+J3QczQWDmQevqhGGG+295m1G7QZ1LDMDiCWaYTUiPpKXCzoTMXiN
wbfRELWQnTJltYKrlWOU0bLSeYtbyd2773iPP9KoFy1OwAePz39xgSSALwDOEIBa+D+1/Q4OPdv8
iUFmQWmqHIP1ApeI2j2foYmloHpwMbRbtdmsoWqiR+YHR3pa0lM6jlObW6gy7QD3XI+K92JyANVj
NB61w1wmgBh4RESujipetm+64Gxvs6P1h77s3oKCcMtVbl6ur9Zz8dCL2x8id8rvDlu+iNKL9HjR
bHkpY/aoBhHO03Uo6+v/fpsEW/JJRa0da2/uilhT2pVll2lFpjYRjSDN/GUUeWax5u39YWLDEjgk
N8sgQ3XzyguCTnJe5opozLZDpaqeXHpB+TG5ej+rwnoqsTpK72GoefKDs7Sz8EDx37GDiObb2dyk
NoubE2D9U/yFYtb2gk+WB34IbXNRF/LKyErDEdiDpDPh3dt+POoPGt+m62XfPByvkoYKXeTXgcG7
pc5N3DsdPxUronCA1zANeXlw82ehywKzqSSIPc5U1S6FW+3IQZ+YEjFSMelxG7lBCw+THgIDxavH
Re+t4lDCjiht92u29MpsPtk8MFde2hhy6FU/fQwQBjWEMePNPP9DbXrMaM22TwHADbQpLSEgnmAB
KxedGtNOw0dv9GFbGxsSIno/JNvhebQVfbv+ellS8+fAvRlUu61NsI6JRBNhswRWj9gB3X9nz8Mp
xxHBzI9l3THYq6V4QgalmsPuK3a1jGwzgIflmc5dWRgZO40ZKdWFH9tJa/Wq/ppnoYjmbalaA3df
geH8tiuzbig60PoWeBnO164n7dCdxUx9NfyshI99br0YXkodeFjmqEHy9ejHl/EcxeMrFNh1n/5t
KOOvVIQl3rfGHXXxUuwgGSnPbmFhZLSgaiNfrjN/I3QyPfvWiKjTaYKGh5JwMp5gNC+SxW5rjWwh
N2Q4zxWUnr3Zy3AIVgWt4I8lwogd69T7aHjOiHHkGCzxknDShu5AliqDlwM46oe+spBSRgj3iye/
YJ25ENDwZIpH92AhVMHwN/+e71eif482pnAJhrkxdmFpHYoqNHRkxuTirdiKy/aDvs6vqS36Wx8y
q5Jq/CCBdPLunDL/PTXjwgURH3lvJOKDuKa0Dg02ZTPTL5xYGJZOyWAHJro2P3SrxPNJ48x+g89b
0hJpiHib7QVNDb7rvZXY5b5Pik3uykwsbwk5Ro9P4RjVTwbMILyjs9jB2TkF+zJCRhuffaKdKsW6
msKg+Ruh+OtDOqG00B/rfuiyX6d7O6RJcW+aqOwLtEHcF9UypPTRIwR6EYdh9ZCn93hiEs9SK5qU
vChQZWnGu9QMeP3FYdA5y/XArnwS1mP7s0xLn45GkxLLPzS+bh9pnACKjp8Wh9/54emiOlymqX1A
dEIdwftQR7Xfty290Fm5Y/owaKmBte4NT/9XhHG7VhTgZ/VcLGjsNPffJjNuufoyxJNqoPT87cqO
4wsHKdh2Ggj+ZdmBkKvNxpDS2cgU7LoBcogDOr0Jv0yyDuz1itSBnL6gnxcAGt2zfBNUbMif43C+
GXkEFwRYFrrVHnDwP7RsFIwH81KtjPUYBvSL52lbKB9M1l7Q5akSMoEQhKQxrpptDFB8XEfs62Ca
2sKgCw9gi51dopFhevkUi/eHF6Om1b3+rtymTumb59cSY+jt3IjUSxmKj0LHxJxgJJSGyAGkzIXY
tSrjbHZvR3f09PkQUpZd4SfUTHETOJIDRJbq9vUTRbkeBBFYoWuYXmVt6hhkZKo0h8V3iNm/bjff
miiKeRVYdCpD4unj4w5B3GpfPnT/IkDEhFcQftKeFpZLxe/PEICtCSiXjqncq2RHgyHfQ5vTEcm5
05rk0UQDwerk43EpH3A1PePHtaGkSd7oHfFvCgoLn92R01iVR8iWJBl4hsiq7tncLOXlqp881WxX
5TcJvGfAHU7X+bWxxZ+jrQ34aGxYX1WZv4p/lU43yxamjh1z+rpS3bAfaWDewKcsnM9Q/bFr9ZlH
O5m9ktQQtWAWwbzzpYvHsV4l/Cb+m9VJduNk0N5Nl/LEuVSrtujhs4nMDtNestFHs4yoZot6BWYx
QajwiIT2b0daSsxepw4DClf+xX2vo4CzJ2LY1wAuMVwpGJS+w3WJHchCL46myE+jnGByOL29805o
sy77jtPN4ZsB5GwrQpm1RBzBZO82D9xJoh868pB+86DbxyO7wxjbr5V2p9tPf1WeSLvV61cathvw
aVElom34JeU9MxHSVdRdm2LgMoQQ36Ea22Am5WUVvZjd5Tby1dU6
`pragma protect end_protected
