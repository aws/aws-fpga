`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
OfnLbSkNJvU+N0FLARMxUmp4FdKSCnNVQpg+fWwku8C4XDDTrEnyDe/tgfyDA0nLuAyWkNmuhQdS
EZ1RZ7RBVrE3kv31CmZRqTqfBDu7l0xJWSZmdhedYIipaRXMNfLT0vMBSjfGuUGFtqhZiZkX/911
V7dpUU7Ft46nJaZdZfz5ZnQeC3siV/qTBV247Dr00rwzBB5MyEKW3FIfR2H2Y3+4SyRvwkhrHY6K
H9nLt42ac3qH4UKQ/XXgbV2oXUdL2PX02Q0mILkiAbbb3TfJ8d0Aox6RwXl4BJhyiga0azEIZtRW
9N2HcUE2t9ssyKnwe0Rx4jL17Gi5uOx5S31ApQ==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
lVhLpHh3CuWTyF/6T5t7P1X3K99JRb2yBGhDxRtht5jqV+ykOfX43qFQrDeJ3ifUwTkokPIiRq7q
0a2T2LqJiDP5MkKTVfUoLmjpYCdBudcQYZoTg1fCsKDa649B8ENossiy3cRiw+ak3r6tjaUXYOSr
1uk52hKA+qZL5M125C8=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
J8he47quSLbiY8zTejOVuCY7HjBp/Pgg28YVzRbZfBFavsGL1FFD5ZQFYiH3gwe06JZDeDKx19W9
IXN01QpN/rJyiHJAmmxzYmRHJxjc4B+YMftUi5kl9KWLVzhVn+sGcbQW7ItufIrohPt/QjCsIltw
5dT9ZPgN/NbVFNWOvpY=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5568)
`pragma protect data_block
YkjjgQTjcHsMJVp+BGRXERUZrdM2EtOEH0hcKxiWpZQuIy3tey6HRalPoRW0JaYdGzi5G6+Xiyd6
eHveD8Kz+rfaFF3EfYU2ubeBODi0HzO2qSRXkTqQooVZjCzMeDAWzJqg5wwr8FXYq7jfcjNh7sIH
CNo+c1x1JLlQJpV5r4vywdEAAHERVg5AGbklXCctMmtSOY8wT/zvNRrumyI0ptjfa2fgu1SdNE0T
Od9LAhy5sQaZRifhlxl5zJrFBcQN5vW/a34P+1WGhAiNt4PvlCQCOIh8Isn1+wWk59hE8L+XzdQO
wMFrqDa/QGyp6NHxCOzEXJvZ6yyBe8Kc7mkWSSoiRnB3wCiyKFyBIqxLdrx4N7b25dKQcOV8EZro
VP5wO5X+rWm4EPUoemaqp8ekeMthQQaYg2NFXgQqqBNpbYuftcBtyZj0RgVebz8oRwyoXeTdWZEe
eEWYeIcStkBZVzoU+WDQ+Wq35WMafyGcUpgxfdUyt5x7LEKjJVrjW18S8Fqcb4RTCse5ojgYLMAo
wR2X/liFxLols8sz5QUZxUp+yxmxiDOGLPcza4H//Wh6G6B5ZUK1RMHNHVB/NcaLnd5ruKPbgPBJ
v67E48iPRYSSTzNAMT5oRTJma9qN9aSXdbdC0jCNLtPAYfWUhU+ykr38kKbNwzvQ72RSsX55UUI7
aVSOl2KxAdKEoAndvf8k7mnUVRO0MdO9MX+HHBDFgCl1zUa67n7PUPj4qW9soy/uBwWlv9NGMFRH
/RY43GssSa+cNG541h2A8M027puXHs8GIYLMoTWHZ+kYUlU9N8HCo54O/K1ecOG3S6X83l21jacl
9DtxJvyVUiVOZK9ibVP2LNKfKXaHi5dh7VOI5w/0HbFGqYf5XOPmRlWgVg1OXKFqRLavqiftjPuH
epqea53wa9Lz0sfJHTktbXxlL7dOZ/9Aj7Ww+Tev9npVTCvhUowI9NJ3u/YcRZVjQMD9l8Jg56if
oh7Ojz5Ffu+j2YdhlNWw1/ZZPeKWAnmZOIqNxqxz3SNSmEnNxJdFSHWAE3gMC+G/aa/zju9DRyyQ
gaf9xegi6gly5qPUSWYnZAq+4vKrdw3SKl/uXrs43hu8ci1t0HCN+1eiLwwomJo3JwOnPPmf5Ybz
90hFUtFvL4UL+qPFVa6Q0n8qw6R5BmPUVciBrZULZEDNGJSu4o6CO8rvfLJpZzoqXtUu/AB9MTWV
HU7xuo3XDXpZxeOrnCkKO4/loerUzY5ZomFRPQUBQ6NXVJqFCQmuBfNw3FdCxo35s3ATyiV+tyvC
fHKn6rUMSSFuFxuGDeJ3SPhT8pNyJXY3yyHaWDwvsfBi32xbTRCVqvBGferbmLtNYX09J6V/iE7i
s+5gibl22XjmYTpywE26ul6R4+DTFnNuV6H1WjzuWXp6lmGhRWgXv+giMNr7PjLYlxx7FxE+iRFi
1OBrr0X9CaDXcODEm6WZGZ2rIKrf9uYS1VpttXK7XsPiKDsCWz2hlMzc5UOudWXJMy1/1jlBFell
oL8G9EEapcyje5sF6qzQBmoRfFyVYvXiNvctNpOixzxSeSHepeixk5XncRIoK/g0YeefqK2eVGYS
Igq7Kjds+s2lSH9rhZSRZiscacCkNyT+fZxRuFlxOOD2qfSXzq1w72yJ176i1j3fNX25gBTG6GpF
ponOV6K3YDhO/YyB/BHe8H7qqeq3prE9jPyLr1ebQj8mulYkGpw6EZJamPX5XWMZwDBVE6JVQMwF
fO1SZzENYoCg3PC+Pnqh4J7nVDvxbczc767gbajTZBaASlAUczwPvPstyD5geOA6qcOB7bHorCy2
5WQK3c5yY88z3FEDYbRT3hmQjy0ZzVEOWIUqonOmBRvYn7o80OrkW5JN7aw/0BXUi52Cgkne0R8f
eo0fhZx1dZ3gXjuoI/fQmAmOFZrUsRic6CSAhqyqXbBxIouOTrWoMm8Tx6DLoFfhC/kIPsJMHbk1
tAphs8CqRjKha9p/5SNGaQh/OTBmFgG8EH6ugG4ncXSrUi3Fa7T6xNnKSGBJoqziLKaro0A5m4M5
4IqATFP5F/TYc7twW4txGlJ9vRPkotyhCkNbNKXYJfUZ/KkH0Oz9fShDzTm8UZRw0E6O2t7olDaJ
Jt7LIrKGFFafNtmSzQKrIQt/xRVQWbVxmYsmbfoctnzNEoz64W1ygh6PufhFAA6/xWb+4tcHIcM1
GXW0DIuTOIDVAGyHeO1PveMvfd4sjuQGseakr4ryyjSzbcB13+89T5y8prWNITzKCWNqAocmUAG7
hIjfMajSYDruopb4j2USeP+B9Ux7hpDnte1xdC7fHmxaIO3gG418+qArr/+se/XqAAgy5SpoU8YT
VBhyDO5w83Aany8OFQWJjduC3YcWuXySM/D/SsMJYlTs1JoiNgThK4y88Zg1rVVTotwt3prAMsHp
3XOMF1yItAGJWEYbum3X7zlawNQtwLfzBIZZ9gDVyRqoQMuapZCTJA6B74JvBVDFFPK59smmm3Du
2c2fqdwpF0uYkZCH7s1vEQ5cZEXEO+RtG7sZzQtYH37mtszopTds7dJU7AQaxquzYkszhSmNY+Uu
5BoDhNAuORD5ncppDEJflmXwyqMNXK2sXB0bkXYEyzKyfN7DVohg7gm0P1dRpPX0cn5sjVQKaCoZ
tUpYq+XGa2OnP8sMmXtbukoNQRr9kHiFAbE9Ds00SbqLD8QLTkeMxmxNbAjtCKo+dUVLbketulGY
39Se/IHU2JrWciXt1LTWSTWcEmDe/G4tEYKwD6VPK0aDPOWRtTZz/HRz5FQOe4AlhU3o+ifZ1maj
Ps2aIt3DNtnO2okryq9/YsnTo5hHTWyGbBtKmfrk+jUFUPd/JWglzqbK8Z+wPF8KfGpF2mNbyS9o
y0lNc8UZuTstgmplieIH8p5wnHbEWQeoMb9qRJe2JPDQqDacB1S0bfZjNVH9DtM6CA6Vp+XZm+G2
f1+88+54IjuM60s244Fqqw4wkNmgcmD9i0+4nQQbuwP0WHZj94D8cNv51eU7N3OffAxCxU286Bc3
QXsNEDGmsl82BV91elhIVw2H/KTJ2+ycc77ZEys7p8IoIC8tX+g8bvthiRDc6slREIkUcvFDe/g2
FNlfvwwfwtwCJV/dSDLyRQ2Omg+X3Nz1oS3biR72Eom5q7jQf82AkM5sZVeTHk5bO45fMylkfghW
anUd5nh6Ch0GkEmlPhIA99YC9ted8GW9ELQruTVMQrX4Fff/c+qDI+I3Ot/vqxlQwD9/2tsT7fgE
1Pke1S/wvaTTzBpbMBCSLJ03lkEKbqJ5/SgGPnlADD6VRfMNh5xh8Vc7dT4edOyDRk1RKtT8vCSc
sGM2o/DTUZzA0u7Gv2VgkHUfDNg2nCfUbBm6SHrP2yW7pMLGZGheRo33KSzZqvQM6aQy32CuA7RS
qWiPxGp/OfPFwNDcFLg+FWb56ifrQq2xL9EFIytcExyxVT0AaC9d9B1XA6M/mQzQd/4pdWsULqYp
K3Dztq0WsbF6KXFJg7sBIL/AcO6FxWo7tuB8COjgCZLVhZ5zJov9HEOUmoT4xv3+sNXpPwcs14vD
FLsNcGeSLMl0TFnN/8g19f+34O/RWuuHSfNUL+Gm1g8HO3vL92kIiZScbhXKnDDxi/qR5Q6p/Yym
iVOa7Kkt21k4Cc13awh/XswrleaybV+9tM2KpnDWZKn9twLwRSP2pD+oj6D7+8JpSDlgOstLM8nL
gSUqcJKuK4WibE9mccrZjhf/QxVFvsGo25pCYKWOjYo14Zg2zBVDC1OBB6VVvULqo9SmEFB6dc3f
9dm6D6bQeuZu/fuzENFpAeG4cbzIlEiCkL9YPFsDYTPIid7WXmzjzDKI727/4cVsQ57RSHeyHLS1
8/EwlB6pbmOt55DyJpOQYyHVyFEK2Ziy4SY6jM61ZE70XS/H0EtqtSvQ3Ig10PXqUCajKGAGc+r5
6zY9LxoVkmA5EklU8h8i/fqdj7bvfGpaklG7o7n3SwVFf/8IVQc0pDIQ7YisLVHHWSzr4FsnYY77
/4Et71XmyHFkIDGtEw/yhGwF7MkdCU2gdjXXaXcHQEkzmqPjbYy0mlf9TuDmWfc1Ot9eYncnE4JI
1E76Jr56s3P5dNGkuXHb5tndAbmsVWoKnsSlAof5Nb/6TdIvm3uDWhgErOAu3m3ZFw4INRl31YFF
b85pLKdrusYN5fs7Vm2qjMR8R8n6FaRp36TUcx1GZS5wRtjpmx64o25PqR1GVxaOd5n1CAL4CCxn
TumfRYpggn7dzbVONhigOU3Bzwi872+gqSf+bIcj/E/Zd1JayCJXuPTEdaHxzWetAZNuS3rypGAY
0rZvlJLH83cfoJsYxSWrsAoYmQzkpy2AiW1V5LtzbN6z8975TYTASUiYEnsW+3SDboYpr4i8BL3C
ogluVvEnuApIGx/d0nhF7dajWA8cbDOKLV3+VBlhKc5K0gRVxv+Pl4HUfA7bSPQB2eyOfls5N0RJ
+xF5iovbFdaPHCsqIVRvQLpyLbWEE9t52xj22/mJQKv14zyZ5Jtq950i2LoEIGItALTwkbJQ2IOr
700F5mE1M+Y26Pl56CP0zFthMjI72PzcGR45ODppCZezKssOyoj6OOl5od5/2ZH5/mZmHSMAQVIH
9+Y2zhvjYRfq+HNU9a2X7xqGi8j93hLJQnfwlqijKo37MpyW3s/ymoNxrX7fxzttvb8YkhqPXj+u
V/mL/r87iE6BWQkgIxE68XxXcXJZP1MIAg02M1ri4o1nva2X7Te3WC2QAZDYSkQMhlocFVk2LUOl
Z695bB0CgKQYNXOA8GJqSO1zuCI7aJ3/wzMQJD49vnRNGVUQZEORkQISLxmLO22Pa17mExTPOtvE
B9HNrUR6ajdijYJWpxr/AZNVwLKiocLWlLGiP3cSLjDHVgBHKOwl9HEX/qMce7tBmmLHVOlaIar6
M/SWB4/AqYR49AKQ16Nb2DS0NwXpvsYbrOTUuKv4O66FC4FfdXaJZHx6W0TVcMzBYGs7FgYsiC++
y+/AYB2oiF1Os3iVz0vWV7YopchsnysUfDSM3f0NWehzM2gIi8ANQmSJUec2aNNSKaogZw74E2L8
w3X+3t0aY7QW3DSr9OIQzZ9mQTfW4vyibcWFlIWoip4ElvpqetqEOS/qcu4nPSVoFLfO2b02T64d
2ANXjseyzcowfmElJKpc1UcxYVvc11SEidBGRsU7ztOiijagnvz7tGgzJoSGhqG0uqtngC6vH/0f
IESd9Xqwx3jHyRF20CGcku0uMG9QsbM7xCiaJCYPdiA4hrOPewYsfwanKJObn0M0hZH5PbQGFRPS
SrcQuLKqbC3FANgrbL+oTnuUE+M8wi3bAk4tpvkrW+mC0uWjVJ7sVVPzDcUNLD6RfyXJE5I3+/ef
cZejUqzQOIQgZ8pToSztulctbN72+xERzmOL7PIJ0006n2LpnKm7c5xjOHXJ6hJ6joAuorNM+zBy
elpOAwtUqhF+Fv9BGEN+/V3THxY3GuHUi76HFLPlts6DIu67EImKwvzC0WUza2K4HaHwC5Wm/hHB
V7bVneSL3+l3H8aS3csMwzk/6OaQMuInDteVt0OKhrw6slc4PAFMxhanGWunydjKbxh2+ReYrFvK
SbGpBDFOALl9VhOGeRj1bWbDPaCBqvCA//2h+Rm2jXP0b5lTZH9jt+jCoeAd4K6fuWKe+v72HReV
iucjN/F2y+WZ3VHC4BGXET1OXG/t5p7O3tMJnBwilGzX6GF9tpGK/dMmTs/FYyxusTTxk7MS8Kru
DI3hVKPwIP0h5QFnmfe3Hv7W68HhGg7HLFdHe0DDTTZakxhzAdjE7bPil+r+ARXxT29SYLu+yrAZ
CIPg27B3kv58B4s20IFKlaZEvNOJ6X17EjZyQJALK/2PU34BxN3xrUe4y/ll1A7OimWzq3E/2j6S
v+886F7g1Us3hzVpv9g6d8haPUXFFjc/y9FsVUcatHF8uyHdLB+Qa7ie6JL4ru0gmPjGK0SRWbJX
0O/l5BkiI+2i2DVQnlqoNW8+ULHfABLQ5zTmfQoRaxWAzJ0dvhSdNTn3y/YfNgUabi4Ph8PcR3v0
/VY75zPuvIn2r5XEfTRlR4/DdGg2sWzlB1SdItsA4A7KfQXMhGOQQvxl+kNagDPb9G8I+XqGPo3M
f+qCQ5wjAQGE7Gh1AZNmcUUOOzvPRu+tjhkwrUW+CQchOjH3KUV0biyt2GG0U/K9sSE1E1h+e5A2
mU1vtItYBY8dhDMl+ziIg7Pz0K9msI19inuT4Ra38PFQ2Rp+OESFBGozfg4ig4vWJmH1B7BCJcim
+TpOO/d4UUhDU/C4vrVfkYTTvVMZTMojjqpe8pCBcLvJq6CzKSq+AN5VglTt7N+7Hd1L/myjI8+h
V62kfMGTrnwRDDlCde3029frGKLG6TFKtToXEGVF3LUFHfu+Sd1qWePaX8IA8SBl9xSwkd+CDgqH
4RXZdUsCPwCqCWccwePd/dRkoaKYiPAdH0u0A68J8RjtvD6CHwImDaaz/Y6TcCxpP+9/t6AOvH1K
MJCQQZcqhn+aGJ+IL2+2Fy4myHtHVi2d41J6WrwvLkO7kfJurBR6T6eLS8PF+DwOnmWVdkaSmDx5
LMWXs39sD9Am9+vg5nIA01/mu+cHaKOP7BKlNIiTbNRQTbRU+HkS0XzDn9KooGGXuiKS7HMEUvRs
PwmMm/6AmB3ZZtt1g1cLOd6z9IbMBZH7d38swlYFcOsY23RQMY3Bj6VH9e0P9bfP8fwF+QDPcztG
mOc5dHQT9C3OGiha9QSyYghjJzpgoF2ncT3kiILVYFFb9+StlYqRj9+hksVJZxd7KpNxsr1J/ahx
78JPy/3xFlfmyJBab1uaY4NTdc+tEJXTnKSbDCjSkffkkJ5KmBBe7/jspfD+2WSUysyGZkyMk7PQ
9YTpzeYLzGraK3u7AZDYYNCjPBaHd1ij2gkf8TSy2weBPqG+eJS/9VJYHS9lZULX/ylfDOKLU3Qx
O400pb9x1H3BT/5MDamVdzqvbLt8yPpRWKWIpfhWBqbh20d+jy2XtobzH1nuqtlRwHykKLX/xyAB
dOYp2o9cEaqkTiLm0ilOoiGdZ2OqPBbJKZlsxeIy4njQSKpLx1GHkBX41PcEQAe8D0NFqVvqB1FT
GhKmePPczZTguqVgRGp+2YMN/4qQbxwKT9gfg3jemqNsOIX8+L64Wl9rc5jroPm2onHOFi7E/+df
nSQ4uw+J3DnsqbNfDOEEPjLpk4aUyoVsCkSGEM99ZIvNopOoM/7v6Sz9EdnLKUdZ64h1f2zXGQ5C
vxVKi0XXWgi8G6G90lgEZTnZd4zzqMcQhbwe/xqBQHPHZhyU2ebXrsWQhX9tJR288fpC9zPAy15d
2Z8fDiF7hVkzdyYkAGpb+DI0xkVz0FgAFKipcHrilKg64R0E6WsZ
`pragma protect end_protected
