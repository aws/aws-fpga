`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
RxZWm+Lu3LiGsyOy4YoCr//Mpec1THnquCUz9Dj4k6rhhKvCBvyHje8cLhAWGqGOcDo9tIJsAGMi
fDD/d4eUpxHLw7kxaXeKYvr3dlHIvEMqCvN0NC8sKyh+V6D3qivBF5VZwfZkPaYIDtxA/IGU8YRw
nmCJ7HwHhcZTw/Ey8OmSEK1Dhsw856h+ggGQGEzg1uzZ+26Xb5wlH+6t9hyB8ktyeYu9vdCrKWfx
932WZ1M1crIpEPJ3jbRUAbbwGm9XEl9EhnsUkY9SaC9YOOgbjOMaOxRbnyiSmYohkFFJQU4qf0Ql
1Brrv9A1h4Zrzzm4R140/tsePLdRUEFdBNk4rw==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
0RvF4XNqKSGIecq8GH72mw9klDA8StidI3xYrGL9Z8aEH/5nvBn18OjsV6oRqX4NQi7KPGsjBxNU
e6vzRIefoe4CgFPHdz6sVHc3y9Mq/z8A3nRpYar3+fDgC7RKW53F/F4FZGFTNoG3gmNW8Oy8y1Pi
Ks+lmDcUpKGzgR+YB20=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
oB1uxWvnpj9cUWMHNGY4+Vl+6ZP7Ea/zhN1SmSch6SvXRP0GM0w0bFk0NEmN6/I71abBjmvTAap4
eN+D7rdsOtfQZarZnDaOxM2KaiBW/IrYJ4AktUi1D7oyzv2UrqMBmjf2hw3vEpgqww765rN9H0qp
kwNIjrVFGhMhzBxMYwk=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3504)
`pragma protect data_block
P7rD5QvoefO07vDM5GxCiXCHSFwvL2X7wozFL7cHR/E4Vs6fDOGNLoVY0H15Sc+jTG7e1tA5FEdn
EMHJEL0GMl6R+Aqiz8+XyAGAAlYT+CtSA4zk1vB4xguSYIRfMz0aINh/2cJqv0P4x0TfMsyF0OIW
Paw/3DyEL/dweldRYsK6rrW35Ba33N0mUXAbhSh/ePyEH7gucM7mg75puRBEjh3ZGbWObYtMQmD2
/OmpRuVU4rqQ8o6XVeTTBI59xbibzruKxfLRAsTLVPzmGOwReRl4w+OdJQO9MoXunTzbN9KG6FC9
clPUxrX902p1mwE32wVabwYNZYXxWl06zx4CmdxyO0ddnIHHHTHxjr4tubCmUsNI2cc/A7jP7lkS
UHdZpkNRodwkWtVVJP0WprJEp+t17iv1+Em8Tyfq0OXxQSwIlcvBdkRevUvZNt2HbWHtSTRFHM5O
aAXjFK0Ez6viFNj4KX+BeYm5QjMHS/SGIjIwFZAMOGvqOsJUGe6gP1M911gmJXMRM5XUsy8PEuMB
h0BDiyazLFP7WBGge3OVejODSDZBQ/QoLuKbQQd5OtMsHZtRhdp6W2UFoCT4Y7w1I5h9Lo/sNYvG
Zsb3B3j/ObfoUy9OImuaom61DopHCjX+537gygQixlrC4UXRWC1A0uy67HVbsCX7tbza/2jVnUOj
W9Rm3mqgVQQPmEqpgeLgaPUhk6VItxL0eg8+Sgu9GY7YSD6v5LMdNJfPdOFqqilIcFBx90LWnRzU
BFuqOxjsT7a5jtIXZrB6csJ0wCKjPScJytEYLbGDA5WUVIzypT3dVlx8/49Fq9kxYUfZW+1CcGFk
vyU0CIGKH/y7xrqzeAXLTJ3uIg3eb68FkgO+vw9GECvJnFSt4DveSp/mVkcoKTDZ9mwh1H/A84Jm
z2oexvbStZUvyIxxk+np4IJnEYMyWRaI5Yk83w6N977nreszMo/hoaM0KsvShxzZ/77TymqRJv24
kq8ITSkc56XNKTCZjza1klwLcPH/261xdTZ/A52uYSHJ/vII2hUf+VD+qRCDiYGq72qGwjNoAreC
5SnImPjfAOX7GlNSn/utDHbYgkapqIi9UvanssW30lGvCxoYmzGii4HR2CJL9bRk61N2h/z0L8MC
hjVIvZERT6ep/hL3m4TDF0jMm26tgIpq2EiOpYPcDdMDl8VoKPs9RORTGhNKvG/HHHbZzJC+ao5s
kXv/DGbAurp9p1Cr1FvbK4aoMnBPmoXMXV+QESneKQBXW8SpKi89p4tqnl7pheeEt/BtwjVkuH+/
WOI2SyJ1TRV6+B1yqoQ1kcfLI4lGTInMcCWaoMnnjJySTOaJLPQq1WtuKdNqBttkYJPZ8/A9bnDc
pXmW5V3FqonZMx/dmhm0HLpQBk3G/JuwDnvJZAj1YZ5hVhY3sJDIJS5YL0ArWYMZYK7AoOT3wn7G
46ALNd4xE7aaSwLpap2XDiYK//M3F4koRo++FGJn9EPsJy/HgSrRRBWRKpSfb9IL3CV1cMn577tH
T5oyBRwd5tnKycSzSJETSppFL4hUUbXmISN8E7QJxJ5mTSvpay2IlKmvERVr9aGsKEk9/TvGM5NQ
khxZXhniB6nPEBdDK3HxPX+s14s1OnoIQdkmWTIt8cCk1dLgtcC5f0rPNVM51j/oz2bvKQ+bV3l6
x2G3KON3r/KQ0owGxGikbnsv8Iw9MhiAF8Ri2RaPG47Zk5FCxqwfJPgus8hWAU3tq8B2RYMlFkaW
CSRycxgliDQ9fDjO0aeqF8DICzN62zWJzmip+fePUkQWia603nvk5k3DSSxanrlXQi1duTprbzpz
ybJ1V35eWxbtbr7hq5JMlwpDApeUGO+cwLwFOy4I5JRt/fROLSYaDXsXBIyYhIp26lbhMdjhVESt
pBKrgJopdZ4h6PwMWdcXbipt8pLzuNyQfcPEnfrQTLyNeegeP65YdVVJOkZLWaVX80p4ElA/GEr7
UKh7N5c/2QhT4Ur5VkhoRonQA3eeLrwBvQSp7rPzDjrTT51UgDZ2AEjlAU8VI/TJE1SHu4j7oijl
zivmEqUkbClRt1SYHewQRv2r2KxPaxAKUtqCR//+cUwovAuPGHdk6NK7IRTVZjQZbJv+5VHkG3xO
+G+iZw2N9aakitZXSOS2ZW2He1VbnZ+rHKb/Yg+UKZ4nsS00HNoFDY2XdIxxdbXlNBSNvGS9A39R
Z+No3j5K3lrawcMh17sU6Pp2NXRtmFldecNNDSAiv05nOEz32JpYxwOG9+7l2dXJrMmjIzpgR6HQ
TjY/srMBUKEsgh4BlESGuztEJdk4GBSH/qFHOD/uGEw34Qf3l5VMJtwa5xeAP7+WcckiCshqwh5V
olifyvgkdkmHqsiJxZfJaYg4WFj+vaL4RM4F5Q+1mZujZnxsekq7OrMgHY/3smmoRkUgSdDGYBp/
97ovRzL8SbSHf4kN3EYhcNeV1WIiL1fo2zqcSKWvtwOpYQ377zFzIQTqvEKZAoWIvB/Y0NzwDaGe
3+OCF59CxoTXdspBiH6BoY+5J2DbJ+8U+T26sjAUH60AyFDgicXQA2aoVA838jC15sok0dX2dzxp
Sk/Xt64Asi1YFRepBN4n5cx5i+C2yLfW5CYplCFVs4sIG5kQYGcgSVywJYfjGzakjtdVbOJbof2G
Gc6tkaYj1ija7/kyH/AlgGxXp+OFY6X2/ow9fpENyw74KmNimXJPWbaVs6FEv/SN33Tnryh/24Tx
l2NR8Ce+2aEUaT/EEe+5abl1DF3p/812U7RygcorJXuiF9d/Hqn7yWCOHp4GF861XCqeXwGj9Ba2
JGEytynfQ95co4rO6YuLq/AVeJ8XXSfJcP+CSPKun6rXGT+myX3SjiwjPPMaSkXzf1PmQcBzMXNn
3Ts+B5MLYqajli0jIMvSlEzAsEKjVYjNKd6xGjrhUcLQA3y7pyNhTD6ox16GYvyEDO+mBfnB18nd
2BKcrLYUWRfJgS6YWLgj4cuikO0+j0xq3WPRYHH951A0dObDrqP+K+ds94mwZ8LY85p3OKeTu3S1
K0vGJWimRU6c622Mc8R5iZ858iKVTupWP5+NWwxmTP5RiFJfH5HYhTiGkfg1a38qO0blTT5nSm1B
LAqqW1idy+5Ryctz9LNTxu6nxG8tXDEOgoJLdijbaOFUl3jeTbXkb7wHmCYcDM+Ff03JMDoPYJpr
ADc6CExFMdEBh/YTO5NCmcBmwi8dl/lNfUoDzKGKRf7UR/7DCIX/N+d6UeiGQ5mrYOsz2Mrqc9Ua
bb9K4LLVOgdvFVc3hev/IxzvK5YhW5EwNVEnEsCxYGfFzjlD7DuX7CYiXL+acRyZ20rY68VPAqH3
pIYT4JWcLfJuAHqDF6+Nvt/G+P7GWaMux6RjJdgYQ1VCkVnk/CZHejY0giw0SaUmBR63bsyhHxre
D/JXyk1FduUucw3tBJl+IzV44eRt1gkK3jWSbmx24zqM5CP21r4NK73Mx+/b3ITa/LVeBtHS8bau
pGqhE9iGqgveIdOTpe1GGstJzlWcrmspSHwSPorbN+XM0AYrH1KGbjzluSCUddy/lNLn2h09+hbx
g5zI/d7m89jk5FgM2bMMCdYQGKZXz6EunMcWAlPkjUw+ZQXA1m1v7KnSB4o0F6jq+2lb0/JE5Vwa
tXld3LuFannkYqfnUL7s/RgLyEZ9iHFbR4IgOJQoNU/aa9bSAcRAcL6j1R9JQgyklbPnXbJ/fj2d
6A/Pu86GUf+dX6oWX7bD4CxvKPJLvFLrOhcZnaOciu3DT7BIxJd6DdWw8EDI4d6Oi4bZAXTzNKtk
Jbn7zoJKVSXsL0WOGQS5Fh7SEWH8BdEKuDqUCijn7e/l6SpN0apUKeKMyeonBef0Bq+Iq69z/SXT
EgQQDO2Jz9Tm0Tbm9hH8pSvRqno0Tzb+nZyhZ+PPutKHvMale+dxEhYVrQAdJ0/r1aXkOLGxcmEe
5cQmqxWa87AMHyAHSd1UnwSYY2ThJ5KzOPAl3gbOCsuaogamv8lln7TQNAXs4f2q+vdfNXt+fzvq
MqoFRQNAHUgJ/0OCCwmQiMVHSH9BW54mXazxQnw+H6hihamvWbWpAGigXo0XED/d1SeUvuI2TTl/
7hYghio7QbVhKbTxK0+20jwSgVaiWeVkuzvAyUi14YHQMWpmPZMNLL7u963es/N0U1E0VfgjTBRQ
1WPwRCDltKlGuqQxVUxyfBLMvK0tfpzGryPm8k2xtxX4qcPfwjeOv6MHyiaROQnbdIkVBWlc+l/o
pBT5TZpppNWcY0AVqY5U+NY6GGGVoz/dPQKeL++qvvq3GTzwXYYnVBMLhGLOCS/42w7JM+/ixWdP
JEi+ddX+0lIddNSkkdSpGGUKDsgT1F7w2e6uVb4EyoxxO0ZIPrRs9kLkxk+0TUh3Vx2rpUqEbD2j
OtTK8B/JxgzaU0Iz85pcU9X055OfxlDxOGSkblBmVUz97UIpzt7bQYAVoHb2JARkAef7BCuHYMyu
bJScz06UjBilwPOEoU6pVv/dZIj/8taAulx3wZmR8FkzVdUUEHVBxq87PjTBp2P0aEaSxTzQyBIw
+QzvW/JRsWvpu0rAaBroYK3SWA1lS/wS9LzzGkx2LvIcnA4g6RYijKM0XJhIQJTAfk6Hyi2hkAYO
eFN366IFa1fMiWqWOaPQpXKxVK/AegRQNK5s
`pragma protect end_protected
