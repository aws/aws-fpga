`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
a32L6jRsmqZIg7YCjPWIo7zUFyri4sFQEsG94CbRiOqqMyqh+/TJGDUDdthWasTDsAxvXmvn04dc
RxWPKS9zZTPTatHeUJHl0EeuBAzKeYizXZToTc851F5pVzzroUFfctbIozbjX8lxBPNcgWgGIZ5T
BPzcvB/dkPKZSqZkjyz5aufD9xHtVMl08Tdrg9VzXupgRN/LZNatNJ3SyKy2xzH2RXwmewqdknUo
vuFjluUJSAjpX4eymD/+si3wTUmz8JszlO4zwbd8ztq/v5k4hExI2dPTbJwFrsVopl39XyQbRR9U
2vLB2S32bWXphXOpkcJbq7Il/dAn4kcbh3RDPA==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
MhGjz3vt4cB442qCni5LwqPSozIpJOrO98jEyF4PVQvyPyYX+H/MaR5yTvsOxbZJGaXqoaut5bGY
H6AyLoVq/aS1LESiZQ1Dyn7BysN+DrHXUZXdR5J0bkmjsrw2AM5CcXGwrLOA0k0lSW+MnW18PCtk
0pJNsQd007LJcqgFq4U=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
aUyq1jIjxAMyb1ipSW3t7iXgXYZiO9B0zgb+cq/YaLu84wKxG1S/I/dAgB3a0oNi2eZih02R4qpH
h2CkeD/iowwhxAmHuSgg1nGim9I46DQ+HakcN/+oEaEtP4T4UHz+c+Cx/Bkr++G6GXSZRvsHr5E7
/kfcMLarZQNfuUpq9Fc=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4080)
`pragma protect data_block
L/2LpVwSBPRNgYkylC9nAWKEQyboEAWMD/HEAS3Ikr5vqeBLw4lLibjz7czVJKjI0cyqvbc3dfAy
sCj53c92NpJv/JV8WuISWG/Zu9RkYsEXOJipQYcfsyCgWddNSenoGzX8SszjBbm7M/YF7JZhvJbX
kQHuTP8Kc9KrUuORBddQUuGvBFM2ejxQSHm8ZeZvHVFwJwtxMwObciCXKifOQNp3wDS1H2XT5inE
c8TmM6vBtIk4syAPJLajD1fAhGI6s+xKIO/10fip430vdXvZZKoV/1IxGZQFiepPNDFxn4tIQE6K
L2keFC5WmbnPzV+xndIjJNhTrvy0sERr6Nctd+ShH7V1IKWrY7h8Ruex57+rYt9fcOcgV9xlmMAk
HXF01k9zfkj2w37x5UsLAmeOEdGQ3BvnIYj93510CH9lCQWGBYXRuaUh2POheOebTyxEkXw8CTOF
q0EHbD3ptufR/rH6x/iEOFuaxwMksE44fi87w9TdiUDGjZD9T++LxajGEk5w1rVLNVroqVoIo7sX
wOEdu7iiK2g+8P2RzNGRDuXIIyZATD1TKnI6fdPvA/8aqvddhsm4FJoDFsL/kb7im+baC6E4LovJ
fg2By4cbC4HLEO80zmy7zTXvM7bcpRwlf1UiMr9UdS0LsuFpgR67rErwBxJyqix+WGAVY05VCUFZ
R2+tw38ZNr6bPQ5byU6ZvIE19/yDWjgLtVMa6UFfu98o/NRhwKH5xD2sL7I467xeF8ujs/wsidII
pV27R4TmUpCXG/0b689UwIcuEvzQ26MPFhr2ftcKpaYB8qyFDTu2gVUv4VOjwgi2Vvo4+Q9wq36u
9DkWpRaC75+IkA49W0/7OQnUNEsgc2PbhTCrlZ/T+uuyI/QO9CTPWrTCJpvN4GReEH6KcftoQpwg
6DcgrAF8V8+kKiXzvlDH4yN3n9uXkempJdT53Zi9q6dI5q43wpBZ6Wixcf/I7UedK+RsHE3HiPRc
arULY3NG27hWHPdOoHk1fvkuagnD2pxw5QiFQmA4SlAPZ9guzrQfgAP8cZEIYJ+4/x7SpdNyV9fM
mIuufAK6BjylvRtBLmDizJM2CULjmAEHfXA7q1IQXXu/B+KC7RPYVNotnUdXmDiVhqxREyP8KM6L
yCeBx1SBMOzyePyPaTdwENuIQdUXGFYSIpL3mDy1J1gLkVlCc89KzzMfxnCA0OPDfyELAk2U7QQw
ONvASzGSAArGStH0tmYGTZll4C8R4yYDmNAtwTytO0WkhuNefhKuDw+N/2y6Rt7wbIdDAcYBY8e4
w89u8koMboVKCrAVlLWd7yWJlaNI1sBh8BvPUdnur1GHT0mrkGft9ScTBcZDwfN2wUCktS6+zf55
A9S7rRawnQRQsjJp075+SA6ykdRAiZva87r5uoQhVOW0hANXxFQb4XMoeF3kQml1js4gCTz313j2
erZ/a1bT7ZwZqHBiQHiyw1AtunXR6zD2fTy0wgatElyHx0DzpQZw5MuUwWEgJel1i3jDTG9yTnOy
FRZRhmV43mz4KHQb/c+zG5YGrH4lM1zo5R6gOYLIQU2lycmBrDwoiv7i/AnfCkzCmv5lpM40zDkO
ijEMFWPPLz+tYkCRXZeXM4fCtgRqwr+PmTSv9HJaw+OqoS00eFPzz3pA36GvczhsvGkWO4mWEuIX
OX4FyFCpfQzI08cuLGA3vCnoLyWnS0O95JIcia4eHzWZ3OTP3NyrUtA/iMcFSrG9Xm3BwFeItM+D
Al/HNF23OSqi+DLrVojirzYiYvRBGoCOqRDvGXOR6mofOcgGYdyIXGcz8GJFmgRUEsNi/O9IUgRn
a9RCD/c72DZ2DYmXCjyp4ReVWBk2Ou/o7QQ/w+93g49v8pUm6VGIYox2e3zGUJaokcz84LPmETGa
qEBlcy9chbvXxuihGdyEXf5BKuliZCUqVKK18RHmjypsv/CHc3AgW1SOqqlBcq+hRD9MLZZYgTqK
X+GfmWbnFWIEawYjx37a6+ki6aS1GQpibEkeP7fw750nAh2DNVBbzfQszJZJjL9HDXRt2ezv9YsN
PWnxUquQDcDa0Zm4SJ6RL/+aAYAdmV25U0lKVtNThHxHaLDuVItIfaP93kqe8DB2+1GRw+aUcrLc
vuI5DPDFDO5LIFeSQGgcbZ2Y2cf1wQt14WQxl/LcQMUWtQIAcbrdb6USwNl2/zd9N7Qr2dbuazCy
Cv8cEaUHI3DTvNvhl/qGxBXxc4GCZSG7XzoHdHjBn0RNCI3SVBTIMO4ptUL3rKDOI7FT7sjn/LEA
pFA1MSrCgWRLftAsBRqTpXipCGUwflD2pLCCL3mFgys3TUDxKYZq5rOaiXweiz+KjjkHI1kkoP8B
ddRiINNS3xSS6YARwFdqHObmHLvsEKy4dcGv1ZCoBDrBjfW+fEMyzC3EpChhPbZSsh90YSR6z+D0
7Lva1zERNt3NN/LOpWq5g4lG4nnGeJdjQPeU8auDuAEZHkzhdQCjhKr3SW6X25SkwIKjlHwC94XM
OvXZM2YNN1byai+GzAmxAncFC3e/G2Cf649mqUhjURhV/1RVjj4i2XoY60uweGIIR9PDgMRawFZL
NTokvEV9vofTbjzAwVfHY/+3f6L+mTX85pUuobirjV6t1UJAk3bP9OAWJXzquxPsJiXt1Zlc/NVL
3xqvBxhNhcM7YRMSV3eZyD/JuiBCYnp18m3o0IqizQKDhhTaG/WN+idyRbLmsPwKio7NPUgUHSkU
udS0b4zWU+B1D4k0zqv6b4y8zSiESWPdFEnesbZpdcjw2iP1nj2stzADDCHc9O7pJ+FcHBQxfXUH
AzzFWwpGHAWoycMSbByyqDgsFY+zaiB41cB7ie3tc5hOGzb9aW+8jjsNfKUGnBzuJV3IsGOxwRXJ
S7fl8fWQkXLMgQGJS/lSW+TfqogLFpbXpi3AgZ1wTN96hNRH6X+wcvzQlBwxnrCURZJkNah4d4/e
01UDL6CBonewxZq/Wd30g/0txoOX2R0vb4kX0X2qTc0NWk9LKiII6yB1JRLU7vyKezQ7OiQFpmFw
iNK4ALFuTyKEpP7+MA+3U9TgBlu/EuOf9yEla5fJXdvldHKlTNJH1NZcko3fvm2eSumtCGZDuz1D
2n32fdj16V6M/12+9hQQsLgTmxXz7bJaqjGUNIcEJmDzRAZ1leMhCwiSFPrFwyVuq9kp8TIk9H/z
PxWQeDSyC22QE4q39gU3X0OzhiOZg2w4miQNaqLFF0nRnUpGPpBzje+xfE9CxSxA6XM6fHCQPa3D
YZQ6dEpSThdxo9UAzCltrqNjyMxEdQfxQSlw2Wck9ozlDf4f0Z/0ED0PEtmnlrK04ffeSiAL/qqZ
hnYoD1sG6xGmxNDVFrNWC649i72Qa41AqH9mcJXggmxWDQ98s9vmKm12iZs478JfldZGb5sWmH3e
KqTz8p64jMrdTwzKGl00VgJ/nZBVpRX98mDv7zXworFleyObpUVQ1xAul//QgKyObwEoaPW6zKyp
o7QUff7xoXpGgkHVLFjFdTwDOW/CWwL8aqc/YE0MpS/GizcFOxEGEy11b+0WAmHv8un96wrv4xUo
2ONRblfKeOLDyswtlpDFPl4kV5BvSWfKQYTrokDFXrINnJR1WZxEr78fs/M7qKfBWw/xnC6rqVn3
TfRK0v7wm+Go+2WrtmT8n/2mDT2tb7kD3oY/IiNHjIZaClGWqFkMrN5zj+1MO7QTRZgQ9WlA8v/2
DHqGfWVazwoWuIJQPPldYFsUMxzJ5g0pJtUqMXeVSZkk1gXj5DsmBDq8JUWDw3y9j63i3/eTplGG
uh27HzT3T2aV6mLnTORuVdNv9XFunTvImoNh/os3JS9vl2YfNNvjyT2h6CCXL0+noNBau+MkSGbs
Jm1M5sQjTUZuCkoUOJ5okEz/felfirXp588d3/yd3qYX6oaGyxcq7JJuaMZBVnjOC58VoikeklG+
5nBcbNTnPXsSkk4/QKHP3IAXUrOEkNinyqfaYv1xzCjkulH+KWRvy+T78xrJZ9+zUis4ah+xAua1
ZEbCmopS2ZuYahwED0Kp9t1E3weHniM0lPlLv98+/XA/aUYWMhspDFpUThlbyrd0/FIWThk3PhgB
6sIcrpW8DJwPlwhpLapvWQAIY58UhHDD1rXRD6qcYLS68i6obHXzF4D4i2qtXTye61x/TR4lavrM
tofOVIfeEt22psDnoLAgpR2X0Y+OKk/2+Dbe2RHz/BBt5sfYrClJ25cC+k83vBuo3FwDJbAdE00Q
IbBxs77ossWTAZFXP4MZsmkLvvo2LMstE42lD1D8dP99/zNS79qdr9BMmBLFrwhCn3rQFuugy/6G
OwrpTrxh58J5kEwYuUDiC5qY3JhNk16zj1gt0SYbj5Vo3Zf5Mp+onyeADUNWtWqt1R+NDc9bDR9M
bx/XizqK5lo6FxA8JgXbwpA8Id1Dzjq7Q4373v7LQcnYI0HIQqaq4o9hRhZAW5uz4w6r4DEgeJ+a
UuysaX/dFwN58pOF1RMslWqG/F0w9TRJjt9vOGqYgUypFs8NTV9WibvMRAKtCFPuklMaPJx3tbOw
q/+jlIN2idEuTV/z4mP2/YwCa+zZjXth/uAO1oEsD+bwc50rYsscSbKmxVqC5bQ/YsbZwhbCXRrm
4IWIy1/C4HGnGFKBbtOa2oFqDL17yRGb+OYZzSGE0oFCX3kwZaVv+1PUTao9ilL2yz4+HOMsYnqS
5d6zgIusKHhnS74Ao5DrLHpNrNUlnEAs7O7EBq/U7JR6agLZAz8xdg17SC6mQqKkoaTxJJZL6b/2
pYeEdMtGHubh8paDJZ8j0l1GOHHKkswUY4bA8XU7I1P6l3WPvHAUhSQATXhbhwYDLGc1RdYIYi9o
pvRKlQqPJHRwV7gqK4KLJMwZ2M2FkqPbHa9jiVvMbL5P2atNfZUrBxzkP8UIZi+YmFuF3KDpZulp
kIb/ORvJB7MrOhI0/saOidstli1pbjFCMUyWDuSDjqi4goxak0ysxcyP9KpF5WCFb5/Ge16ebi2J
Knu1Hgs2YbMRUkw08zLR708nnV/5dROOTzSbl7MSaHPqn/LevCrGqOhXnUmFHIZXefXWJuXcbfKM
jtVnA/OISm/gTnFdL+GuI/9Qfi7wNpdvCag5JFuo6Thv270XL4SHWziLoMfj2kTh3e7k7rMVU+5/
jIge1SEMO2qJeM8rcmQCW+4xn/5NdWCWDb6L+440OOQJERhBAOLzv3h1jjApthg8qux0iw5rXPH2
dKCDnRSePvrjOKj7KNCZOI562MgTxyYyP87zCInTISOor3SOv4IR/ntXJSWh+kYllB/xtM+8SlVs
jrUU5DvS8FmDmDNgZLC/RvrY/3Kk+Bob7fg3jSoVlVPAN27wHO3MtjGFZgRP/YYDhU5xyEXV0dPR
oXs3qSt5Dz2hXXe6q9XErbKd/Qvl8E67cMeijahYy5V1
`pragma protect end_protected
