`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
aH4WLdGmo0c74wSq+ByEcKN0AHrF1/OD5g7utJql4yMFR1kC7F+GAV7QKe57yLrNv5yR2J4KK+Aa
aSh89IKjbaTXtrVeQj8zvNXniN1eEBvYLxKqOTQ2R4xYzI6Q0RLvgd4oxkYL6E2nTXv4eWMUs4WO
QFxorgJBkTRvO6lHmX+eP0DZ+SczhrsliPqMklVrJljM0/RgRn7yUGbZhKfl0VQgN9Lo8dumHsAt
4gQEtQeYxP871emYPpa8mwhzje//OrXDQ4OOQRbREctPIqwroQvgUj8Fa2vgu6XwKB6a3Q41/GrA
1eYg+Km8N9W3bL5RssWJliM6Dm/QnEdwcyK/JQ==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
uyplYCQWt2fvObx/t0roUegqs4K+qrzGty28X0RTvfxXaAK5adpd+euYmaSYlSaJ7NLmDZEH+q36
UKGusbgVAAX4/5ZGYIHg2KUz+C31tShvhO6cRXVpcfyvG0jBPqhn0hVuqcgb8xkVMfUPIAeTEa9U
KQmjNpE639QIl0qgv/g=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
MFp+ZoS7urdvBQyCwW202Q52D5Gr5rR/fTyYMzcA9v48hiqGG7QPJ7kqkWXVjUNgEr1blUcZ0HfV
7dbRPabZnIgsVL0jd5TgcSlE3OXbHhqlqKO60DRVLu+14pDB/dYHl42hBUgOQEijsUtF2cqrsKJ8
As2Eco0IKMNKr5gbVS0=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5008)
`pragma protect data_block
Ufk5ixIeRWUuSt+MOyyAvbkXByyRxuFIqVBPdaY2duvzuChbYYaSDnKFn0OnxsKobZ1aYYnjgc9m
hi7uNWEVJrauSDzFJzU3z0spRNtO7PniXdKA5JLdPs3unKI1QbZGfZeDNIq4xjJd+53J3/Ve1C5o
hxBlUQgQBR3ox+0nMBWMIB4/NVQMAonp1IEBOCkaabKZx2RgjDAsE8htshqt5ur/mht/v4I0te7/
Fe5pbE6SZ2H3TfUL3h+EYEn2lfI3fbUOK3YULuE1lkV3YuEUxZef3EcJWkbYY3yx4lQxexUA95tw
seAM3SHSISR7TlIn6eK5RyaqbgN8YVzDm8YVtbJxYQBR50cE6vQ7OB6XWwECv0xjGhsQz15x1b3X
CR8Tz73mHgA+Vgbr15An431iKP/Piz4uhGnShbDOz3rX2Q3Ky6oXdC8no1n1DCjsaFDlRl2XUg3h
xMLupu4n6JfRqMVzblsFmi/qCtqAE6CLG6x4zAYZAMV2/5kgDxGIBzIR45kbP8jN+6IuxS2Ey3qY
FFu5Kua3vqH9XW9Erbsr1TURgwbc4cXfQtheKTbbkUMoF/JQtrIU54s+2SCtz9SvCjzi4+AWc6bj
LtMY6Vr/nDtj0kmJ9lBXtrcg2GymVm/FCBCcSPkzlJ4PQGpWgVzR5hwXtWjagkV5Ey8dbS95b0Zm
xac5wbwZyiZPNcxeBiql22lIQCDJhfOjTUhmBq1NyCv7sXsO48OeSVfvhNjQ+PSP+3sYmlTN9CKr
LzDkcanweN5C+jMT+gk0xg/repBB/SVj+IlIWsj9N7uCXsJjM0RjSmTQKocc40jrNTFQ8P/kpqZO
JSrzoxHegGqlSzpSmWqzmlVjIEHsQd2jOojx/E2Ryf0OSvhvMDaRL8sVtp60ByAM+ytIHwuBzKB5
q5mvNm1dSCxqZsLZiqTAVJUVMvNBDmMnveG1bP1MikEiKAcmgiDuju3MnAeKe01c2PuXSbu+k7jB
5MMRO8Xkf0/FqKNOGh8VmGhQ0+KhcVt6E84QyQbWm29PkAhvl2AIwiEuiAX3ZrobWrsVC+tTXctH
RoekNdJtFRR+cFnFEtYdxabgKtierAM6AL+sJkTdGbWexAG04geDXd+kxBZwprLfATk3yeu3Z4wa
vTU5xNx8ImdfW/FSbgLmdGFLCcqqwwOZj5fSdq+7e27IOzOZO0CVMZKl+uuaGFuBpDNyamBKrjVx
pKQAFJm08EH0eqDDnGNsvQL9+EnJzOJPtnCaelYQXK/XlU8tgLMBF/0I0lycKgnDyZdPyZaRC0ms
68aYJq1liuV4AGGbr6ZtMyOszoh0zBcd3DsmXcxxiHLx+71+whRdKgC1It/KnrW9CJZU3cW+8Lo6
z1hZW+OU8UfB1BZnBVbYArf1F+rvsipK9zPYiKmyk5QLJRegQ6zO0kEqCppTWCPdzH+lyaZ4fxGN
fQzt4E91D3W0qB1GumH8Ed1bakJBZECYvstq3+tM7czf6/LVZuXKPUJMRw327BZjx5c58A2QD5xS
jFTMni5tKxH7fq3dDgqkO4yq/WjrZ5bjBTixCY1uWqJZhoO3PIHdxOYLsRu/s/rL+BsbLJzGK098
Mer+wGqq0tb7+AFFMIIF0cbilqbflft2k9BiYx5l0VoNT+cHSXw5Ho+0Dm6cz1BVC90HZT1BrjJf
iJYGMpU/dyoRuUgt7z5+Lc4Cg56vXmjX8N5VU58NEfrvR0FgCOKqGbmqVuDJ2uEeZrB/x/Gz5IGZ
DzIolxIKWxXPjfvtsXDyL6kA1tEIEYGRejvLaMXYAUyPpcDowzKAREbO+/XQOvkQd1nudLiza8Us
6dfAWxntecRnopp6sg5cFlW3D4DDaONW9qEPFGKyi6ikYyaEfAVwIdwt1tfbLT2EM/Ebq8sft9kO
fC0ducosKwnL5mAEAlP37r3n8joc3iItK0/yU+BuDJhsyXdT67AvF61JqihW2dY3A2dTn+B2pGQ7
+3oe4MsWj1/9O1y4bJoRmpEZVAm/xfk4WRLTiRRdLMu8YQu9mN0/v2CQy8uOiXkn5fRccTn01aD+
F8e8qjQpsldsn7R6knuDGHBQrJBqUp6XxuzfPKVbQ88L6NsFIfneRZCEZ/zv+74bzERSOdm1135o
3VMFDyZgXUJ8dWdW7JgyaPK6AY3HXEzyFyobs2gFvXJ+kVFfTDuFHdkIhQbNrTHESJnNeXpPvW7f
2UBwRxHa5t+BXwCGPcq+I7uFjZDQuthBjrnSWQKvIRy3UUvn6kN0a2gqr2QW+rQqOuDk3OwgaQmU
3ZPCg1hCKF+hjGWEAXYf2/eQ6Df/MW5ukWbdORtv83Bg2+kXC5r9j5DnCOBp1sJ8IXitTMsUj7I5
wSOlmsSrgSuRYibuikLMOQlZEhA77kMa6//GTfz3W/ILygmfDbUh5QWcrjUNG6IQmFjmyc3Qq13x
/tz7ThAh2ZPCuIe3FUI0Zhn/GqfRINUR31ZUg4gC/S5ZofTKXBiiYrab5SrMUJhYk7bWTHBPI2LI
gqpPtdzzruZCy5CB3tF6dbii2TfobGCRfW2H4hSgEW/4Gp6kyCuRQdFsSVe85kP9nzU6bmFTmAbO
8THgvRqwNgMIaUG2AplBY+ur0XuQFYhy1X2sUH/qqS1QmCs+h5C1b8QvioRgFQTUAzdf8CvW0x4X
KCMwC8gV4F3F9eHar/QfcHjYKMWsh1aTiZqkzQTZK/AGSiqSi6JsS53InpS/R+TQKbnIEZMu1ZOC
HArXVfbp3AgEFzlrhaRuGFmW4EWipTbDQbcDLAc+LWI4jsf/Sp+YlqsJ2wCW0sc6URi4qzdp8w5u
1WtJGr2tkFX2jWlYGYKJFkoQr5+hPGZZIKL1UJ5iMJirhJoDygNRRFaBbZfaPXD9+GK97A/XlwBj
lfPy6O+fKqDaHCo8jfIvmaSWlG0B39ZUaZx4lpEaXehoJM5Gcokm1MpRwyvlDpVPNwBR5AXiefbb
PcfJZhbrobM2x0qgO1XPjXHtT7j2V+GIhWFato1W1ktVj8WUPsFRI7zAwTPxudhWecOpbZ+Hz4eO
aahKuDsJwNFVtPbaLkCsxxCG5mn6RVB29QlotWdWZoN9ZIztMnGeBcICt7og0NiwHlLG2VBFADTZ
yU07M/GMT5wuwYtDEHx4lU1vaFlg7OUZeaXCYueisY7HG0bdKzYjnHqdLQop4RoDWRMKP3AViLjr
VxGgIKehav79+hFi659zD92E15L1Ip8hNW0RX1N/2/a8HcVWN/+AzZ6yCMNbKNrhBXkqmOYukNTz
gyb3EtU+YhgEnrcchWmQtFq+mVNrxRc0CNzir7wnwMAZGIsQdaBvpi77R4uwuoQuev9KWHZPHq57
8uKy4SsAOXWAmJlMx0sA04BHLn90YcRxO+4wP4v0ONuJp1h83GrnmbRPg4erArTphAfl9OFZT9si
U74f9GUrfhimrucxhPNWqypwFBHYxUgTAy0fJ63W9lhBO3YTmSE0dBvbfUqEL9z0bQrriBVhkRVG
SqGmH/0/TlBbWwmTB8TTj78apNV99totX87Do+sK8exvdTX5jupYwNGrhnCjtm3yHziiPsRNNsJL
ZjHS2daSXEt9s7Rl7xAvo6kQadoA7aujgdUtiHZe5QRL4SjZe5dz9/ePwagF2Dvk4eOT4vcj2MtZ
wxy1Qca+XPgPSZQhUdjZJh4bsDqhV3/hzooGcW9GJdZhnFEla6CL7PKPb7eBW0qNZjeorQ5Wk6fa
E0ca+ytXM2Rn/uJO0JKwHt8ccnPM/5t6WcQdLm8WUSNeBJbqOynHjorSjVMA0upQm7xeXOLu7QzG
7mZUJvWFjHizkkzSWrDFhIL/zi+7tcgpn1jbfrzaKtNheNNqCrDzUZtJ9rUdts8gso6Q+k7AWkI4
pToAkDM3DHKBU3zEDz3CvnrLu/X/NsbLXT+HT39DpiwBrcqqOs+kjIpnQxhX2DSKpQQavHfe4hUz
1t8Plfms/vwljghv1abEvUZtpgIXQfWNDr+WQ8oW1MyyHRp2Utc8AbLARwuEVm4cPlOAoJH+Pb+T
uMMbu35IXAALJ+iOfAGXck97TggRE8umAWsDJhQwfEAJ9du7UuevfAyDZ/YY7ZDZLn0BPfkv7a4/
8tl51xV3flEv4b29/JKsB9UJr0hpcQZIsMAtTVk2F/0ij8cvIyVyW/YE2ulGbLHtAv1f9n4gqC/o
dhsE9ir/B6elNVFDALGG5Uj8a4bASeQH4+mOk4PpDhtZZg4H/guTvIa4NkdxXxMLdDinPNY+PEnh
DOl+95/YaEHkG0qS/rYjuiRe9O9q5LaoHQ/tEdK8EIYwfzFEY0yD+yOwFaybS84ksgHArY38SHl3
i2deOgOoGD6ZSpuJs1Px0yM5SImvBFKtv4suRrmpOG6yhidUXNBZHi+KSDBFdIVaaYA99sKBbrvb
Nmv/v2sIu2QSSMGU6uEv8li/5GKvCxD8OWNGf0UaYVuOI2bauDBq+9glGwG6TGt3xiHFgxhKH3w2
sv+IFm6e+NpMpwrE6nKXpBwyZeWEcQlDYloUzxdtbsotXyLzsgAhLgJ3S0Xr4wb/dafBgXL6T1jx
NfzG3bpxXZfe0yrj+VdGqcEUG6FJzagtAnn9q9UdREiTSPFWXXTPye4RFr5pJu2Cz9wY5uVXtNLk
05Rui+YJuFvfdpREDWjhUlFsr2I6taC6ecu5fIy3HTIdejUIat3TniSOMIdsPFEhEvHaW/F3S9n0
UiNEYwNgTvSUPXNMjRsQu9jB0UVWqXLk1dHlTUil4VoFc0SLdTPCqiStD0y2cXqkEYMsQmqUvgPl
RhVXvrFRQ0H9eMiqJjjbun+f6YTI7sRiZHUiMPo+8/bkeXFKOP06VMQT6+722NCog9oa76EhCao1
H4wjeWDhusydW99aTHCGilemKiwnB+245ZJg93Jthx4jl0T29dfPPDMUCVXBknjiJlAThu50CJTL
OC1xQEMgQQ4H5+t9CrsNdQ6LoH+EMP9AnEGqoJF6uCQ5QkDL8+8aMOlKEAATWuSI+/a4kDitg13I
dFygFGTX6mzaf21gFe1DoWdFE0s4pReR1W93MB2D9biNAqx35iusH0nsrXdo8EtPGO1DYXE4cF8V
hH0d2KV4178ZePoMaOM301eTPP4ZGzFXVA57YnSol9BROWBt7RCcDxcAZVQIRMqX88nIQ5iTBIk8
3UmlFDBmTj+7HDgDbPiB/ftHjlTsjyhVettaSJIS3LZ7bGh85A2ZiwukvdbIAXC0pfuESuDef25N
zZEMzfNhNtkFEfsoqAq3Y2ze9VST70Uhxf+YYua5Ith/iRRbcnkzInsPlULdCMHYaUvVmDxQPEQy
wHtSkw4IM3yN9HZBdsBXYCiQbx458iwLpEBy2viCELiGnyLk9zyx9RiQ9EBy4n4tOVx/4gJ2O8Et
nrU/3gesksKSikNbXoe+kADZFcODa3KkjvnPaIPqg+ZMUeJdHk7L/cm1ae9ycKiie4hFOvKhEMlp
sv409WpbHmF0MY/B2Eu7z1dzF/V2780WzixIYu5CFplMxOdh/H5TmD1qoiKdk94rq8dxu1cYsYpi
/pinx55iTSmzlepZZ/sQ47ArPNc8VJ4M9Ieyd7fsO3v6AnfT3Th6MoZel0NkxUm0hN7TRZ/B3pWd
qGg/CA+y/xSonBAHQlm9r94X410eELeja01vPU5ilsrfsi9L+kc/cvo+9IwRnSBK6cUaEmUTvMw+
6Ph1eMIiQ0+O41h8js8KPG3PTbUhrxmt/D/Y8bT+VPkQmx9UszSXT7ptzwIpmwt2+YRM0urrhrA5
2UhvvA5FSms7Zg3I+J4D5PLdGzsMsXkf/K1qTUQL4yoEgPKpsFMJ/8wibhyD/RdocV7Zx0wcMJyQ
qEe1/kfs6unWMkvLyZ7HmMmHEi4ghrl5Zom9OanJw26zAIJn+10s0DSKzImELBi2g/hnIP+mgGeY
hIyjnDrWX55pAoYCQ/9IJoVItAD+YQXqOeJhK/ITzVKJ7/+GV13dEewnXlNJB0/44TkHV4VecVby
x6ZA7BIP2T8BnlIL4/PUQ2PxaZ1e5+oC9no3RYUD7hvFFJ1XOTB0cuAMJ61am4BZ35xDQ9NDm20f
7iS0gRJES1DQDSX4RFZ4cCn9pLWeiMFHvTbCUfKQzFq/IwMBpdxEDBxpxTrF2HZCEUqj6vcWh2CR
4iy7opTHSpibFrn+NOAklyrKcDf8VkPROlN7s8g5fd2oOW/TKXlXPxes91BZKRScqatpanwHxkpC
7Ibe5eBYBCTTT5PvSSz0f1RlitfY+H+AxloykHUhY+2d58xtn2zIlCHDgToP/9WvAkn2ewM/74iO
+NF45lSD6RWjvG99vSsdJ5vrAHOvfg+BUu1BNtsMGUZ7686u7wc31OcK0zBk+YCgI8TSGeAj5v06
coK2gNJDBo1vCpyKMLtrrUjEvMwxvwbuPAn38wq50u3WPa1KQhHW63uvrKmPiTPmc/suZoWYf4kg
NWdW41VzDkIQ8UVGqmcDeWMyYz0McVDlINkx4IxBzLAVrRJoMHgbWGrxoDMyHV2rxHEqUZwbXHou
oto0WPDg63/Jk7xNbhianesTv+fR6cAv9WXUOeUriA45T06kngKr6NUvt8mYX6DKAwDzY9KNsyao
E8hJZhWbeZDXG6uRJbjxNeYZGoghrXtW6mY+6pHMEX1StnDc1+v+t5wCZ83kpBx+3Q==
`pragma protect end_protected
