`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
kccS7LGRiYCWXsvGn5BDuuWFedcj2xj8qy/7gMN5F9XPq/HtzapgmEj+j2wLTwKDz48saUtHYkf4
Ce+s/riBtbPQOrVngvOcMr0qU38KruMs2r8IlGUZd77NG9JXBgI3CBHdkHSEpNO5t/3DyvNSuJ5U
Ie07WqWaJH27484VQT1D6qNffCeZG60H94MYEsuerkvqkqxrtw0l3JLXUAoofS9pudbQyUVyLZKa
NHiZN3AE5m+GfrAGgP/ou4dU6ZAvGLRz/a757tMygDx02KuWJze/dwU++e8LOPnC8FrbaGeeNAxk
bOxrXj3hhnrT5fDZto6dN8IlLUOGV0dVv8PwVg==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
vPqin7igm7dJrbcg2MRWPxsRjxOFJJMe6i39G4b7KQN6rcOZSHdZBMbI22t3F/GL4TuD3a70N+Qi
i2A6iqSIrmirkqvIc9fcXvjWsPFPAtKlZd2u+02A+6pv9KIZf15OMNHUXk+sQ/9fELDsvy/QbtTJ
NRP8xdgF0TZlToM/+fk=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
oAJPtiPDZXamckLv+awlNUkPogH6su4sC8rh9Xgm1Z6cVfSvBrlLzl7wYNiUy6nY5Tpq9IkjYwch
lHryFXgseqA1KtBW4HSi9PypTPJqy5Anf+bGuIjFqanq/kDUpUBFBgY+AyWfVIBfMrxG+RiWZGqa
fVtRofUEiWC2mjzfY9M=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2688)
`pragma protect data_block
UCVHrpN0PpSSuCa5X5VzjKgCd/sB/dY0eUzzKYw59OMLrJab4ghOnlEbXok3z76v2hU/TaZw1lAu
x48RWy7lf68P1Xdk+ENMotryRxOBDY9fNJFYxOxE+lylVudC8qdiSWPmd8FEG3MkRt4G7S5Eq3kR
O036al8WKdHI+CKtNfbsSyO9tqCspQhonCDtPwb5ldXZdPRWr1rl3se+4XziAy6KHYzmmYvqXqyM
WuqkufseEIN7kMjSZKsjon9wl4lfWdMuksBWPkLR7nY4WxWQB+TBWyiussSGYzdt/Erf4+CZ7X2u
fdf8O+ybnExUVXNqVf75KLoXbyz56uZrjXARoJM+R1ft/bh8NYyMnxrQSL99eOWxwoxiUFomMghv
61V6NdaPE4UHpDrnfhblQtfbL4t4usAkGpyKPtzNNYp5VFnlMaYE8QtsqIik/ko8IHKIFKR013EK
kkaqmhhFpD8q/EiI6pkZs6KI6iv0Lih8yNj8+ubDYxLnzU4M2pSeP8UHf2d3xGTwfIxV9nR4N40N
Yxr+bnrosEsAfMW+keX58osFocXQXFAacJ1Dlk3MEFQT7RJ7kDQbOh16v+T5I7S46S74M/HbsPit
11mZrTIJCLMt57uCtHIBcTQooR9oU3FZbMMB9J5A6XBu+Wfgosc/AkmyD6C2SLOXffgXgYKCBNHi
WgbEWb+krIqaqQcC26fRdBFmkQIPSXXaBJQ+cMfuI7yFigQAtl/z3uSzFsyn9XNNEZR07VVLTdDP
cDyae7yGVwgVvyMh229UZfqkxytMAdnoGul9EQKWOhrJzObI3z/a+SThnJpvS9RJolrT2CHL/6Kl
v+tEwwpnUrM75DAsNMXXgX0/q+pdinxiiy9DjZ5+EHwkfN85Nrv1aOKRZTVJPsEHTIeW8I/tvF5g
OHBc+6z1/1y9Qmoxjo8wpPhgKFZxOfKn/mNcAMa5X+VwhliwQafpzAYvqaHKBzdVGb0RcPXN2Z+u
hHPfsoxTt7IVtO5MEoVu3sufy6Pv0inbidCdA0c4MfXoO52H8AV07I7vNrVmP4zXHDZdnmikBQcE
KHUV++hew3Ok3GLzWKEXCOCIpNScNHSO5usLKbDU5KJba/xGSaBZHBLQctk1fiwrEa+HRasuLrHC
YrLs8cA+0ZkdEG/0o++Yorb0g5ABthRJS5ajNvcLUAA2MLjliqu8Jg5cWqHHA0rVOp5rTrFI75In
0Jp1A6BWaCaFHk/NJfYKcEX8BsSrYaAAoWtBPXLnoov7NhmyWwvgf4ZB58lvuAq2osyaQrW8dnhS
2h8z9HIzldNXNgQ3M0yp/jqjwdGJXCwUwLk9+r+6pBE2s20/STA/cnYx4qEWLa00AyHHkkAW99rB
K1UvAnzH82FGWPid+8DHkQGws65Bwy9jdLvD9zgY+QBVsjwjTxs3q+T5QDEeet3WoaQNYb5MIUVL
eDWkxWGm+zEgVaOoIKohkhdpJ7ANqrJFmO2rIDrcXNXLg2wXjA2svZLQadsftL3FM8Xyko72vHpr
flKPDrezcqhcJGLzHWJ5+VY95oqgJqIJsABLOFimXV4iR3/SiLEq0qM1LJ2JvMVVknT1YFR3xFLx
6/CHzKynEOCkO1Pvf6tui0PmFkfRFC58eOtkSObea8Con9W8jVaDhxV0fXr0gc8dpx7aZF6GeOy2
fUaXueodIx5kOgem8dAaE90hYE6MQKSQkY29sQ+lpeNzhMDVcAO+f6DdZCPA7DLd6XlpWNhTBYgq
9zgyFfkvNCKxe92gGPpaeDOlyLBq3PfLsV3590+t93dG4o1eOuAfOKXSjXkV/LFsaDxxISXCiJ25
HJs2e4TyHwBZ48y9YVFNA49twxsUyiWCorNiKX1XCb8yz9Zca7Ieiww0JppGUfQ2+8C5FdWinBYL
V+tVw50OJvlfyI+TaqHtntKaIQsuvNfcrdYr9nq55PJ14MJmFwBtViqLoO+m2HMZ9A8h0sKdkGBf
rEu1ZQre4E2izyHr9JK77DVZ2AFewIVAN86z6Zwo9Xh1vj8zsYxs4fRVoYL8hlnoVSPox6uI/tus
iQL0rCOiG4A0n6iDc1zHkIdGTQrwhSR2irhOZzwKP8mhgN2WCpzaPMNsszhljB4cqWbwU6BUqN4I
uc7IfyrjuUw6CmFt/hAg48I+3s1qHvh5rA1jUOZxJmzZ0nsHE3xyuIJzs7hGw5p9YRcgmwB//0tv
I6s+kbw1XMcme3mhOXS3nvSbtXrrS6VN1i86lerHEEEFaQeY6LOni3YwTk8CxzlIjSoF5pkl+eRB
EQa/YOlPGuwYLMhTlEHwW9aQ8qt4YasgYDEweVwqJw8/yFs2zS6rlVuKLZpZlVPa1DxMJzrATUMA
eykBHuoNAVL3cBYSHuaDHMaHIsUgObDhtR/zxByt2febF/0gvea9FvGnPbk/mAIMmvA7SzD2hZ3Z
L9eBY7QEE27IlmB9bjjdPzBxYzT9wBfK9PLWTHr+k6Sgje3VQTkOqu3a0f9IH2ilddsUEWcNHFzd
im3KvUrE2ilJuLHX0LidZtXdUKRysL5Whb18vDjzagi/43dDPGob9/hIVoWQLbJ871q8UNMti5Pn
YdvhOIULCDJCp70bmexrOI3biVhyRMrgDeWYoRaf6cHcGZEoo1vFOV7an5tbwK0re89j5+3Lslcv
YR7RMyjuXdX52whWY9UBs3CNA+DNgVVTgRzP2KsY+wktKpq525ZA/NxEcPYpS5ro53ZjtFBWPpfZ
XnijIpLF2Iw5sv1lG3uNr60H0chVWtGw12zYxfryDvIXCRSAd2mLTad9NY4XL4BADRgB3IOP+w9S
GaUiDqv4G66wbk9n/7OxZgGOb+cnBVugUpQAB4v0uZMwUquFDPA3gWO0/WGaHIXh23k0/32AVOEI
24RwMIlyVhOmyS2j3Z4joaEF8uATupfjrd2wc7iTjbCAwXsHPQlSUT2IXu81JyfdeCAN+avbnM4k
qzm3G1vefNH+01j/FWxgngj/ZHI4heaBDL0kOwDaShufVB5TbHauXXi8ugHNugUdwBQ1muDEkBDx
nyH6YyRqo5NvL0PdZE9fdXImSyMtRFCTXnUiHs6x926VfBthzPqscL5E5TU+VbI1DyAn4mdIrf7E
uX2LxojJ8Jvj7Fw46tFFJkzg9i5FrdysfoeMaAwBJtMo9nTzv9lVoc+Btif4uA+4lUwiz96dBkQ5
+OV9yCrcCS1NBTbjgc+vPs2PX311TswyFCd/soyINDf1D5sHLnDXgCdRXyvQdmocPHZrlaui+6F2
vrHTmhcuilYJptIqlgPSRPyASStKI5EkPVZkvQUnFrCyUzKilCKNKY9Mt9RHmFU5DqmPv7zar6iM
HKvu1UAGSOc7UnrQlpF6WYBnthtRSzEilKXG8UTFSnkuXG6lgYQRsTjyBlqh/NmFC6r5D3rRG4p3
rgcW6xjBzj2C9gdG76c7LOYLmSJxMzmbsaP7CxxhYS3Id+/sp3UKg4s302CUjT1fBTd0NXcRBAKc
z0Dzw+AonjeOt7pm9j3DemQqYfHatv8FA13sljvpVsZM3rbDERodOhScp+b5EjxlhVXy8JJjlFH/
c2sAQ6IQVsKk
`pragma protect end_protected
