`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
k+KlIjK+YNsxX9OmD3j3+qHhlVBF0wyTgXADacV1dJBpyTMErUyvx5CSsosg4cEUo+50msNV2jq7
1T0pPia0WFk79sqhtJIV3QKQtY1L40/uZyORk1nXIm3DmmImfUnsRgu919huWw8pRTPHDgUWoLBO
75seUsmBOeB5PEDXHQKXGjJ8MWQgQRjLg32BtuV/nHEnjBBwybqLOJuCIhJby39V3ALUpNYLpLwp
sJH+2QDa4Nqh7v26kbn/mpPOaPLUEIO19M1GaItxHNexkM778SJgittAKxBUPiCN3A6r1U+RKXm4
T5ttPKMrXnlFQi2zgKZht85WJzg/K/mikh2YlQ==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
qfMEWqHG0iEpQbkFY6P5TNAktVx9MkWXp6OuJcIPeGekKOG9IdcgJCg+f5uXHSVfYQLpwCuCVhWq
iklWSqmx9EVzqtm+efcZEqiKkbymWL4VuvNpUIXvI4ef2C9tvuPtPK1zZXpqcO6ORtx4yht6EkS2
j5BqNCRIYwkbJ5C4Ji4=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
gxys3cZI6HcygPTCFeIf1k3SsSxclOPJ2VOeqyYh47nd4qnXXjf3SyBlel+JulWZE6IvtJdqJiy1
GMm3S/192Zwiw/r97r/9CVY6UJp6joaHwnq7pGv8RY0he76N5g9wTj+lnSc6Ke+EGpnGOvN1vtJq
XD9SGTu8K5Cpa7Xzv9A=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1600)
`pragma protect data_block
djK1OMDx32nOoUA5lX41Nl7xidTl8uFcZpfij8mGgKJGpp8sInnJlaZ2zP+BWpg/JOuyVucbASas
cqmNhosMZmY/jORsxUGKJwwggEYemqabawMdLyaj4vL7AZ9wI0QxlJ4jBr+y8lOi95Hc+Nrtbp2Z
oZQWB1wSGwQAdu34iyL+tMdGS2eWEColHXrThQEoNHNUcIz9M2qgDpI5CsFwx+TL18QAtk4zN5A9
yYgjEGFSFT8w6cXx3L42slZ8HKaoWn84di8fKPptyZXhlVcvXJXBLqQH2bRy15Ss7ldiOC53hx90
UYfGu7W3utcaJjWQmJXcF4L4i1sWYqGWlhRjyPxZMMhnmzTLzK0GK4Vp4ZM2so1d6t+JdIda4BvR
OKfY7i3TNNmi7rF5HKIJvjMY69MJh8s+MeVrL+hYCoXC7XXNgqZjdQ4fl9c5BXJ8nCp6mM13Wt26
gTua7tOr0XMfBuui6jvEbabsNa+hSqcrSiuCqkpOSeXSwktfsVEi3P3ftPFMBFfcCzfWOEaxC2vV
2D3lL8m59gteIvzb3zFQhkxDqAFbPtOT1LB7WD5F+epoqp0G7GddGzoaGBpL9FOIZtj28CXVUA/U
ERnBte7LOiLakUYb5qloIcDtL034s0Q1bc2JBpXOI7y3p49UveFDLBkhpxIL+uZ0X20V/nOGwCSB
vVNN8vBXQmQL+6oIW8wyDxMQSD9sSA/R4JfcNpPvgo2fZ8dZorenNnhkKu1d/espU9QOVuYZ57xY
G0OzZ1FIBn0BGQQXpg60E8xriKrqY4cfjvx3qNu96DvL3NsUdEL4Cqxrx7l7yoOBuNKNPXlfwqxb
+wcb47+6xzOBWMr1Zry7py4G5WWhZDI0IEMRwjm6Ay5UThLFGIY9XlrcBq4i7x7+G2eppaFBMAzR
Ctgxd5zEhKtlwfscHXvm4a/KBHvVQj14AMv0KxdxyfC/WrRjPE6i0s9SBNZb9ZpHxHI87BtvJDIQ
skyaea609Glg1iZLOnmQ7/76F37/b9TRkrbXCs/K/O5lSnqPh/7GGaOL4B1wxZAUxqT7D8YhA+UP
75sbi/s5ZK+Jhsm8NTRIju6BmG51Fr4PGLYvyQVx022ICSLvJsK+Qq7dnmZlVmND0rZ7JnPQanaE
TClWz3blHFWmsMyzvEduk1k43IfkZMCiSLsqb2OSt2sObyWiPFBs7y2DewluIPi4YEHXq4tpRTrv
cKyyBUsu0eZDw58e9X4M4zjDKUMG7qMBAp11tjO7nTqdGQD3JtJUjxkdFinJ1g2xZ2UMnJzenZKf
sIK5dWcC7AwxvXVWsSgoUWZryCzVPfR9wkONMgWOmCnrm/Az5jsU39GCN62RCCydZ2+feljY+CII
NYMVxiRN8BgmwI/v3maRUcKfZPmQZEIvMyuVi1aXKEgOwM8Qkqp7TxXWRVJoBl2ckdsho34qXdSt
GwfxD8RAx7BO298Fg8Q7nIxTV9oSgQKoLtXL4c/PXtkBBQmSz0uSlKlvpyV1iYIHxnJXjVzYWAMd
yygOEuxTcdHr6qRuzWp59FumWtvTMVlgt8n3+oFtuGN1mvLeOX+w20m2Tp04IyIch5cd69kMHGrm
bMp0qFK74TSc3O7T48ruFQAuFz7oo3eVg+HUMX3InxWYhyOHzeiRkDfvkkIHpW3MCL1Rz2upn/Y0
VDCWEgFOTNe/T75bmrtwOi3xhrLD9yGz4A2IBlfvnGhk3+AsA7Q2tfwywqrpgdoNuID+LyeCoa+z
I5EQb3wOTONXeY2ffpKtgZIF+PoaUVgnQW7CNYTR3dwA7SlRUaAyXqo7yeikNDHbZ+6qBYrQ1FPN
6VtwYNMuj8PQ9UCd4nG/VKMeEURuydSrMJfVsEQDiCv+oF09UjOWYl+iqYhkxLx3WBTVZgVyDojI
qaLmu4aWvCMkXdqud+jEhvo5bpTymhKsQ7Kw1OhhzwXcy1NZgANrr1kwVwh1KevlNIiVTKOFrO0X
xhXgHtuaGmg0QcIZwmbROx5OyxYdYA95Thfq15Tyw91XN6/VhlizsAjd2lNHd8wEkOLwzxUGefvA
Rzw/DNKTsFWQPNklwScdwFg9wIvBzBw100SexDW29s/NKOszUNEoHimt5nEKjatgPBa9s8tV0Vdy
4ikMEA==
`pragma protect end_protected
