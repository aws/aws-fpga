./../../../cl_dram_hbm_dma/verif/tests/test_dma_pcim_concurrent.sv