`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
hWF55EtsHThLlaQdLsn2L9P4Jr7mTFckYIh7J8kEYzHlT/w1F+xKW2mIjRFqUW1WOs6kOdC/tH3X
tVg6xMkGU4RWtnIyEB5Sr1KCuS/OhQmk4DsoKr73uSq44B5V1KK3Wd1s1QyUJ9DqA9rAE7b0iA8U
TGVsybm/LQqWY/Cim6mB+dCpkmzxrfDFIjVOkjGN9xo+8+UimyqipfkmFb/n9wiBApyMoEJhYYG0
YQkbNDEdVsQjUn16zMW0r7QZEhbfw0Vt9WJu4S6PjVxScbD00GWZy6sZE1o5NC6NpAR/OB1I61Ry
riIYURoa/sVPpkVQodXd6sKOA0qmdkISxAMY2A==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
FmgNAHPjpMPNcisSiXn66EMr+Rli1y7r6chkICAgN2DGyXZ5cLZwillS/m9ft+zPcGK8FKeJs30G
JYIkLAEq+Mehuv1MgMNkSL05yJNnuXMwsfozb/p2jDBo8bBvqJfoA/xOoa6C+/2t+nARD2pleg1Q
6eZIsf/vizrFNkTX10U=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
DAeiyYexuG/9L5bErS0J9ic20AToCzg5/9pvFpviuemJkn1MltTD6NGCAIcsaXZPKpdZZY6dALHq
cS2fHSur8BNpnfyFqafS1+uG99/cMqhrs+BabqJLb0CzxxNFg/1N2/cQxDaTCKQR3Na5Km9Lbvr7
KT9inafBADvYHYpsQww=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11968)
`pragma protect data_block
oLg+0YukDgJd4HzHfN0yp7lzwTDqkYQB9JL7lw6teSB+1GOG3/+LLvhvw9dZNNUuAxqNtYDjQCsL
3jFo1sSVUMs8PePFhLAjeprcrkuCkmir3UfyHHqW+Q3UdrR1YvcAtBW5va1TikLjJyAW3SbaSgIk
uB48fg+8tC7jkfdkN3aJYW8lnA8C6WHCIQUrpMWhCQ49QouM/QodYuka5zjoz0ZhG2F351XM3xhU
CFCNAetBqz+1uDpezObQShg8oLAZF5kHm88ii6wqQsLi8rnuBF4TYATzwCg6xI/IM980B7lwGTMh
0lEnrvg82ypu1tnQAVKdp9x6tXi44GXuWxsen3/drhTXaBc8p3bS5JR3icgT3HoNbnERyug0cYGD
5rT6CG+uH2Hg4lX1FjxKi5QOUEP0AbXWKNi9/+6TTeX2mb+xVxv9CtMTxtQi0AS1nzH4yYYaiJ+v
Sh1ai3AILyRjShOGco+VOsmAaNLzJHlKf0Yl2TyPIALl45bMBs3y3GdnTiHss2MNKPQuefHb8UzL
tgZ/xxINxg49n+N2pWNYegz1kxPdPynLgJ+ArjIiiZ+IKXRGuqsKTidH73S6Kwj+nWd3+Dv4aoY4
b5zKbhxT3RZ24TCqoBJmqv5R/CJREEHqugKeReMaUO41pWePpEUj6qDya4dBhZQfN/kC8SwzSqMn
zS0KWAiLgEAWSbjwAYMMvtlSZaAFepOKTzLwS2nv+7gSUKdFlg86Gpl7kBRFbsTytH4Gp0vXi/iC
B6KMeYzuAPij6piE5EyjqGoR2rPiy4ly/VVev3CX9Csde6qk6VtYEe8smihJRqV+b4kQy6+RApEl
3i5kBwAGiH05Lp7gkR8Rbds4nNiZXuLB2Wi/ld2ZYY7O7RDc9RwKrEeqAkkfIkndKFaKDgmNhIMC
Ia5cDA4lnz3ueLxVpRSf64BPNe5hrDVNL7u3w/4oagjDyA4vsKp3KIm1oV92PXQFVmlroFZLuNR4
EVSZKdWT/vUd6UEGY5hAAqTxtW/8kJxtSN39Tn3SF/KSXhS88RT079FhXIRBFOit3WyMzS3Ona2t
2ZKTdEm7vu/kbbOKdExxiEumcbXKMqt+nmQlLCe+RNE/67JZ2JGlpy99WyHSvRmXj+VKhzEWiNff
3bVlygpWHJogy/4e9TiOFaCCYX6B9piMtnJOInccslO8eT3KUeEkfKQfH7ySwCC07QBZ4KdzSf1l
eEJSPFBtwNDU16/U76Yj3rl463ZW/7q0LjaPqOkFZ5zpZn9x8GVo/OjDDGRtk2KMMEa6w6C/Dn1B
igPbGI4zVb9R+qCFiD6OmB0gS5ApSeIE0D5uTFfFbnnBEiqW8dqE7E5gQHDf+NjpCB7X9x5pm6ZE
GToyn8QydxfQddkmTvVnkJmHBGXIf51qm+SK4ULpX6N03NXSPLgqWH2+kbW+6Gs+SCiqw3mIpy2C
z9ha3oi5klHAugCphkfsoNsPZ+tcwxAN5AHU91VaZGku9XnnD36VaL4tM2AjBZvbLW1YCT8rRGUI
XHxLn+3ta6pg2z/n8wun6CbsEXR5ErUPlw+eDiz+U/FGdupsX3uOWR7v/kjFzkLpU+xs7UEWBOya
/pabyAPJG8k1vPd/HeknNtGWx+pEUFt6YpjSazrXbYHbu47XSHGLO8HD71vFEoHm6UYva54yfwQN
i/bmXZ4Mjyn3t84ZdxqSZqEY/5kvL0nvVQXovPeH02gsdMy63DppKs2Rzyd/N069u3HASjJY+hRC
8PscLf0ryNBM6q4IB3/gHqIf9FJQzTQzCTYHxOlnNMDEt7EXJLAG0TljYWJYt+m/Tcf67Y1qb/rG
YXoJ05OIiHP8SLHkSSoZU5kt0ooR4qER94NpAhbzN3WJbF2LNMLlNWyPnY1amK/v1E4mpm/bhIwX
V/mu+iVaCdNNImri4qIhbDF0m09ax2PKOlgY5dxJdG9EhDvIpJoMmIGLFk5CS/jW9ffJfB+eP6/s
9cKFAharBhsK/jWSuWRQRMM6eSkyDJ2Sd+VISEbbeUu3niPUhmOYTegTxSA4stpJsxlfvkm/OVVK
JlxzPPS3Rug8pnCovulJf/QKMvjCJsVe08Jk+lxzRhPtJtFgP7vh799y4/rX5JQno3lSOrB14syi
cIf1Gd0BFAkc96Y1HC+WIONMYlrNoHe2JksjuQncqOp2TTi2GGj0wWuxTEZ0LlSP52/260FAL/6u
tfEXMMqM5pVF+eOo+ZNusJkf7XGb6yaftEBz4iMNg67WzCHc0zCQrQtXOdIyFUgJWLVKn74kW3WQ
0yZEv1XeiV3TpD4QuNdANxjeUe53kT4vmromDxqk01H4fF/D/b7lr/b6anfK65ITRgM/dgGRbUJi
bBmAjNdGtArNBgfBnIcXUvCiJZj1YXPBOKe4W2mjDYkt5pY9T18Iui+KkbHrHx/xEAmIcoovnwve
lorGmSDoMz4uzdoQaMND+XDNf9lUTrUW3H6KNeAhqAZ2bpg8qAj1qxzsywsV2wX7uTIIxypvuN9v
GsVAQPF9niYsbJrSZXdp0r/07YQcgdPl7/W2jDE7uIBSLf/eX4APQsQSjGkxs6Fsxy76NQH05MUj
O2w6lHpwY+5/G9EJZSxg+1lHK6Vp1LmdeHdA4zMZd7wkdMAieV5mVvs8uEL/+SuESWPFj1S90WOL
gcm5hv68RgwH3ATXMyDDLpJrJyDkWM3RB2xzpWvQdPMmx+9Hao41i2m6TAAFvEh2Qsz2GBRIWtht
Tf5eTJvzIvswot3gKl/ySxWFTR3Z/4UYRvRfpC+bEBdF5xfnSPz20A7uj1cLwVq8S3PNz+oQZE7q
TaKPvPiRORtenrW/G0CDbYNk6TvOlhsYcdq/DRouFkDYUIfM2Hgv0PBWBjyy36g45VtJuXUdOmG2
yygMmmQzsMdoaWDCIvd6oQM1R0Aq1dTkvh7kl1KgcM71tyDkYezdmaK9IZcm6OJgJwt637Ay+3PC
bSQdELCNH7453Ei8a6WOXTMXosAkROBe51PJoqI8IOOwv8LdGeBg+Yu7ueyEXa3rhQnTqFvzfuSc
SVJHHmbt5z3fwwQlpC5VNoXgl5IgjtH93wZj+B7fKHCYFfa26gHf8ArGz1+3TWv37JAUZxxOCBoH
EdxCbkPgF28WehhLEN7h5QVq2C+bjQmHdC0V8AD8JB4xNYH84bPdhMyeskAmV8WJN5707seo5IFC
HL75ua4r1aQb+DAqt5h/jn/et3ym2URNdF/Cz/nhYtt3tI18J1pMPB59w7p7VzZEFFIBa071chOF
s0L3sQaXROw418MdiHpvwwllg0sjPaJMCDhZMMtpaZrOHAp4Mro0SSeV5uxQKZcpHeg5ka6obREd
D15KL+RfHuLvBtSuQVBoizmfrhMEfWhs9czTMxhY2FfhVKi8AwvsYdpDGwQLKkZzDY8/+yHoaPOS
zGtB9TwvxUnwqciSdOglbDjh+ulXGrgPbJ9cpRIP4CQNFWL+7s158DIZpWRDoFRbs5/LGD3+ge1j
0cCfJYLw9Nr7erfvI0Yawblw5+jmjNgTRrCjECqpkPqcf8DkiaUQ1aOHJk3/tbQooDiwtmYnbVvh
02chh9xFwMWxiuXTCI6bz1AcbP9dS2BBoqiy2IBzVtI6j0+K5AormrgfwRgoVuj9qcHdYHnMRIy+
PE7FDNEEXGivelzJHneYbgZTghSaBnlA76UNlaHxic8dyHtJPLRJR+ibgOIfIMowm6hTgqwARm+E
CWlUiRvBdm3RRCfFyNi6/PZyXMT7IarVsy1fxMAtqe4SLq0mIbbgfOhMmmK3eWsThftzvy/4lECp
EcfV75nJIavAOniDJynunK6mQ4WSYnblcF2SJmhH980otkiHVW/t0aBmKIQ3PkknY5DXglOOAg8u
uSgSJHYe2b/npfskLxxHqSlOH4csOXnqs1rN3xmZ0dqYmB3FFy/uanIwsvmF/mm+QRmokIjb5V4l
4/Kq9yfvUGT8QrqR67TC10nYMSzTG4UWfD3E979rHBJnDMY14Gj/iFm3C5AEzHlSx0RBqQ3sbU0c
niL2NP4euLXCxQH9S0Axfq8ArejnwtHl5gXH2SQw6eHb3B/WtJaw9uVEHGIZVd0Uu8aXenDwbssO
sf3Wzzgoskh+jJGcZGRMtwpOVY5qvPHjwI3LI0lVWXGSJTumCIEKacXmKIIMJ2HLQwerM73s+aen
RQ1dCCklgIQq99fOSAdKlwpPKNmQ59gR3gtCi/Z6D44HQt9PmnOmVuSeyLltGh0sNYwJqeGMOeP2
2wYSm15L/xIF2pXzhbc6xQz+Qs7FEDaKf6vInFl/ET51nX8lu2/BgiK6bKFkshj5VI0OOZ5LASoN
/RwpFM8PeQuJ6xelaNccQWmmkEzQfzKL0S7yeZBCMLb/FrtHNVZhYf7QOE4+GWbGYM1up05xic8x
YX2xjhNKnFB0tR/yXRfSGBKNw7Dk2x2/Qtl76avl04pOieLBnZ6p1Xai2buBdEP1laSWMC4MHkHE
8iZqKU1FpqdGcJdXXE4be7j5w2KVxOamXI3JeLWJzrwDx4cQdnkxOypKaFrMFu/JCs3MqpTZF1ds
At266fFHCy0aaoNd/oIcbfN6abM4MpveBGDHb/tRnA5qdUc09VqVOel26f/MrMlpHUS0abk0kdeP
jhTQR9Xv+6xSRoFUUS/zxgddy4VqUIDDIPe9j9weyTJY0VtnSARbFHznemZkBEvU0cvYez+juAtU
MFOjj+tHwQXfPREBYvolOrAOmFDp/Xd7XF3Tln9F+hwEDbXf2ubc98VeXmLqVrmoGW1+vijh4nTx
M98N4NqDu9DwzDY4uo7IPzSA0MQUqYVetV356tZtfJMs71zBDm0vsILtqDSoR4kGTTP4wAMN24X4
z1wKChqDNJGowBs57BeuvfzFWVOCOwruzrsAKwm/wTJC/Q3D69S13iBdG6kAstfY2gyghr/V+QQm
WRboqHnXed5NPzUp3fLVAKcrK8a6+WUcMzHsVz1ocybI+rQJMdxttCfCVqjisXUl6D4fTpu151KO
sLp/kvuEZlCk4ulnPQ+xTnXckO8dzoSZUYhG2bdrNSXEllPbQ0YAsXiHHb/0eA6BDCFoqbBYrveL
SXdMl1I7JtklGhkFPsvyIJmIe6hO/2h7Ory3LW1pv8DwvajoDiqKnCrjUSQK66o8Zzr0Jje3P9Ia
mFPiINqb4LAHHFfFhuNKVvUsAXUVJO79rPPO0WdXxSJEbB0EzY3o083ntSxuetiwXIrDFj5IvI05
kbqGhpQr9vMHO1JyjF9f91LC8X70fn8T/dK0ElNZINBKcHuDxSvZftP4H0KvMwBjrq+3jg1+P5zG
iiaPWOy/PKauJ1bekf7ANlunD9+Q9RiTcoI4ul4yNa6ZLnaRlBeU0E3ctEUfqyZqxbjyNHEB0LQF
DGpoJCKZ5amQmzS/oeCQUKRalvs4b383c4NEZ1LYN7xxDeVWQWHkq6H3OdAYr0EfTvPLn3UBCFbx
wtyk0SlBiOl80TB54wr5VZxbq82InO02ov73JhAyg+jgXeJTCnG2lkrmGrh6QDpdi+SehGc1fUJq
VGNhJ7PhjsJ14x5tyZv3ETCgqXYd/wQnfQ/wxX5DQwy7Wg98n2BSIWoHYJS99121UJtxX3vmL/qT
HYuOaDtrSiSx5ZX59RFla1ulPnh1LdolAzPUGmJPwheb3RKV0t1UDvS2kr12u7w9tauUBLOYC9yr
wEiN2qgtSWUNs4QtcuT8CnOF7Pu/86BJftoyyfMC8fhrOlzXAeo4Sex8A6pFqbZwDo2oTDnKT/py
9to9SWogflc603QhEerM3FjYr2Fg2LQ8w/glONdAR20wv67vEpvy2xe32yXfVwcazX0AjMkUtEul
tS6rlrSZ25hIen8TXrmKFbrARtNfy+UtT0W/ntuwi1MSkntafWvFGa4X8arJIg3q3i9mszEwPQoB
yMrLb0mjEXDjKzlxiB+gZlThVz+V2kN7jqmPLLdCJjIhmlwPvT0lDt2hCUmM9D/wkMCQ2/4vCM+o
vEXlxyC46CZVAzuTtKgZF5wr08OYgmvHlAcBg9Mt2FxPC9s5MDjaFQw2Fko85/KHnbXSBcw8RlFI
tz4fVvoPbkxc9nXI3rMXAmNJ/Ycfe3alr2wx/hphrl+UzZDQErpgt9/i0M2iS0YETeDW3Xn7NCni
VoorZbS1ThQ6ldbcTGS95ZYdTu+eMc4twEBRfoXQO9JcbXGc/4cObHz72csBZ76RBViZ3RAOIsjZ
oDh9PwgvE8QTKO2N45186QRjELgN0KtOf8/nUQnTcba6d3ZoA8TnuRyVHNFWNHz6vSa4fR9NHpIA
axWPNyw4+fXus6mZAyyESYVJhO4BC4NzHpRPZWABAg2vDSCTzkUP4PxxpyKvjP6CnnEJLJvInyld
wkL/cC61w26tUM7G980Rh8HnG+gS8rE/x7fC3hrln732YNmiGcPcDwg0fbsFxnEBAUzPjzpIndrD
6taHyFfXGWI5B+oMSuurZkBDfZtCZKAYzFUvot5u4YxsFD0lUc4JwCI4FuUuAo5V/UfZK3XmECCd
nU9SFwY/5IlIQQZwlpcoYIfAPrbhfEUvInaltnfvCr1mJlZqcn+ToA6Gi2BL4LnP4Gt78Oi2zdwo
aQvWjU+LFXQ45OHZBI3ctyiigicglKmwHneoQbGV5yy1Xl3IsC/DpuZ7vlo4CdMlTj0ETxC/H9FV
UZwAhmGLNOCqY6VsV6GR+bjxL2JkBg2kxAs3x+5SUJGbmN/kCtlii6BWD2q15wkMp2pUpg4+AMAO
4yTlIOsyUsCDn6TrCmjPPBU2wNHRqZp0B02Bk+Wxr+mvZkAdJQBSJ41pr3CTK29rZBvFVj6jdJrF
1NsP8cjm91qP4V3KMFdos2dx2e3wCrUjXItdZbRgtZ52csSQhRwGOWbjC4MvcEtlb3ya7X4kWq08
JBefugOytxjA/K97xSNAc8+7SJZMCOWmaWJwY8X6w2/MR/Y6iTQELGEFogRijsWMBH48R6d5kVvs
8rEnpRwfW338o5ZCT/kbNHjhFjvSCzQN+QosTWs1AID1TjGPfvaCQrd3wXDJyyQBSBM68R9j1k75
zr5DgwFhYwGtmX7tl2OpJ4ecHwDigMoxYiYPsYYpq+rQaxG14zchT/Bxn2rVlftMmSnBXNxGRTkS
E7BGFPKgzyto1Mec75RJ1+HPdfJLhWtWse8GVeH4OA27Kc2vFlm+wxFt3k6L8FW/wcveciVQD22J
5GIZB8s65v7IJZlQrUXqWKBSHISUcbkNgSqcocowJVHmB4Sn5ALyIRVmQQvAquFtzrV6BRJI21OY
1VDv/9uFE+05H1ljQ9xox6cYqoUBZbkpzz3yqPjV8xe2W0fyFG3Ezu1XJfWaThG++hIuyE9J1+Rq
L+rmxtLoLkKoq8Be32/KMTxW4zDEg8esS7PATgf7z2J4P/NwCUXVau4UvxN9Qpr8DbiYOLIV0QVL
EhgE5/LZ4tddGRVUMc+fKgwNjnAoIyEH2FWSo5YmH/HSkwsguHCC9E34pLjbiN1sOHQ0L9dFCHKv
QfLNIIHpLchmzUckClOfp8SeT2FyVZSkkvmLQFCeGyuxYNkzybT2YRGv4rgQHeyXqw6JfEGk51g/
dyIl5sOYP3ltOt5ZCE/02B4C7BQuY1xIA3JGCEVtoXh1L8NQmqx+MSgmA7Om1tELhs5IqkSdo9TN
zzx+WBRPjX0syPq1943axD8PwosDu8FB/WDRzjcHFkuVJoMYJ7W2WKy805F60qIWSKIfPWAhbemX
APoHuEh7Y127TizXuGB5lFxVDqPRNZ49Edhdhm1RmRcxcGQuztuxK2avRDrK4jlsf7h7a7QU6/0M
icfDRtKxvyOCfzo6dTBAiepEQrBOahSGb+5D8tJISkPJSVDKwUVVvPq/63JjD5X49gRy1BfAGdUi
5Pc8YhNwXB+ej9vX0XhEjotYj3SGJOf7T4bKKLWgm3a633LCWG3lHDK1XQzDAm7LvmXcrE98Wx91
0vAp53CNFpPpN0oAq8ZIBvnvRCwgsvycvH8Z9X9Z2BFhp9ReBOPRkxv3lIA5x3IRaAaT474Rpg66
teeu+YK4mcGUjFWO47OXt5Dq1IjkDijyfR+y/rTRNP/TqS5O6eDtP4ZxN6qfiyHnIJ/Ktp0/2X63
ZOhVs1wEXdVWEMxs4l1LWXHi6FC1WwxRsLY75wAo416H5fj7tF7a9U89I0mhyKEBscdfV+PTA9Dg
/IMKOFz1WaLMjyPgqPhO+4sp6NV9gNtIQ/QhrnvMdcu+z+zkadFN/2PV3d9X08jNt+NL6ZaHOJPy
OngM9X5dHqg0SLI320BN/ojsMrB+ZvCO0Q/1XauczXkxPS2aLpdDTY0DgJhSbL3VXRoyVbqHlwHM
JxD+5gxzUjmfjWjMpKtc7y+o4kXQxTscMn30X66e8AvpvmNLsOOK2YI3YQGiWhFDFTZd1jgSfCKI
iQ+mwP67w7U4kpY6dwwPXWtD7B2/PUICc8elOW46LB9YQagjp9LzQ3OAR3QV6jDFu1eHy1F1/TKv
TqyDxLrLBdvzzSdFRLSy1hlrGmL2V1rtrlXmEz+0+uIO8k+j4bD04LciguxqdbYYQPdC+enmRftD
1zUBl673GF36cYadJTnKNH69k27HteI0qS60dNqwY7KCa94f35nmaUwvryjaLShGzYmBCb2vAV1n
7Oj9QSEzraiy2eKqv1zsmPjCcXUx9nNUS5mHqOQq5/HZJyvtYGJwgGvJH6FqYmAW9hJotjZkRawY
oefY39whHZeWxoGH5d/pgitvf3CGuxLY6X5708lZxv6NEQv72e0kqaIn71pzCok/1zhaavCLmLte
HohDwiBXdF3qF7HbPNdOobK1w6qFwuTsotFJvECdJDe7f5FKpNQsWteZavZyNa1Z6HmJLVgI50sP
V6FagQo9fsakXLLck70KgCMTt2nJbb7VwMIxZA23JTY7XFGTccDJtsypE7xPfKHFSdvnaEdbPdqP
jF608wz1nlHZjlnmiKsJTsXjXn5n7Bc2pK9yRD/oz74ucuglWBRFhQrS3yMpZ+MZYZ+AaFjoPa/q
NJ+eSHQNmh7U9JyPwHVLSpXROsbHA8Mm20/w3q8M9bh4yP9g9De0p/09hMeFYALv1V8SDW+9+Tgw
hA0wTzYKUCSBt1uVPRx3s7AqBxBI51/jj/GTlc0Woq7vDnOWXVCxddqPx4CGF2qq2DNocdZKlD4k
Ds28HPi1T4TyDoMMG/9B+DG6wc6RDHAJsEf7hqMR0tzNfEggglBAGz9gbS+osq1eHVwuy27WjsYn
pW8OG5axvkT5kh+qvYEW8lKF9UNQc6kkqOFK/RurctVzAslsNGXqg3KuflitiScSmRaeFdKtUY2s
a0xMKEmdc8soeVaCXzX4Gj+CBR9OWP6o+Cez/+Yfp+ZJsrfaU/8lqM1+Zom8bLx639DhdkT8nrdm
hZaI5s+e5prx4iFnkXnIe1tIsxaeDgP2R4oQUwcqEisOVV+dQqzP9LNRqZXp2h8Px4zzRbjjaKNS
dYA4eORYNLbf7GmI9s7r53eA7kTg8UfArwZ0Enen/07T+jQa6nq+7DJmBHUf2ceEK2mC0j9e8xLo
+AbE25Hjw7M8QgQVjV83JMsb8XTKyINQf12nqfeGJA8ItZR56OB9fWvTEujr8N5ZdpYacPGan9lA
UTu0U0b8cqMyi4HuShZK4zAYu4zp563tSAZWqjiIERVDFkw2a7/92sNFpE0x9P/KT7n5CPCNSU9i
/4iZ4S7UwfNU6V/2A6+h5xFH0uaG9CobX6bE/zPqZqH3U4sB2OVZRNzFD56JiDxvEb+BqbYx30e+
vnY6Rstl+3Qbq19j5p1afhl41yGYTDoE8YiqMuM3BB+Rm1iIxuhq6aMXceNWZLSdHIV4tzvLuTXH
7WlzxOoPFmIlKGWklmCw8TXywyGtuvK3lsQV9/nPsKa5HwEpQDED5dnSmNGy8VPRY/txe3mfoYUm
joJvjRvnRfrsCuEjxSxH+4HoCCagBp8jR2fG3lLIT0Qv3JEH7jkACGkAFeVO/okJ7KBTEEwv1G8U
k+lFgxfgM9JqJ5jwF8VpmzF4kMqnxilNCYYqL8qyx7ZwylfPL/w3iCKbCeHb7BBWnKGAK4dMVwc/
pKVeMVwixmEES3ZlucAgOkGZVewyCCTanEpTWCb+Ogc0RpA5yWmdlzaERPtm3vmEbaTYzhA2Af9G
tHSo48gRAwkGGoqNVr4F8JcaVOFg75njR14fQR/b9joy03tHjAue1fWiyabJJIBdofSrVLWgC8bg
m7eogSkeEHXnYFRDF/d20KPRF8eQneKfUhAxVs+zANqc7Y35/msNpQgQPAuulxbmh5Uub+W+m2wX
e0r1gTNjbAY7o1whs5fD82OIR7aC8ppOCQnev8lu76PBRymHa4X7alIGY+lQky/3z9mHhAA5vGJE
Hdl7dwH9vLcAKwoJ8ZY1EELMFOw9JcxX1QhE4l8WGNnvu1tjy1uKZ+3urYrvmKvZWR7HvpxWJ0Pl
kuxsSdRHgXt9v3JvQcf5NsYq8zGW5or0oeFxfs9hiKuMMRBYMWknjckufy/4imExdiUMQ4UygwOJ
KHpKxv2vFWD2NM+A6f22tzPHaMCLFVgL/zEmfgtuj7sHbsiS3gRADFsYz/fG0X5kJpitpWaCwbht
Z0LQtZJGFCk5/vsudlnb+S76hCdbWl1R9fwk5K6vOF8AUcEJ0UiRwRsWzDm4uNsNmncYIDj48p5R
STfNFGZdNSUBcevbiHYIzWUYdl5T7pWlnrXXJ9/mY9OyZC8f39luP+6rXSmU+Yb2hB4UUDpMiz5T
5C5AmFr3rOCqmjvsrmmRGfdQ/syfiPBGoA3977bbEhvtKgHG+2PByeV71hXojyR+g/cqj19pZd3+
WVK4RJWV167BVXgy8Me5zuEjl/QZYfoIyVcRgpNpV+xErpZeLAUPQzAFzJkPACZriWJrhWfXX4/t
G42Q77Oa3fomh6ZjL3zPGvoiTwm1L+jbkdcirVd30+m2CItIpjFtsyBz1V1wU3duOhKvMkn910F0
L/NTZY/94FroZDokWos82BoGEB8tCPBiep5emQ3lVtQ9lINYXA3I+4NLKteyLmdiApoInRcFUouB
e/hKQXavllKl4+E0oSZQseVInXt8/MYXp6aVidU4vofmiZkFJKjChNToPC5SLDAp4FgjVdXrn2lY
E1u7D1cP+nZEaSHVD/lxh+irFTbnb9SccXTJknSP/g17aHDaJrtIuDLFNSCU2W1BK2Y5P/TLnE65
nhXarTiusBcR6Nm9jozvPrAOuxdt2f89x7L3jLHmzoTaY13duXf+QKB8bY9boFFn8ZpXK+oM6gTv
8BFNJfnM8OG+e4Aj7WoPYcHpYC10hef8fHxyzfH8kPoNg5E/1I1jxhJ7WKWTut5//bvfGWdJ4u9Z
/xiGQFVt5npd4KqgS9X5P91yXm/+0Kary05H8JIlRaXBGB1DY0y+TU67OAjV1jFHmfMQDqydiTbb
R4tLb/EoxT6R41ppoy1apK2Wmv1VUWGMXGzgM+Ge6fJIbCsPbnwEem0wo9jaek5z4Ax3VVWJssRj
/4j3rwHIFhEfxl7IMqwQHgpktrrTkAfnF8FX2ApnwXUJKVKmk8Hmr3iXsfJPFLv4t5AHVzrqa9Pl
01ontdA4eH3opdDlbUVV811OcpSZVkUuFqmM0b/HGvyxQXfBXZbxtHou+xL9QWq4Vk4SCEte9P+h
yp+G4KC98a1XiE7NeUlFVUvm2BE+OgH/sg9ePjp2aOgpOVRUToDhq0bJIVbNFRJwQTr1XzAs9vzm
JTnY/CUA4/tC0O7GB393E6v9OlOFKSBqpmhGn5CoNVfNX2w3PUQpb4tKYIGnX9uMZ61abjRci6Uw
F2STBJAOe1SgcrdCXl9oEs6nGr0S7CJZC1mgOccV1zHCR4m9V/675Jz34wYUf0EE8PFM9jAy+f7B
6mqUGIXsin0u5h3FdBOHurtZn7YSJc9EVvnh/W+i8PJHf9Gfewkqi3BjJCoGUo4llrPvhSy8RmYR
bBIVVIN5ZXbc7vSaLUIiWMI17yd606fKICxnsrxvkxJhCftnvWxGIsUuo/9TdKMJ0pH59J49JPhQ
oPPHEpjaBYqnGQVrojW3vPz9P0FhjRrYt9MV7TPBxfrV+iqqLfwcUgFy+Mt/2giuZrNqg/sFp+PV
jlLg2aE6Tq5xEALCQINIYKljPgd94kelAn2Qi2OiPPNyQ10P7StDksXbWpNBbxijTbdm1iEAlBda
auv0nVts24rWLIloR+hetwKaQutOrHrjomLArrOn0K3ei4mG8D8bf3/8eqewmnFq0mGsifGJPK46
r857AUiZ9HZyHiakinhZUKC7gV5yQJ6Rdld5kuUXeNEmnReEyOek0FVmtdr2HW4J101csBiwKMRs
32mCvIaTp0OFzh3ZkqM2vnfN/HirBW4/VCBUH4rMoIZ7SUucrP1wP6KYYykSSH5M8bJqnruNbttc
tDhl0N7QcBz6MNY/Rjy4YwgElccpgtlV7oB04VVFnBjnU79flKOf7JUmA/HkBMEYcFtYkBKwy94t
VfROXplSUXg+WCRzoOTsq8QM90lJnjzuNk3pzxZaBg/6gZ2EvMe5C3xWQ+ZuUtC7yxoZTSm+7cTh
WIewu+7jYBRjuFS2gkeWWcrUMuTOFdt8+O1DsTqRUBNSNLVMb30kwCa91lm64cb5Iy7EM4WHPjmo
Bilp3KObIVISYkdJj9ZAZg20CIdctxzk2YKKFV2eZ74uWDYzOTAFL9bfLuV2u6y3VKncZfRsa4fA
27Ea9l8MhMTWmybknSvcQYKtAWd10vjUpMgF0cvdaLZx966wVYkUJLP7117JC8tFgSUWlkurL35R
DRwaAQ5jsVZSJOIj97tCqQeIL0GC0BemsPY8xcFvlwuA8aQyt98RjxCrM/xFwklyH/DkjvGCUD6V
iOI5K6lZ1SFAFsBuLP74f3LP41sw6N0dfYr5/w7J0NOGgcxvPKaR4QKeKRwm2wsng5BTvmAXEtco
au5WYV5kuGpve2+q1c/RSYIahMv7FRVI+ysK/hdIl1MSdNMWfIm2OOuMOQ2XCNfLQCFAhl47eIZc
gz5WL/nNF1iqGzwrqFGZudHRhLDWsjAzLCjtTm9b0Xuv6N/mBaoXUplHWQdHA46XCSPKf5EZDXGw
K28n7KMrxpLYiwqcGPRD10k5/dcb5QlRi8JPCllJ1scffNVHAhuFJ+MQFSWM20+eeEzpqoI3PBIf
LhpfIGqyRYgCank6yqU6xFJFuvefZjzm2/JtrQYA/86xUq3N/j3avJiUY54vfTLp28KNWJsyonbQ
rLUV1e494UOQLz8UY2XqziNP8lqfpfO7OcVTu/cyBjoYnBtzgFwupZvYth/V//Ek8Ivx1ajqKlxr
bLybXTWP0QBXNBzxfNM6JE/m4/NNP65ubwBexo7ks+1ygoh1qeyWndzQQ6/aN5mS2ZWDDl82MGF4
goHFu3C0qniWPyjjt5r/sTpQx/qdT0IpJABewR1HtHaZ+EdbDArbKEeMv/LBZu561c+zQp0fDioZ
+JqV9DAELFS3yR3KS74IP2AabSdYI90M8W9F55s+KCbMhkfXxJqx+FX0gzvmU95kp59HuSKfbjBB
ZyjwQqpdzuDmCMqcIJCJNH0lo1phxu5L1uKv05bqEu0RhBSU/pnDfjwmWy0eJIEpn3rsrVHQFFnH
4xuYVk9p5IOCizcM0S06ehylqdMQdr2id0WgMXAAo1nyiI4KflPO8puTHFJ8rNqoG9RACqhD6DDj
gnEsn9mhyMz9/3yDGYDSGd34potinP1a7tpQZBcyraSDwew1r/Mb/Qr7Qr9Fx5NLS7bsTpzGfMUU
WIytT0Y6et63RjHtnfTYL5dfh/VORLOYM8VUx1ugXzc1UZhpYh6dwTlGEXMUZEMNPrlqRFTrqODs
EiVeMf0+qmOj3r1pp/qyDFvK4jkoH1npM8K2FXTcAGq8PKXo4VwIjD5onZLJjPPWNTaipQEo6j06
IRWKWL1QVZXvc2avOi6MeBHwa8vgIlDKXOMzgKDz8I+JxLRgPzRZpb0xOA+adrQvAAsmMVABGhQf
5V7K0JTC8HjB4YlSwcXLx7nGeXXLBUUD5Er/c4czlKdFjGsSwIHJRBa6mVj+mkQpwvRi8bVHO2rp
fUuLdAjIRCVboTzTPLHLTJA9VNO7l/z5ZLbfoX1SIDAAjjGoUyCqAoe9w306QqaXyqC9sozhyQKw
y1tSJbsH8QA+DZbTJ1cBAtos5jaq0IWYz8fPBT5RFHP10umqp1UR8Da2h2KXoQEV44rI7meAsxBG
QwFku0zY/mE4VaEo+V0EIXvn3epE4qAyGt9t8fYrNU4OUKFhqZbgAPdttYWfDMBW1rwNbPOVcx8c
UkyRYuXigCCzWwxYb1PmASEyx/eJFW2/VyQBBHb9lRFO+NEk9qkIC8NweKEfFbKzt5zMbDxauHNQ
e7SZiiO/Hv0eG6h7lq1e8v5+UggByVW9SlgfCH66SV6XTmlfQYwJ3q/52chsB+F4anjV8ym7Hkoa
ZeRq2W/aoY3/6r+nk8lmr9YqkqXy+xM+b4rZkOBRQUxCnp29FvUYPaK9AquAtPWptuPrWzKWjWpa
GmlAAkdjpRb0wLCrqPq9Zl9770cN6zTeQ7cW9qZO+rusFriJeB3ke8atdvZlnuh9gViEh2+RUtIj
9AXRx9zLxezrZLmZApcleKQFth3ais8zSUrX+m/DlzLlihmfcygqy7pZPyExVPl8gsnBcsueOEBi
RCK085hqRjsgR2sEAd2oGWxX1iYR9gMfp8G2FTz9YHI7fuUr/i47JPkZjuVtsaH57Ic5GJ4vjPgR
CXvLLpCPTIbZMghRMLcswpLjjcEgvcCKMN65WAzMmrggkRRyOP8aRP18ISRJy3xW2Vdz1nYi3Dda
WJUk6bASbjohTNAxyZVX6jO8uRYlsbFCr/WTMwb2Nv9Ydc5mN51JKz6vszQST0fYL8k1Ox+QI2yS
Xp81tC0/CJhk9VaG0wCKBAtezLEK/UkJTaQgSauAI94Erg78rEg4dvz8wAbf7smzhpdQzGQHPRWO
zWzH4cmSY8vy4R9pwcPlGJgNWLXuhMhYOWQKeSrDGjHshpigGe/bbgoB3NNhWX60187Se5jgVeWk
9/7zKP2Uk/txALWx76jOnhUfLsJKH1JpUnyKwTV6dbgjEwfIADAdyyaKDQUPRXio/oJKyKFeH+/p
UgRQdlb6Prb1XtnIS/P2iBULafwZX1uDMgueuN1mPGsqiIiwGwJN0hIiE8ITlmvCU+DhsFERcHv4
G3qnhC09wEtxBe7jKm0HBEmzHdJ3FLwnHq47p95UXYeUhcAkOXLfV4O0dd639ETqjTD2tlvkHWKD
ukuGdtzDEPu3tKZLcim1i4tlOn66d/uCu6dBUi003RK90ap1UktS5ddYY2nTWQQdUA3LROw6L5P9
YJuYgjThxofnwzCxocAhX5sYglNB+j6phYfaS8R1I+3WNLZjbe39w1aJDz9VNOlUdIp9yDNH0F17
7sRfIL+x1hJXUhA0nNvLWYjR9UtismNgDkNGa/dCxpc+clLp6aBeYAddDqQGdpkIFwvYkYi1lOtM
6aYFB9XwrpcJci8+bKuv8AckbfLKoSU6AQy4HAe1W0xFviC2h0/cy9fWqi0yWxOgTZuoOnjpRFXj
52yHYNn0xFq4EIjEXktqt8TUh6Cht5bVVh/oCLxqXqPJQcSWw8Xt94Jl0B4C6xPvfOk2Jt7hxv1F
LkrqY5V0EsWBNU54winbllyPjYziWDu21g3PsS/gRgitDRGb4r2YTkdDU9FZK8dn0mh9qpJM1xoM
cU5yAaQbj2L45ug6ErnU8hvtjQnOSxCs9g997MRxg7QSkWa9wLOZVlOsCa+wAa9X86m1OqlvyoMh
JSjm3AtAjEBcvzG1zeMqqdoOwsAu/n2a3myF+YnkG3TnzK4nmFkXz0p296VyXOrgNEORDWMAlg==
`pragma protect end_protected
