`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
OvlwvZLpkXPpI8t1pX+dhixMP70+lHoy9pQ+N/HqvxrY83Gm4XpEtApO9TF9qHOUjyC81/81cwVU
NacawZNZF8Slej4BnoI/3usrN9thEH257K10Cxu+FQ9lhmqyJ6LF3yb/+igjYDo1tXmgJ3Ilyujp
WK5MAxGMtMOE71x17YMFYWymz7wDxUqIC9Ke06hsZPRDbWA7r1gmmfG2w4tKPvEiptNd2W+yzQmZ
ryaYWiQFmue6/kjq+tmgiG2xO5KDHw0VZeCv9xvrJKwHSS87/NhtZnPWY3STms8kj3BeUQFu+4sT
6QOFmNNS7xY17U3mwzZffXRsSoaqjp8HohIGjg==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
1e3KQp6EnbzF7WnDxt/j/Nlmi1J3crnwdZ+pGgK5H3IqkADFyx2dV4g0wxd0ym5cfS05bRc1V7jA
rGbFT+T5eBP7MrXyFYOMzqe+jIinM8I2QJtZknqYvfzCtI035WE7c5HIr1SYyeTndjgZhM5ovRse
nOQpNhppm+Q0KJeQeEQ=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
e+PcKQ2sWJr0laIu8+R0ebfZXtAdZ54qUIjg2An8kKAd/C7KdiXOzb96RHsVA67S3VenPOec0LCh
fq8AlYOMAw993JSaKfqmIYWZcyNGMw0gPNumMSX6+8i3WMO7Tt/e0JWGYjM2LYP26doP1OVBGOC+
2We/Sc7MrQnE9zkpjKA=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11520)
`pragma protect data_block
1yuynMGRhbZJyVjDv5Fst71LCP919AvfWPeCb39JdL3ODu66yLB1K8MmGqIsBsqJIPD5ddtT78XS
6QUIz4ofellTKGwhpwniu+iOYDQ4lNacXgrlaKoV7tKo+6l2RZ+J8kL5wLLDmBEf86tk17S213wV
mU6AIOPfm1MDcMJl2BC4UlAxvRnEurxJr4LnBUVi8T3M8KYenM9Bu1jDOLU0lhsBptckfoSmYz3M
U0hDvce4OWmxur7nlhIqhkrawhR8WtSImkQSrUmtqkM5jHok0XmzywpgdXtAroYnAyBiryfUdITs
GeWy17NcaP9cDobjpcU/MJmP+JEe+0ElHuzARWuvfe7rBWLL8AZ8VdkJXMl1oqmnTiKMIHufNGiE
FOGtZ16xOl+QLZhQ2486oLfNb65xRMseKjiu3DXQmsNUMRHRillgKE/hmjIdB8yMM58ecmvFEpZM
MywtfvFygHVp9ebsycTDVTyfc5CTXE/cfr4PvanDhoejmqGUfd8sVgVpj2nUMI52ydm+/XyxQ/0V
PB45KB39ueY4B8MgSvmbRfLmzOZlLWIYi5E+vLeAfZJ2Sa4khLJqS9o+0IrrcPXwdNTaua2XKLlW
hJi5tHLRm/XIaGDa+HADOPJ72B9221BUDXzqVkhd4c7KKKTmDHenWOxLpcuTb3eH2y/r7X3Hxihg
1A6cby1lZ4kznDB7OWVE0+Uqtzm7at6O7Ii+CUC62W88Jk0teyzvW8Rv3JC8J+a3ke/5IO7AUjpe
10T6bGYmqVUQpVe+Abt7UAhvzC9PFSHedsjstme23xmK1dQaBceaK0me6xwg0jusiUMaKQlfIDDP
FCaNv+MYc7DqcbQsfGFjxIqiD1GRvdGqLzRxd7m2a1cv7Mq0IFOmhRq8hRUuU/nS43SXH7NO+hHb
HgcwDms6QmetsylKs/FK3LN58fiFjCsBlLsawnWX0jxCdsUG0YhtVxzU+7Z5pne6IWWoT0vP1UQV
TIeTJpUNXpv86q3UWKjEjqqH3kb5vscFGyOdM7O7nzpL9IMDM917jzmady2O60qyLBLmIsYEL/St
3qqtzEfqpNRDN06D2iQ3M5jE8YCuRN5uZ8tINxSENa7RjfgDIDJj3Vc1jSALwclLamGyM8Ou5PDp
PptVIEvrdR52xgFBoOrK8qLOu/0fCn8gb1ppPnTqcMcoN3daS97XXFMsPNnGbmjGr9MqkmphNGVy
y2JfdWjWVREOBYVCrMIqPTbvEKnreFA9cgu65lMR4BHVQAG+EnBmbwIY0+cwpGhQvPkLG6I3i0C/
ybf348GpCd+z5mqJMRGTdTcSaw/es5MTzvtwbjU3bceNj70/h6CMVIX/nEduim22L1xAiPGJhjfc
Ns1SY2yRKFk6WTc/Gd78FZUnSjBFK3GEU1J/bY4hPGK1Elb5h5LDUwUtdmBZgpLk1zu1alo/4QIj
8h84uA12MjM2a4VcDq/bTIr9njn1ZCrlrdfCSFgUpSowkbojNZkekgEX+KfWOwnaGI6Ah2RrjEyH
XZd19e8tobI4R2/xwFKzVaJXq7MI01Vj0u6mkGrmTmsPZbDT6B1tKri+ptaFgWxFbEaj2GsvRORa
azs8T98QwiiuQpJ87r5dwrPsM3XPMKXljPuMfsbUxFEPLpvkF6NJJn+8/O2QEYaCRq4P2wlA7w7k
+X4HKk9k49KGGSD+l0847MOS+a9Rmlp5JFklrHFE8zgXrpU9S716+RqyyyXRLePleODjtRpYWC5/
J8dKaGuFP3paIGwPJpXend4zlGHrn5bSZPBW0AzKC39Gi4YoWPrfPElvu9Pkncs+3y8uh401Pf99
NXEL8MRfnNOcWNGJladBjKzP3bMwmD4CdqyaBKpq90iEe7UmUvFimFfZRvCPyVrFSUPSINWlmnjx
9ONttJcTkyiM32HvBeyoRDP8Bk2HWihUXGN22BJt8cGLcl2qWdpPL22EpHzebQKgEU3A9X8lYLKQ
s3eJXYB57oqrAt8o17ExrJ5961dJS7OLPH4g2ChrY2yXjJ2BvQvrBWGp/mpZ1amYJmyT2tTOa5Eg
9loOWmSq69XugGjdDl+AsG4RH4xcaANnrIgI2c6SugyCL3b5X4tKhPai1uHWI23Gj9616zIEt4LY
WZAcjETKJTr9j/iO9iPsBDZH9iEMO09oLMy/2qViKNfu3xMcai/kSLMgcFnBjNtD3VVlm+aUMLTu
duW47ITeCHkeNyiohXitwkok/9aYIOec4R6AkUZocYZP3r6QnIdFCUrK7ldO0PBi3lieLxrSxwXm
obmLecBXAIJH9oTRpD45kRxcF7YOGxyl7I2VOgNW1mlm93J1+VeGq19J9u53bYzD0h06VBho2CWC
J/5zGa2EIhm5qFTrhpvhw8N0mPnQtc+ljjqH3ZdnUlWX3k5qb+HOqsm3tyiWooAeOrwqCaTzkC8L
pijokRY86uBtENKDzcEt+WREYfWfaCTvEA/OoM2UvgTFWbjppXq2mSl0KAEa7RhTPkJ76Zegh3Kx
2mQX7mIdTGiga7GZpYYpGwCJDZ2GbsLWi8EyCEsf9VFSa67LYwSZIq33V3q8bffgBQUeaeZ1Gd/p
dwDJQDuhGlxi6r2ZqfiL89LnbEtpyJPPhwczx5a0CRQ+fS1868X8iV5soz6Bo3Om4p8Xr0+5D9UX
kODBd8A1mxY4bmtmPxa+5MaLjXS5inPTlokl2BEfST8dT657wrE0Ql2e5fiA6lNBj6utyP+ZSD1M
QuiUUOJRBJOGCuoSpwfQTdcRgBa1dWIpmmRUa98FOW0vs64bco9Aifw6nEmMRFuXnaNy/wkzWGet
bBERs8BmwO+FjhhVfGOVolBhueAWWjXG/dSpgn5itJZajoeqXJSCskyo/7b0xFv46CGJYRz4Njmr
rD7YmWPuBmoxu8icNQvRfqzI+gPuI0FczXX+OpeXU0qoOmyfkUSF30xA8LXZrszs48LXwO6Noe+o
/xyvODBeymkS1bJiVki91276Eei7RveDoBZZrjt/2BYlI7vukImkk2kZv7xpoA2CIJz+cySRCvto
xHu4KtgPMxiGuxg1G7xl0Y7r7lOXazygi1TKCuVZoJbPC1els7k1d5uEfPI9+xExuuXG39+B3IEb
nRnvWX+qfTUY5EIGVXNdna3Zu+S9YwFbAc5Dj8RTbD4olFFjHwxcN3CoqbNplWUQfc5wsKlpv8eD
neVFSpdAltOXXbXXCPSjfSr0p9Y8/s25fEUMfhesDBn0OK+QJWtcTn06f4gIaCaTXTUmVr4prhII
6tdT5/lvOH78pGzm5mhcUQU19UlE3mwMtWByh3AFJ2z9F6/otyr1SAYw0S1nlIDagDbKwQrdLWXx
jFokW1odUj2OKRO8WIxos5TnHPfEWmhXJSUlwa/B1p8nLKnQwevofXd7WEJymbST0ZKPt7kA6rnT
IVrRQJ3nFVpBhfukJVrMq/XuO7+8OEq98COE60+8OvLx9yrfqsvNhVj7z8fliloEyqgG65NynFkJ
Vc96olA3BRDNyPL+UIP77OwAqosVRYemj5uPau0KjcqFD/3Kxaw4TWjhkJi+CrWGPETd4VeuUbE2
bB6yBWbvfPJUrJh25p1IDj4bdGwIPqpA6Rx3+DMH0otc1uc7owQ5umV5cQHp2uFAa0AwJatnNKev
MlujsakfSy4s1DHDBmCNeFS5fjPck1ZL74ydHiwAbw0iQSowbmTsMoAgmMaWIamXpCOd7sIbDrJH
CgJv61Y8Pu1aYfMMskr1YE/88ZvnmCUIet2jeY8sS+c/Qj9m84U0RsHC1NrgLj1I7ZDNHVy6kboQ
S5gs0xblg7QQ+lK8RJiouLCT0IZWddsiRc8qCXeqhs8l5/3WB5A9KhZntqecK13NTU+7FHky0nqo
ZQUktChGJi1XaplHB8JKD3Q6XkuGnVUWGvzryg3Shmw6tSNod3VMBlND0skiQ32EDPp7ud8LtkuU
UehUhxEX/FK+oXhtI99yLBKNv3Mzm1UVp5kDUfZzKFAOBk61m69fGMNZR1XZ79kPT6RsHaiRm8ZC
cgnRPOEo+pihCKYNy6jbZYJOmhp0ir2uvmsVyVuQKUNrT6cDJi93HAhawNF6joBBJADzGwQ6uxU5
f3PI3utDek2P6EIrlHBmpdhCcEwVxnrd9auQcJFa3dg1hRlVPZBZWXjwanqOLdJLiiGxS86Yt/X6
Y8KP3nSS54LteLygCGHjJAnHGS6n4dyr6f4YFqq/kqYbN3606LJaI/2NJud7VZpcAWQdKo8/54or
vW+KCJsbT47lzmw3EVWNqhjeYTKgGGKVHJiFutSJBQH+Rr3NeEy4WSZVegzujAPv5sX4N3FQthPW
Blh/sfd+To+jgC9yPELuys4CJt+Uedo8VjxqU8oHCIN8V/8mZU+FWngBPpN9ZhZH0kpQc0/3w042
9gX2jYXYW/hHOP4vS9d4ba84SPCw6RbGaWLr2xIeDR+v0VRlqTklnfs6gEuWbxvj2YLwPL77IGq/
xCZceeZmzNICyWMnXSpqqXGvRaKDW2yI5E1c5Wfpr7qzHwNkDAE1VsNgoRFjI611tyovR868OBjE
Ditsuzl8PfnIQFzJlSCYugX7nF9oVIgKYSpxwOazuZLoqeTlUuYEgJQ0I+ASr5dr27rwRKx/Xjp7
ADKP6TvjL5essLazX+0jlVlvNLjjm9r54VRe3GbW9gST+YaVvB9+5WJGSs/DyyD6BAlEdQpNpJwn
dqJTcZPXHi81uC6l55p5UYONJ6e1D0JZID+Cg+HZd+RFr2AS8Q+bzYzokKI4drk2SjRkqGv0FZxw
DqWobRdxtYkYyTMX+qxL5NNNXhcZhX+ZI75FcmEQloOvjHBrsJt/pXwz2MKZYK9obF8P+GrVmijb
8Ka5gG6nt52ezAI0Z+zoQuQyOFBfQrOFyeqqyGz8iPVM86AjJMhSO+QVKYbDTWgRK4OBROi/APX2
g+azRD5TuUWBCPkoanHmtuXuuEbyA2P3hQqfuHBq0X4zO3ykEqtXIrXLiQSTd5unN/G3nUhCvw1C
R/qEKr4lwN+G/ZBmm9nbca8RgrW3gxitaLIbdIOiTpC80JGtfE4dyLMkX9Cuhjt4GFn5g5q8nxPO
pAWsuU/HwbGdek35m5nFSzFHY7z44hJOL07NGN7VXOGj83K6tjVbCPCHdCbM3i0+dj/nlFD41yho
5hnXiQvclONk1THCWqlqyuhPLtFNtBOFcrV1iGvZC1ptg8TDJSI+WMuzN9o5h/jkk7ot3JYXLtpE
FsmXLVYc5pUPZw/7lb0p4UFeoNe0ON5rPobudf2yV7L3mP/BzOPJIe57cZBxLLmqlyn1AiwToSLY
3KWZ/1R1CLVZcsNVBM0RTvlcj2q9OZExWc8IElDbPgzfcl9I2ZFZFoR4W2tnolwys1sOSo8Kri0N
LWXoMjwNqdVrr1H/mEHhEMqA9H/9hKc3TvynNWpVYdqHED79RLZM1e/an3MoTXe75YmvAQOdkQfZ
whRsmDz2JIas/JTmfzxnpgeknGVRiXZ8izMMmduXRLaK1ZvV9j/fn7b2Wd6U7lRWqB4XvQDWqxqX
4Vqien6kA7qQ9FOOeSlTmDeoJgctB+bqY3vhxEfp4FfZORNflTzjbgWgP5oHh8cRcSVB02FMSFee
m4EpUYrJqXBxDb7NNn9ebiI8E293AUq69Xd2GGrppPuuwSTnsS2kYejjYUA1zTofKtaJzKmeDDOb
nyePFpkaowFUDZlD575lyUWzsX11iKHEbce/WIMO2gyS95dBPFxdY+vDWt1o5EFg2KSPwMozsGit
Kx4I3u6UwfJsoMFBuyoROJqbxS5TZxBPT8k2b77BOG8rff88isGl6TjF/D65q59vsVGFPMUyjzex
3f3RFduDYQ1WH0zjDvvpWOZ0XEm/MpgPGyxy2etukvnKdUzLgv6tKlv032HXzg8LrRwYTCUwcbzw
+C+V9jYC20KsdUcdy/xyfxRbayKvXvorng7+t5FEFHdIh5u8f/oUr9IXF76z8R/ZadhZs+RnVZkR
7s5WZbOL+anqTZbWP57kSaXaNYTxtJ97Aq1a/t2E6+50XuPJCq5obEyOpYJL8vIVdoS2gL6BpKQT
g5QhtiJ0tqfqiwMJe0obl5NbvuE4GviLGbDRSRwBmsn9MwfitDHxbnjAVtdBVxvi9EJNwOdntodQ
/JrQg+7/5wzFLBPbADYKaUHrh+kcFCZBZYS32/oTFAodpjVRCFopzD8WxfBc7cFc5bX5nqazwgi0
iCUTUE0GJDHOaHPhBZCL5W0q2s2fdAUfjZDGOlEBGZptUvDcAYxHpwzsF8mRjU6wZhpRYtxKMAeC
jeMJVzNnbDm0RTgVbATQbE3kJPBlt3cEggGmmaecbXF2tQuOnaQCFLEQuD+X2UP7/zRUwr3e8/hb
rilf/+IUpI2qZjvnHPpVbm80j+XVRLVyH/cxi9YNQ4VXGOHg3Qbm/gEgSgNQgYYov5vVhe/A9g8P
ZOWUZpvBKMHoZHJ4C12+WjtXk+VJTrNrvZ4n8aMtQKzqLU7ze8J4nW3bcwJM5kHvqTrYXbi4djSN
phYYg5nS2XLcE/YC8WwtCFejZwNJkGCci0TiGI5aek+IstUF2G7l+bq3O+yrvv3stUL07cJOKcR8
8CLZNMkVyhLvg/gzTUG4sEQOrQFcZLI04FOgRsX6Kx8tw/zV7USZeV8TWfkTaasZtHPapmGBpCsH
ZAJRLT1s+n//PSnTy+fsAkmUYscfdJFUpYxFmQp7aNGg5yzSa/iSfjE73eOA7XRChqvXos1wHYaJ
FT6rnovvLn1/IkPqlbMBt3JfMJxApx2rGXWNGi8OHSJaHccpGgljZfNvAnD+LnBfJMGKcDoQ/+bM
gz6AHacOSr6pq0tXDuDUilMXwJiZmCgspGxfhCf2fJm2EDe2KZ5JFH9gPOQIMXOBhboCUQCKU0hk
HskVd71OElG4sMpgNFLwRKEP2KVYG5lLpPT89khfSbt00R8WsmlproQrgs1N/J9Ju/64AxMpaLpZ
vtUTbMPEmDjpWebK4+Ofq0H/SKrbHdPR4L5tLq3X7+U2DIlREKLj5NK9OBx5b2xEpqB5ASTwXfQL
TlYDcgba/CurAKR8sJprjyVkHcWkAtCw6uWbVc97ZF3/X2Bdo9u+mpHyfmUqjuV8DDaPxcb5yRWF
xY9LEXL9yY6D5u8jnOIMwJXRrMwed5ItVsVTupa6duGvPWGDUk5s1bgDRMrslJ8YWjVAOjIV7/xV
Q7p0Eyl9y9mULF3SA0l2FE2QvMR9gnc3koGYrOxlt13zTyIZMJ6lpJPe5WibF55Nmxqq4yum4OuR
wXf1uqYRgAFNIng/WEfTT9yJ3EtxMd33uZqn44CI3YM0uUJIIWO2wk+zdolMCR/U3I6fxjIlRQGv
8fvXPzOfLOc3rdJyJM4w5azBDZUosJ41nzdYKaWPLzHI7uwwcyihJrJA8zUmcNGL8TA8TwqdY6s/
/ggmx/o8Qj5VnjmyrkveSqMOxqSxD5OhHxFKBhDMqgW1N6cWDHgT0+10dB6kQ49OgGk3eSJrJvSS
lHosqvUAQ+BCMMhkPAGDtD+hEl4UOo6L2nn6J0QoRnuXcyuccvXOpEg125ufiyO8k3rJy6aDUfNG
sU6OfZZP/KKazFr+ImJyR1lVajwlr8mbx2JcL4i7OwJVib1kxf2DDNm3RLBH+lEvJ25DpYyCfy0T
0E64uX+YyKgyhMoD7rvUVrq92+9e9PzQGhLGuSP5nHuc186IR0yVFfKElUg9dbfZDzH2UqzZ6I1x
MDpGniGnN5uiKZYO0hLdxgYrsdvFyMvUWh7n9Q54Yra8eS1OFBZIxlpSUF57SK2vlYtBmh40/7NW
qX8WZs4HoxHJzLFDQr4r9Jx/5/kso6gCB36S8YAWMJATNqxZlQCSrbHiQgQ8PQh+H2w+HB1MEhLs
L+E13F05oQDPL38Vuw9UKU+lbZ/mKUVi5m+QCXQy6+DdJHs2p6zfKj/vUlpuOjMF4l4LCIuxXMFi
npj3iwnrD02JA1ZeFK/3Bu3bsWz5M2T9PT1gW6xjzSwf67+yu18x36nNYUPCeX6WSX9odB/RWxqp
0lgol7xRnekqhpNs0/G/igSc9BPgH5sNGZ2wk+0BvKxbDzzU2n+tubi5cV/3cyqoWWqU4yrSkJkG
fvgyb24uSk+/LZYXNkvJ4lRdMtU8chZsVRboRRx9wOzzaWhfAQLCz+6r/HMp2ef1MKLrbAlKZ+CL
A9Tsdg1HdlSx5VTKPIBoFlz21XbpKYtnZggi+DJH/jjJ8NQUIq9IdsM2fuBOuqGH17M36BZvJD7t
iMuE8Oe3WpHXtPW4hdtjORaDQ/BEy0/Dwm8YQ4jYKAYes2iH2x2SVlX17noorii8GMReBbfYX48S
mLQqlmgmXk1g1smct4h1Xzh1kCpVyDqeHXORO95S1Z1kaTB6GKauPdcTVvHxjRbBus+WN9FKdl+D
s8fwyUWCdc+dMrwNkCCM6nmXkQ3aMUJWdDErtkUaY8GCXWDbbRik9Hf+0N7PLCCfHwXo8OTg0zOd
MX8RBLr+VUkp2/xGW67mToozsnpR0lnqRztycCdZQsqKofzSAOSaPkpG+mvzcc2oDXL1uRkfOisi
cjjbzD7p5DTc355y/dqW4GfDr2AM4nnfCyIHgQMQK6xbfgEbWoEOVQAoP4647TzQOeBVUvoFqq+I
vhHrt4AosCkRCBh9CmgPHXSe1j5IXyqY1neUpBD/Ub90ss6Zmtfg7LZxcKG0Bo4GHqd9waQgkGD3
a0RRNAI14xq0Vs2JKXoBAW3Io5Ixn5C2suumt/XRU+qtlZ744WCxM/o2c2plPuPxJN0Myq5MWaU2
KiQwfCbAaw5e0KDUlC3YBYz+3AVq87kdTsC1kf+xa94+g6eqXbyxs0EX4XH0qSdsF2YEewYFCnFO
ofhs5mu2IFqOkMmjeD0sBPPkoYWaCmXP+ufEUFE2H1VamiX30+DOfH/KXBoPwxqE56fMxm/jG1GI
dE5GguZpmMl7H6bUGGFQSjGQzRI8Fxc8KrqU1LFJIpDeiN+/bIPhTA21nRobXAvZuqbe96dpliRc
rKQzRhJq5HUrAZfp33LBr/5Ls5kFzq+YAy+gGs+bq1x8hjvAoTqBVVB19cwPHK5YJWQIINhTNfSF
E+82i6DJ6FJaErEI99q/yvn5ERvuM6Ws9ffSRZ1sOsmcjmI8qh/ZNy9hmyGLgx8ooQ1y38GAsWEL
ZXfhvn4xF2EH6/yT+lrC+9Mp2ZLyERbPCR060JvcSNrYSDEtWJhV79iJF3KV8AA2ZsMYqkOjCLHm
selP8MRbkNa+yLCqEPkJ7bYKu49yb1V1n8/kBWKWhd6mGdfoU1wVzRux3/VOOG0NgbfEd42rIblm
KQorffk/ovlv0x+phaL7+fJ3Et/eAOEQECSwI/OK4BuE6ahoFVCb05N/xIw599sSlsf48q3uN8R9
uiI8TiKgY93jYn6VN6gKWLW230suKxS82a43qOpXuKVsJabyOyI+512j7kPVfg6ikfWw5QD1c2L+
BwBIRVBlgFePlAx1IUmwqGVoPgb6duxQmmLWPk7hfnmix1+HRzzf+fgotoi7ayegN9xJFt7aBqkn
9EOvdEOK8eXN83cKP0lz9torigksaBdxbJq2TcUchX5VMVmlmymhEG0oVEEObY2TDME2tZ6ORWpu
QisT6D3eEvT2e1+2JQjrr4hwVf7tt/LrU4yvgEJdnmV1R7tFQsjAmRPGPUlw4+selG8TKoKtuidY
DfrOiqSaWr7Ln9WbalQ2N2VeJ9rYjO41sQzST5KVuDnCURjO2+yFbSjDV3ff0eWxjygejsXAsM0i
TyIa/YbUOvfhCdsKAgGst4jPlEVyYtH/oUo6Ey1Lj9WW/SqB3ERjfg9a7IaG2cQwVGNWvAwLEdL9
cVpXUj05pXktjBiKbljYJZV0j3uRJmCALoWgcT4ARgS/rk7+sD1W3QNS9Cv5I1OFcmLdJev1rhwF
+PD9ZFk2whgHmTCJBHCrBXo42bZkwnsXWlqiJhdrWsOXoj5y6+pt+Rn0eiN+pkCiQjMg6J2DFHBg
vGRpQFIoqiHxN4qGX7KkbGEOkobdZEGJCRBF1+MS3XH8L/jXWFy3UiVMlrZPsC8TKM1n4GSs/Djp
aNaRqqFr1x7ldccPcLfTxG5bXikSrazkU8cBfGD56HyWFNgLUjgjZb3n8pn2Pv2WpGJDYYs6mYsY
81wReCwfv2hgTvHjHZjfq08v6dYJTSR+8xKrDCUn9nByFR6PaBWZJxm3pvBT3IlWACBq3SvVjOuG
kk8XQ1lyjUIncTI9LQQtpwoWojXTU2+19EMULg/1lM0S+7DyAlDy72aagXJ62snCelYOIVyXwG3c
xcwwIpFq4gpXsSuLALtxvHQ/arOUcC7kvCctCGTJ2jEWHXd+7TC6wkgC1TfoqUenqXyR99a3SlOJ
s8igKMLkVNB7fS1TuEAnmX9iF5XpmkcwnKxT5OyyIrpoqS7yHbtQNSgRYyA/tJvkvKEViaIb9JgC
PHFTAqXfhqR4jzfltAoiD7nTrNeTDvq+5ZYzKuNoFHs++GInqXaPKCLMyJFxo0UwPy23QxHybJTo
r3G7px2H78dzMwrLMvtckB945/MjnO+7QD2galRaTII8uFzYahYz8tkgRvpS+nIwrDlVuEMeuVby
0eT5WknZOmZz8WJ4ccSlVo0sz3Tw8aYW0uPwVtE0m5zTCnnVBVrhY1MTLArfjpmnuo6C0n2+1+Zo
rZNa/585qR4OnMzM6mgXEtajP9luuykLrQy7VIkIR7bu6KNkcr2Y6i5zYjmqg60mge83ixfrfs2c
HlbC0tVdNp5W/H0/EbuYXWi3fiLgb9q5d/nyBhU6o5PBzTeNI2bHujNEN0dXiUViYGffRGzPQYzS
bn5sqFPDXsE2+srN/mYUzlPMH8cY4zORyXMgRjepVJ3BhUc8l3PT0mFqTvuTELLBLkm7TC8hvOMT
wzOhTIpgr0nFWyMwnwXYG0gkkJygiAIei97vNEcGL+VlfyxAbSqqsqmwSvkCRhZHYZTKz1kozwQB
IZrZxlc6+/8h1tMigX2bpvz7Wte9VBRH9FQOkLtUU6LmJ9CGoB/cFxd3U//Z4JxSRJg/LswHinkj
aFLecsmf5fXREooXh4ePtKZhqkQJSzQi9qUE6pwj9zAtj4gkRZXsBJS6Gm1ZRgXfGmWeGEjqfGzP
ZL2KjIkXJSZHtM2Pwofqi+i0pUgnjhqGOyKyq1kd4F6IjwtYqNZAiQxJ0jsrLPbLwpaSvu2aQB0a
gMcPFtNB3kZpqB6rwbSioN24FJd4udtnZvMZAMvPysSwwZTdZJQBinGFCaRtW450HFy9rIFWPRfH
x1cz/gGwfxHIx1gSq/dc4PU2C7K8AKLV3M6MEl1VfZkYLzJjdzt5sQX4WEHYgwrw/+rkg0rKtSwj
TU3YpbPmqk+Yc2AsAmE39URW9DpO+dBTQQ8U1hLWkFgSYpHW4IHCvY29xVG01yL3AsFn1poyfcT/
xnkY5Nd8AIgUGiKikFDy+06MrIGnkDBUum+nFXd6cXaAjHiN6xZPB5GgveIG6yXcR2CobqjcNTXc
ZcqPVXjbjL5tfdWxFOxjq5cceLTa3orYac94B5R6psilpfwxOm3vrYUV9NMF2APulAsFhH+Ls8Yp
sGA9an3c6NA9Y0hBs+q/PSOqsoUlCT9JgIZZO+yBz5FV5EQBzviM6sR+gDnRQfm/4yB4DXrqAwQe
LDLfcLv1c+GALyQQWND/6tFBioRqfiYTBdpLDdhhum7YCy677aXGoooE1E7eM2W6bp5tADWuShqZ
qUeWh3Eb0iWIXlD+wMmLspZ4q9BbzbIsA9kztT922gEjeXLsDYZVrleQxgjgxVfyxTdDqnBrGkg0
ykAbILMRKcx9dQmhy1UZtTZs6hFvQNTsSwx/gcXuojk6KWKtmhSkQqWUxbNG/lRDwt6lDAfMPZMe
92IB1voPud6XP/Em/nt5N5bGtb8iGhpOmvV4v9SmfFm6TKFOHitQlWZLB4Sm+v1lWR0eKdEnuJFG
PEZesAaXxUI18VoJH1yeDKTXVbz/nC194uTElvieNnmCMT/EXMfKSz/8ymudk3YlWiS7gWMd97gj
X/IoKemMXa9niubocFzzKeZmr81eKB67lWpD8RrP/lO9DmZsmQv1ns1kL5SdmCNfzRamvBWKQtwc
5iHNAErNQSpbNA6RkZXch3dEx0lgSRBRMl8NPBaSkhV0vV2qkY1tgbkfqfLwd38C++gvBCrFahLf
CmB99UrwhkiCbG/ZIKAeCjqDCTekyI+NFvq7mBbnmPy+0CPHH6Hl2CQD/w3hww40WVW9hsAE1rj1
ST7IW2jR8FIDC4JdzjeURjn9xuVHA7KukTu/eEIkvmfOM/ksqo3i2u3wNCJ/Nq1iCwWotiE/BvdY
QlTXjqKnmf0gWQb5BwAMUR149Z0sVe8TzywyF1IIreM9d/OOQOLeGenSSpIX1ebR6MjFpaGq3NNT
KH6x203alcv3yOZkuO32qGhC76hSGg/N9CSAEFFkOp/NAWs2eBibYSyublEEpQRQGPrPGz2uYnGL
PXHWSOHI63VCdjwh2IJsgBYJFQOshorRtcLx9O2/RIUfHcuaHHAmyW89tmSDF9z4NBfpNpPERnN5
NUjNMdAWqxS5TnHwMDiPLJJ9fJh+2pTWOve4FJPqfHvVouybj7YSdSP/lpRWabSGloEVxpd2kyLv
BqGxBfYtCMEINsUd7sjXeS1HV+Z+yp3IFUVW/15JVWhDYAcPxUg8ni0q7WxoR7j/vfa5MPFxwOOP
I+Ccm28cdw2uxBQb7dRHeel7GcyrDcyBAZ/kHOj3BrBo4hnWjyFBe61rPI37el3MFsJET4ROZ1Jj
V2roN7C4vHq0ChYiuM+3qc6Ddk3lI7UmBgx5DZE/3h+V5J236E/X620gXWe9gk4/ShvOkMSFtj+5
TqEoVsWo7thSiKjdg1vr1CdqCwfOWXkJ5NwtCpi6Tm7UjgvC80OdTQ9JmAKex0UuPhDgsVs3AsHr
Bb4K9PV1KGC27o0/a6vHzTV7ok/ENJmxK6sCp/FWBIaq36VRyF6rGZ5SpW9QAYEILzMBwxTuL1ka
Cbw8ACod4v2t5YswnKQwbT38kvg6vJNHG+FgZ+GElz2j/SDdb14F0od/Enpu8k2v3uHKT2ZfCPKu
l1nOnDC4+aZzGk9uQSvpwRp4GxlkCrUzPyuC1F6dg4fwp65shdOMemi3Qs6Pc0WyVhpTxERk61jd
dJ6fFQApNNuJT9QNM9COJEfJRLIAXcoUqecBbDLtJJLLxg4oNbQTIEv7j07CVQqqOlDWJJE2mT/V
Ln8yXjcUInX5OsPQrIrDn5tznRuKGHARuFtpGGbVedRd3X/Ou9bS7Ql0hYEIdpiTL13LM8kwxpI2
vKwqypx/iWLzayF4T4tyNe7d+p7/rs6YKjtDlR2rbivbJM+SkFE/IYIStL552S9wxNKbO5BcXyNw
w6zpbGZfWbiOO9sIYwgKHcNUam1E1fHj62RvBXkRjhuu4vOPytmKSGmgQsobFJfqVsaohO7VfXfi
rkPjXheEACzVcWnIaeUNcqH/a5PKjLRoGBn0ZZOdf+ZxK6Q7SY39YTaPSQV/Epuv8UQenXZVER7X
gHgiyHgWOpPiBIzyxMoW02rnjblzmJpVnBqPonaLwH4EfVK/lSc91eEBCTlGGU/DTBgSXKjebNY2
bdr3LL/3eHz7HfyMqpuXSBvFjEh23XimMd4c5v8aJb2BAF5lHZ0/hE2cRwlWA/NWIaHousPz+hbf
NC40H7+uHJwFi14oCW6M4uxRB6+3Ppav0GM2YtbI2VLwxlkgRXRY3M7/C3kUZ3dlIYxXCuhHgWYl
e3gno8Cm0ShG7sxsFJsxpE6B/8DSp1iODuOonhMORvNWkJT5HqkhaYqMrFyBk2s/SriTEdi80YfK
O7RiWsLacTA4EYhvBxgfbRJaRqqx6ZO0s3k5g2DUHsp2Htcz4WLGb60vkyDrXF0TogkCpTFdGDPT
MGKQsB5Hc1vOSvLngCpQChh7De7QwS85B5syotdgqfY8W6ma4cbnRqBXHTTGoa3EmOSasZxO+ASx
tiVwhkPeH38ccBZhvSkFLDAVOZU/iMjpNVh0O5z8kNklstzfJiq653lcBFNNhgALZe2IsbEDgJ1w
WLWOFhr9aJfk0eBO0TJSzOk0j0hmfDKilS+3U5irGIpWZNNZbQ1usfgJx9kIwEKtgTlXhz946viA
NYix2TdHQC9RtDr6NKTyFCxV9K4699YfTppqZvP9ymIE8r1HsD5HhHMW6qJEmecqieiG8HfV+o8g
4OA6NutKZl2Z1VWiHjRFgXsQp+CJI5KyjN8ksQ7MBo0cNb5r7LP+4QSKb/5kH9ZxKpeDolmn8bG3
wEczxUpwWnf1d+8TFF8qS7OkOj2ypBGzF0cacxTvvIdil7E22uC1Phn77Xu+pDQ/7+TCy7518flg
cwgfqj7ZrfmSERL0aacXJV9oRGbpC3VkolNe16xig43HvDFc4kR8U8DWImGw/Cko0nN1R3WaWPM6
VG8dvs9Ip9cfXm4rLhO3t7jG2kBYknhv+C5UrfpdCgBFwoOCBtU9xuDiuXiIr9BVIyKob97foDps
ZAdIehuv9BjBjQMeKLWtgc8ouXvEitiPCRJE88i9vG9Q5mYlg6/RSlklxEgWmVUAYAtT4qsqaFr7
m478nPSy5R/c+gCGdx7+Q0iYmCD5LcMn66MMCIlhFrsu+u1OwETuaeufHhjIxD/Sw34fpGETPt4O
cEdQHEbcB2vQAi8JFOYQOSST0+0d+fGKd1n7ME2dzEkVbCNP3t+hH1vAS6GexIliGvVe6M9nxIRg
8arHank8GMOPulB8gAiJKgQ30zcoeDxVlHStQWK10BNxPARv820ruum1lEDallzIpgxT5lBz6zfv
UPLwp4INCSdo5OuEDUIaU48iO3WzVfN42uE9G/6IR0Ez8W0vCDyTaEOVV3GJW43mcSD71sJAjohY
V2Qn1ehEoKPGfhhiQJQrlM+UaTIHNNk4/g/woE3r8TXVlO8riwuAfHLXz3zlktQcXzrE6dZO7rky
AH9or5m6HbB2EgwqnRg37qLyQ2b0xB/lMFGPMFp4tc2c4yyq18eE/w1MHfm+eHGdkhmLz2Y0CZ5b
ums7hqllzflBSWJjePfY0JpaNA+ngh8FWM49J+B7XJvfUG2NTIpBz+Yk8CNb7W/2ZyCs/qNtQzNx
dqpeleZF1djr/YseIVT32tav4cakSpipPPgSFz2WBp9tq7xXHArZK5bscA0OUF0Y7JBIYgpbbs/D
w1ccNmI224TgDXoXxn8L2SFMeml1EEHPN0VFu1KS20l0ptjPK9WtkHSvetGDN/EiKFJNpAxiPRrP
WDo3tY7w
`pragma protect end_protected
