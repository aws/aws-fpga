`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect begin_commonblock
`pragma protect control error_handling="delegated"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa", key_block
XSsTGNGtJgHES/2ibVRfmOC+TJ+NcI66C8EXdFNnkLq8ZaEZcS6wTOi2OVHij0a3Jfd7QEG9C7Ww
7LHpCKpPB+lzQix2DX9JGwYtipFQEwnzwS4R52NMpHYmtOm+DHcgSPq/CBa6hXg9zVVQNHzCN4bA
ll3GciYcI6Fg0q4L5j0q6DNEshte6jVwIUgfv8JfcHOY7IBrLyWL0elYND/SFVToydoLLRMZvhDL
96QCXrGdM6VNguTWzF7eGZiGQ9m71TPxlLFW1id6pZ/HilvHm2n7zCZ4cZNQ6a5zW8eiaTnb86W7
1dRD4DatNRzQ1bmBU/vZpyKtPw9QK2J/sHo88g==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect end_toolblock="TLJlajGRGtfqxVHY7I18YjQo3AgqA2+MGrE5L46wXLw="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 22560)
`pragma protect data_block
Zfg/kKeVj1J7Dp9TMQbfz6dnkuDLWmqPPdGRTILGxxD7+Qnc1L85NEo4x9N7lPYdxFsMJ36LnOAN
uCf5KjSQ1MO6aS01j+9m1ZyXj/Z55tOcdiRfJOL3Woyt5jgTpujwxLsMJ00eWAs9RWCrpLzoZTBj
M9vedDxy11H24N9XHPwL5Q0PsOmdJb5djscBv+QN1EBdHLXhVWNIXDuQeXaS+P/67rzBmCFolUVT
ou5fivg3LaE18rlS4JEp1G6MKIFEIBpNyYj9kGt8zR2BEK4WvTxLioSzdo46ZwHP5f6s5Ck4lqFk
YvOlRDuvDdOKnJBfgxR+P1rY2yBS9xgtj7dteCNjHj6d60j+ivHMGL/C8MuC8q8QQ2pI4r3jVJdG
T1th+QUyiSvPoctw//brAIV08wwwQlAwahglN6/3rRQ6GSEdo29YVoYipeAICSnqQaEz7qtObMpf
RxA6/9iV5yHxly7rMMosgjEiMK4EJPz+cEqsyj7rKlno94I26cP/EkxCVixXMUz67dflnSXvgyEH
6HRUXdRpLtACZ3fEiO1DSOsdDtn4bwRz0TlX69l1W0h2VTex4qXRI8miWUzjWOSRExypN5sDDuxn
on4MTM4l6MiK/D8wdt2qm9ph5tucslUZqQVHS0kf2wyAdj011YOwDyHQx8uaZNpMmfp7xPqBx7U4
R8MICzPOZK3tZfQcFFLQoIVoHGTN6I1ere7RiqN+fXlmp/pMDrtyM39e639jhw/RxCfOU7moPc9d
qT/e514J23gNZhvhP8i3+4XJSZS8DCDfetp38KA9dQX3DrxXQaT3lM66vn3n5CwOBtB83Htvc3Rd
yIHFrv20A+Op30vc21S+3GKOb25PgU55jhacg+kESh/frsXtHPvJZzBSmgjAB+wQv4e1tIDBbrbc
J3dzA5aA4aH0EGVJUHqEguNS9D42se/qkdwdP9A4kV+x4SG4mraMlqU4JXB6P/lcnwHPF+x++yi/
SzD92cMhmVx6ktk8Wb9CVFP7fhs4IUMODskZCKjkSO0lWkwWvd+Hw1TIjSoaTlqIE+fg4qDUkF09
Fo0OguXa3BrPOKYd4BzFa37ZYMop8vsGqDhoFKDZ4a/Q1ejQLX5Ldl2dCugcSkndQ+lkCwd64GkH
BZHKuS686h4TIkHiNeacEgnAaVv2hYqn09/gG9QhX65h9mZ8mLx2K+DhKlKq+2wJKOZkA7J+yoSv
yP8F4+pCD9anCxUJLFIB9hFkf/OsU6fNqBRFDDCWJ/wTC1Zh1VJUMmiA1Yf2+T+wPk8PceyoJdMi
nmygaq7RTdEfMKSooC/IKcGuPqlV6jFXt5xRUpNJHpHfmsTcF5Acl/dCz8ykwTEabv2xErc+ytZz
DqkFnSpxqf9/5itBVXFaxGPzYT+1XJ3P1c1b99xIET14wsmDMwVRDytgclOacaxtf18JSTV3P91t
MU3jE8j+wpsnRnLwHpVVuTcnpwHPtrVmmxAAWHhwNRsuaV+lWd2H441lUDLM8uu8Cf8cw+i+aoTF
EXgiY8QQ1gJ1zCa3F3BRFdn7/yBe2oVcgDdE9N/n+SdiCaHam1WMEjKAG2ZseKT7A4Uw6XbpA0FG
znEycCcAkbZZyX7Smx8cDx4+2G9UL9BL0T++eewfBqWox8HQsL0wJKBLObQCgjM2nvdVpF3vtBoS
/NnEH7AyJfQwBp8TR2F8I4BmCVLy8mBhGwWByurHSAq4Y8Kmpk3J3K8a/AnhNQS0mbayUj7aSDcV
8jauRnFhtXiwiZYYYQW5t1/senb9wilAw7sMphgK3bG8r8E/otRYRkRi8MyIvZ//yvph8rEBC9sw
GE2tKp5BECGCJUGaQeJfPLfzAyCG46gPxroO+tK+uPBO63XEBQeMsF8znm9cPSh0H4RDF3aRYqbp
KvAmbSIzW2pqqPv9lvM8Ldtk7rkpSixpbeRM07/blQBHNA7vBIpIN1dRjxlUuSrQowZcdXEwtqAj
Lw5x3yL+Kf2OKFrDHj9W83kcFywrTPzcYhq5E7uAAfOpp6VxBkcrGEYz1Aqg0Zo6wLoqbx5LL0Ny
3W5w3BbhQMFfCJr4Dp15chR3Nzp4GA8IXBjktieO/P3imQfk/7EAgdsxyRPpVzWDTX3qkW62d7sY
yCg9zfcf1l4Z51L14WaQ4KIXp4d5TQKO9nIz6P+4MYlmJuCD4oLQS32KcF/Wwm8SskwZWK2fB9T1
vNxCUHwfoTlchJVj6HfCadm50fGieurlLMS6u0V4RpbjjgZYG3A0uqhd70+5iQEoSTcRYAyMmr3f
xONmFsEUxZuFxJ4rH1GR4waCgnSSVPah0QpA0LJ8jc7i4dRVgHxnJ4HUioAuV1fw+GkhEXBtVZah
Qycr4LKbVwVBjSNN5okqbsQbZUxQJlETgDMZIIWQuwpnjnZW7VGPN5ML46yT8uha6zl9Apeap+Yp
zCkfshhKEOH9h5f5Bf6S4gvQu64zpYUeiPyVVvoKWKUZciu7oo1n8kUtxye0UWYAk3PByyvTGiD+
UP2aYyG1sO5hjvkyooGTu78z0OOJQeu2nSWtl3sC++HNyKkmnoHbGqzjEeTsvd1oIk/zzsAkF85d
zfljNRkjQOJMZ/BtUt0a3/hV27oWQzpwJdBC0MkfybCIrrjYYQU7BvqBd6eFjYDtEvq4ZrrLIbQN
nS05ga/4CuoiVpsEVIK7S3Vvdcrshbx1lKgqcOVe+9S874A22yle60wam+tPqOamD6cr8gZBaLiv
DdicIcdEYQSsSVZk1j7gEDyssYCdsrlAAD8HUzG1BWz7eQngOApD5/manY4+VbxnFoaVEHzECb3e
GtH6+s/Wy1nfbKOx8tXch2UUBDXFlCglUgJIrScwlcNxvUgyw0T9+woVlAzY531Mf8x3QgQtN07A
OPqUoVGSGPsXfrFgLmy6cIDGKjv0MT7OvIDsosGH0AR4MnrRMgnOzn9ns5MzrBerCDpR0JXu/cmK
bR7Db4G7OBa5vW26Vgt6kMwdFD9OGrLdUeJqukvOnA71ZJESZEAPJdSO/cUyMm7OychzO63QSHXJ
fEJMCE3q4Msi5BOOR75BPQj0ZvClcTphJhLD9PF7/lss/wmECwkRaGA01PyFzVIEtWlyUZ2pLuC0
eyhUA/t1QlQDuRZBvHNqTgCnNBV03byvB0k+HEH99IkecI8uiNmLOXnjeAdg3eKYUSTm2aTdc9hB
30Spi+0JQcLJrHAVUuRfwLXsn3/+QSGOVLzk+1xFTWlA6CqOh6HCUD+u4bUaHPa99yKzx5jr/dGc
avoj8LUJiCfZMFuCOgSeINboEQusOt80mPvMxfonMsMle3ZdFeNBPFOBM8AuNhOhf6091MgmzUtx
l16wEhn71Y/+UwzKFBWtczS7e/1qPnGuEsXa6DgixLtOJXKV7mPi9lIyWMQoDZN1mL/PC4BfBMn8
cPtw4hHffyVKvELZhQ/JqVgOoHMZITuwZFSur02186qEXu2Y6udt/O6ceqmr3vC6dW2JoeJJ64Xi
szxvhRfOYZJ7QBXk+vWNHJ7FfKA4cwEI44lOnGz4hDenzPoNio16cc20YHJSQnX4hFa3Pb12KSva
fZPVLwR/KFjx7vRvHLyl2204X3QN6MkNCPqTEDQOPkGXzgUCdqUmv7ld7/53VynNa+Sh06aRe6Tw
bGsBgaMeu+p1XQr1oy5/uCvmUZTG7mzgzLTMrjSKdDV7ENpZmTPna5Y1iq9NKYZoleJAxLup+G4w
4Ss3di5d3WVJ9m5MSLerog6NdkWAMBnS9EZcCHhGAn4VvyrlLgXlvfIDeGqt8485oSfZrEp93kdT
WX8eH1H2D6UWUu/MNkw3scaVIHKtLzkGY1Uqq+LaDO0fm1257RehbDAJzkqGooCYCgZoSQ6YpWBa
KT3PCzhS/Nqrr9rHCM4g1rIkrqq0tL2Nco4FhTj2RMSm2KVK8WBRnnmUPUPIdrO6hBY44LOSrBAL
hFTMtrrdSbZJ5NneVKNoh1VN1eJ1K9WaTZsEA9RG6HMXNVbIQ8rrYVep0SBJHYHwlnCATVkvDlLC
fdLLpsZuxhYviezoAiy2QXI2mX0LPcJSyD7ND3jrSiDIa/h1nYm3sTuN63n9LXbaZeOXY9CeYEJm
kM7z2W9HArYaNc66Dj+aO0aN1wLGxz6LsHcMwYf+A+TpdfckB1VAkM5mMxa94q/u2qtO48TWwhJa
xlsrF6Tg5uqp8mqEo2nANw1l88e6knLDEvwHPydDO5wkAqOJOHvIxxQeQUEdLWy8UwHeiapJmch2
MPzeO2zgPnTKajlNT05F6E5NcPGOW1gzcjqCXLvZXU3seWKww5FJApsVSlQK7JXjHtT/l5bqNSJp
sRr3M2k/sjN+HjEflcevDklMwbUsbpVa0/GPX1a50iSjskhKMu/lBxDOWt4Sh4T5YFpg1BX0SdXx
58zNIvzsQbK9cQNM3clCxfyyf8GGhE7+5BGS3N7l0nkzshmBUTdqw1GEi1abwqklUd0j0sa567iL
s/5ZOPpbl5LHLO8Deggeyh8KhuZtYicLTW5FNyGgYJUbI7GvX234dSIw4WVoPNT5gRMFZ9rdHH4c
8B3nUVWC2Q5ty1pno3UIi0rJmdE8aHZvkiO/vhpTQRrX1ubVxdjFcIGTgQNWtffahxSGjaLDQwkW
DZ1oDeY2UaTVfxcv6SWJBtldKiofd7ZaG6YTE9YevulXOkGPe4JgC6kSkjaXyqUB9qGJZ2I02z5T
5D4Nak2dOF0cLB4pZa3dMYkAgANBAYurhT1W7uDB7XtSPcjaGMO0zOCs1Noh5UkkbMY/H+qweRUD
6yBu7BX/Y7T7z7rWi11GoBoeadNjw0DBsTtAznfO4Afh3bw5kviF8OGg1AjkHcM3atwJhzOeap6j
37/eWHopJz2mQ1g/J9LLf4656u17b47vUrzeQ7+etsEVmxwPsPu8FFFuh4itDzDGSXYoQ40JowVk
dfS2oFhkfw6HAIUGqRVgVz9eJObnxL6sXoWiwlTuJBpZvzakitMrQsiFGOO5iEQlPMc00t2m+/qA
hOqkdVePdNOUZ5wbZhHu8q+d+8Vh8Isu9417Z3Tbv/stCFl40uYAWiWlf29Apattoylid8IumDPm
HMSlUI7nr4NDgVoj9zRPXwiXnDlyEBEo9Rd4ckkBMLhHyq7kKSdFlKgLt2TmFtYaEN7HiYvbQuye
FcyXrE8I4mv1YQVAFN+nhErv03nhxL0HYRusBR6ZYPBPkYVqH85ZtZWmb81FudVL1B085wllRemc
sTZcsnIztxgi16+B3/onXPVD1Y7iHCWsiHv8T/WfNAIJziaaStpUqLy9dTxWmYKNbD+rTAFPIK3p
mDobqo1x5vJM1/JEsFTn0GmnIDqhJEipj4KWgHaLczNjqF3v9SF7PmU3GNcQqGmXNAlH4biAa68M
nYqF37QdlxgSSrDRL+UyGRPf4tMxSw9euhv28DKBkBMmTp7p4YMz/E3IeIZ9FpZ2ypfkt0IPTYf/
R3NXHJhawicEVhPZzdxpyOyrg2qgyb9mzk0+VWHu1nj9VbRce5gRbaKqkUyCfZzX9GPvmW+U8dK5
Y3VEz+TgQAhxgUhpp5wZRwDO26Ou95zwz0sWUqlE+1r80sfZdhUyhRfKRfVCsS+l0hwk5LCAq9hf
87LzfHAubuwohHCTKLYxL2mL5cTyjHsCp7Fj+ByENGxokah5IDEUdX+JKFybmSUKi5wedwK2Y3Kb
p76ddMwmUTbU69CQrwknsTR//g8XOoKlvIRJFu6YCh4OE8NKw8qtkBz79L0JgBTqycfa+ThBgWPr
Db35LzAHy48rp57L/SplGtOFn3CZTTZtR/DHEjWAsnAkLoQb/t0ZnLxk+idSK3HsdXUu0kewVfdI
4mZ9m6gVpXmAj7ue4IQudRawUSfnomrUGjazEpfPz/re21DwPRi5mWkbnP9IvtmAD8lXpEdCsHVB
O1BuNXm7Q2UJy8a7lNsvGaP8dCq1hncD90t/ay3edJa4bCuesg0JqzMS4w8TNv6FzV3J857BTJ/h
vucKry3/Ro43X0piCBEKU5CTUi03EW29oAMzpv3yJeb6NyHTRg8B939hSTSdf1UmSLLDdtiVRlAD
89MtCF4Djyt854pzn8EgANHjfKaVrfL9nGArN1THL+2vNvMIod6J6uKfwi+wfBLA+cE385xmDg6o
5jR3qjDNSKCseOn8J56xGeQnz0XZHm70jyuEy0xXpmyRsjauLvQf48qmpafXPUXwlg9Yu3SwEVAK
Z/kqZ/lq9vzvJ3igrUrfUPxHFEz8Y03hTIqJGAlC93/t+v+x0bgUf8/8l9z3mZEB7SIQneyTg2JQ
L1y37LlGpA1qH/bWmB9Df/bCiJnKLXk/aUwU4jyW4Ha5k8SXKoHbAq8M5yPu91yyE2A89Fyh1qwz
fok0rA9mRfa06RGEisLLY7feNvkYutsIW3L1iNhsd/Ry9cmBNyfu1fY0D/flZG1VPLisAthIkFJQ
ti3hPpO1wPddIrR31E/yNGy6IQiIjqUULiR+e77l4gTgAcw9UCGSoHP30Hn/r7lxz+MxqhN9+yxL
YrqG/2HWWOrGFfCGGc2bYj34gb+79jb8483XsgYUC/cNk9iFM/Md+rdpZk6D0nCjyeTIRh92Il8J
COfxvTMiVWy/4wND5l1MrryT4DHODM4JSGLs3Kx1HxDFqaErnvlItD8UdnsDmATgWdehgzrougoC
ZlIxy2IlVO5gAJPwjDPf5RB5Hghk9U8ftQsl8yKwgqghvlxJJh5+LZDLzDJX0f/jaJt3oLgPcvf8
y4y/qGyT2gSY1/kY3nOK1KeXkGy+24i6Om/BP/QcE9YE7I+PHb45EUZVdQFXBy8EowshLCN/lXZ3
Lnd+ll2s7+gbYQIfYUNyM6qCYWIjdSg1TM2oSk84gzplrMgV/bb6VH49v9MDGCRHdqDbQmjUyBT0
CS/zYVAcRn6/TRrrTtAf0Lu3kqlxCm9M3IuaaKzoP5zf0QpaFaBa1EswjUJ849AGSb84XZxu0yeW
gQ9p7rqwxYjwGRuLXViJZXNyeY1AqxO1CM9BxwwHV5YtJax+Lpzw3H5/TUUd8Qy72R0kHX1ajHIQ
Ml4iBoO8b+3XggSOfVB0ZNxseJt+RxWrAgOzo647e8U7bkGFT+ERt4zlCFaV3U3ZwLE7tUJAtAE4
DL7SuQ81qp3DhgRUBe7wyGz0imBUTdfXdVy7UKWj4ipOsNMK/LUkxDbsS6hO3y3RPrC7GVcF9+aB
VHOMI6FP9ySkR0b+HhFNBGzIXrV2SYZYIQgBoN2pingnYFt8QnjgKsjO+f8kw689cBXa3q4GQCTK
0ksja9YVhFwN502tm1uGFRmNAeCqqyb8+g64XTw8Qu16tUsGn2ENqLN0Zw0dBJJTTrKD/qEBjag0
M8sXgfnGb6Kd3U4XSxLn5MDDAqBOQXzrZiYoMnHXqRScfrKm56gtHt8e6711hm9F2Y4TCluYJr8u
hbasgTb97ChJAt0VUr5XBICo3e/58ghUOLdCJqXUAeudt887p8dmtUxdSNFBA6tIbqF29J5A5tCt
VdafuHylfa0NvBei47/0E5PeXrs4QyzukeGEL6hiOzptYbMYba9OcE/NfMl+iFWVeYReBDf8bT1G
DNLjZZ73sMsT+YwyrP/1RkmCuvqC38gLDnFLeFLKvIVr45W/nb8HHkN4wYPYkDABIL0/f5oyVmGp
ELSnhyz4kkvaVL7enm6pP6Qc6J37SJ9hUV7wpe2CvwORL7uWJ0KQDiL+iyJqkh/fmhl3Re1DWzF2
KJ7LCAQ0ZFz3lMeeu0BNoxeTG+s9nLUwF/sySpZvf+nnA/bXqzEBlYSWRj0mdBaquVtqedq8QFFe
jPnKh/SgaIhIlB0XD4Xvj5RjLii+Q7BBwyafF813i0YDnb4Yej60v1dkYzB7WsiFnBxavE75rrdt
+1mfeugQ6MCs0wjlyq50Sa71fDT27OyoveudYGiY4Dux74TNN45+QQ7SYPi5XtJ6Y2b+A+52u1AK
0HtLlS2DGl145B8xNwC4NXq7BsS1N4XPeeRD6yRhx1wtFoWcwr6ccGmkhHyMkn6AInA88vn8BzNF
lim7flBewck67GlR+l5S8tUx71iczzv3ThQmL46f4CBfeI2caXZcbp7s0Mlxyd41O3lXI5ChIIqV
IhwFFJ0vRgHvgz1EsXKcE5ER3/QTHzJ17NHSKkAuNy8RYGv6ni1N9u4AnC4WnrC11U6R4VcMW6OL
pzlm1/YqnA+UduIMCZOJs4wxcaiQv7MQuGTQlh5+cQmZIreGpQSD3SC5WcmMTfuYnGtDcwuC2gpM
znNjUBRoiYQcZXcSyH7oY2OSXeMgrVmMHcD8Rm19gBgfULmG+XPUs1uOLpk+7+rviMZZkxX87bcx
ulI3ASPirhdSb7lzffhC5Q09Eg8QRrXuSJK8j8ZJxlUK7/t8S7xKUMLd1UZ77admoDmb2QsL4ZrU
36eeJzjPqvKSCp5EfkvtPv47ew89Fb707TTI51IZN7LhgiY1zVggy1uJUz+8dAKTfR4uINP9w4T8
W7+DhNNtAcd+ANM3LqckCMUzSjDk8xDspwzcBlK+neeg92jzCdNyoBrZ7lbi031axc3rUwmPlAj2
/HC54LrRuO1zi8Y5UFwW/03csirucWQeSpS6R4NH71FBnI+OxW1D3RHCKDxKMc4E1in5hKrx0aB0
5Qx0QKcLTHskrYWmboBVytS8QwCHTrlw3N7CgtGPgPeYGn82WC90MwmWliUl6Og59h58FdXvrdc+
AqxQJOW0qdZgU1PaCi0iT0xCGQNaDeY1TWFYPoxObB2OEiWR2MglNARp655Lqrp7sdhR8SDPkMFo
325OZZeEWkOBoSaggGnMzUeSDv/Cx46ATUXQzbIQdlUvBMjZQlyRmGJeqynx3V15KXU4uPfjSUnU
vc71YftzmP45o2U7Zq08cSNMNk5f3587V8pYedd4S/XYqWQEY0g2g47YaIgfT5k/SrJabO/ylJdw
mu2If24A0dztuCCZOBiZmofZCHOI5cjm7POalRwoQ96+TuiavwcWXfbR8pOPpaI9UN87wdvTaw1Z
6BJMWdt2lZrmviCcaG1Be8zoA8R1OP0RlDljFnSzoHjyGP+FMxu+yI8JJqJNbb8qOjqjbPEV/IK7
29S78Lr4X83FQ6h1fqmDRThgFV4zGcQMU4tces8Z0c/SlfIT0Qj8WrquUcVbEpvO/roJH5wRUurX
klsgmXO9TQ6GEJZNXaLGvfjOLn/zKjz8CGtxYN/JZtc18RD4pgGS4IOeT7glE39h95Kyu5oKHqv7
9I2TQs7AxgLLaSVLMi9kBmn0oSbUDtA4PjkKmcCLCkce+C2JNSdb3IoqJAk9ZUhhnl+uupKV3sPN
JSY+H8/pELA4OT17SLGkai53P8agXSxL49lvglml06UmU3Uj6TCxNr12+hoa5Ew4dkdEQpo70aae
9aDVbDqy1EQotxVq5j1qtT1iy+v0yJXkeNgmepJAi70Lm5/II6LLzYxKWo2rfKM7pFOK3vzqgD41
QWGuvzhKgkzYtYP72pbj490J4gxbwYLoCZ8O6mPnAh1NXnrmJrcBmTw7FFjd/FQ7sfDiBkOe9aEr
F5zz3ESo9YW+7WW/JvMmHu4KYUoF9njP+DUXqdxBJqm1UqOfvLCfHqqaHWBUv9rFX0IwVfGcx4nE
jgVE2zuNxTtLHnVnPXrsA9CMmmeo7UAUlWrpSKuwSm/SmPBpl3XHGM86AIjCy4hIYA6syxF6LeIq
w1njJ2Kzv6mgp1oamrjLsEq/i0aADnFaqXagc3BA2DwcIwCujjXv+X1lnH9w2u0A/aBht3oJPMxj
cBAiwhwLliDpAVxUzKyQfarjerImUvBZ2rK3gPmPBlj39q1dgTqjjOSFddhNWOCVfJ+Mxz5Jg+/s
eID7vICAqa42CHK1XN1rYAEjmyUZU6KNGZiGSZKVuqovyg2X4nIcpisF0SDoMjzL0LIUuCWI05tv
bgf9YteviPaRqasj/imf2gqnJim02Z8FwY1KZWqvf7NeeWuelUFifyKIr7UiboYiV8xYM/hoNC5u
OJ8BHFS1WhXLktUIi+kR4/sfJd5XMrHNFuPyPmya/WVY83p4VyyitgMCH+TTA1POh2TsY3TvTW/L
kPXbOU/MUu9r4tQBHTuxsQicI5VWaHoLrZEXGbGhAPOX/UxSz3n0kwvLqlkKu7RCpDdQLoTydbxo
lK4ej9H30b5BDk8MnEGO3FzeJTVyfBFm3j5m24Vl+b4X1eBTcX3FgSEFMwUBsFqDNhB/h1v728ZM
ZpbJpSyr6u9h9bm1O9CS0D7V7PZIy4q7rT48gN8p9rXRkMZrRJdZpXNnYzY3XeAQNXaJxnftJd0S
w0watLcLbcVQa5fjgPIUHdQRVQiQDgrLYVTo+eP1evrAVZ1pupcMPdJjLGUR1wOuVJtmWV1+hhIN
ogHwbWp4rzW4lTbNFcacTH40/3E5XHF/8BaRjX2ecY5GAmvxODArcZDmzQLFGxEzhR0kdQJJsvl0
RP7tgIOhHiAgG5nEeqorDdRWfJHptAS/+86aKu24v+ah9GgFh71AdlNJedd73ORy+nvrTKxUQzyH
DZbRLhIjcE+b1C1ZIOWsZ6Wg1eqHa9xBAoQRETCWEN1Wvmo/HNokQ01LuoHwN70ekMJcg6RWjmrk
mhzF5nBqsOEHZx7Vmtf8//M3cXQ/fI8jspt172tyYpCuhEbG0lwC209jNcyaVzkFLc3wGMYU+cus
h3ssSlr2DkTr8rttreUYAN3+aStZZP1kV9FqwjM/iQDN17TO/1tBwfz/xyOcbReZB3SK5dvdgll+
k4yEO2Zmq8pnsvu3agmY9vGXJtLMkFQu55vBwI1NvkEKULqfzePx67FZudt+e04gpLp/aF43DSuK
4KDB8teBQrjRk4fTAWBmkkJ5/FlC7QMuAVEHUINQVMEoJ4L9sv07jmgpZqhlGofXel0ENttDDR9F
bu7/AwHkenHv4OMDl4xTIgnRNbdLR9voXuF/O0nLBIA4NCcGA5Ywhq4LdJ9wZCatpj+NpWVwIDnF
uW/dxLjFnWRATskYYvZj4XrdKURG004vzjc6QZ0+yRexI7Xwxhq5hjfX+V0ZpQQ2OkDi3ixTqmxe
vOPccxWdp41yBWyL0lGn4RWygK4i53fwzEnu8tex8T7Y1V84smu14ic7+zSnrwb0pvWhwVn0qptO
ZrVVc9OGHN4YnXozBX/jLCKyFl1LKfagrI2zFyje+c+FzMTcqFp9XaEBYdk8KIyv25+8qwjjTJQl
d5FxsR1wQHKAtKQ3CBCztrTM/ZgFqiC0hlvFRVhrvhJiT1ghxXp6dfXCEeichZMNo3DL2i2l+n4D
QGQ088HJ7+YvMLtbmzFhk/UrY36dffAEWcDsowQC+D2kkGGjKq+SLq4Fku5IypvALEMjGoNsSx3U
MIFtjqqVzy1oyflma7JF2k6cmlNGpIwAQrMKrMwnkNXmIu8QtFxMMRItwyT806IEIPSts40GQ9Fj
TJMknqVOp/rfWIZJ3xbo6+fitcZQqEDpQZGMave7PrBYMVxdtNjtrY05wO8+G+mrAMny9wJj83RZ
PTE1SvUVKGsn/5VsHFXJstCJ5OzctgbFFZznhTN1RFbc5P1OQZsXGRjPHFGc8kcDmEAfX+hMqS6I
jBffWCSEEZbF+fISvOFmw64VgJKS5YqxmRo+vb0OPN/x07p+S2FAvq8ZxCaoKGvQHe/wSU5kaZuv
KdR8cAAl/rsHKJv+m61H2hiR5qlUEm6zPhSnX7a9JQSv9Ss6F3b7KT4dKigeIQLKDFPuztwpPGN2
hl3hZfdQqViXPBMWIUxo4DOpHKNJUT+0auc/HUCtz+9KqhFFz09kzZUz5A4MijOq1kKmFADNPEyi
ETaeWIwDLzegL1Io7rWKmV+kZIyQZGVr0ZWi+vum7ec/tdmomIZ3h09ICU7ywHwbqbELP00IEXfA
1e+dlhnIusJD55HSbs+NG8pM7oSQd3Vlwzh3PMLBc6azBLTv9/F6qMV29Lq5u5jQHVdAgvX8fPHR
IDN1tqPc0Puvy0FG/mri0BgrTrr9f+9UcsIQslqy6fMM+52kzo1Pc06gUOQkP/2RNvHOBNM9Yw56
xhjYI+8c1DAJ3QmUr9WW6LZC4C7BDUDAsKd3I6vd88zmBsp6qYlZMnlnxaAkgX5qL75dJgo5+SLQ
RAT3rxPuyR6Q46TQ8RS2M5/G1gOGxKutay1QT9WT37RczE0fbxqw2zqjlZwkJLhb+tigq3S6gSUW
7KS+11V6AQFT/+i0FthrLqD3rLyKP4YrMNOWXHuh+ff2B0ax8CLg/z9FVuMGcjkZ6dB5FAVbJG2c
qR6Dktm3/G6QQXph1gjAvFa1oLiHznDa50tzyDBLT3RDqlWdTUWo8q0aakyVWcTxNgcPZT3Slobi
/rixuRzQ9ZT2ISQdJm93419f7GMTA/PUUTB637YsSyhMSvGfga3wecEaY7oXStDiYb9qF5xsHr9K
WQGHK96mOOuST0HrbU390JTzGkXYe+RMY0evKaQ72hn1rr5yAQHahIqaYUpV0F0Nv5WzzZXM5SwD
DFsRmsNSiop9Sblz44BZHX7q+BXuIXYOwGclS3VfTrpFiRgjeE/vCrbgWiYG6B64TDyHkplgpqza
TwFgno2R+Kl0K1RFnc9xWjqb3xrVhpGsi6DMzVYGqYf/sM5itebAdM57D08gAJRckbk9lVUcMtvQ
9TbaogVxMWIc5rV8VGRqu7dw+2br+QBwhvqa9er/vyIEP7zUMIokrJBxQyjeIIndR72gkatHctsM
xuhTRDdReMwv8gvQ5DvcOU4w/5iKZTKsEijbihSqzboZw54xujs/+GluC8fbezkhSjfOn2ZZZY2Z
RXoe+fhQmPWLACr4vCQcq4GvAncCYJuSI5l/ZNWnGJ9kjzOrsc2oP6l8z0nm/Pecu3ra1AcwmZaw
VIWgrAfdVDChi+YDb31ODdTYKUkH/HRX5jS9kKsv/3LmWjlvoPwqh2+Gt807qb4kbfTPYfrLi5F9
mV76/ZqoflmJdeULjznHCMnCE3FC0ptubIvCqBxyCU/f13b9GGsTVXawyZ4tUJuwD4GP5qmhxOfQ
1IqR9ZJbrGupw/rMOIm8El57PI/yFMuTL5JoqH/D5AjgCp53d68mO7HKEYNwW4lOjw1f9beC8nrP
9lU4xQt4C7AMkRczRfHKzQlg1FYWf+nKaVgkFHJZJ+9PdJVrK1nuh+WB5R9L0IUXD1Z9dmBhSrMa
4OdhxapmkTVGfSDOlWCBwgYv51heG3GCpQsPplolhXdriddO2b8BE5Xa1a06GJoc4ZYBloZkGQc/
hCWMTGk0pl9rjthAJFx3EEXfjN0G+yTM+lAXIb0nQY6MUv8UolQfXEMTEz6UfhDgFqNXHNZNKfhA
NQYm71mCumI7fGT5UFQOD5ZscLhtJ/izmeBH7ldbacB2zBMZoclELLgNPVIceLbzTLbx96PAh8zF
2XSWHIfBCh5rgxTeH00HT23NMj+dA+Ia902nYrTspbHpdzmrqhE6chVARDDdC/4t+Pv0SwVd2XL3
hqRVEY3tGwg9+7iOARY2G2KZ518taxwo7FX8EeCCm+7TDJ7XxzSF10lojdWM8ETdJDGULyShRy/U
VNgAVbd5gPbxOGZV96Y87+b2xBjbsJ05J7tzOJctznsrxOYyKTthiafqTqEH9BMmND3ozjUaL5FM
gTiezQkaNXZqdqszMxCREvjDi+ZW/L2aIvlFBF2An00b0ZauIZaxsCh7fJ8spyKXyH3J7ezK8d3K
iGMDcy0XR4g1oTrVtLow5+jr24Q6zYBJeQ3vsx1bsccRgBIB5xeshvUR2SFJ23YSYh3tnKLCmeU7
zAAi/DtXsZ57yH1kkc8knG9VZYUyAmzBXZEMcgibVuz6QfHLQoLgJN5dAaEZoGY01PtpWgIFaR7P
4agcX5qpPCA+ttnwNCa1HqiM61vgCrAx5zjA31hW3TfJkyM/actjZXevZ0tfcr5egR8Oq9SzSmmw
s90mxgvKlYhOtFIGAerTVdDvILRDONpsd4h20ddkerERaeq6Q6p66+Q82UQADKs0HWxb3ipDdYfY
dG02kG6CZLd2NPmqLOF3Q0BsUP8g2GWPmg//FjHWgGgcEpR2+2RM9W8vLEChb0SzBjYccEQPJ5sd
2C7waUzbOQJnoPfz+tTYSGOf4eQ+f4jMmjM30xhauIASgPVnL1XdsgpG8I20m3Vs+O9QFFSzj3hR
HoY8I4iEZFtG3o1i1NZ769pHotqj853nQWgVUA2dPuTzzIVitmOC3pEqwhOIpOrNXYiZtFVfK/Xe
I+15S/ATYKnwK9Ln+NwWIbhHqyKoLlcHhKSYF1sE6xL06dwKky6LdeEUsMR5p/gY3Ozp3wbeyPn3
T2sReoOENFjGHwBZTErXrX72y53HcvXhpt+VEMhlt+LX0EtXnEm7FIi8qAv0N/qXH7o+gJzm7Ks8
oKs1I/Un6ji4FMb/CaLDTlszI6LYRNlsv3sq0n/X7jkZf8CI22xyItbtIlX74JBcdjkgx4lnZKby
IXqanaCLOJCSzTi3qTVBrFAAo+e5siT0/+pdgIaXESjsce/GIhy+0jPrfvvlVO7PsO/7vtqNfHoK
Mo1E1WClRyyT70AVfmF4Ia23d8RnhwTbUm8VmYwiOxxNph4cScRHfjxBXD/TsvqWLARgC/Zitzff
fe56obcDMrxA0HV7P+IaQWe361QsnIm+2dZMGkdw9qLufPirzDANWgW1UMT0im7LVztqAhqKNvs9
jqJiqy6At2LkvvQlzqYEcVKpt+/rZ2okYh9SCQCi5aK5XMBd4zH3kTAW+jcbu0TO29qc+Tq1YlkI
NnUWAgo5ioJKC1bFCf8MWlvu+za/9XOfQ5x0bhluJAKlvCOPEPuig+ag/O3hCOthXVmKGtgltR57
LazEtzC1iAL2ZBsji7YdT1VSJS9v360L3oLza8qAeedGMZvisK3bn6Lxl9V7NENIhfE7ig8CvTvN
gnNR0rFRbh/IxjZM81Y4RpLKm/0iS/YD4fcBrWlxSdJdh4eRbp3uBMeKJL/3DPeUyPAKFz9Ha+i2
qqZT3zhtta+bak9o97Vk3BYsWG3GxTgSZC17wrZ84JkPY3HWGW2JKB+2GndR+aJ3Af4EL4ScGJQ5
5DtSwi90mS3BAV3u8L41hEbgPNffH9UOo+kulVCzP3mmjZlfqbe6H6vkMn5gJwK9NqAkLHyCOx5Z
nHXnSO1BWISri3+iId+LsVz8bGipililvM6X85MZ2HlX9G2ULlp4XGnFRtbcwdUXo5YGye3ExjKk
yp9x0+KQrIsw5MJxDR+58TJ2EFwSx0XElPhEjHrgeJL6mE07aPiJ+5naMgyrzvRouHP22JK2wus/
9BTItQivE5MyeTZnpQb+S+WgiiEF+YZwnCGtiEuIxUT7rQ0CcS3HF7ZhXNu6+T+TeUW1SBApYfA2
KGUsHdqQManc94kz6xM2RpefQZyF4PkNx6hCMAg6+Erp5bgz8Ud8ilol8rFvpRhlmNEhjXRZHm6i
wI6yrbgJZhZSvmuRI1CBiCbnFE2wXKNK15h1TxbdWaoPEvC7tuPudd01UCpMMHOTgTCLWxmuHHm1
lVsPiVcWzCv4pI65VfpZGLORMIncGKzLX9/scF9iTYYg52/X6NC6nJolh0Hl2/IS9LQpFgD6TFvS
OuHMhEIS0EOJr1i2ZMGhkSDW3DGfOy2bbLHoorkvxAoZcIa85emUfkKxYxTEClMvyFoRJ0d5evTZ
Z6tfYPFTiGuE3I0NcIQKROdbBJbOc5gZcOXjIdyUJQm7X1ZN/xTgFuhrPsjuvXTO+bmlZ32SOVWp
zae4Lr1kIV7sfSR7L3JQ121VbyrqoHpBaXtTPIYiGBzll4V5Uu8/c5kFqxPAYnCkiyypea+hdWCv
rJRGdOcnXEEMEm9bJ885DPYzCvkYScmCvC/iSue9DJXtN6n/gwHycy2IrLKQRAXuK02AVu7Dkm/2
2q9H/OpLuNiPYeUv+vu+WUhhkAKxONptGIBqX3bSSbl78w0G5cJvrEm113Kaa4RAqmXcNNiKZ/Ox
i687Q+RP5j3twNgU5y1rOv39DjVqdMczBDvvDDVGNAlyjeVxNA8fm0MFDcnLV/oHKfla6TqsyS9r
hcXcxRUUsNt+CZ+0OKLz1UBsNJsHj47jBCQz59vlUK24wG21OzyuOkhsv/mXKF5RsY7xx2awNNMt
WcFy4Xe2CzZJh4/IGDEGso9a0fJF4OpfDitwFpiUkGWedBnW4NSHKDas+1WRy+ZKUCFD346zNQxP
fNLGrUvSke2Y9DAq867bI0pAwa8ccKxdeQRlPus0VEVUIlF/Q4tCBnnYHzCifBnxpn9Wfo0ki3VN
TXmEfYHlTYMV5TOMiZAw/MRbuaPWwk0zII+JCWNaDqJxhe1NFPRiaD1Bm1sxynzYn1ZA0DvlF/09
bFXTxAGj3VG4rQWlCDu48XyPyAIfuCaHUw/IQIu49SiTEkn9wtt3SYj93vxpCpQ64lPtm2OVG8w6
VmWAvANr+TzqVS49pw1VjxRaU1hVsf9X9O72g7oY/gyajwziyUORtNJ+mSvirNHf9l0ka6wV532x
egpw907MorVw+Bix65XQFkT0Jgrkq4MIuJAZv79BrUPoBM4ITfj9ztyoWUND04VB9hUr8t52bP5k
wkSuy9XNtOeagFwfnRqYMYvR2NYfwPg67655Pt9kx6oD2p0gSF7PeHD/bbwGJpSxV0WVeo49tSKn
5GVstTZxvLHdfbusbrpjbfdqiD9KnGkQZEzwDXfCKOhOTJ0cLI0AIDF4MJ33B/FDXfOaUxxtAD3l
L0w9bBAs6SwgsI/1dMGyfKuWsAf/yIBi6TgRvfSc64Ljx3b4lWT9pAEQX/1dLgDu70LfCjSaUWeQ
7iWteE+eom5locEItldutSKDPjmV6QtZ8F5nD9jjXzZgkkgIQrSyaFjVmataFUHw07Y17c1TKEuu
ULOCqCvLzET6jiS9Ml2Am3KCeaa4EqIbsMAy/971sifkq2q/sT6ClEf0i9EkXHS91x71up94Qdl7
Qy0ALQ3huoguTn0G3dbCuzuC37YiV8xII2z2ZIEBQm+ISCLs3gGQM/+BbfXwaQBMldL7QEat0pkP
HBTbv+HuuXGhJiciHWVeTOEXAmEvlN2BBuB97AQ0he2TBMle4A0FTIYQo2oEuTJs+5Ay2nzEwsQb
u1+71m3CdEYRqF/YNAd1TK2EfnppIPVS7oeHBzV5pnEm21NcB6AebADsRjxnyQYafBmxzpyCTCsd
y24kMo1kOhAreupH5mRar0RNdvkzEEu/BtYBYEWqvnme/RhyU12fnW1/nowsednvah7IsdD1wGj2
Ozf3s+Vdg7vQ1T7N/RxSRhkL9y0R8K5tWnaH8plDno4cBQF/vBRlLbP14TnFdBMqrRY0wH5Vy+4y
X96nPtD6J1XDEa5DIsX9ZxiGzZ9oTNRa4f1L0hKniquo25KUzaOtUy5BRSbtQ65nQTmYhNPuiLCy
DR4KnowCWihXVHcUYNF3STIfwLUfSjooJmiX+qqSJqj6TZD6+Un4OrS1XDX50QEWnYcoEegwjOQu
V/fNB5NjfDiPCCn5LYxPcnkypsJM85oNCjF2f5VommAsRA+vtOxO3A1DlIo4nH+/CCBc3mUJZVTb
/9+sjWpLIsJL/TPc5fxYmi3QXu7lfDV7+PjSAnO6/Tx2H2PbAqdXclCJKYVuP1oTfAu/CkR3xvAU
GZvERhpO5ov2UZ9EsDnZESmbpVO2kCcxfQBxdlq0/pr1c8ZqzQJxVwZoqPPMjF5upIEgIXy0cZIV
CAkfIRTltd5c2uCUTrVPa47fZJHUur5kEseLdirM7wP40gpYtPqz1NQt6R2T6HAeDspmlkK1jOw+
8LY3oOrQvILxq2PqVot5aQRawwn55RkbT/V4dERkdO7HyVEK0LABPtwFNEZdlWmDt6CF663p8oXd
eK+86TDnb8viuop0XPirPbTmeOZ1Nydd09J50HKJk1KEEkLloFbVOq7aqYyF1GmmSEe00yNxBYou
2Ad0sIrPboCOJv5lfJLhYHRBG4kzaQ+Yvoid0cKQg+CoobwQAt8EU4cWKP09UfKQfVwHdPnCll/l
z4dDIvQJRulqPYzgmR6TgrpH3c30bEFFarSPs3zcxkrjM+jRAgv8LFFNGP3cWmwhgQYs5nFqAQl1
kCR2YGhfGbx4LcqJ0ojhi2q92st/Ji/U9Wl9Z7weKBax3QU7/JoFHyWCDwwPSm+MTCARRAhSAgGr
wAl7LwaYW3MYPoOOec0x8yLsI/TClhuOkp8QwgsfzVBYqxcPdEtKg/lZ5wPwR7p0nTMOgde/PbFZ
2+YEccVN4ZLGiywHkEj0jL38QFVjecAJDF97Ime3jbCUAXK3VRzf2k4NbGSSTFwyMNSqWLLKfjiz
aJOn6k/DI2TkfEhRjmBcLojc9MSztWw+06bdYqPUgYxAJNkP/41helxfxXWYp6wZ/JKaNreagYWk
0BM6t33DWtMwh9lZGh45gyQ9xUCA/vNXoq2ABT37LKqW2OHguJ1c1OozZyfuMVVde5hiLH1qSgE+
YHCLe1oSyBH0qFyuO4IUPhxuoFmg3GZLZN7Qf1Ld4I6XAjZyVddIcfMx7feiHNSSneq+NaGbpIay
6Vka/5n21MyIu/IpAP6B1n6L3QH02l1FHj+9fs2jgE8klObFU0gQKS9O0VAH7fBKDb2c3qx2S8qT
CNw/8TuwO5wc0FkfkJZQhY8JxFfoNC/MNzFxszT0XX2ktqFNHOAKn+keX5NB1bJ2iPj5GP3G5972
qPpSAevGO/Wn3B7f9RThYoZFosuWc5E039zmfzT0kzInkzKfBFGFK1X2kaw8WgnPtpuAk0cjou9O
sG5pOrnqWI7QtRkpUCm3yUcV/CN9h6pDuJKweubXJjtJifyLeJdPrzYhH6dLT6POII9G25XH/UHh
8zhGS9MIg/YnSaf7J5H2Ap7dGrslraFpalgT6II9OGFdZMqIjpGBfFFW1EwI1F6MkRj0fhjqa4Xf
cOcIkfWb+1Ic3XgP53mn+Xyv3ddOT5ESZACnA74vPGfL8YOCYYHa3JQBmVEsMH3hzvwcUMy2Xou3
+VOJ1qEKZoSumfTMo+34bGeiFnuegHHtw3Ea/ymzZPKRjToa/wNBlopBEu/UM1OKk+X4Pktw+mql
+VwY4j+UP/Q+tCHVajluyTn4YW3XrZMOT6zX2RIvQGhdj6mAhbsMmOVa7EZmzlY7wVtGhhrKQ2um
R+/7D8XH6ncT1bJfYNosuvG31+tcABoUU4Th01Ofz/U3BWuIjWSLUFl6mbzldCDNvzYI+FOrr1gu
JcT5LrzuUI8NPgb8qVDyXz2sZANbBA4snkNuDf3ii97GllUU5S2U+Qk2EnKDX/35QNoVko/djYyX
2K0E53rsgVr8lj6CUgHs9/68KUFPBs6eFLvHEIFUW+21yf1dQlVwNySPNLl0u0RcNzRVUgvIlFH6
PYDEqjSmq5O5q0Rsw6e/rwqA0jwDnlAm/+EPPjTowVCTIzN5VxyLYwspicWFIc9WxhAWOtcalSwC
dl1mIvhQqiJbSHdKSzwQrBF+MHAGiqtCyASi/JufXmgOSipgbnrKFZ04v1U31y5mNL+oQR/KkUG8
nvhBDPcTwFMUvS3UzGZkJx2Z87HhqW0PaPO/33WpWm5BeZKuUfoYvBtKwbA22yzsBuPlBuiJi0go
Uh1x6rTyl0x7AotKmyur75roiVldKUTMFkv+1h6dQiTfaNxdXNK3OrFGijCCRUPsNe+eTfT3ev3B
ZAR62grLqXQESSW6HOaphXXNX9zOgZXXth3ZSAi53AozX5E3G62lKkbKX91vALemKWY+lecV5GPl
7pVHQgx4tJKjJ9Yhk1UHjbrlzi5eTjEdo5xalSWxnl0JQ06oz8LPQlpvJL9axTE6mB7OkCZossw8
TERORirVnZ6EQQxU0TaaTyEUSzlzPObUzuDvWNd0D6GHM6lXbdI+RCkj35sCQ+i5n7I1kDjAoLPs
kArT46Q5r51DElMaiQLcShOISquzGr+emsZ3+FSO0yoPUh/Bkh1c/MYIofVjo2F0XBahRbJ8C+Cj
dNvQ8UOI9hrSioNRbHDLtVz+4p0tth3dZ5UNuMdjCGfDe9qMHzCkQXEHBJx8StsYYDv9WKUlm9y6
xYFAPkHGiuidgLtjoQyl1Hb3zIEUFmZhgx/4kXN5QUdfKcsMsRDceJwGuYgGdGo75j8yglbHkOCC
JvQxzLHEL3oYqEhwowPGvaS2itO2vFQ6TTBk7I/H62226PgA+balEdxkK4cHjIHUbwLP7TgU75+2
OxzyOGdD4NyWP3kuYNpoMbVt4gM3Gd5jHcbt+TKdl7+i3StHS0IaXOw+LeoYQV2sJr5j8c4vzeT0
8lKYvYvu92Z3/XGTFQgm1AdQOeUOJ9XhZvP3zEn7Ub7MIzRzvbM7u7azSnBXk0WHrzD//MzPC3Fr
Esag3TuS1H151zW/acmAKyqkKVHuEIDzEd9svgt2j5QtMTEI8Rrb8iX93id+IQNGOW+UkmA1+qom
0uxX4TvsR17982jQTisIa6x2VwwCTJDC5AqI7RiDkS8nabTi6KIjUMoGX0Xwv/mEED8XU1QFwM2P
FfDKXH6LOIW1FA4SGU+Q4Ozly2YiJhja5QjgjtmS3WmUxU10b7a4P1g+1xBXlmObulZ2I6dqtSMp
L6gpvQu1+FgEvuNiEViHYcPmer2pPEKIXGMuKkm76unKOS2C+K+9TNhbqGmg4M1zmvfKW44/Tu5T
/8yWCdmCLjBt9AsCUFvAfu5S3nwJhFHUgz4mKk4Enl7Jw5blg14JI86J9RZqawuVtQiBb0mJkRUL
T2qyiWDHukGFiXJOL665yVv+4WgPD9D35n+o5iJQ/Ph/7XmiudKe4XTO4J7kMPK9X2C9F4AMveaw
D/maRWcTrB8YWCNTUO26bp2vnx33kR/Tylj1RNrT3JLrS/QqxXg8yVpSvqELa+cJsAwYATbDVbyD
2dHDq/VBmRr/UDgctiPN/NFquCWqcp4Xl1fODKt3IRhNJfmgrN2LS6yGJl91lWoF4StKB0mtn2l4
nF+/igs0GVI5pa1wFMIXuStAbc32qEOOg7WYPqZT9GBxQRv7/aVigwtItwzB1Ql2klA7YuzLB/98
BjO+xei008dJ/EQbpkd+YUyuCgwPNlVmmocv1jRwAzUMemB2+d5LhWttb4wKObNnHaGFhgFFLkqD
zoHp9p5W5hrMX08nxESDK42vSNB+Eoh9P995SmbPcOgauJl0fD6vVrvtGq1kt/QYt+1Hyusbt2sU
E4yjf9ospYQo2pbJCWD/1ArrM41jpsybXgpRy7FdHJwf59BxwhKXnxtTJyqUYWTqx+sSBDO5spkY
cdAQ09JUDbJGjrGyapm2RhaibIKs6797igG5fSRvaeXq5y4D56VAzQj50EQS1iQfTjxB+xzE87X1
KlKY/G95OCc8WsKHDBXzHPS9nDSJ8xgaOJIcAAAeyhN9QCAAJaMfbERR7FDL0x42AjXEefj0zogF
OiwbLTilISlfbqkp89+bdG2jupXUaoCnN2xv2kN3HLi62SBBUBdbiZhE26Kr1rc/SW33elPU5ax8
W2sijXDY7KAbBgr3hSaWJ/MMHzwvNmat7dSR5E/EY67HMn5RCAdSpk2/JDHZ2F/cFQ0rdJ7ZHMr+
B+mv37lSCsr5zipiR6z0wnxapsxnZV0QP3FvbWNSxBMwQtSd7R7AjoHP/sOJYUorcBIS46LcqvOi
DffT4mIZUwpoXfEDiCjCPtuUSVP3QpL6NxySbG7s/4YWrF+w9/ndSpRGmw9SChb5Xm7gt5c4L2U4
ROf2pUVRvxcxC7ZgKmW0E+stYhs7FU/HF27R9sSZIOWl6Z/AdmPEEO3VeLUWPdnOb8xPn1PBvta+
8ehb0X5mNRirCMFkGOuSEhcQZvqHa5kYdcHdeIWQxlamBl3Q6cSCkkhl901P+AlN084oNrPzF49S
2ttxYJ8dkxYOYlU+6XvWA8XZjbgAd3f0ZXq3ml//lmtpFtRAFle2Ml7Ign7udlqrCy46AWJfep3I
/AmZkui2CW1qb5Z3Z7loYMsJ2dlSt81DxAnkWA5uZbohbrJbMOvyO3HxJ1MopcNwdEnJjBuYT5JB
AAY+vGIcUyH/BiuCaKoG0TBTciEC+N8uysFc/FOkTJc8VT5eHBAw5GqqBhGwGadT6PDEelji0KCV
h5Lb1ZLEPM5fHrzCEsecqxIWjRtcd6J/esIQ0eJYzkGmIwYKLP4j4stjyP2dSMAkdxzk04ZPprvJ
tC7SyWtUnV3RbHkRM+MYbWiB/Cn352GF+0ixtLGY7DrGegGMgSZsP4MjPhbVjKRNl9dl0bBSmf+Z
y3XsIf14imOhQ5b9LciEWBpZBlTUjwGozao9P8VUZEyIF5jmUpFBdEEF8uEWkHOC0yC2QZY7hsfh
9+aKZgzhoU0MLHlqdesB1AMK0EFrUuj7u9fk2puL3i/8HMu/BW4kYJGyYb3Ng/zg434lBjcc0uJZ
0jd6PzoMg10FYACY+Dr7ZUmRJSqv5yFWyuPwSXgUNWDXDFDPS87mYfV0565SsQzHQa1Rwq6Pq4BC
9OHLS79XZwvXXgLNG5VzfljpWfAot+XieLp5qv0my7S2J5RcJGXudUazwDxhfKECU/9nm7JO8TmC
cRJB7BKMfvDbk8n8QPtlI6KBAT+0WgwE854n1jz2Kdg1/WSTSogpJy+fZr99TXnXgJH2/bTuy1h1
m8iCvo4SK2QfbXbD+vNTiJHz0RyK/kf/q5HQAxet3jT9Dp/wGKS1D8yvAwyAlQJ4zeZ1zoWr8CX6
hUgZSONyF/EH+vWfOX+1iQSfjSEuCLRs5ZkxPOgdsCesez18b1tvz2JwVAwQLwJ1eQLypBkjgjXD
BPgfg75FHW360FCMW/HYFQ508U/10aVLn2LfzzG3ZxrmGe8wsINH3iQgKx0XiaZdfMeghbRbGS6a
AU3aFs7cTF+2zke64cH11BjqzNl42yLNO6lqaRJsEPIBHaU52qmVt3ab3ocXXAEGunQhclfpcCCe
BEAW+kysqBQ+7v/HCBUFKZyDshGUi9EAhLg0/iqKM6gJ3Pz7Be8VM0ySDGieDDyPH2qRa/VFMmRN
ryex4ejryVduj/Qq6EJfV2VwTeLkcu/Ov5WDThD6duSc2XulCCHNwcy8eAXf9XeNpL0psDBcqSSQ
TenL8S26YvrdGb3paUoRjxr7+iEKWOphFNWf7XP6BgDnEbMdE803i2zitspzz+eRksHWQJ9sc2Y7
AKUiZ1zP+cKl6mxNR2rH2FR+X+WJqvxkxcVrQTtQNYF1RpyS6qM9h/KYxzH/a0UrS1vRdaAO3x9Q
vYCps+s8UPNH13hVe+xcXcqXH+nA4/wsIRRQGevbdGjpiYJOyaEDt5kdZqMcewuZIrj/ri+rJ2oU
dyAlw/5tncHF8MwsH1408khJ5Wv2/41HoH40NoNFdNl41zveifRuxPiP+2jSetMvnpnM5sxqJPG9
lFuw9vEjbQVpvnmhNe7q13HikoPS9vTcyfh9YV/QF5fd5ukblazyDElHonkmbYb5BGM1nx5n7yfQ
eiP2WPd+TW+9+DFpJ20bLvgIN/H06asOXAJkKXj3RTdyubQqMD1wUGPIEYnc/bX9+BInJk6Qvwuu
yiDYjOdL78AphdmaPKKqWUh5mDtbQcJTJP+/zhyPJD/DnROln90sHivAybKYmEpdD5uKyM5+blH3
Bfl+eiDOiiXSQxiTG9bgn0FXOnDVgl0pHQb4D0VG6v1E2EhyQBFIAKB8ikeVjN961WKSB05OZJh5
+F/Tb3F4DAfy7jznRp2Y13EzaNeRcRrJ4XMhlJvUTDjpyzoOSqCeW/Cyf9LeM+1udPJVJpvRwJzc
pRftg/UdyLi+F3NFGpi1po1/rCx2wFn3o3A+29NxowXMwDSkYQ7AeFoZymTF+RCfK6xUYVX3PKC2
VtVZtfyq0eq5tOilATP+P06u0RS5weBvidyJVl2UtQ4LD+lZxIOYCDhSXz24/xYE8TwMklXKxd7F
756s2BHbhKfMFLIhEU8aEo3/WG7z7vi9xEtlIqAIxmyI3LjbpFL3zqonFv1urOMtt2mj3ID47ytb
+mCSAxmVb0EZHJCz1ihC9JBu0VauEqZNApSDiuE2INUNcYFTUlFfXm0pQopx+WjPw+6sgkhatrPP
cisv4Qwge60Yt4j4eOulVR7Y0LpYitAug2FpZnkbBRurVVJnNcNHSOqRh+mpCsE9LvbyRL9mOzSC
0APQ9Rh7bN+dSAM/+EqYmVgiE/p9iIeACV/pG2iPr/aej3nhmjWXIJpfxDtQczlMI8iDbTzvttNh
7FpM0/w/MCTY6pN6QE0Z42HKDmKLkBcaJ9J+mPFjqoSu/20gks8RpO/HAivIEZJVufRueurMi0jX
DrCzhcDZSeaqiPx2Dzi0Kk0b59vl9jGc80M98Fdj27BPQLqEPyORM4q6kpXXrixnFKragWM7q7PT
bGpFN4Hxh0SqW9QPlol4hXoRgX07gAu5Bms1+m778aGepCU0MAEKnlSXKnu9CHwJRnjUG+68ISRe
d45H5ekhaL7n7PkBGLAdBle3tmVSc/FnW38I0hEHrACZzVkbJqrYi4hYh0A/Nlar9euj3jKOdxR5
NBkxq59FSU7uq+ODlzvQwU4vBdJqSNssuypm9h7ydy5Wn+tiz8eXxu/q/HOvjALrED/Vae2HPGLl
6/q36reFtUrzUTnbvlbfN4b4uUyR96Tp9jTfnpe1utOj52VlHrqLyvjof3JxWbf63TpsvATmZ3pN
s2atj5VvuzPiBw/41hZqB9SCfBcGWEqgcAuE/GusZzxnzCDC6cDizRA7EVBXY8Q4RCwsp0Jr0QKA
+DnnBHUskDhGhXr6FpceHoXlB5CK20eyew2vaQYH57hasO4ZCRrhRGWxlpQmqiuiJkH7PTORc1Pf
RhtwuBuewgYfXgARcND3mKM52U7GwYP8x0Dh2LNcS0/mAPhyYKkBgAoHHKXoaBijC1gsYxrdMCf5
6Jc/setu5oZd6mpd5UGiZivDpTExHrU67S/CKnUMAG8gx3eySskiW/6d8DYk0GKDNNtubIOMYz7+
iH1dsFBnw9LmiPpKIAc93Tv3jnneDZ+wtVYB69D01nlZA7m/ohSPKJ0C3dtd3Oden6sa+0hZCxGm
pgPHvd/rfSmHZbKSWPSmcTdaLCmU5TLMRBvjXTA1YI2stJdPrAZ2j/5Vcpkegz3JDVuogdZ9eAzP
I2xO+LQIKra9BC2gTnv6kHyoqAWLgWJhx6u+qdJlXPnIVUjplS7H/vcD6XMQ6coBG7S9yrDEN2PU
qvVpy8C7B7P1E4TFRM4XyvuZDfdC+bN1b1t0bNvpNC8mqv2WRfr4gqhMrzCIsSRKlVI1YaLWoWUO
ezpmfB4flJfbM6CK20BrTvh/S/pz59QvfZwRIahW02lFl7d4TodV36rjt7pga6ooX5WrFRJFfDMr
ffcSH3w4Het4AJUJREyGpuAB7CuoCu76kcCkqEH0XHmi/l+KMVg44Ba2edTt0cWGonvHr6TMekKW
5MEqogVqsI75Me2imVnwN+ZUiTdUStQlC8sAVC7K00H1UfM3A52i3cFRxCWL3cJ1d43jbw0ncMBp
VUANqafR8APhkLwfzfMPkit4lTU4TI1DnGRr60xdAwMjJ97szOBs+OstWZTLroc0UDHqSh0jKyBS
QGdCgT2OXqbkW1cbGBuWeIrRdHg8yayLUbr7mnaiYOag9arxQsXaPMrysqWEaHHwZCCSmda0N4nn
R49wv0dvrcwfFtYX6QNWcMzlaYws37CNUT5q+7ryqQapb/Zn9OnPyFofpGrtTxcHr8krQk9OLRIP
ViN6OQaSP6/tCKGBwWtRpNBRzjYaHSdFSeaBhoP/rZG21SvNl9rMi3l5xFX/JWScV5/PcH0JyW/K
+zMh90Pmd7MsG/dbR75RWg5vTOXlx9lB8iU6TF2eMCQa3zdS7g6e2w8gio7gQzsj41BSciU4/VvJ
BXeAOKMkT/6OFawlsQEQYZi1uxFWxaLQp04FqBBSyUXdIbgosI0nZxDxOxPp2kgW0+2M/2h93F01
QlcSgIU0515CKvuGnDrCfqNWTc3VzD8mnqDFsl1oB4UxbvrXGJv3+0pYPmmxHWmcHIHvZ2zt6dUe
7vuxgw6loom9qw8rzXWuZVNdywt0oe6wDqTLcws+vJIt7cxHoA45NHTIohgyXDEWStxuHs8SPLfJ
kVgzQN71jyH5Njc11u9bh2SxwSij4XLvBdoGYqSIpneB1/1NGe07dKDxfW5C4QiwsjM9M5P8KbR3
ER6YiXr2ZCVYuYXu+H9QGzyeyUpU5Ga9x622/sSEFmcFPhPSBvY05yoNwtnxkNsLZaBhLXDzAtqw
wC/xGASOB8he7rDOW4nQpjj5R3njS+dacAM5cr9ozyXdRi6SYIjJwR11q0E3KdhWyfrJ7Ryfl8Tn
VTK8awn0qtaVHxDP9a65VNadA3RnYL9im0iQF+jGnN09nb4ToTOVJrG+jNNDojpOvLThTsvouH8t
uHBnQPwhAIqALMh/W/ZpdTPl5IB7zG6pIpOSiyAs+eLTGzEpkMBSyC4z1Uk5oH8Pu6FfVky9tfBb
1yOPrXIVZPpPjcCrmBe5PJo3y2pwns9Pna6vBS3/Bj0sOvF60CkqatEMt7ZQVa+QOtnGgn28rLoj
nkgkJXQT1xbpPbgCHph2grUTCNIDJo9K31iN0E03worR0oOBZQyMwiYgyACEi00ObrMOj+aW9RB5
7bdiJXvGRW2BaFs8kNZH6Tz8h1sfgT78NieAd7pZsa7Qc66zjj4BNAVSWZtqVRyNEpgDjDzluYJN
xh8oN6zgKOtD+JasOlowit3ZwpEmeWAsJZtp07pMKrBZ5gI7lMqYDhs8kC2C6MlDxlvyedbAG+ze
yeXMMyWJgQOcFqarlpNZp4L3JZat5btUa+J5PQ7W0hnEhjYYINTMPD6AAXlVSeVXIWAeFAwayc6o
ty1eTGZHPa1FDe25Ya4hIHrJ3Iv1vNPP/grGpskwPZu+vdHjxBI+lFWffcT1bUu+M1xI099U3iZi
7R4EBZCZYkq+S8coVEY2gkle2mhHe1MwgFNR/T8cdA/m86TxcISuq0dWKtXooVogBziH/a5h9B+R
PuHC/C4w+8BPbMH7zOiLet7yXiEI+uv0vnHw2AtwUWyCMr/E7kGY/L8JiJqRk6W9kmnD3Q6RZKIu
R2ADffwazi6kF82WRm7QJWXl0rJmJsSbrirIYKq8oKwyQbCAWA01kmKjnDw2VDn3RYG5IN8bYN7B
xJD0ROFsJsDcsxcAngEnIeNEeJ4cnr/AINMRKSyxA3G+Tx3HBgSUI3dWyjuxnmGYjfQKNKZeBaLO
PHxsQUaHLigcq2T29w2i3qNrslROSpel6DDuOO5OzGRkPRw1nQWtkPKqjH51R7+RqyaXIONgDfsl
OvQQrPiKNexUEs1p0n+slyKi9oCewOMerg9mA6F4m+VrxZhHw6brEAJdMsLSIUKvCC6VPvB2XCb1
a9bdmr2F8e/qipqGM2/IAAT/o2ZTK0YloV8Ho6u6GRsajAU2c0w0PKOq/ejoDgMKdz1QyHUMfook
q+wdMM/h5MlFy1qsFOhbkTOBKnjF0f9pwOfVxGED3k+PYInLJpHfJYzMEZwABJv6tASMqbHRQYFt
TaTCXcDLGUcujddau4v0oTyAvbfKIPiyz/IsooUsj5L8wqgAn/FwG+N6biNnac+786awD5usA7c0
kRRT8QWXIh6LZlo+SpKFJ9IdI6X57/vXAmLy29n/WmVecLfEwa3pxRpW2ZnefuT1Je5CM3mEk/2o
Bbfl9GgHd6IXpa6BSuhXWdFQ+OR1h7MuvRI81y4oQkDg7wCptLg77GFJQzHAvRtcXXhLi9SHcL4j
Qe18Wjj7HOhaGM2BGpnHoj6XC780cHZpdUg/Kc3nQOzg6d/n0I7j6WnRn+ujgBU2x7Qy7aMwWxKy
kmljOvopEpbh5KFj4FaeLBNe9a3gydR2n2R1A7ucWFwj9PGv8uSCHZEc2K30/G1vlwVBh3gb3dfw
qaVio482ECerhIZepPZXbm9wT8to/SrvOTiBY/peA/kphjzoMe0x1b78njUJM74DYHs+WpIjYHBu
kkyuDspQyge/104k4p62H5MMU0F2zNMN+70yYBzlkafd4eecMU3PEihSSCAUYIouVBypC+TFEHut
e51h2lphVC16H2Aoiji6c8n+hZ3m+9C/7dxnTYvFwp/ieKEqKNYwLiIyzhvYGcBiHbmjmlQYVimh
POWmixSwu9hFzIPsn/8qBCprGLIj5QythGOlLFSjFYmVHyKigQ6lDnVoH6Kk7z5JCz7NmcnuzkY+
0R3iDuhNHlSDiLnDpYOwTCQ35jCsnPWNiZfZhKrgeK6UN2Dj7LhrOUsPCN1RBCd2YTdbxbvphUk1
jfFvb8KsVwxEhNQV+xUQ7gNxjGNivNqGBurly0iR/gl+kqXq0vaa23Frp8e4VVJ9zRZhTNOgJRav
UwLzs4SUkTLnk4+7Zayi2rM2T0pSe/GOHPonJi+bJDLBt1IlJjLLbLYZ+XGIS+s3HGcUN/HZK4JI
YpDZfCfDEc6MDpQXTON284zLXcsNtQO6h39svfowp+Czt5yIxRZbWO4g0pAL57YSS4NOQGsDy8zI
gHXNP/Rdq7iYvBIzlm8MWJ16fSOHL2zVf3jygRYzclDf2pWL0rB1k8yYZMj5AANdlmoOSz5XUuow
drQoMrP/hOUOjBhzHtlCKRAKKIrcFAol2HeqJungEYt/CFmU/IhjE1dee89LzR1wcd61/jr3LFaI
TaEoZNL7pMymkfLV/Y6jKt1fljoGnFfpXWvkeDYlCme+ajb2clV5tA7kGyIWbise+7FFFdezmRqn
DBaIN4kh8HYugpT3p0mBVC2QmCwrtiIYOuaxV9Kvu2jWK5tBQlDrePpoYNHdDZDo+WwG1i5q2el2
YnOdxC69bTqnWD9A+3DHWKi2KzLkcRu+k1c1gNSXKUPuut43l5wHIRTaOYvUoskarjSl1159G3Jt
0mg29KY6MZASZdv8DJVYHnRkYApTnLPoWJIz5nlSpFluSZ9vBjNeWN8PysagwlITlG9qurev+NHk
kUnTritK9NOWIHoKcQ5MuqWImB5zkcisYyhD7D8RTxv8ZAyj6ECjuWN+3e9UYexNf9PoFZb8cxu2
qrg1sI2NaLKmST4MFCoGeRUcEQ+3YWQ/eLN2lCAhI/eNXcVJHX85BCi36RqkleTQsWlfTHWFtttC
D99IZJ9uIPo+C+CGzFIRMSa3GL2ZtOGLLpSp3VGre2cqZN7Q7BbvGqMBP4zHDoLaK+E8Gp+he0tn
BZb9AQB4i2E+e2L9aIa7q28saA9ODsf+SaUvEi2IalMn3iLACCvshfuWbMLMpUPgnW4F3yv0+Uar
0BiSE0B4QYRo+l4nOXHZapwZuLAYF12y9TYfRpRJV94HQ2YuqW2Kj/trsiFjc6mdqf2GZX7glrUr
GYFFZuAymIfR9GHou7bG/scIILr/5O17YN+exAEyyFJWJkx0pFVvev0r0yT4u0JHR0m7wU24KpoR
Uf3mS44vyt4bKKJZivyPbf3tRxzUltnbafmd2qV6zhTOFcUS+V/cX9zk0McI6P0BbCFlFcPl50sj
PoSIFP7DWFpDPm7yhMFNE4xN9RfT5kKhkmhQsp47wfHViVkLqJ7hxslTW8jPP2YFy4D7PcDy+DM/
F0Avq+G5lFo2thrYKKjMBRrgIwDg33lExBnGNaehvkU8ly7762zURDwygo/MFEIRZ5d0CCtg9fZZ
MiGpgRF6AP/3UIHwGh/O3hp49RnJk3jUhGVEl9sISybz9TEbeGvn33H3L6VnCB89kxHkFRf7yv6l
7gdlAQMZmbDolRlXSLGrFl4rRkMznLOgBqrfnXJyOhnmj5aWR6OxRDNnN2oNG6oJCMU2eJZGjQrO
UOb9n7aOcaBbozasleF1ShQInZ56SH3+sSdO34r4KJtfFEH3/KmtSgawRGPXbkdS8GtLors2AaKb
yzA6JFj40+h7lYrayidnIDaUTnsexb1BpTUPxHDSIwN8qNat19M9W6WcmhOK
`pragma protect end_protected
