`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
G5iF7uHN6uixJmVNsQzPYWIV2bMMe07tRcG1WRKLdabMQR1amZWDIrDvqpa6jT5+aLz3mspzCX8r
yCQMB25OMAd81SdqvohTP/UCFuD/XxjEwJAKeVzKdfQ3IRnvCKk8ID37RDKMZCJMiXTTezSvhDDN
mcr1qtpCw2OjbrifPnSQ0rO+xnYbIWu/0Xg6KYVdeUAkLQ3vno/DEllGLr7gJ9ee9wZr/lec1SNG
WEu1KzFdfDSlCywgvm0x9i6lkszXBmP4/4nfzwQyKpaG2qE2t9QziDuEztthuHOUajsZwcwLBiML
34ODEp4NkIMaNsVFLmLQm96sps7SsZNuhpS83Q==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
bZBNLRsV0lLSd0y3au2q2SFk9st0qs5Xw37wAFqVrSEGK7f5s31W8cDhwxNnjO2VDvUPMsONvkxi
pjgnhTjvrRa+rb8Ps4bI848RaD8e1qE3EVMJpvRty1WUyik4DDyC7ffMvZdHWiyDh9At7CEO10mZ
Xo+FIwPzjzoy4u3z0ww=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
NM6ltWTSLLcCTqVC5g6y3cq/g5DYGSxNDR14Ge+WDkWrVax3QDEaFUfcnmFV6/2UToqwlOBs/qjK
VKaS+SGmA3ptbiMZ/s5oNnigNyInrfklDcdG+qxsv9bf8d43TwPeEPNAEs8Gvn5uxVioZMUJtTcH
QLyxpMuU7G4nwXIdwrA=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3024)
`pragma protect data_block
pkWYWH55J3CRbdmI+nyIilj+LV2sSxSew4tBNIU/PCTOvM8MiwyuXCJZjOS30ENTbfPY/MDZzb1Y
z6wvxJv2KlGWI8O175HZBDEqEPP3ZBBM9lVz9Zl4WwLq9spOfy/R+oQhFsM+unUkr34tFFeSVb9l
ZxV3kkgDEbpZntlT/Og1hE4M1V3zoANnegH0htTqumnxQSmT/RGnXPegkEbT7Vs5dykVMj1rnIjw
elEdqhddr5wnjL8H3WUR5Y/XkBrhGtGTPd9uHGtQ7yWIPd8ve017Fqj6qnAuz83VYDXZIMPFsw3g
sRZtm9I2pmVoeZzgJzsVlhBfJGnaBpObSR6tLUKqqiMWcmJhDy8LNtWvQO4XvtYFZ9hgdKahlgY9
H+5NEwRo1OlvlsCg6p3CffCZsfphmC6i7LsQVyJOx1VL7h8Sn05FZ+tfzenYrh9MbKle7lV915o/
mZN6WV39aRfqh1TK9ex3q/gT4gSg3peNkznqnI+9yvuKjGtng5aKnADDYqHldqrDKr9M44wfbWYm
/cCmVOfQHkxd61kwwumUz/HnTRMnN77JT+PEhzGgclNv+FxlxB4sIYjchjc5HIEDJONHv8SR76rZ
arfJx9fLgf+4RtQo13jp3jg3M9VYe5JbdDkkinDyNCrGgcmdbIOyWO6ZCXPXEiUaxvMU33ZZAvnw
KacBb2m+aabZQUyae/2iMx8m7vzISbeOJdlMZj1bSWIxrIGYschCnrzv/ymgWhZIXONdI9J4D5oH
0XpRCfyMvTJMuh9+0li/F3Rg5L+HHCsV4KXb92ztBsYFR8zPWgyWqARcNehOC7o7uZyg8rIaiM5W
RaJkpl2UjAJzXWILcn4I3CRfV4ILI83xWOQkyk2klmn74xQ3CeFtvp479g7/bGAQj3WQUWbzhJD0
4qVtbxsr8XXAsS4Y4bTFe7gqGfyAc4QjzhWegQ5tbsCTtLN+f430cVwqlvRrxXbeFfmEC9lA34Q1
ceUXfdl+fLTplS3qPk3Or3LtNeo6qAUm/ob12UbZtQqv7Kt1EGPz+WXl5amTWnleWJqSyIPWLn/m
lN457xcHO00gde1aStKriCp5GNSPZbl7Q6BXBXbKL2yTgqd4vbLCK+AqpFNeipwA9w7dxp4q2/By
3xBIlxblRY/33NJawiR56eVnnn1R3QIfaGid8Rj80GjXaM6isShzZP9D9/gysQrOMkTrIT/VD0WZ
avfBcJKv5qWIEwqaQK3nWclQs/aE/o2Nw7tWyPeElJEuo/Cl7x1iSqDQbq9YGXUWHA1Aq4XS/6eK
6055l2ZznaWqSBr2tEjcosdTxts2pkx+Ctj/NBLA+cD0dHbVKJ2v3iTqk/9M/GL0evDjt/7k2kw3
4Bk5baYBzO7ucYoA/g5zRyPJydkSJSmN7ovyDWcbh1k+rExxSU9oIloPBUv5HVVGuMtTqppC2Z+Y
uPsN2TeU4D7g1EG12yEXltmN10CYNM5+R6w8B1GkMDgKQ49KLbQ/13UyNJ95965wx3+UbI9+WOk9
BnUOtwVzMQlhHvcLae2D0CXlnZtiYAokktkUAvEgcErXUqUvWAigydtVO35ZQOmUQ/DHYFZGDUjv
sk7p98mssW2G9JmvpnPAONPJXNucXEnFOw1EmDDteP1l45bXK91Gr506wO2KfK1DCVcHn73BwBmu
R2+QgRyLl3kBxM4LJjkHvRGFu7eM0NvWJ6V8Jghb9utfBUYOz/07j4AaRQ379HD1R5Lj6M0MUwyn
bBrzxGDuXlRZwoyurHlnWZlr7uyGMBPuzSyPIG5K1yP12aYr/nee8DrCz2d5h3GOsVgl89RX2pKA
Kq2P3aoSIAnKFNdWeBhUIJ+TA7lopBXBDy0uQTsW6vcrk+YAPMQ/U3+CiuaOrcg53OvErbAdpSr4
bgJ8K0qj2unF4HQBhwA9g4A33jlX07/vK42LfoqyJNQRbFwnRDnWY/fgMYWa+l4C6tK11z5HPnKk
eCvycbanZNOEvh679XjFk5xTXPLo29tFGzo9MZUtYeOtKMX7Sxfw1yLbVUip2qq5V77xm80G4D3P
AUJFXI6d0TrC7uNCRsGqBftCjrYKPnYZA+4IuSmtsoYvK3oYkjWvzB7aZkdoC3CH0PrmgaOsb3aQ
EhYLhCwvrUGt953sfNkHzCiNtwDc8FWFxlOl0LxqB3GvtGYeaEKt8iaDXU21HZJ6sgxuwDigBMJu
+lRiuKoq9nQeistu6wvSFmZbgSovFjH+JbKm7n0eI4TS9EoktB5FyQibcZfwk3ICLQEqSTXjk5tt
mtygqZwd9trrdiFcEUISxbszvinvEydMbtdvic6vNnfl1xFD6OMOL4UT+uOkQUPR+uDN+Dwt3/1m
ksqZhG8YaW9Tm01qKjO942HyzjBpPgau8Ah2kv0X9P/YeiXcYEWUtSEAQSXnu65ld4eUePyYdUNa
mYKzHwTBCT89vwMpEl3ELpq7NIuxLy4Iht5Kf8ieArMsRagdMhU46gkfCB77hUQOT88PEvRiQ2Ef
yUm/mELxys07G4cbUa4FRvRjy9GnG/i1EWFaEODX/nJIa6Se1rHlxfQohG89qHqepFp0UoJDvLj4
CK8wY9Aee+PxT9+QKjDZnh2aA9zVj1dwGqCtIWneJzePoPGPO0oKACzODliTHpqPw6H2MW5eiifC
fQIHpZzwjgmlJH7DqL9N5nS+/O3m4/37hjL+N/P3Jy4DxEy527XR2d1cQFA3/aGfwW4pgJc+oAEp
DGAxhro5+nbA8mle+LfFqCc7SZfU1KYv3UNUYEWWreMke7PxewbeXln7SToeQzDFZdJYxvqLxb9o
KhBW4aCf4ms10Aea9IpSOVGNnVtad/u4SezKqdEjk1g8ndfOYxNw2LO291ZMvMLExQiT0Ym7Adve
eewNksYUPFIaITsQmdZlwlpXhKATskeYyv/RrG2TVyw7HDE9bYBhLF0YzJLJr/QDonE3WnSAJHeo
Y08RWrEcq6U9EkNxDsPswJCoStgyOCz7jlgDzfSem8du7NBPwTFaDcbaCsnKHLrEJ8dPPfof6Y/L
TVCD3OEt0AYfPt+fg48jxGX/RaRhCInZwNlr673+iGFnQcgHbL3yZO65vqf8PBu3yv29Nb2/0KgK
R2NR7DTPplQFBKBtcqXFTDGDhvgf0b4BAeVEX+MTFqbtRbagIhFgVmz4mu9BuPEy+q5Ywi395Yc1
/jgswulwLKnLwmc65pAL5LeIpINRtypkdERS4CSJOW/II/0UupNn1dX9MFsDUyL1bacAnshHC8JW
fc6DaH4iZqkNO3IslOIhzrliqDfaf4q4d+5PQkApRKHYDwv2YBNd8euWUsZWOIRGx43dIUlgk3aM
XY+tiXmZYAbpBWuN6Cgeb9ok7Glsx1tM5E3PlAROsi0Ppr17Pn5CzsDqrZMdjpwDLTJ+EFhVV4AK
64jar3eJ5V6SAzRxPtnGk5435bIR/h2l+BpoMxr1/DnbVGptVTdlIX+U2Y3liErJTCRz8s/DtQik
TAkRptAFpSxBlt+N00x/BUrsDwQ0tndVFV8+y0NFB4ukiFPxfZSDGhO7qqe/YllQWSMxUslhsOi3
6hhi0nEPVDPpDGUwItNSYKXGqRy3LKAIIYZr+OCtRuI+3vI/Px93p7Pp30tPDthnrYNYstUmW48x
bN3KBt+1K89YwkF9YzttCXlt0k8MWNGlIpkXbKlAyKZJMOCpfjHilVpbQl5H3I26+G5jvRnOOR++
tUs3n8UK5N+EjacyM3vP0u1e1nd4JfY3L5QCAlfLbWdoKD14Bq85fTKvL2IGdDi6I91zn5DVnVH5
MWoNDWhOWBfpzBbczjX6xyz1boHimGhMb3+P4gP5gSviGWc6vKT1vn+2DS34+pj0iCz+z7QQk/NP
RtdzAJyb6m082OtHK7v++7DjpoxaKOo7ICEnhNYCRq2XWRNz3kYKoCpHsrwqyhrtcmH0tQJg2ag4
Fm4THIJffS/uSATNNXNzOisVuaDjEnDk1yAeBL6VqKkNoLigEYuYLqb83fqONh+HQDH8ST1+Qts6
d5kO
`pragma protect end_protected
