// Amazon FPGA Hardware Development Kit
//
// Copyright 2016 Amazon.com, Inc. or its affiliates. All Rights Reserved.
//
// Licensed under the Amazon Software License (the "License"). You may not use
// this file except in compliance with the License. A copy of the License is
// located at
//
//    http://aws.amazon.com/asl/
//
// or in the "license" file accompanying this file. This file is distributed on
// an "AS IS" BASIS, WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, express or
// implied. See the License for the specific language governing permissions and
// limitations under the License.


`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Cc8WUvuxbRcmC7gvgCkNhTYvcxATjawVEir45SJG3WAFFxTTofKqX9sCqDBAE6IiJRaYh/MMJRjh
r4x7SVoMzJ8TwOlhwY95ru+KrxrpTXB7Pbw2cNSNHtuIF2g/hb2AKDsyEaUqQEuhVxg5FPyDVFge
/eWOXgOfBHAGMPBXQIrTjEXwJ87NcnMB/7tDxlqSzWltcf79aGGe/CV+A/4779/orCEAMr5UYMHj
3Vn4avqofWmGNw/sj52tBzSsfS7Ulu+HjiNQBbMoWAortSpZdTNbj0SvH9D5rC2C0mPIByUwlrjU
x1NzdGFe1FEcyYLRO92JtcucyH9M//yDGRGHiQ==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
UzyKnsQa7GNjyS48gwj4FCnQv0r9p/owVRUxr1KT50APEOzpggVAI3dxfzDTe33AKwVQkBdJNYaX
q2DdCGNRk5VJVV9GGrGxF3Xtp/R4TSJx2CHJi0xIrHnejwp/jWMz8yQbOCLJ5eIWTxGBy5B41kAJ
il9IjhBxdB6Psb/SDQY=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
PFRf2PFKraV7XyszIl7ff7SqtJCHrv1sxHDeBKpJycFT1Rw5ay+eT70WdDiJKP1OdJANjCS5D/d0
iFw3lHWSK60dOfJLahamuln58BYxeRrQKRu+0anRFPFWOmAiaX2wvSTusqHB4Zi85XSOc7mmqd7g
kFFxpBFvamqKHNDsbyU=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3248)
`pragma protect data_block
nhnA4QRxQ3OS/pFgwISNUFfc1e1F/pCec01kQGY79uLoIODwGIUB7YfMVibaHtL5xJU/niLVsLUo
rQgpMrRY1GbCSuA5bbIE6QDUYl1HCgB6+PimRoG5ji0ndTmoi4Hy8Pu8/91Q3yoMdLgx2fDOgyMk
sHgIHi1ORg7AlzLD4hqg68l5NlHL4A/f95zH4/x9vDfll6wOmoM/7KLCLkJl+brgNsnavoybp5C8
0JK1kVQ1qKu334wtPLMVv1lmctHqT7nHzpCn+2JrtNqM+rq2EtZvyjXq9qmEqnG4bmYcUrDYSG0A
nCJBeCy5N+iYDEvGb+Pn9o+qI/+6d0xf6ziErvbtkau37Ey0FZT3WnQokmS19oX6dfT+LpLzTiib
+I/HwLmotpDLVYfUI/jbncjOqpJBmaW0QBGYUrVhkFshfuzYlIRaw+nr7+WcZLl3JmQkGAXO4gy6
D2xcV5rqlGUaoC1ICcrXiAxYkyHOpMSBSfchs/wLFKYzpzZAo8I5wuSqZUS4qTGPY1imd+u6GdfX
m32Gg55jKXLI3sHYMeWpe3WHVvEvlEcP0Lty2rh+x3DbHivrnpliqZanR8gb4BeQfkfIK/EiqInM
X0esI00OuFZXeeG3/3Ll7gbM6Vst3zbjlcJ0oFQ97/ZVlStL2wMVCZqIpbReMgMIjWXWP9iOR0u4
LEKhbmMn1Rxp5fyANSzHqnlEjPxyxgmvIDy6+BokqdLSKoSJ+W91bYLSb35SiJOZ7Jgo+fZkGiC5
ify1s04fk5kZqxD2DtEQEYkr1I7/CDbsr6rrqYHy+3V1+I5qH42fS0ZZts1sZNWUnQmTSU++w5Jc
3BT/ltnIexi86amOnF1Xwfl9moDYUTfDuRbJTwVKKmcceNrAT5nVBhD+9ASX6t+wFWjMs3nVBdYC
WOefrNguyDh4o7ZxwL/sD5g+dWComHGMGS1iawL9TTF9OSsIVhGE617vp/fAOYganpTnmmdFbk5S
PwbLbFO6M+gL85AbfF9X6OUezHRcwtEXybn+HI982SM3x0QRznS12uvLwcF5bR8f8+ew3tO9v86O
tmqjKa7uBvmvRePD1okT3sRI56GT3W0K5TliGeEfHwJDXv2WV+ihGbj/MFWu1gOByYJBwNI3DFqy
BYvB2ryEQvdHK8LpIL4CKbU11drTb7a9o3646XAtzT355GoSXrqJRcqQ1OZWRkglzCHc+a5SZLhA
NJ5GWdSHBFs+S2lhgtbb3Syw4H7TFVPHT0KHZcMWg4d4lMVEJ16tFl+MrTHTZNc+iOhMMHw7SLT2
Bqr9T7Zyq4Z8DT5x0+vCRmaUCJ5f7R5Vqq3hXdUtEJtpWOHnIIjtFbEaUUIfd9S4iylIv4tw8/Dg
qpV5kRXxVc/0xsS60u2/m3zwI2Vw9mJq1WJ6YiBO7o6Ik9a0G2ZTKLPVctiXycDZB/z3ASI4f9wL
BZKoWF+e0VlqgMsda/+O+i8Y+dAMHu2oMvyS7zIZLjvVH3Ry5JWNUAjLPO6WAn1cTqk+/6wbYA+b
BXclkTOVYNKgR+oeJH+UBbdaLo1rF+l2fQ2HbbibkgznI3z7vUgPq6RGoYve1uU/ZZqnVuvNichb
70JOkJ5LCaRzet+rELF76GTwjGFnyQjQb2KQ6XnCXKFoN9X3pJ9UfJ7fBB2uoxWQB54rwRU0807d
ZineT+9NlEKC2ccalP1pLOWL4N20VAAGEb+fsj8uYw165TfnG3i1u9HkF9XYjcv09P9+9DjYzHhL
Ve11tyB1O4Ba2zpETuFGB74QtgUe+NC5KVKi7YKRRHdjTS2hvjbn0wOafb3mjF9lJXVPaJGBMXpe
pOrR3tbdUsORgGoL3PSXBM9hSQDErz0d8rNJYzt0rmXU3E4U4k/j02V1PoRYo/MqUmjjasVRde37
Iru8DRA1+vJZMLkmh3fWQqhfbo65siiojLX/8hsnrPAYAD34e7B/dgKmhDqSyQqbbXED1ijsBKWO
5Ywk6BRPqeHTtRdU1TfmnQawJSzFqs/OyL7sYsPOevO4rmQ/g8RIIcmao5N2xaNdIKut24nnT2yD
t+eC2UJwrhi2w/Y4b3kN05H2njjp7OV8pgksJMJPyfMg+FU5camuvAkj07P2RfCAj7EpjwUpizp3
VIsXzE/MNV4K0C/kxlv+i2r/OnYxZZ+xWP+nK4X1RuOBNTbmtSw4pyfRMg4kcCTKiyV+02qbcdd4
aESgMD0HkR0RKSwB8l8qa76bANxV8EkeDs5hwa/O/wGrsqYnDnuonYQ8BQYUYhUd6AnQVAD19sAH
kTpaVLc+Xq2k39ZUlbVIUj2wH+TKdmVep1KKKIPUuBopAS5lUT8f/rc5ZlovbJIo/xFNXO0FOvPn
FIb2epQyqGqtHuJXszqrGZ+nK/Qsv7rZijku3mff2PbFYUpf96GM9B2Qh4bG7QPnjwqDEVeuCR9C
kW3/OBfmRhSphx3xxvRbEYM/oChgPGC9VIWVEIgaEjGsAqvoQU7JPuXXtESqGNVlQaHSSiEWiTwj
br+B/iCcAzAtPFG6qIqI4+EJLvTylVDRhXP/r3iK0lWNShQQIOPQk0bY5MGl9pKXsErC4oY1aMdr
joRYvs29UDRE4grB8J0RqMmDjDeAA8x56sk6mOa/smtufjQxKfhlCjHQXJvRTd8tyScGZMaJSvCl
UR5tQhlJlQBfZYMyMLtySIga35mfe7HwLvqhVRhJIYU0zZl6kfTfd+Nd/sCQuhCsT/8alvrV5+IW
iemU3AAIeRnD7OnSmJiwsFJgx6VDsUsPf+z9GynfheYsL7swpdU7mlBqnGQ3dS3h0oX7+BtJFR+u
IhjxepWjH2/ncSoC9bDaw32F3T0scA9HGLyHFrFmJx23H7QyADmwTVSaHOFiJpbf8Y0xM11JBoWf
bKs89hYMYKLNtCdi8hTcv2YsZNlYfESF1jPT9TKOUX6xeko756asCGQHBcnp8S/XC/g5v1L/OPN3
0iTctaXtEUJiranEN6ozjMV+gxCi7/75FtufsKWgoAhemXjbKI7G7Upk8TRI+jP+bNGTbv6y8pTv
V4ufjq9aPcbns9PDhUO8qALGlDIMr5hD90ZTk03kfYEvsb/2hlieALEWr8vJTU/wOj0orC2u64O9
fKPMxESq45aDeBecfaEqycDr93ERVgyQ03+v/Z5q01Wr1sVtg/iQD/uB6mQjWFhJAJyoVb/SbpjT
mlqJVBSMHCQXvKINqjSbfz6iw+hNU5wvs+Kre0+ULAYfuJG0sX8FHKnWBJlQ/AwIkzWSwoqJj/fZ
VNBjA1GvdF+LR80uRlOfgpuvMNekwSIsVKzHqXXILTFXSmlKJG0N53dXxYMVNmXXd8xUrmYVkH9Q
7ZkJ7OOQ28epQdeO/AlINlwXAWdgnJMRYrSqC64FLXZBoDW32sJ//pS1w8sQ5nrM0lDLtNMOKjMG
AUFqaDKuyRAhfEPUc2/FssunNI9I7yDFXFNESjMgV5dMiv8RVPx2wjiSI/lmftwRwrmc8cY1FqqV
dmvS8Fo6/bzv+HySbRx8G2w1TDRUpjICUTCdBUBXhwtgwNa4p+kuV5OpM1lnq6uQD0f7lA0t5td2
kgHplgbWQwtr5NjNIUIlHGMAqaA0dhGhkeCiryv0ARUsbEWzFzVniP+0SqIgbZqKkIIsD+KOHdEh
D0C8xCz5qoBtQB+OE90AdyQPmuWjYAAseapA1EKGcrU8CX5aWtlc9onJnzEGpkIuuDtlBEzDynr0
FbIHtdb3mYzBogp+9XjwmRYsmpG+u04uVbD0zoto/+AuAdVC2hRHpVoN9oduBqra2A6Wtxn/CFZp
78z+fG+jlPzXBEOUzHTj5PH+kwifG1pnswi4vcdHf0wotNkkvP9uIiF7h9dcHaXCkiTrp2Ymy35+
BHQdczNffQFGTSpUpd8vIrDZIJrdB9+f+ydpK8gpxfS7C7Aa42DSrji/LkPr8DmlQDesiQX13Ksa
d6bUc9JyCfjf82T7FzSLtyzHDGXWemEP9VeU07g0r4qkoVLFAfSwPqtgL8o5TgL81uQFPMPKZnnO
3mUQktx5jruVcF/2ulx3FDl7BYoX9oYP0+4wPHoC26VjC9E6WJA+sXtWVZ2cAymO/SxYRNRlZMLA
sd+I8J7QRT06u2RJBa13jjyMoL0kGcZ3Vsdl/Yv6sEikOIp+W72k06OPuLpWwR7EIX061EEtNOUl
uU6E3OKbZkoLWaKwSQ3tISiR6d78/5jhJsHhNgjoKGZfHJ6WuBEA+1OfM3PXYVvIXttGfnH00aGH
6ZFwm5KT6TggK77hW/dvr5LEIhY2uRDB0TWldhIzL3xEq74kbVKibRhedXun66plZVsDbYySQWg=
`pragma protect end_protected
