// Amazon FPGA Hardware Development Kit
//
// Copyright 2016 Amazon.com, Inc. or its affiliates. All Rights Reserved.
//
// Licensed under the Amazon Software License (the "License"). You may not use
// this file except in compliance with the License. A copy of the License is
// located at
//
//    http://aws.amazon.com/asl/
//
// or in the "license" file accompanying this file. This file is distributed on
// an "AS IS" BASIS, WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, express or
// implied. See the License for the specific language governing permissions and
// limitations under the License.

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
lOcjuXbKbpAAW3Jkjca1YSn8tMN5HWCsBBDdSzVURUzdkiVKfkpuWLYRJHvoXE8/zZWmn1p06YkB
V7yDZR88oS0PoiopAROHWHUxGU4a4e1wATtqwQNsC3HR+w09pBPSehorSz0QlDB7ylbpaMbQD3qe
o8yMHKUDuhjQCzcor7eR2dGThAtFXJ1ISgD1bW5GcDgB/V4R72IOu35p+4bqITk6w7Pcpe/u6llt
8wpsSTeh33NYc5+tos8h6SJKqwCN0trOyT27wy2soI84DDFYrTRqFiMf6LS8jCzRnYBz8vrAOoY3
aeEVStXKO5jTSUSa6jevObuIc9/kjBz7P1cTgg==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
YjkyAQ7p7nNnPawRGh/i89LENXvli+N7S7q9VHaMJI+2rTyAMw54tpuoDzs+UEGH4MhYejzinDVD
Gr+rh9wVIRRlNmN7P7QENUZRkjuwItzlnTvIm/rKJbCVZ1kjd/MKGasLE7fs9gUZtJRvGcfxYpYE
KNamIQytSk+XfL0s8OE=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
SNgV9MNGybYhYrNaGpDFBPXc4aDKRl4tHOqbiaxv5ESqOVnFoq4pxGQV8zE4/rwUft9JEdEDVpeR
JIzEv/JyCP9ypwgw6QZ2f9QEIgmRKdZVptEow+X13huxNh+iIPTavxejZYSM1iJaYos2rQ3UADXG
uU6lwqxHs524RCoLoFU=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3056)
`pragma protect data_block
VypC1CLWG9eVXucQ4KNSYm4eCmXp038Ak1Zb6G26lm2hTsJOMahhuD8ccSJJRHcvTS8fAKVq1Fn/
cgT2+V6cvllrCRimwTqUbFTXIt7Ta+egWmejWE23YTYkiduQiU4izn4CqN/vxF6J4VZWRgjGo8VF
iJPBZI85pvcthzDj8TLBjv2/j8pq8D5jjGoXMMXnhbXMOJSPystSy6n5SzRxmp3+FefoNWeIC7OS
bZxmzmvWS3rtSq7LoVkjmQnSZbyNhSZjQj6oYWyafaqyrfjVAQRaW3ejFjQLR5Gc5nKXYSn9ytH4
fO8wpdmpabEuh6UeDoA3orEDVCqsp4vsH6lx5E+WGbowDgb59Pg+l8q+i6zfnr26qKAWTZREm0L9
6INoLIxL0Fm9T3mu2boD1xuk9Pd9k2/UNPZ7A0Az/PBdIliwbjcveTF/c3zh7ISvye22fN+3BiSS
FWXA+2WG7J77Fpek2xc923Az+Uur92sRGXmY3eNNA4IA8k08Epi6ENDI67sCbHwlMQ7eZcoTNPiN
+rsoE88hmajGequyV8GCMAW6FIqXZYbElgrcVF0cYUrLzbsRegZRXUgjhBRC5cU8ezIu5FFatV40
yIxrSDRK1DNlaIg3BGf9J0/x0GVw2sZ7FlEoRSqv24VkrV97753zR4EatCsiaaLh1cUlj9MQ7N38
MJ7z5R7SEOwYiga1mZNEgLtZB/MXXswmUFupZehC1TZue5gzozav0DIY4bWg38rSnbDr9K41zQXn
B6o9kRwNyTcZc1GE6BP5rBvUrx5h1O+dDuwNjV1Vb6zF9xfXia632xVd/LBSSwoj/KIn+TxuH+/b
2Lo4eakcEARcnW1LxYh+QL4Gh0ewLtnnNuKrZ0kRqlZVbP9Tc1FS4Umq5e5gJx376cwLcSQoKz8x
ApycP0mtMDpycOmMIM0oPM2MAwVU0YUnXOByvDykq8eGAFhb/sgV4rizaXpYPgmXnhl8o+eaXHla
HivLoRkTQYEn0/mFaJyRdcbjNg1/r0afQLC/suql/AzMF0Y5p9H6DAiOHdoPZKux449HTnQ90KJz
7vm+NGtJk9hsZFUQYG1luV4BXmSkHi03hgU9LzxBNFOcKiwS+ewO86FyNb3GkmlM0YyKcwI45eR6
IPz/o0cTQMpz4sSjjzsqbZGtRNYsIwdCUrpPW9MWAByMi4uHCtzE7u9hOv3axq2Ao0PC7Vd0kdCl
b/SC6Kk4wkrYUvIG+3DJJPr7wybS4IpcJBCTsWKrU/TBCfaoP1iuATVklyO89rtxEH3OiOtDuYuU
vkcOG2R5gRT3wgHhhZnudbV9s6ZMNwbEfUGyWhF0/HKeVG8MKBVPnslv7Mgp2lR4fS66ufKdnXr2
sT+VHf/Ksu6WPrFMcHa39j8fXzJcdcb1GjoAPVpJw6EoIy6rURu/2keyeohKyxJ79zeaWKAPJyWE
CFLnStB5s2lXUn5yFU8WffYy0dp6kUa7UnViB82AHnnfaUHip8GzmySHiIRERrbl+8/eo5+ygF0t
/tNV0DFfwD0On0EFPUxf3gKoCzxSTXp6EEhyC3Z51hW2nRb5MiqLjfrYnzxUKh4qYE7OsZTko5Np
xgv5FZN/Z2EeZrP5wu9jd58gCozXJmDl19jXi8YZ2ajH7h3O8Cl0uY5TQmUcS/9pxYZ+LKdmVo8m
sBXTlv4SqyinHuVw2ZOfEU5WIaJhRt6REtU15oMQLQprQCD9ZHy987K6pUUuIKlb28adZAhCcT56
iM6IIBSegkdwUIgFrYCjggBCa2bYdgdWZN051CNfZlNnp6PyvXJ1TfCTxn2b4KbuD/XvNqzXN5xh
YwmFljh25TnKXYEmuG0CitCj5oQ+7SDQNxtl9zngcU3qMqOWW+2FMGCYsABWOseeye+srRCqYHSt
piLuCT3v/ukJzVwyAT2Dp5abQQIKcIFFxjTmLbBgiExf3nSX/y0skFzBcNDN41VOVsAOKXlETaxd
KU/8wyQN2OE89Ve8qiLtEviS1f4WQ9qWrTAeqfm0qX9TrEeztm5Qy76zkj15cY4NT9++zJDKXoYq
4y5rNpffIbnUm4px/pofHT/JJd0KjnijD8+r7p0FWyQYrScYoX8HddTQvkVIlDTgzpxgQKTJ9ipv
MKW+OHF4gl7NS+DuLWRdBTW1i8WF6MxILO8mYseLQkbJcx87K2DRMBORwte0p2loQ9gLBysVE23A
VeHoTNtIAnaI9QMj4kk3pTxcos2GWKy+CwcJigKtvh/N/61+2wSFbBXUpeUjcnY8j4o99HD+wQnU
O61KiIyWb0xeMZus3DA0NAJ0kqTZQ7UUPqj5+teZ/q9BWpdIx8aDy2WzQ0rAOGZXR3Quj81Os1Qr
75OIPqLS0V0HYS6bLoBhZsP3EmA4wjMvwbALmwWdDBWZAwR9jHItnE/uel9vhZ9uwxukbL8f5FBa
2LLLF6DN/iGQrozaFxp4bm5gzri2hAtZbiVyNLNqioipNZ0qGzmU+FU+GduQF+a9qcijLf9kEse4
5AoBzIKW6J3vj/OO4+dBlFCjrwsOQ9D1qKmg8hK6yZ0un5wXPjBS+aDz7LZ6YESozd0nyxKOK1lC
VGRJ9fDd92KjZLgIUj9DcPYMsrD6THAF/hte9JmCzFg/PeSmYdBy4vQBiltba1LDBl0go9DokCDV
bGGstyteA7DPANG9guuU1TR/VfmC2A1wXtwUOM/uZtC4//K79Ij2ehY9jmKBUIDWfjqwlkSH2g4b
FaK5F51+KEnN9pg15p1VkF7MdN0gMJk5Jw0qUghVbeIg9hzl+gS8XP6svY19qf6C+DmOA3H4H8tl
DmlKg4fyDBuV8lWEpRjitPbxuMhdrJ8tdYk3lcAtAJDBJvrBch+43z7C15lnqE5tUMAg758jOnHi
FGfG7Q5EsHvxQLTRueIQSCQDzK4L3grmo7gRkmGqZVCy+YQVP58fBjNQ2fFPcwAeSqQbc/7r8dVT
kagVVg7iAOcgu2DhoNDXa1h8CEROwgdSLC25MV8bw+cYGeDRbtvqma1oterp3UxrfrluAZQUbnHD
hw0voUOvo6k/xxfSEjw+YcjC1ZiIu+Zh57E/sPeX8LFz9WH3FO3IxvGsLKDdfY2dtUYJQ4s1GPpn
nvXwDh/7jnIhWzQYbh4ggPOCl0ZTjrTcVlE1UF0iQ5jZVyaN4OPS7YyvZYdB51u1hiUYX/9ny27Q
g5P/7tFHCJ2Pc7Lk5b1bbQr+E2AWsTWQpzwYU8S3zF6nNgf1OG+u3BCCDoPNTUNtNkcimOHC6xbj
CtQBXm/FKeG1rMXqqxdK6v2pftH9p213xFREMFy4e4GzOMiIEtdmj25RY3TG/p/6eauW+M56Epsx
QUHleZAAd9XPZd4TA6cAhgC+/6K1eUO4Jnt9wZUAqRNyT4OWva36iI3Ca1SDYwaxPzqw/14ui3g8
L+1H+wWOyOg6yAEYhitnDcLCH14zHG7EJiKj6txRMkjwGDHETMY2zl5BAkBmGqop+3spz5zyC0GW
2cmUUpCWVnFFCr6Y+Rx7nO/zSLVM+ww6cNksW9mMlPPmmsfochR+Who3GUNeGgWMO8xQnvrByjJP
hNLN8y4Z3OfEEVWiwJ6Owc9NFylWRbVwQGBv5fVOKt1laQ88Ylh+e6f7EGNE61uHCwgRABLOj1Qs
nGjgxf7INtLHO9/HksBvflA5irDezvDPyQFTzR7ZaBZJDVgRhd9kZF+8z3veFMZ5zN4QVCvEsVsq
OOpChPGPSnc7B2Gi9HchyBxRIs2Xv/WfxNUseKniPAQOMo0ER5tnBLUT3W1VVHj6k/EJD4f2Eri/
WVhdTL1du+QeUr4dbjP+wMG3g6g4I3NAM1hiFN3K7miO7VIJporzwXmULIn3Alz7qU0aAuK7f9Wt
LJpMUrQjT7KFQpgwBscuuNneMyIpc1ptZ1S7Bx0abAcinYfQbli6r2Zi7C2M/FBoukKcyCOVMElW
Nb3jZOFTXIfGYr4CkM9Op0J1xKRE/NlGBW9KAjBKsFnKAbmgAlKU0WPbCRBkBKVDLP3TjUR2vxKj
6MHFib+lecUC40rr65CpD7LWRGXhKHBcuw0S/4Pab8BWFRA=
`pragma protect end_protected
