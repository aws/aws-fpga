`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
imULVMT9sTBrgQv8myPwYgI3DVRNOqwvOOQykGcUKMpx3Sq3nWW7NooxD5OGXzqcemx0NbjD71sy
UG7hoalSSL81FR8Zk0XCgE/0gXGENW0S2kV/0QZ9wFArGlvj7ccPQ4qde+165Idma4Q8yTOhlJdg
29K+Bz1OUSx4YGF3nFzlLLhOOYxLdOzcaHidN5OIUKdlckvbAznMInTFN0I45KeLiDmTPpHOhjlA
a/fJVdb/zT3j7sr09UrwAGG6GY9p4T1B604VDYIE2V8EUp2xdjY6daadXuLM2yn9vNN19yatq1d7
Hk+Y9PEXG/HjUSyphcNbwfn/wIWtcxBT/8eVWA==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
pjQUceqJ+v0suzO7zUt891DCrei0A6bsSDr4UtP3lKTaHTqJ94d3dbklxl+BnTDfenI7XaHahdxl
SFMwoZG5cVgbkaeTe+CKepaWfiLS3EoQ6xvBvN7NI8L8Z2lUWTLwedaZcaAOU3NRN+/gU3m6HogB
33nSfAh1sUK80ECSge4=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
BFBJi8i7Eq2F8xNxJOeiQdbDUN2pSuAj5h83Xq0wQVvhA/UmneNf3vDs86IPznuNEqVfrLtngw9u
MHfp5RVqj/u1IWEV3qHI9ecqGp/fQ54F16JvJgfQ22ovsVWAm8D3NI/rl8Yjt+qYpDgSPFhgsHT5
D8nXgruJ1sn2J6npr2E=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2160)
`pragma protect data_block
vmBAbK4ZRfOj7nBFhvkrnwN2dbGsVxw8chJlTz46cNQjseDMrsPglhWxy3UxKoGrrewUOGDMbLkE
oVN9TZv0Pjrf8sOGYPMJ1RHotunQr7bh6UFP3jDrfOjek67xh8GuEljGr5/0kBHjc+HJeyYajAWt
U0ftX0Eulv6Dj/1NsSKd2qsfWo+2F2IbOg5Tp82/ArrlfSa1Yv+0XWndGoqine0/TZOjMHc6HkyG
GLwFg63i6Za6LUxbZi9tpmSyJPglkFf6ZHv8jC3p8FQzI5hemTtCUcqAnl6trkIPRgT/CgAVR5k3
0CsMpjGgsZRVlqwx/QKlf+HN6fs9ijfqYPk/lWu5VI9ZOC1oo9NMct02ABjhj9XFDYKje2lVz15n
nYd1C2G6GjA+BU4qr11keVEo076djQ8ZqJztKfrGCyMqofKyjGS/m2KAfz2LBmLuOe3yUVL6AVAO
RRWWPzTb3F5C6yK+Ob79OfBLuMQdPPoo/y2kQHwoQIc3exzy6ciS6zNUPAG+Lz723MMGAZAA/SVA
KiFavakbFjvUudF0eQ+yaEMRcg5F15njjXdEnYK3/hJZkva7BM9js2YowcsYwJfRQZrrkAlnpXiu
4FdcFoYb600wMqlVdo3N8qBy8hHhnbnWpaKixSl/02+cMwp7CKyvYUPhHZmgJgpb4YFxLf1WumFn
r3zBLSiZwbUOVS/0H8MWOCgIsZzTV42IHaIOA9ZT6CwWPz9LdVzI25oYBm7EDme+31gzHiTtAO8T
C4CHeOCVRELbVGv2a6/PmNdvGMrkl8gFrY80TejjzXzzAXkOt0AWpJZK1Q0VMBax5/dqjPA5l1nT
6RzB2InnofduEuUDNw6v0FPh5q74ixmB3SsGSRDjg0lu8loGYuDhQsq2miG71uszH35q4PK42VGV
6xn5KLrXC5qdnLdmYUCOOyzTL8P1necaVTKs/uo2EjwOA6QlxczYSx/TGLf3YgUZ+A9VtjnDF9Fo
05WS1fgSvSL5dtZvcH1rCjWyDkOm7cSmiZ+2U4tXIV06YjwXpWUBaEPkBwo3SLlxP94bjvdHa5FX
Jc+HGnj6ZjFRZsI2nPKDc9ri3flxWbpLeAlaFx1jUtCBkPK0F6UsUWMslI76EU6T23zhXwGXT7UH
/+mJjJb4bhdjuotv0KLMelBq+TDykLCLZFqCySFpheOXA8Zn/7d4AfcbdqN9Mqb7yA3IYm08ZbyC
KyXwjzC/kdkz7qbip5xPAP0qKb+v5wOTI/Qv/OwUdKV8KOhH8d79106HM3PpFr/0kUhMqJAJveOf
Czl7FliHBrPsy12xu3xzU/us26z2oLzIYhqtdr2mbUUQS8Yb6MmkXQcPbR7VYUJdc/MYP0Q1J3Wp
olj1/lZuwViJpI+9Byclw8GlNCbZoGjpxEOjPgdaBvRa2Nw+sWelTFGkjP3wR/Z15fSh1oHhwHiE
X5Ft+K2wHG5+BgIjhQNIfZSN3ogPbW7MXvC2/s6YJ1Swq0r0eouuNWsAosbIGO6tIzYTEHXNclWb
oCF7y+qT9NtCpUMbW7fHZtS/Upy8+s1IJFaHKh1G0l5kSApM+stfnP2SPeW9/o5Baj/m+PR0o+PN
eJbkd1fgD880dAs/aiH/57s9suhYnSBWPqrpJVNu6wriYRxJpdrBKK4ZODFAxqI3obC3FdsleLex
HrE7g8guQf6GJRI4kz2STvhIbirdYPQmDnqYkMxhPL+9kDxuMU0VCxyYB7eIpDNv7bxTPNjkFHzw
wSGil2gv52MFGZdV1Ao9MKd7A74w/IQAXBeVC4QT5nRwbQeNgOscGyMvsxPedcjmOeojT+6kXiM2
hNk9MxUmG3OrWgV0fTHPeP7qxNdnt0bv8A38JmvDz5eLp7mtxZ9AXKMuwHMJZf4gTQ1M69Yy/uTI
+v27dd0ym/+d3hC4Hn7ZyYt9e8yHXDXXijYD6BWQkfw2PL0PRUjGPJtBVDFUhAB9oKvIMYzDr/bc
C8T6E+iS3bmEgeu7avz8LjeYlo6cM1UTBhKzz2D8L/AWBTzwlQgOuVblx00tO57ojkHw8LgAvsvu
VkGALVrx7wJJpPfy+Lpgzo5pn20WRTX9f8Djot5k5EryotoGwi1yIUFvkx5USsegkuE/V/spI1GS
ev7OFujHPrC8TrE47EtpyE6+WCjAR5TgQy0OiUhMboQglLyt50YHPx3vR/FkE7vmTIynCXe60uDf
d51UDBhIKJbpqlezTeB/RpHkinN/fZLNPNy2/KoNrRdAuFRX/XieKFz/mTG/JkE7dYtEgagl6rRK
600J2Bz5mZ/9P/RQOyXOA9ZTeXBlR/zQCaR09bliJikIRyHcXg+4KnNBc19Ecwan9WJblxCNbNjE
2hRXExmcDCy5arOsJofpuCTS0q50IOb6LJllXd+A1VtdAB8yOH3LXDB7TxDLZzTrK2liI5hQ4xbk
e8Bf5tJGcNlm9kc9AWmEMoOzWJONPJCwlv8QTPcO890a+9GGafwsLTq7hGie2xtifFJ5Yw3SBUTK
0BNqak8WAMy2N+uS1QGY3AJP2tS3KVCp2KLIRjYAj8Qk+WIcc+vXQkvX90UPvAsgM0aF8AEOzIk3
ub/OUm+xWm/OIQr4cfaH+RbYCZ85KQMQsEEkzm6v1PzL8ghZpsyKBW+n0mx6uWZFYT1N5jPRkbBX
Y/B7n4lqRrJkMdbnte567Rn3+MmmqMVDVxdD1HDMyeoVYeb/SOpgKaj7CUIe8mbZHx49wadTxqTD
doKzQqzuSQJ8yUjJ0oUM5eZ8N4AiWb+nvfp/JEPk8JHjsLOhvIiqfhBWFC2ps1oAg5fcPaeliYMo
DCKImfzJ56Q9oPRu05FdhT9IVFkxf1Xhse7MWds2h2UNgJ0oPeBS9Pshhows8V8XNLBT
`pragma protect end_protected
