`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
E8iQRlzGr9F/g6co9M+VkxHyP1M7l/1wle92uLbT9yEQMFAG72az5nzEDxQQ0FfYOdnHgZGl2dvD
NljKsz0+Bdpqbiu3TPmVLllssjwGqD2s1ATREJiBmQLOv70A8RF07NQTS1Niq8BSl1M0pBg6rDSR
HXVcjlcuoOPTnQ9a7O19Otbf7UYXsYeR/mMyO3nLwK1JbUTHt4O4tfWcEyJd/Y8vJdgodQfcxTd4
RZuWNckt5YAtvDclsmVDVB9FjPix1k3vfHgqFP5HSHSPT55pgpw7duz08wM6G/6uhEwWr5aAKVx+
faO3asiF9yBHteqBn+VpCo1MdHKadmeTYS+6rQ==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
W8UcGY/zshtQjFqhQ7VLzNHqDvwypvYPntCNREWoHEqFdnrx0TUPKhpCb+aiiPOvBLwVZXS7AaEO
/8u9JL+kMtZVrBQgPmxMitQcMFiRYcMUR+FQqAyAnZD3ic4zfOyswE7OlrA09GlCj5j6eDQsFojA
SdTkGJnfTPnoGBut+Dw=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
QnLFrmPFJ0dsvoy5pX1DXGiUHgIjSkThk2C3SGkHUrjqPaFA1rnJfcfVINlSuPL8G2yTP/5rc+ii
LTQmrD95/3v43ngjp7xkKdZt1BKsYmSiE7nFM+Vx0J8r1nA/c14MNf26tek9yEYM2iwAfYvvlIeF
w3NCGK9YgPIjqXXdi/0=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2720)
`pragma protect data_block
vSNQtwnfuKeYoosRThCcDR76joQ/0/zeS89InGhh2Ykaq7HDy0dWr3JxPBjzk90Uz+9g58bdRjFH
k+MgEWZF9+W+dnS3na4SYKxDqhphjzCeWduBuQSs/85JuhLjD/lWlS8JxsrukXwZID+n8QS0m9pi
TU7BXHFUxoQTj3dWRdlK6fmcuWKDVI4YAl3k9rdvkE+GqMuAcwTqIO4505VkQyBEb/x1ntJXRmlm
ODQvETWYHwEYMnvfJBKajU6db4y9PGuCVk0TVGOzlTMuzL77en2q0IPEcHaxUsbabIYEAPOEH01c
lxvTm+u+bBuEgVwM3NMWxHNBQ1Nu54z8+EDHacF+nWXf8Ja13LoMQTkYl+k6lhTK+rogySuWl1ek
Yy27pXARPW2bOT/6lQEJPBK3PcK81DhmmJbGZtw+dH5jflPMJ9CMFIS5cVYHP9QjP2u/Mh29ev7/
n+VJguLQ+ndhnuZi7sc9ZRiXR/NPXHSRemYcH0ljJEN7z8aEHvFeeTE8IRFzOsu9CqmGvLpqtitI
Dj0geBLSQ9Gl8eGNmnlBkfXkFiNt55QcSG+au96Iv10a/WqH1dW3UwEuWUnhcdUsOTmfvyirxsvH
/O0Zk0TeUdDiaC1QA27tBl8gEMAa9rZMsdaaodZ6bDneGljijtb+XicMnJ4gZXXgnkY0gz4IfHaw
4r3thfcVziwbVuOqyPV2nGJUeowL9kIKhDqnWAcMtmvR3PRafg4GCgdvsGv6kUQqWAam4CZqAYz+
0EzwaxvxPDicuMI9CRvBPrXTHtcaiiMGYlpFhsDLVLik6k97Vj7F9cM+mCUXvBvJH1jsg29BVl9T
7Iz1Eg2GXnQfjAZyCKIx8uV0XBkNHv+dmvlFk3K1GYAD/qAfUZWbkm2ZxZHRoyxjhZ0czgrTNiJb
4Q2LtyWQelQNLhdalK5KDWCzzvpw5owCrMuVXCLA8qdkp4cv6eMgmY0f5YCWhFwPfwlwZukTjl1R
A9Icyz8ndmoOxYJ1rOQ3OKK6/4kdGhCmWxfRY2+9XvppFjuJzxQklAQlRyCFSLsf7dTOPLG+hTWR
AMjCc39sorgCB3LnoX0p2wI60CBkQ/0Hgg3fMbUPj2v/doRjA9Gl1Pyo59vsw184kOOyyNZCNyuN
QzqbRA1tcl+GBwVkJw0T4EQPtxZInpse1RftUAA2qh551GU6nD3nlxDIbwaZS1O+Pbbn/O/eTZqk
b4+uroG24eSpteOR+GlugBcdy4GJGhQW8s0t2DRDk0hOVdW75oogU6q7a1IOiigE0A2kwvtonDjb
Ffm5ApgDA66067JUks4BRvcmPa69bEo7FJsjeViGPTzSgbAdj9pECmtNdu8L7exvbg6kO62FSysK
qbd3zFYV+vIiW7Pfa3c1CGhn/M5aEUAOkfxCIwV61mCwFEohQTQbty3jW1VDEmndQtxgaAI1nUGs
Iehz+Wb10HoyduscCTqSQ0JJpgmoZMoO0oyoBBRP06ZlEKXp3J+cEXXsCB2yz20p/QJ7AekKdNyR
7qdicb7wr1KwyMXsNXPqTqSVja+ygIs7NGnqUvWw1+M0MlLiKhNm0icKMNrv0KATBNbXqjYCyA3W
HUFo3nisFg+9QytH+Z8olYj6vXEMG0PxHpVfvJ1EsnGte5uNn8XDdZR4fJZSJms8Em3xdKBCI6+m
GoMfR9/dXni9aDfuvV6xVtTvPwdOnS7PAsltj0gCfAkHtEeGHr2gwVPlSG2QN6r4qRHYR29xK54G
GA0mOBPzInEjPqSxaN6K5qMo8zSbT9UvMJ7B34BsOqsuzDCT0SYbR2gMVUHa5NH5XvfwCuDpJWHC
DohdnI0lVCoqWIb1PX+jayY29+56QCPC2mIe2CqhlWpj9BUqE2f9p8o2Yhkhg4K7OVsVw5tsOwDY
didheS7sYQVWmzLfDtDVL4tYZIPzk0SzIw98L6Wce+XkWnS2Q/IIhGSHWdhwj+GfynZR3u2Ljc4Z
THEIySXINgH3LmDZLzwzI25J2qr2vaNdya4MLE7P9fczCqUm9UekRuJgoNTO4Xp6WebxJp2noE1n
LRvwIVpgqjhA4qeIlHZEpZSLqCfP2NjJKfpG9APLxmDMPGlkYMYIaF24tiA+sOIzUi80tDYrAq9G
VsQCXej0n49AQDzxjBqJM3SoXpsWZpSOAfQwwtYIwfr2GT30IG9eEN6eGbZQVLNms/B1Hg6E10gI
6qKG19j7yyiMSitZZUtRm/+IO6Q9wZ9zxpEbXC14hwcDnTUrUuvW26MCZZlfoX3bJH4sQVd5eCxp
uZb8RS2YgYmDsn5gcBQYnOt7AGbTf6KwRCn2LKwjNTajxFyIhX3d6HzL0WWF6aEmlYsB+X9IMHEK
sl2Keo8//4+pZ7yvLE7bcTl5CpBw3xTF4fB8eRD4nblomRfhh1G7EOT21To2ncJlfRb8AJijFwT4
HcgvcEtBWatavP+wH1nSHf+Qkaf3UAK9gyX0dLFUTb+rz/O4kq7aW7toNPQcOErs+EU5WAqrgxs6
paoHlacYAMOt8qCNQ+CFKG0DBEXebAxtxX4AtPTsA1K6YFyD/UjJP52Q3nvx3qtoCbIT+Icnqz10
zAdFjpwCMlm5aKLLSjboF9EpaDXzsomaavmr4xNiYm2H4cEI17z02elKs/xiapacAt8QYAh/QFnJ
ZsnDMlwzvDpVVE30sMAVPqBHliYcV9jY6AC3JzIQLwgJdm+DDbsJ+8RT8sf5IQohcr64GBWIOhW1
LswRKesaHLUDWGD8e76F1Pwe0dIjwt2qIz+1KKq1mQWnZku/HZhcMq4YRgAWxTzu1TBPDxObw8Zc
JxcseZwmcXyKufMjq0gOAMeeqnAiavwoytYA+KFHE8pkrJgdk6YVNSXB6uHQadd2ABs4pGVkIY5x
vXg8da/OpyBWdnzb+jDAOduzf5actJqCQisvUDHnjftL4M47h195U0JyU5yCCPHrHU7LE18ypNZw
bcqNtTrFpJMh7c9QKjnwgOW7/9ORXi1pqeLrqbHcXwL3qKfdSpcDjbVRKVHr8A6Zqacy9tEknlDa
H1mDQfJKda1KG4hdIKuY8oFDHLt27oeZIHStRydjR9EBhx251PgU7IQQPlKC8QT0pmyxJ4BP+gIN
ueNl358SBKNqaWBwRwkm96EZJSpIr1BuEB5rGJonGRXQraGTAl4AiwJm7fSRLW5QwyCtvTtIGw2y
RZtghkCTELVsN41rVOnuqGE/fnKklLhfs0sC8qXc7wAba53c6GWxdqwfDX3tl9HC8vqBp/boRM7L
o+NtfxeUVBgw2wSSkREb7tfJTmwcHbGKrsO92AWfG9Slse/fSytDJ8K9JRAEICENAnn6F7wmQEVS
EwBlGAJDOZn73nd2/rmRCT4j9D/AoB2klLRJH2iKXx44+RHbbY4flzY4dyAuT3lWzxe1zc1Ap0ud
bfIxBM8CdoANO8Rdf30dPvZdtQF9iwK75dFZ20RULrE8U0i9H/6FmjqJa3pZPQhEHIfY1iSxJUjB
KwwHQ9+Hg6o5EMFR0Zl9rghqQIPx2oWtS5KwtoUghRKBKhQ/UbSoZU6gubvpXrCwDUNPLErE63fi
G/ycuW1XZTMzSMtyWk//Wigs4REJYf8qg9ZF6oTR/6mwbWxbh/STcWo=
`pragma protect end_protected
