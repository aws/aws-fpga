`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
M3zW1tp6SfekI4BfdhYdEJ7IwFON1tROpXbSRdcKG2KTF9rIdJrcuIR4FJNBi81E4pwxL9xWcL8L
PiePiBddiCxXoe1zwgpvAoB3DgJu6mSlNig+r8e3f0BnrbQI/nVFQrUMmP0MXdNUAHTwP8vgxUKN
2flOkKkzRApRFTS3oxDKqu9w5dFhPvnUvlnYzfNRGPfMhvEM8LY/oJlbYbiAjEyl+WeY3XTActzq
sYxZw5/+RdOl4JkgaqA5LFn8GwQwjJEjBppNnzRjTQ0QoOUJ5yh7zjLpTeZCa9GKpefmrnVF/qWq
POMix1yF/a7k29J2ibUSQVAIRt/7OESJf21pDQ==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
w3pNw4ZL43tPW9rf4eyrIeqFd5D26hvpPFFGM+a2bmOb1DlPYqZBgnXWOpajnq+QTaQerx8BX5P+
K55rzN0lx/Bak0fpW/zm8UkDcicdbxjp90K6+OBILnNtvmGRtH+oaJZ89pImdn7HZkOluqBQt0ci
oTzuzyXajZ10tqg+Abo=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
EsQ5UZ1Cl5AN0+lhnHGXZ9IMmjqyh6+ki9/wG9eEp6zz87hL2YWhrf69S/zeXF0hCgSXB32R/MMi
M4k53P8gPClORWX/l/uvLEioRhOpsxMQxAnqRAd9RS90b0Snsqx5T3MXNLAcbsDa5zWmDW71Dx1E
1KcD5yaa283JpdCC5SQ=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1600)
`pragma protect data_block
u8K9bQTO1QorrIJZ4CTKetF5sa5tx3nyfLVT/VTZMGbI9nQe/VqwckGszU37g5eqAHV4BnfrpY0p
BcbvNRzszbJR99Xkq3+I2BWEM7Mg7ZgFLN1BmDHbtdvurogrUeyJoNfs9g45gAe4OLillTj9HjIG
Y7UBjd1jm/Of0ax+HskiJvJEivobADQLHhBvKY7rLuvR06Ona7EA5Qeg+OX1jf7GBrLXHhp0uB8E
F/KydnIGH9lGBbWxNIRQV4UXA1a/u7BE62pspkL0SoIrPsdfyS7Cj8wyyNtJYy5VHIu6y8dNlfn5
nVeWc845D9o3KQ0COAZ4wvrq0xgzOazrVIIYsVg58NeIt8g1cZpFOHJHjxunxsllRYiW7nL/b0T4
6ilvHl2qYuDUu+XH0Ta+LW1C5yiU1gQISGrx4ZYBpzb9+xLAAcErAQ1PzD9n+611Ns0WfU7d0hA2
tYzwV0kP5Gk9CNes2EYOv7v6fAZHDLUO5Zx9PfFETs2slTmq04gMc1aUQv0Csrg7PCnOJXy/wWcw
ZVznJZB4k3gElNdIBEzyk6wFuzUIY5doKk7NZkwLi5VAMz6XbqZT+8fOkWNBlFmHzo94VIFvImFr
Emf2Zzf6cSRYMI6cjCyt2aj+fLzpz7nYsyKCFXAsytg76G45v1wvnxqe0rMcf7AZN1/taokJhQrF
DJNZD6195xVJPVgJybr3F0jQod2oLHvn30JqD2xLk8mxA/fjYROnkODCcmcTcLlHOWBGFmIPYHxl
YME8cFqf2FmoUYNF0gbyIimGW/gDKjvg2fNygUlFbG/XyjQk3cAtDHcVEN8xOPujctokN8/SsScX
aSJE10ii4C6rGQ5scvME9LDOCtD8Qt6skRFSdcyA6ozNV0mCD3lwb7XirFjh9K4f+Mmg9wU2hcb7
FzzwcJL4OBv0SMYQmHG1LRj7VoKzV4pfwbBGxUPscocrD8tyJOVyh4RzJc067z6zbpMbkeJdRzt1
KuDcmZuUpjxosFBo0vRw+cJZGIjgkgoh/icgYWvaiTkmlH2R3gygqtU+jwIjZoyWhSyHNEaqe0iP
Lk3r29Ve3jbZpTnXPNk40SKXkM89LjjefoqMuN7XaeTn8XiB1DC0fPwNNLwjhQxJAFicdav24J4P
x3AnSUW+WuuT478JBVuCEMWWGA8QW1NEAb2/uIt/7+ep8wcNW1kIgzipuWUXKkuf5Xxe5iwnhrTy
ykGIgLIxNc+AfdXCp5Ko4bNZdvAJ8nCBM8TAbmEbAEDa1BwobEYaT6UAxm3M6rj9x0Bvn4/DuYER
9sV0M68zqJjaTd7iD5cUHHDZ/sc3HOOdN/C9Nhxv+gXGvL1Yfhg9Zc+WFWFpYimTQ0I5gexDSMWu
sJtRGHKXDYy+vctk95txiIZiGA4RfB3uSVU2wdkdqtw4ZWMcTQ95WIs8Mh6WpPGUIGyPrzTySMG8
8MaauzUUIfQqglVPWdfe5RWgzqTJFP/PharkDBhLomKq1wqQCt2quiT3oheFkWVMyy6rFgmrbaxF
n6LiaJVS3nMRzji63/8FeSHbGkZwWzY7onR+eZ3AMqyOz1H6K8oMAzqprpqCjSQ6Rn5FbP2AVuJR
vkd+wg/BEOSNnzZ750F6NaZ37nt1H6qMSf0WOmnFh4FEFhXkBPUU8y8xQFyOAKZpMfCSZ+K2vGVl
ZHlGu3mHHHbuu/JLYEhiryb9hQmbJbjNocHMsEPWZOU0Oi2oR9AZ9HPzgRAum8ScsFTAO03iGHtI
zDwTHjYW5yWJy6q9I7x3ZTyyNSUsbYUrUeN/K7BvSSzbI73cPs7H9dRpKLDpm34ggCDgJ9TTC1iu
RQOaCD3Nzz5CFkEfrutAiCgh4s5cKGYGnpHaLL8ff99UYeqSL2UPBZ8cctzR/RUeOX4WDQVTkbZu
d2RYMUxiwh+j4+C3xirrCDllCN7caaF/OTzChRpF6OT5bWEuzqy7T5K6s5VSgI+1q8FjthgYZHXA
HjTX7Etx6+HzW7iuHySvNcN7Z5+NuURI4OGYPAwrNd1OxEps/Q0Ehdc526Zlcu/ReCl1cAnQ3BYc
paVsov2No3D4YhIIhA6efR9CaC6UAa1QwqR29ziMaY04E2ibhyE8J7MGKZwvXbbXSW9IpBpJ29dN
ySSN3g==
`pragma protect end_protected
