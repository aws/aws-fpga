`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect begin_commonblock
`pragma protect control error_handling="delegated"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa", key_block
meJsVHy7Gy3rYY75NH9wT/T4lU6JojVuBnqilfSz9cfBLcX7zgZENGlc1niM6hw9UnoijYJtk5jr
yylF8GgF7zg1+INUyfRrTpbq+KYNehInPgFHHvmrOugO+Afn0/Vny6qW3TwbAIJTcFPpuUXxwrxB
0AYPUfh3tFgGADQ4MmRw+Pzv/fekzl1+cEtqBApiDEhiBJlHcf7SR/s5X6CbcAHrYYqELhGIs1W+
wrJKoC2YUj3i5zMOK8/RkCn1CfdKMN8fhj46e57b3l+XEmpSZWimRB+HTTERAPy/vJ1gW0wipcKh
GOXHm1VUAFwaYcHtqKJdKhqiCAXccQ0eL2CecA==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect end_toolblock="CcHN/kTualhIHkvRUPrPqBcobcf0l2k5TavBGHOoZMY="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2368)
`pragma protect data_block
ycSU27/VRZdB89TBcLF+FA7ch++GBOoSP8+NxBZgU9PO783Z1Ale/Q1DGDsfg6VJmJ6Sw2mCQDHw
C1/i2KoOwvkOwNBG+77/9n7HsBKC7BgzNJuEYzh42B3XHk752FbLoP4bKyeE3FzheluflkZl2Av3
7Gc/vRUa9VojwP7UugzzpQlDjkxBP9SGplQDAEzsV+aw+7ttLAsTPpNkYvosrsolhqhgX++B451p
Tiggp6RlxcQt1WnrcUHjAJObA510l+0+AqrvnoRl0H7nD49WT3A0/VgMHSg9ZOpcB1TKHzBpVDfl
boTbxWg5l1Y4EQToE9HUMvjwRMu/7OZokO5SXKIDDZYzoPw1gOvLU4rxWgphyk0S44WMdvitscax
Wrk0wlLO98bO1zLalWhkGn5dD48EBPSa9HmJ9ybmdZVSDgkn7Q6xEFC+X84icon7WhbHgEVszR4U
ASORjWp/V/agMD/+rBfVAU/kvRS0frH1OhqX+FdkPcafVUeWHO26mpoK6JV4mO3pXgwLYI/hkit5
Sr+AybzyEuj7Nd1sl1z4gLumQe//ubybMeVeacI5QNaUxkBBfDBeOXEL5jlA31ZXv8O9aUz9SKS4
CISkMkHAC+W+qTX1YKJFB0FiJQyR88s6e6PayULiayGB/3Tn6yk1yJST1vi5W53WUZQYu1spBFwz
GXhjzxG8LRbbWVDpR4r21Zr3guaapkAzSwiKgdZK+BRT95P0OcN6SgHyvPpQeI36NwTcjjt3SDAG
aoDiJx8P9YsF0yxh0FlQxG5R3kfkyreu1hy4FMbvV7kxnI73hmePLmGbJeENAoCiBAURdYDM8icO
W9Flek8geZC4kTtBauJ1/pTDIMoVjyfx7vVCWreAnVMgGmFJRsonUw/9A4wBpNiSuz14ot2kdBK6
uzIbNu/k1PiOL7zhkLafongo0MdEph+UqtSlYyPg78GFMtFokVE72Xt/pPOJpJWIDRqiqOeFu/7x
7j36B9Gl3U2ru7JoJQZ3zSzoZk/FqWprDsXPg6BtN40pUbQAn1ytptOTUemn6xOJ02IHBps9XiNA
9i/PXqssB8zR34z3Q63iCfi/u9/9FgWHowFf1Fptsgnk6a51eXzWEdXmd7nIW+oNqguXSYsfuqXQ
+zHDiNlh6X8O1bbP5miP/CmY7tUlbwMTf35a+rOOM3czuHWiPoQQ9pGBfW9VdlNqYZzOJJt7Jq8M
LS4Pyen00n1RVtMTPH3SZT8K01cVzRLT95VRXtrz+yDIODBHM5iiwoYL2bB9PfmI1xu/onuNx8VW
8WiWciVN1AATL+JQZrcB2nE8Mo38Q8b2POfDY6deRG41V3/PMYYBCbAqvgp+KODvStuWB/CFhAp1
AA+GEz8UrQfZq/qKA02o9rG1Dq0Fq/BLQg8e+Eisxf6yJ7JxfxDAOJfQZeM0vuV1ffSOIq8X9jeO
ouUascRuXV9lFODzGRVdwEBL1aAIGenhtemvhh6d2Ls1baYF7TA236HiHSAibHboXIfuYglBTJRp
JRVxvSMnmnsYEivZ7h/0Xvaf4Bp/Ox9zlBoK/9q6lMDdUzr1hZHfZf9ALP3zy4Nurahf86NIh8/z
zNJpgH39EhiC5U+KDrkB4L1hb4NsVX+alE5NspgkuKn2u7YKCby/PSXvsl2XG1W1F6KlzXhqSWhw
PwADppn8tUh+7Vg7+ySbD2UWtKXjnCRYCjF12eUtymvAxNNAckjSG81I7W38Ty8tnHOP0GqTnrxC
uh8aLuioA3TETjl8bh4QL8BIHsqp2mVKfoDowDSrA8PRGVbn/hx6uOd28zFFD816zBHdhclwnV0G
7j0WZmeAWAXQsg8abSw0D9mbI0ZA3nYFzPBbZceNo2BFzH5CTEU4273AFYP0Gma43P2W4lAnnV9H
VYgzOI63Sl2cW//AHu1HjtT6bwmc+oISmnMxZCaYng1DEKSRPUMrMCxTsSbmxJ9jnVqNDOTMzHwT
0ftL8kaZoyMOu1SAHqDDNc81Y2xe1+u9pwRRen6Z6bup7eSYDoNqQCDksTsN0e8UJM+YLd866ObJ
Eruu2w3lQhhFcwMWtai1nBp9okGeS3nimERME4aTQsVKdWzxKXkXqATKnjq+kedvSpLsTKVxpBdD
5+yp0p9nV/l9PZhoZ267ZznEIn7ENPo+r3iyVwQM/Qa0rTjreJXUdgiWEakFbxD39zD6FJCnHZPD
Xi/mdhDXN05/ehhPJOyCFpUCq/Am8bYMVvajzV9vcEPpze6gqsnnyWigS8hcmHDzSSojTEaN+tvr
2mR+4ZmlLlMiHF/jEdEw2Fs3yBtooEGF6HggCNkssZZ5ANqukWO6dUcT7S6DnNAVsH0NzjJzl48Q
2BSQJymlFUVTP0Lp/N89OC8XnAcgohehf0MqzPLn19Tb62vWeCSyMjExf+DuKy91TX351FlHDUU7
U4JKUUZtO3bZcngLiPsZHeSqX4Zw+jwwKZ0yBBU+/6rUlXooRIGRwhSpX+SlApS8Q00P5VMtEcAq
ag4vVkSlFrUeU0fjLujCuzDOERoFEhcoVd7JYUDUWdFvm6683qgr3P73wxvRBrlxvov1Ia+fFoKs
vYWWT01z3RUlqc0K+6MlqGqixBPB90HhgK6mzOfo6KG5465CoggUnPDXblOyXgTwmhdXHIAt5CHf
P5QexojtoK1DHSIALmVPNCylpQAlna+t91UL8972ZlyIwNRmhxUZGefUbeKkJPVvYF3Zzcolfeff
vtdhDsunEAJaWbHc6XdLuSYIGKUb/7rk6kO1ilgbUdRJtas+GnoqQ34gGXJJMVdN2hHTvjXOC1aZ
mcEmw3gu8ICvq8cvpioiSQtYCxc+WTifqDJXX7yLal07oH4hg9eDoPhQLivYc14aAFLPwXnq9lup
ov0rDTgLA5WrNVBO+ygXjkxEeBlHqP3kuDUkKdSN7oceHAW1lwSnYSkcsqKSSlufZD3nN534DkFQ
08TQj2fqJNuGTY4H3uYa5awJ6HhT4lyNkFZzYmPEYVZFnxfxbI8v3eHhrJoGXDCVzfKAh0w0W/Kj
c7afKdIWB2R+lvQ/bqUglIEs4ugZ86QxgoAez1EQOl5N+VfqaM5ZndJel3QP+n6YbsindPTC7l//
VrpWfmT9uS7ZjXZv2VgxTbhANIHCfzy8OJcsNxrTkA==
`pragma protect end_protected
