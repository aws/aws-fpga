./../../../cl_dram_hbm_dma/verif/tests/test_sda.sv