`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
jlRPg/sUE3Rzrjxk8m0VwGIpGnCmZcmvi+xb/1wgAre5+XaEz3pwehoCA74ddnzysXz5k0oYPxnK
dFsDdAc5DIXVDUc9V5ugRTwF/TvXxpVzaJPD8EgmxxCX19MrN1oaO9scwMP3MhVbD7b6nR35o28Z
L3v7HjzMuCe969tkjKr5aQuDHiZAFDox+8Mx/GIwBnLlwe9Xb/8GqaxY4JbY1/CqB/04As+2/ZJy
caM2S81woGeAmYJFqJ6Uo4zjKz4cdGmCJSsLOnKFNGWT2/AT1nyBOYAOwNKNJtOhbSrgDaCCnFMg
2AV2JRdtHRJgrvWDlPv5LwN93xu0NnL/U53w+Q==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
pVWB/UWbarx0kknIiFgMbidXqeQySZ3W8RzqspL42er1CnFBaUSd0axA6MEwv9GdS/fv58UeRRyK
RwQuS/MzOCbHS1Ap6KsKnrbCd1Df8IL1RKKMSp7Tciw56CQiq09McTB573he8DevnLUnXp7upXxG
/ZfiMo4X13xicWWumfc=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
phgj6mB2wVvo1huw1ANy0Uh5z4P15MRpN0q5W1059Z/Npi4u69B8TISYmBDLOIbzd/efZ/oYJMrI
2WapuJhwoobAbIk5Jv/wu0Smk1GhXbh7UBDmKoUyAu7ek6eoj2n1E9CgqkZTRnrGx7GDTdSt4k7O
prvZ/WEkGI3U3xT0hSI=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 35824)
`pragma protect data_block
N3MKk3w4YJpIh/VoRdvqXqFAIu0yhyd4M55k9PpmFWV8nYcBB29z6ACS6fGOOYm6hiNUhiO5Earq
cq00jQXO1iyCQm91Laf7atw2r3HnpIR3ivHLE0rwXcPIllVfB2BXU9jw3sXoQNxzwibXt9ILFe/h
htDZrwSz6rpGzPcb86GpyS/8x7um0/qX0DURd4MV338m8fljV6ayLZAHvq1fIXnB8gCHhHT4uV+f
sCOzgwaPdc844nP5hrVq8LM7MOaI1KDRikD+lNE5aaC2VF/NQDYTiJ9AdQJNA97BvBcHINwqKs0I
hmKGi4JPrR4a4CtuE9hamkmkh6zrPELvWOc4LIA9pfPhutgBF84q4SZOryhrOfzNZXKy8+M4eGOJ
HFxs/1jQk6yU1CbtCHiy+on2UO4T+Txgi1FSTE9bU7nbu3LJ4pLOMc9QZAMdPGoHBtVypyJFuUAR
y63PtHxw9F/6lLLbYX5PvRN2QrMQKh8eX6VwNju8IS5qfRcF4Hvs1oalf8j62lNrRObYoPtMMhjA
7mNGU86/zVPjvypOWYsJ2avkayH6T+wjahOLcl/Vbg6mYUb0vby/ZjGnqAAD71nNluSA5cwqDeEK
Wn5cV4AoUNvSsxM5wyRL3kNq26MI9cvzABjH7KCAfWjthvScGaCKjp1/yKjNid0B+gHTMV7S2dgk
kHF0dTCLbHUtUf70dQK1k8TFR6xL60nI1JExlt9NU5der2Ay4Lmaujk8KAN/e1ovl7sOlxn9cGFM
3T+GWlOa78PylhVoDq9JTKqn+TEA3pehK2jOmQuIdBJFe9g2McQfKeO7Kuuj4ikiRKi24ZsQNzum
6IoNhUjJqFbLGUrIL7c+p8vJYX3N1JQQ4xzGvGODQh1Z9uTZsHg9jmYCPMpm8qNYlbWy68+cOgcw
UAuyWfGHecetFrmfZO51qu4NN18sx5gUUssK/Q2mgK63bVBqm0jxonsqhpux1pIbzFc7FqLBL7MJ
XS2dSRII+DiK+BNi+fhKCl9SiNDysGKiiTqhHmONZggMuhREIfwOHQab7/Ecxq1dHg779cXInKY3
Uc2Zjztajl5GUmhK7qdXKPgtUVtKFvmqR884NTVxkokpmMng8PuDq76Fey5Nn4Z6hBwHpMpn/zE+
me4qda0pYtTLmKj9gP0FH66+uR2FpDP6HuUlfojknaDqx4pLXAcztXrqrGoz0wwzEShyre5Ls/sX
dnmwQ3u0joedanlFl2FCvaiVSkSEc/HzKcHGcv39Krqulh61FG2QKss139prWFbgLGmEi9s0O9SQ
hO/tGezrIKhW02+NBRvoDejJPq58n3C1PwtJMZcAOweN1yOePiUWeOKazP4EiNCeXC4Qvu25tHjd
fCplKvur0+CBQ8ss6A2+Ql+63JLLmPpj5eBeRsT54vhlRLt1HzXVHF5oKkiy70s3RcxUzRWCGUCN
PoggL+pJe8q5HaI3lOlkiRhOft0/HWswi9ecoYSpDVsoaHgT67korqFWF5MdEvTxTDe5meJjzYFm
PPWoVVB7Sov+AuP/oAqYq5+rgLavqZS7v0f4gB2Hy0bWXOwvcwxd7Au1YLNY4MvHHHgLZ0T2Cmgd
T4RIvEi8EkGAL4+ltC41X/e3CFVkxVoZP7fG9EDbTdKH3hwUjtJHQ403mm/64h/A+1dcXfFC+HZb
yYHifbcsKHFfVDEs1iUy9SsXA5sd38jKnbRd7U1UafhDsoM7CV9N7jcZaVDhSyj/Ozd8lPQcz6h9
gjMr8DrxpoUWJ+FKocfz23XB8AJblptQtXIBaQKn6OhFdEwxL9YoWtTneELIlXavg3A8BP8ADCWT
02M4LegSXFS8wzEEc8LthJg48AG2Hkgg6r7kQOoA/be5mwxQqoum68+vBzzsgULMlJrwnzxIeReS
l7/5xGSxe+j1cgDVCj81h2HcQ0wl4/ZrSilkkCSMpCCcWwmdVx66X9EeAJ77MPeF0x2b0HYLHiSD
V1JIeiRDQPrUtXS8X0ckWEaIHHoAQ9oBqXqc33XcHZikxK/tHTuf8icD96sPcrCOfeb7ChXB2qIF
BM802OTXJvOYPwogozavwuDHYsW1/cPVOMtU4BImOm0LWH1sORI8o2co3tsILDSOtjXtndrZiVIl
UVjRj9rX+SonmuR1oFzqPrRr7xV7OiGVg2QP+4ZdsZwNpFLXrg2BnmCGvehEOl44oUneD/ZWomJX
hM5Aw6tgp5Hra2yy2OScwWcP0+37E/YUtqqwyD8viRYDt/7dxMwg9OmicMFpRiz0RDPZmXhwaSR+
ZfaV8Qz2J6hacf/lwCuf5s1G1X1wubrU/HKxYQeoyMudRTSbermyQ/dYlhghsw2rY+WgpzABtevF
4/XfpJpDCmk19JvKTOUfRv09ViiMttdffCsmsbdQUaMhMfHeYZj1Kcm4iS/uKLjoblhRQtg27+x0
cLiBMDOD/b0msoUmDX76tv1M5zLXil57aWemgeougMAYvV0gpwNrk7GjrE4dnOysZhhp0fzZih1d
dDidQn/hhftAbqzMHswatd3RzcjTpFCemfsW2YbawEFeB5+eqon2k0j7UyNWUHpBG0ZRbk0Zup/p
EAgpz2wdAO4Y6Q623QJPyD6Ijl6k4IYMDWDwGwfxk5e8Q570JVUrsvOj8tr+Tzqi2nLqX8sBbM/M
ij3vAPwuoDR0TKgoDRSYUbHz9J9G2RfIhofBgKX1XWynSPLwtcOqRmQg8mTlsaYtBiR8iu7WMDDt
+SUyNhhVIZXObsuaH3GLhpG3jllQEcst+M5PSugWkXmxiRqHBq1AiYj9dH+oubEYh254PlMLXt4+
Mznx+sUY00H0+m6LgZAa3mc7T1//Q+qu49tZbuifDZXpEgxmXGRyUetGbHUituFJcfCr+GPcgqxk
LWjPOopQFInisAjq1ZO9b4vYxulfOBTRp4K5+qseKOI3bK/mry33WVkA9ARfKtnlKyMNBiiXp5t7
DkF03VVqPFScDTue8sRdI+l9ku3Wi52jGNCAVIpl8J7W2IEqjaeFbIriLPDJscHvGN17EDXFlDo5
/AByMgyIuruDPHFVWyD1WaJTLbhb/T0NaNXCM/eM0fks5T85zsV2/J7lWJKGGgOcqhJL2vpPXUED
8ls+9pZMM9y9DzTBtY3/TnFaf7358lMXQNXtqaOzLbjXGxmloRCEFFuxJ0GojW1qDCTH0iP8UU9A
XaKnJWAYko08uh4gf/sBBD1djo67ZPNaUfZ5QXFQW9gI71bArnWp1r8Fxs8hG3i546K2HJn7Xkxc
iQvkf1OgtIxAPmLZyYdq3jLsN2lVABiC6XPStRLum89Pqj20xJYam4sb74+Jm+IE/KUvQ3AGxqeR
yTx1J0CGBP6PT3eRoA+DY8XSbcLgLRkLJ3EfNvruP6n0z9R9ciXpE5fi+SNeug/OSgIC9FKN2FIe
ChpGs275vB4/p+eqJW6srRrrQBPEZWj+t1MkzYYXSMi2Y4V4KEaXguPfWxW5U+Ided1Rejfx2fcY
ShtfhrC1218Ahj9tYCAheucIB/9hkcIvKj29l8P4Hn+HRwJjq+0zsOXgbz3g0LlgrpCmUiwchGVp
qb3JEQOcicy5VhMpSI5MUaChOq+kq5UmP3yLAtJRs1PDnkjEs23F1geD1nHxgOf7wu3jEF8KL/L4
aKOAf5553pQe0VoZDxgVI3+4W/IRdM67vpVDtb2f5Jg8Ru+IB+3HSeGSXPVmcMyle4ZYOW8gcTo2
PMev+le9tVGeKgiy+sngJd7fxGw/olMRBbJnvC+9uQfFm8c88Z60zGCGXLbPyGdBMDnOe4u3l93t
vOE3ZhQhBH4amg1WxwWoY6ozoRBfag1XSiTXlyuUE0GPvOGaDvocCmPqKOXFvPnl7f8IKB3p1GGG
i6j2Vcs8bGBlPfQW7i803stA9YfPDnwhdWMaxWq6aXd/RuGqCOLqfjb9XQQEX8rsECqHUJ0qSdnw
uqdgCiemEoXsoWKeCA6yo4o5Z/kXgDRKIfApudtN1Ah8I0pTyHtt/gfAZaLP6VfXuk8iY5gtGSWk
W+ERZjcM6WxauMKrYd0joJZ2pa3SioP3Typp41fy5SLsSa6wPt4L8cCXmFYjXeWN0QiOLCPj9hfc
IynSoMFUjspNGO8Vi/9T7KW86eGQuXdpFJnTVDoU5TGKpXYr6FSOqLT+PCbqH82yyoN/BoeF3Hgq
JJXNO8cK4K38p9epztvFbQytiZsipUMNWL0XYsAP9wY8mIwEdPw/lSjUpc8YVnJMWCgW6iHVs27o
ruNcpR9Bti3JRVlwep9Fg5IbKDCMSEAdzcDYMf0cEeooL4QEs7YHRVIG93FduKWeWwDleyEoJe2G
yBYfQZg6WfFxd53pwyo5gl3hAqBJ9tDK47z/xGOMidCh8+eU7ftKZUJNMotxCroM7NNkZ1K3tdnR
cbMbMeHfoa2uSxwfeGAOfjnmjISUciJIr975YFx3xgWcQ3EnfYQ3UPqVnn57GBqkAxjbwgKSAAhd
d/CjWxByHgu0QZ9QHRdU7m4RnzCF7dUdhIZhFgLPRlA5gdXFvaXkXqiC5Kzh1ORoMAhmWTQmIbrQ
3KcYqGJK2j5yaapypQyiPvnERMANikEnb/2bHYfma7uFlW/uISpiDlHEh0GNBc53kIVOwXmc9/1a
6FDLE3tpXblevHSjOXAT3vkSY4RVhZJGNRim8dx6324+M1ZRGCJ31R+dQLyRQTyvSWLHq7mnP/dm
cNb5Y5Dco3aBaRwFxI6LldSBsSYvh47lD2dIgio773PB8MmDwqlj8x3pfEnkR9S0DkoOVtPQsA/z
7ILSdcn7mvIMxyz5uDg3cgf1IkeGzy1uGvV3vPmnQ2B7LEfTzVTvXGGt41U/n2Gb3LmfNRtBz8ID
BPbB/QTjUsU+mdz60vlGZYClNgZOn8LRaVrAw2+8LAa97EALSlCXwyc6X9BYKnSa7fyyIr+VI4w1
5jvVCgeur6lb5U4Xn8i88AhYLe2AAI1y/BIpS0mP2em4KDdgEmtfwjaV7dePtPBpjYSVu9GoOxAP
oQrQ8oXyv/rU0E68cqs0KmWfSgg5SfB99xdoR6voVSPk80sQJDJbDk0v3adMblsEXexJMSJmyrxn
iHZAqROdJYhUozcVf3ghUDdgVltkdd9HZGhU5kkC4DpehVg+RgAsp4NiNZ3Kzq4tLjLU9prQO4c9
5C1t/Ol2nJ/dpImDxq3DU+LZdrABGJ/ib2us+fb+JTa6/zgeUVNEpLGSl7NhxGFNmA73O82G3hdp
o40MaUPG1CBmXtsHlqAqtMUiI4vzq2Izz/LndxM0yIhZjVhjRKsPhRs3TRWU8wRE+Y9bd/vJq2lO
Mn6Gr7hfGaXu12cyg14jw38smW06pwKGywVnuaVO8wT+d46hpsEuNgy95GcgjkGhRF5dqsDo0aFU
hW1YliP0DWEW2t83nmD2cgr+I96k94GYtJIfVSC6+iIi0Lvrq9/zOx+UJt1fdTUI34IaKxyf9HsB
2r9CeEjIIC+al7FLKtC1Ehxo8aSIlMldu9WSEW/J6Xxkl3MLE/AQkr3y9UXBt37jIeULoEpBpq9W
yeDr1i5gheuhXD2t/dqHh8Ld1kHylQYBMaL2PnjB4ni+feND0E1RFKcbeWh+hgzVRJvGCysY9HUs
Dw4vZf5Dicl5PhfTSVUYC+f1Q3eVWchr7YKSfxtAEqMwlniRlHRwSGCVRZskhdyhYH+5hrFE3Um8
FGK2pRbm0ZvnvsdZn1g0tPDoTJQBjyFV6pkSSx/heAJ9xlYWW8yWU4k/kAsLiUxn4CslqspTYZ31
+gTRG8yUdScvHzxx8WbKPunPQQ4uGBmdVvKdaXmJK12Fr7tuCweM/3X85/cJ3E21QqfFTWwdyDxa
Y5EQhIxoqV7xy9U58OzELT5fuNpxAU6y1eKnYg9X5lI9wBVW62pzgonM17t32vvzzWw+lRiQnJIK
VMcvumwQu32wJaPT/igAN9xKWwPEO3ntFCgUnf9BtsOyS82Ilt84iU62GZDgFwnBLdY7fEIl53Lq
siHI5zALU5OH59bAyL3SZVOmvGbs/Mw8/DAlIaH016z8RJoNYtEGgt2tpfiSUPHn4mxVFcD/Dc9N
k27ISfzmpfeBW49dHb8TXyjCRJvyDppodGZoBQqcnUNWdvbhSrw8tre72i8xPPkv4bmijf1HUKP8
Jx1wgE409DxmKKy6yQGFqLKanbiDWQprF/pX3VeZxBPCgcgbl7XWCUhU5M7OPnvpBUwVl75/F3Mf
rL9i/8AZyRnxv+RX8ZAMUUlGhLZR5517SSjckFknQJKni9FuwnXlYLLRu4G90jYXWLQMxpBXpETG
Y4vDsy/gnnhD0kF8CHhq7jGHh3k/AQzdOfXgcVvte8MmSSIEtTvKxiCT/6XNRhc4C/GELDiOk1xH
2lihACVlYoVRkbX9ZUYrhncU4tOuisFK90lrkOiL1v0UAuHPeqrzcYnvTRZv3qReh3mmJ6waFqcz
rrwRji2t4i7eplgIuQLXnHRVHb3tdUs9R9dTqboQpr5LKdmvERByrVWSUH52jyfzFj2mpWH4QD8g
sAlNkpgdp2wdGw8mpqollvuL4nQ20Of2CzHtYPE+GFNJoTsaNxeNLTO4G7NzuQ+ZcXJr4+7CjSsc
gb5hda8Cmbsj6yD1vifpNz5g/xKovcEabq+GyKWDMdY7Wp+izV5CmDikYIkD10xc1Q7BkC+2lKV6
di6njW903SNpWFYzNGL6Ty3lJ2ABotBktfLjl1fAb99aF11OLvVDWhDaJXdaLRzZWU+0iQyo6MLJ
SYsukxlAQQxX/VJTaeVMegNedQ7M62KqznUuP6fZanFmiykQ7PUfKwQgjDtx43ncaMdjN7UWn6rr
LZhqv5U+nzgQrvHSZ4aMp3DPaYHZ3lUn7oZoAugCpeLql9XUtgVvmqg9oSkxZ+w97AxfDlVPNHlN
uGHtdIo/dLFM4uwteDvipp7niZ0pg8EfPQej0XkEszioqY2B/1UFEt0T0N1g95m7wBHpm3aZc9V0
zGe5a7HguGjqh/UVqG8AmHySgoubCP7RVgCI1NiyfewuY704mM92FnrwhYVKOy4m21d8zHpaj+zq
+a8CXQk/rWNUE+7lEggJSWXYdYdicvrtMQ/DNCKomoi6D5mjhY438LF3zgJmVDiasdYi/Q68K8DC
397GHbGgG65ilVoq/cy0soXiFCnXL2aUN6Tf/UynD9aAm/PbtnrK1m7YI6s04QDnBY+LPDehotfg
KVOcoqvJtR9m4eajnW2xbhNX9qJQgYBDHEFBj5p/ZhHxXdcszhgkF8gcyZOW95YbDqycm46f3e9B
VIXuQ7z43mmEabzFtqMUWyEWKADuLqeCEdWLUhUHSvo98wnlr4YTuALKZJx+iLjFIgZEBqscriUL
eJg+aTj/57Uum6rbOADTpcUPjsWC6eIQXIUJ2zF0FKX2LaqZvrJLzH2N/hfqH9/7aBZvocUunO6o
q+k0d9LrvedGG1DQnHzJt5SotOCZ8e4m8vCa4i/v/T8Rnu1UQ8kbn6FKJV3U109/Hew0ngO070iB
Qt5f8bVW1Oy88CGiWFFhoujC8yodiQUAPehpzuTMr/ZP007tHf9OWejZaLKRdhVYuECfDa+7hrxh
uwPP5AQCJ/uSQtXobn0p9hsF7JTpg2CmXZH7W/LM+OHpnlrzvcg/cgjnTJy+NcKVyghHjbm21IUl
aQ2yrPjyTDWaV2RvmQJCrb78lokF2yxtsQeFp7kpnIRijoUgn7OgYPfDXB7SbgJ1jyDAoq4Bmp6Y
o3AF5034tKWr0NVp4qn3tuXoAslGk1Q+pG1OXXVOLNcwS9Vuyz37sq5+LGarX/n6RTkjRpWi9xRY
Qj1l9Fm/uHDCFr2oeR4+Frb4zH25P1gZspFqF6KDhRW5eR79Y/SkYGSEMSto7XEgEmAmypp3MZbs
x+0YUEO+4rGSCxX71dSlWmAB52ZoHp4pU5eAWB8VH2NuNewKeVOfkyL00C9t9jlWrGZFdDMqDDxm
wjfP+bIPf+4zRO6dtrCzM4lrRBHD0n+81RH+67+bPV2AopPjhyQVz8tfEGwCIMl3Gp2t+t2b0B2V
SX3BrbHs/xj7VvPiT3WuFhviGaaZNjM+fEOw2/D1wnokJfSdk+hIT82AUipiB8c1we2C8QhPz2V5
b4n17JJN+GGFQE1HDx7bzlyJlGKky9fsJgLcIeHQw21a8dxkf4It6I7klrFrxsV3AnogxMB0s3Q6
smfS9PJKdmM2na7DR6b7S6sQbuyMKtDmV0zKZ0GS0k/uph8cTHDccMKSVySZOhuOSVnMuIGjE2Gx
JqePGmg8cmGhbxpg9nRtz1fiC/fnhRM+GVOHz1Lf28PJZedqs54GETe6z4PpK1GQuoCrjdEzXtKP
S2WlDzTl3RDc7xcaj8N//lxdPtyy/lYOCi3g3ZDxPKWctCICd8cBedGu+Ptptu0Kg0uixQKecRt5
2HSfpNfr8tbvGPXwfHw8Whx3KQWKy5uqvFNtUBFoTqWMzWUC8KH33dmskAA/62V2IG+/CuusmPJK
XmuIm5iJPKkrFLl4gRTmJwHskA1XRkK5CgN3B6PjQK5MwHoFsszSRfqSfhRXJ9VJMXyyKExRVJBL
MDNLDtEG6eOsTMzb7NAYH+rbWBe5lbuKmtK572lLG0cchYsV4PoiZvf2bGcQQx3fk5vdi8QPYZTZ
+qrc3oTt3wsGq6vV+0wJQzYv5EQYU40wGamocWE0y2vKe1HoWwvcmZoF1QtZXwWX7QeGv9POe5Nu
VbBKNXeeM/PrwPUYM6CbkyPeH86OqothMeXgdmVYRHVNtGjrqo+6fGPVK4AM06ZyGnrQFoBJwp9s
faZhBIAqZS4m4JyKluoiSyRynRJmw84lciBZ9ve/fLXQoZQ0LIs0hoWww8T+xYmt4yBNZZp/+ibc
o1mMv7mSGNdyc+WOihDBaAXi8b0Zd7T67zrRahFr8RWMJvreILAQmlDthPIvQPmClcVMyC7i6Mra
X0HCbQO809MH9vQgEhaXG++2gwbhCfqewXoEGbNJxXdVjzxsoLdgyg27Oo8ZLAGMkPG2VEtFTHvv
sSDkvMM72VE+NEk6OqF0ypxuvY79Y/xIGKM/meJvA97TLytIdMWg3DCGyFDAnU0If4EOtd1R1m5K
vcjrmstsnXpq/H+IC4FvtjqrWSmdR9ooKJT6fMHjdp/CCiGDhAEL9rTHKWeQOyPHb7GIR8ID/7Ej
C9c1sY7lg2XkinFgNidF4HqoGq3bt+vvkOPZxWMG82KC10dgdRlXBp489pLcPHbhSUKZlKMyiTZ3
ISOTppMd4fW/3kQddK/f6e75VIjKxlzGwQ0m1AdAjjU0d31Gxv52XG3XFV4/D4kCt7AYGqBELhNF
CtObhUVWYZ4Zji+xldJR924aAwoJ3RHVHSvijeIJlZLNPkIn3osB7vwaWprrT65HZKYwdcJX9Nek
pu823vd4pThMcFnaB0KsrFns0ojwTbkpqb96apO7A0hdeJH1Kcj4GVwQKizVuQESrqCK5QfKeK+W
5dknxj2mW7YQTzLjeuC4Y8/L2vblswVHOWUKvDB0spVpzHrVqBg+ItqjFH1HkG+4xsi9n1dNYbeu
In4CjeBoBvF82gI9mBIW/YyECFNtmIfDda7avPs/P/pyPEoOLy9GEM1fFr/3Cn3ol9qu5lNg//j/
5p7QoNNV7LUWxVChtBImp4UeqCwmdqi6Gs9hC3XaNPha+f56hlzPygiW+1W86XDR+LhExTIqR3dO
9BxuLIQFg9//2H+WdKXSCBJU9rAcMaFPvBNp1IJsCpwyZPdHNOxO+M30RpbXk2VrRCR+bznX5Wuq
veerqNoVgskYEJ2LLxEjDBEOp3Hjl8AUvvdl0srdoxKXXz6ov7l/xIMH3k9cYWeZkDGJiO3VirgK
F223Ki6doW4lYOvv6u8obBzULPoA0U44qywStJzAd9GNbSbtxiYijGjN3CQDdBGhGqkqLK1HGmM4
Juj2bIy0F3vuIKcZEqj+OZ4EhzWMRQ+pWEJPOlGOm1gVxmxZQFPKjRn04V1TcEEiJW5xoCStXJaY
O0VbWacBQ01hLHh1UZCnP2HEye7GNISVkcHuhQWS7nd1mEuUgl9jiIls7tsX/5TzJ9QzQzQx59VP
sWDX5ZNnD6JviwWpYtAE7FO6+2rCpXnwEXLTja9DqMMd3poEol3rPdivlt++Kuv7vsQq5CEglKhK
becqkef8KLR5yvNhzU+USK835c2uVMY+SLS4FeKTJhCFbOXoa7o8mf6+xge1Oll5tiTugYNWn6PP
V0NSbqoAXmxWjHKxim3MtvjPoJQn7Pl+dBEDkPG++Ic3eEu4CeTKKX+pNDzet8DIOkgXh9lrh5Hd
MXlg346hYfqn/WF4CwUIKbH2e3w+dd4R9+dalPMUDc6ETtPc0pWNi/1oW15xSap9/WOm4f0DA1C5
WTDu0Cc2uBNRvodMDK7jCfAouwcYHGjGVtOt37Ff2wXzALJhDNiywYo0I55hwDHcepuU5sTd6yU5
09zPzB87yvBjMX5BceixQCCA8taRLUOpVEI/dZw4KhIZKu+bSaZqpjiaXgUWdbb7P6WQMXW0hUsl
0qfmynKURVfBiT9wETC+nsgods/kLgYS11NYpi5MxM9o/DznWXNdzA7j0cL3SKaE9EWBYu2lQf8M
8imaArtFkaH+vUrFj1ZvcVlndLrlVBcM+ypxNCPk3SgDgQps9znfKK50vl+1w6+s4PZb7rVEZZ+E
fSfHvJYPzlcXAwCHEt8ESrClzaonn+v9VmStWA++Ujq2GPnuqjSQH3L9tXSDCIXttoUf+LyxACpl
tT+WrOMOGdn3q/QavGh87jsGtn4RNojMmwFM9V/GMGzf8ZZ54tUxu5Ofms/v1bOnHjhVMbeM5mi7
0oWb/u6WxmYh1M9A3KqQQ4SYpOGxTmNv8sEoBkmDbpISCQmzu2waG8mkb5OBoofQlV2pGLFtccek
NYbaX5KUn1D6BEHpCaxnfYVU1PcuX1ijneTZePhc52vIIdnoxAxBEl48lUkkzkYUfmaVz9J9WRr9
yOf0yPans0tWHh8p3fMDWPwybkCoqeXbp+xIgDxnYeUvHD2aXQsSfaHEthCXqs4VB1GZNMdSPsrN
/DRe/EcU9GFzkisYDnLz/fjwHy1mTmikidseI2CmwaI3G73fcJf4U8bOJHi/sQX/bbFHFxZVeZSW
QdTMKMAywWpyO3DFb2wGnWNWDhoh66okUaDAPjMAsWRG5D+NwIuyuTEeGxb6mptp7vVHFfldhtXh
cVjlbwGNq+ToWsemvwQntxUzvhuTNThof2F5HRJR/BLlPG9oIeOZOJQ9eSPfTd+3tBqUmc+7Sl8q
dafCkRQf2VU0sflFh2gI0tYsvtglJ71BvJnmhrkQzuFkjDph7fnsWvZfsFTCA8zk10pY/8YSiWPW
DPFKbDRfpFcjqg5klGvaWXfSjIA2Jtd5RO5my8bg4kaE112tMx5j6tcFcF1/srxJtbyWY2RhJ2Oj
I00cqCjAyj+YDRyiT9BX3+VCw6SmgbQENXdLU1gg7JqKaFuSwKpBoh+dmbaX/5FmXUUzJFieQhVO
512bzkXWPFToba3kK2FqmIVcw9L1c6k2u8FM7Cuy4YwTow8CXy4dpcSLBUFXVKmO0DDy7eLdCEUm
qmRjGuYmWbV1PyNTmOjlQtoD6P3PeiQocX8h9fLvx4EJyafNHIklKH+aA8AIKq+gop5nc+22Q8kL
P+QF3ZMi1ACmyU9Z7IvV1xWasPNX6Oo80GvAxhUToPPeEqgtTvllC2tpWaqKj4tVzOT2oDTU6b8W
JmOBwmEguyeLgefebNgvZEbR7F+AU9xMMYvLFi9G5RfmqbAkaFTwiTKGy4GOb7pnPYEmaeNIAMmA
I107n9ECs/XtgXfY8hoakcqNDEL7rI+Hf7OgvHgTXZhjXXXK+ek95JrIhaLGyq2kKSFmLmZ/j4SA
sT11IE4p3MfkPhaHGhQrOA7K5wZk16inBuHbUq6DxPvn7DNriY1bElEG/yOy3xjRVwWoaacNMTSI
WShKcIFTLM21yxCFjBAuBQ7TrKehT1MATssT9GF9Sy4zhqwDBHc12XLWgA+pyw30Fam8QNwRxE0k
Rw30+cN5j9hy18yh25xMbE5XY/Q2VHVsn3XEqkxLBga0qN5m8ugeQhGB0mrxKMiwI7pidNyQAvQq
g0iIjXu9YGK848y8dEdgrxdReOFZSYuIDlsL6q0MpMkRIUGVbta9npDmGbCNFneMfja5peOTXBkf
utA+NzSdxxkswWMhdB3kzBKUGHrKnRrP04oenbra0CkHJX+NXvrB2gSK65NOe3A8ymBANu4MmtOV
wSdRr0r/Agb2FzyGcgbtBZSyKKVh9/IFUSackQ23Ag6TjAI6Rz6k8xeoGolwL77zC9MMmSEs0aAI
O3VzvomPdKRkSOvyUbPX+ODz1sOZ7x1Ytpo2+jNm3wnzK/PbtGrTjFi92Kwzd4MqTwKxBMnSsXuf
9KfkctfF+AqWmyoz9SR9Vj3SBBAAHS19XVtbn7T+FoI4qCIHGzVD6mvt6GiRhWFNZF8vp1bB7+I1
Ri7DMMQlfSO2SqHEd2kKuE9wTtG5R79g2/OoSxHKozMJUn4tm3z0rrmKt3jdCcGjLfRRN0kMFglA
vipKmNj5RezryvaUe+3huTqdQ6XQU+xYcEVGrmnq9GCVPeQXkEirxt0bRCYG7KJzflI13WBo8oMM
td2yXaR+RIRpeuXHpQkoEax4ipTo7ZXOYTSgZJeF4h+PlSKJxVIPpGzjvvYikdDG5skzGATrhotw
kSOCENfzC/1DPes+rRs1KxSw2kymiSh73n/iS4snw+/3ouArwTrqUFJRdW7mCq2ZRgHI5cM70/uK
I2O4X/ha2hH1C2VtsWs8IqA0ZaXkrIBrxvfYj/7OTXJ0wumQCajncgrUPZQrkYkDkjZcZawa6QVY
IYp4glOyWxDL63klIEb6eFZub19XhfeECw5+e0tcQ/Vncy3Mx6R9XMwrOJj0Mfktdgt/5IZDV56J
SrMv6wNu/6dtlYsPDbK6AmXn4WAL6/Vhe2yluSjgH/ourlNrR/h9uxRIVfKf8qZpHuMQSUx3tw8O
9LmVQaC1IhbKNaG8Wb8/bLyeOPrzlWZvZfZRBgHulu5xbNddmhyXLlmdTwQ3DQcVZ0Qeb7zcWYlI
OfZEpMy1Pbblm6XzMcIcQjX9NqjrZkvIjWEQpacn3M3RkzCPit5DWbqEImY1aEeiEtGkLXhmYalZ
VBvoGXOPDnZGzW+biyvU2V9GmyEIqjATSui5F7Hw+XEqZqgshpE6PpU/9bEc/MNl+gppX1VtaXCj
uF2tklcUpYTjRPgQVIDJ9jes+7EXijR9897DVDcX/PV9luRwoUC7xrvnX8vwFhHEStozw2MUJ59g
KNWC3zoNnR96UdB+StTltZRScbBW/GqqP8T5im4cW8HbKNYsF7fOn+NhMLUIKFdIpIEshwY/ezHz
TDLB9cMMvalYEueyfD3wULXSx+RIY0fR9y1EqAZgQNntN16GHVgpzGRg8EdCdHC9UW747asrpjPZ
Fdzz01TSiH1rIdNapDMh1vQaqesOOdNNF824Vd7Y8xsGAFIoY6Zk77zdTGg9/pNB3o0XBpFsTduX
V645asdLqXYND1UqNNwY4lJ066QlkpChVv/Pqofexi9DbjzvG/lQMXPXBFqalRA7uAUkbr1/7KqO
qx+K7EiDRKI7YTGMN9Vf5u7uL5R+DLNo8vueZ8V17CyViehVHdFHMX3IOl+bVOBpwBZia3N9rXxf
6po0lR3QZYkQJ//ln0ZU71rwDAzo7O0jEn6weoC70X3OaQ58UxAoe6nv4tEh3DLUC8MNnztto18z
W4uaHHDZs5b4MctirBROufok/MHuJLBlcLTBSAVSRNArSWECUY0TiytZ9kV2vi4EYrheWI0AlkZJ
wF5QwoBLMGA7DaV7kTgOdYpnTJ7BL7fT1d3p043DfFgs4L92uVZ5kyuyXptHxyQavmvSgOa1h5bj
s0i9/guyCT2kbt8COoyhhhzrkVGVhWfPOg22T21ri4yZQvHEhybhkb4Jq1Rp/adqAXSv/636+Zmr
XuLpFLmH0cmR0of4EsCKBnNna6WWdUh+/nU2wvpOELdAnJXD3bantvkpLghPRZ4YxODCXGkWETcI
nHD9IVXIaWXzNCn7WjMVfjdhTSixcFm3g6McfDh+4+GjaG8cCXmkNEX5W0fv+btOUNUtNdNX1d3N
poVCwMh56OKkVeA+zoS6ETseovw+FIUZKmJaSOAooaECKI3Euy5UGhK1lG3oE8XD3x/nv4/9kMOG
nPS6fYibOOoxGNvCIHxIlKkisP42pRpBhtYI01EwxwX7A3ojrO4wnAhAPzQQ2rkO+e8rnoUXY5K3
yaqt9Xnd6oaqCOOX7CSI8viCJWa7VbXEhoU3ZL1AaTi/chcxbPoGCdZs708Nrl53wqw5Ztd8Y5+O
hq0jaB/781e0h9Ast4DZy3ZHFdlu8XcmDOqClCa1beOh2m8WEQ6qlyaaGi+h/l4YGiTNJXhk/sBM
swHty32iDeF81HHd+MRzqiSpCoOeHRfVQSDfXrSqqFgo8sT9RncAIE2b4wB2e4fyHUAeMnCE8kwf
56EIdnqXNFEgQdjI///Repi2T0Ceno7k6WkSHeRE4OzCgbwBhtstyCwck2+avlT7BdWWsGyDapW8
5JHbzOotScOGk7dBr+aHYrikEbdL6G/2FMixneNxeuRoOgpIBz/njv/BDys2heIc85G66RjGkqrH
zTWDM0qRYS2BGL/P5PL+/ieae41y6t/lS00eU4MPoC7RQvtezmm/OnmWVV0iBRfVYCe1ARenBTEH
j+Hxx/zCr1k6ATWt++MP4xgIYGWbGV7p5ODPfRKETezetpCKlRYjTvhCVIw+dbpjiwUND9G520A4
22j2GCysMuRO1jzQUXnOFZ0gh99X7vAJzAB7fNwyqdbt0itP27dzRoH62uJSkSVTWkQpgZxJfNLt
HfohX84Wu4j1S6cIYjUD09XA/u4EjlrTZcs818i2Vdu2h94BE1bxXztiD9meN/PR58puvwhLV+QJ
zmgXc/dcmapfPm4bo1q5LMD71xnxL4VVUhQs01UOb2ap298bqZOEw9x0K2s1TvalYLM8qX0nWNd6
QwpdjjpjS0pRPon8K8uePHP8AJdFAIpcsJc8nWNISw3725U9HvAh26Q3FUMHPaQmTE0rOcw1XfgN
eT6m5pT7vxQ2a7kKvfkYAlUBTvOUT/qPkHRHf4m8Q/ae/KMo0nFZboLRVwf1pLmnKNXcxMdUq8hY
9UZlbzo6amEY8eI9w1GxxUSuVztUFrDN7fGIOgTjcNzZZ70UEUAAXXho1s81/O76nbP6z8UFyz5T
Ar7EottJT2DOX27QrPHf70+uZ4UqaaHZLMTsg8uRFCTRz88WCPH6qH1cgnlLYlKhBolNekOOLeh3
Ub5bd2DNcczO1lQ/No7lprnqViS5g/5FL5WzLvfIWtFRsJgEDP/fPWgg/zs9XSXgGLecHDzV7jyV
mBCtfMvwl6jrY6M+NTi/kuldyEzuCsaK51T1FVM2wmnCXXeBUiZSMYsbbW8b/ITYIbIGNbhTUa3B
jFiE4HS0B3X63tpdAzQ/L22ZD4HpUsyr5cVPEFn1Lt5JFXGNg8mtTZcnuLgUKeGUcvs10+WcCk74
88pqprrpHI8RXA+0wEL0mBnZdZKkmzcDPZtTZN5Jt3hFbaWSfvkGrq6843yfg6bpm0KwEIdg1Od3
QkAB+7FYDG5E5JvGDqDwwT5oQlO7NIIMkd22gow5XpZ2KtpqlK0ioRc1GBgYSM+mOF+Wy8UVLmT5
Cph0i2nYlTEbGZiVOQx98jVPqdcrHdIfe8tF57JkE1FIU3ECls0WCY0qbaAfkleSxJW6dXuQzgOT
bFH9sLuov2DvhoGXHiD/aMKSkgF6vt2qqvSxSwBu3+ueCr85kqeGVVUkGBFGQxtk1HQBa4N6/z0e
XaVGpa6/SdgfASSIZg6BhuCBLXjRg/yyRTssBLiR0tCIMpBj+fsR7QfcCCVCKsEUW3dwVVKcD8hG
4fWCXWxamUc1udmE+MIWbOQwl1olvX/5ucqlR2GUnbjF2GCOc1u9LkqELaqiWUCAjdYfbefLkGtl
JaMPl2lMw0VEnpzpRu/AF7j21GgQkthL09/U803yjSe1X09y0llT8jkzZvDKkgwHy+W1U4ZJWFpP
S4j6yYmrJUO2mt//ZGf5W8pTlHxf/dMVihFAJNfEKZlB24ILUnlVs6mhuPmME1NlSnbMen6RW0nz
CLVTirPSO8+s0kQoat7pN/yIQ2paWIT3UmRTqKquddhJPA+HGf17+zwa274y+gjFIXpajTA0iT7O
20tUohObM2IAaOeF9HYfJTNNiqS2iYG1FdGZjH1xIQEnGodQ50heodqXxXZVzh0Bsz9S1Qxsoz5R
dnQZFhNvKempcN0n4MYOvs70tkkY38FKKr4FowWGyNyRjxKR3qep+9uLTSV2Ix9pmWWZaWGfgLWm
AB3CZl1uRP878l3GFcMgVr/qgPyAQdYLTSDqEHgDTbalMtRhl/YOv0dVun1ioWZW1/JYloTcyZlH
2kwJAzDLgrMZUvil3Q+Ky9+qwI1P/4tET8DUZcT+DOeJfPVwqymEOp/qDh8Ldgg/4wnHV3GRSA7f
k/L73Loi8CJB3YvgKLOUixLIAJhl2wn9hTB5T4hpNg+zFjkvIsYZS+TcnjRI8igz/HADSX5zPx3X
lzXeRa4fWmdk+yD7wxEnm1F2FMj4WHTq6TZ4OTN1nHMVOspsA7ZKkyBDg/59i//z/YwsZ4S9SDYt
PwUHXVBXlbnyx4FGnMieAYEPv4fWEaA2GcHZqHkBntPZEzvfV2GJRTDaMovwiG0GtEcdkGCA67sv
lXL8GrF7eRgERHgQuRlGQBH/fU0MUxtAMOlkx9j5TRvExShLZSiF6l4N9L3xsTZLfp+LlXFGGqP3
CaszryCn68jKXdlRPgXTgAXDJIjXKENe7cz+ThzvuQpI7FTH8Y3xrwOBVfVG1cu1IieqoeyoHcCD
oToHv5iHutUodHIrLuKa2FVA3amXUZQVIWXIWhQ2KiyeZIPL14IrsVtVEVqxD48MOffpuujytH7i
n7kTOQcX6AqFU3CFMOxYK5RSzYq3US393Ax0rxwfFjrTw7Ky126+4TBRP4mtxifQQaFaWtNdhQWm
tWg3+sh03cxXzY5ZIGJJBCknvdLndtyf1Lw5raFQYetBIJXcaexZBT3PjyCWenUCweeaiLAaCDoy
mw5DPr3jbPEz34gR9+1zQ8jlea5qbkOHK1ZkdJmZQG4DrQ6hLtysv84VF9hEBRXXgYmQNtoZDtas
hvzTu6tEfeowwjooa11Cn1WBECY/zjZKBoZlfGTlj4ICIQwmT3dDCnYisdC0+xO6a+a61mO7hmuL
x2r6hZaWvHmgDk7wroVep5UU0mfHipePide1CI572J5gVQT0hkLmQvsw2I0ZyUEuUDWV6U9Xpq45
IxzhWQaARzE1rCYijxatbEpkbAkeoXg/whNkbcKNDNifVFekRKCZSRKwyhDucHKhX4wnIxqMtN0r
sfEn/nrK6HWFD+9UNcZp40u7DMcieRijrnfY7V7TgrvDsI7yVW+HFBlh6DStRTPooOK6CQro3QVD
NIcGADnK3c83P+4syLW+ynRW5WEJ+z3etmhxLSgz7O+UipIKP9AMuOh+Siq9FCnVkyIqemPOkhUF
394iTOtfF9mTjfIQMeUGGGv9xg65YnpewPP36cTyupcOr+SGDF4OPjoCDalBpACqKvUJAzmOZj1s
x1DuFi11skUtGlZ4He9kGVQAoDEJ9LwiP0iTJJOce4LoUrcZf3kpWPGDEqO+4BYBwpmGFnp8/f92
C3MU0ToRA3dHoR9UpSBItqmsS0vDvnahTUpHFYGTCZDPDQm0HCEC/fmp1py4zqpdXV2lBfCIHozn
qOM2EzBv/OV+4kiDjEyymY3XmfthMeuUy/6SeGTWNXhZkslklQJ6He0fT07ie2YX5xIQ9PSy9QwI
Zys+n9v25fQiW9J2rubQ7ha2spKxDmIYLR80IX0tnA3txR7g5idQ5Q4hc+Tea/vTbPwQ2/hqr2tu
4r4yuEQCS19O1rhRdgf/NtVjImn/V4XQFAAcrxtYQD7FQMnin9leDk67FEsYPc7k2bm5jKVuDR9F
0nz63yzm3In00PiGb/BGowi9RjhxpWT3RNdKRtGcmLtaU0BD5RzVZ6VqPfX1IhGmwI/8Y+KzQBtz
8Fy5VKVFzbNC2tnFm0bwFoRlj9R0F36hOzwT5M6NY0cshn3Hyws5q6lYO9VdjjUbBTzsacU4CTn9
+1jrfdvaRHPQIjGWnIrUV2H7mSTMtXasCw8l3Si7lEl8a2mE7Mk2c+FLXteDdaaZOIGPA6QSe6zD
trOEbAwheFZxR06y4lwLoZrZoAMOI14DQHN71ygF5gy6az3Swd/JHYkg9wr5OgzLXoWNKJHU2i8A
Xx0svjLtpI3sdcc18tdMuRPe50jXaWmZO8WE0pyNH0U92cevF1M6bl+SK14TjccgHi/m956PgycE
tGyZkiv1uAVNStZr504u6rz0QFAEoSr+TaGFF0avxXZKdeIBgVm7uPXpc7kBKkSTa2NhVMN+uiye
3yJXM6kpt8uAxrnytcurkN9YMm9iQtrmjBV0eL6byua5bDrNk6X4n48i4yBxpP2hoEcrgbJ3sD5e
qryYfnMrzDux9/fPs4PZncltvBOeJRaOe3tPxUWBVhgiNS3btY0V/ffCdCkJc7z2FCTq9FUFjS0d
W6HgrPcfFTfhSsPrDoSvea5GUZGq31fAiXrYBobmEZmsv00bLgK3VTmliRe7M28jKGd88PhTvFlj
MpFubOrehTxt4iSEJO/d8wLXkNK96TeosLZBh1RagStjQpMPJlOneUm7O+QLFxWrt0GA39j03zbk
oxGJgK2phQOcAG0l89OGpQDfR0D+2LZF9XiKJ2B3/sA8H2GJMNf014fD8KoEzUUdlaazPBFkYWyP
ReCi7+zOIgwd6AiKcK7GSMm1GXODE27hxvgMYMmEETtMOgrKKwVRFPLG9d6Hp1uBEi1mzT9oi6AD
BPSIeZy1/mzoxO8m6fPGKdL/FqwG7bMXeDUFrPoRJWfnxWbjenQM9ixlft0pJkG3X0WP9jiBeVkP
DWbjMOh7mV2eFsFzc9+t/intM34zJfL8WTNDfkDGZ0fUMGfGx+OU5+y4sKRB4mewx0PHQiIqoZY4
xDTGuboiLvMLfwvgArqZDPyTjoiXYoQW7vsO+RMS8k9Ap02X8f00wib5VNtXfxeNzb0gfBE5ATUj
eCZ5Ev1hNIYb6+OEQQxK0Mr5EXuzrrP/AkmpNRC5jZvKZQmp3zwYKWMEaqTFXVUORbRpily7J9SH
5UddqXz0fX+t99WUgNdAXd61Yo4ff16O2X9NvSborwjU6XVS1Axk3inyyo/Lc2dgtHTTQyAovfJ+
ylPZbYAxzpPSfjJgo04jQRDGhTU1zWx3auibapgw6Wo9xp4mWGdnnuScUBa+dGHqBAIn77sCurqj
KBitH2/D++sy4eaj3bqvKvaRn2mey1gKmIoURuye+l23ElaMKJfHvmHVc8IEWA1F+dcTX1d9G20H
3d3z5OwTKefPB23aZ97Agddzzi5nReYbFyn0AVL/RV++CL+o9+oNANb+gAAxSZwEfhNeKKtQiccb
Gln3QRkNTOzxhvreR2jEdKMIuHCybU1un4pWxgUw50ngSD6tM8VfKsVP/5icCoPkcjHuWbauIA5e
azf7CsCfqLdmAS+Ta4Wh64RXzGwMpC7G+spJdDaEsFZT7CtdiLT3VEwUE1ABujkN22clgItF8ZZg
pI8/nOq/dXPWf2jynDTwrIDxl3kfEbTglUPbq8GS+mRbQAcvNEcglwf0OiozbR6eemkv/etZBfV0
62vI1L8M+qfpuCFVTKnUzzl+6ikpomhqWXmbCUtV8TXFwg+4cAu6Mp3ifuqbXt3b2hGawHIHDMgB
ltb8rOvKGJdjTqwUmGxVdaJa7qa2R4A+2Y9ZbJ5GQnQ16WfiyvysQxI3/Ac4gtPS/5coxkVzh5Hh
uOc5ZlvTIA2I+KdTJeHZcwKwUmQE7BG4MfsnBnUhvOPHR6SntONqvb9433gJLL+MVP6GKR/UM9cN
gsFlu+zC7fslZxCaTAEcBk/GBScqaSyxtsxEyIsDlsPac38wM3NZq2+azAmC+/PBvlX3zdRgDhM6
A9zBe7SJENYMARLmuRTPlV+Z+TtmG5ZlAMX2vlxfW2HsUJfBWlzEbQvnReuHrOkFJ47PH8GUizQw
czbjX7jJvwYY0lBOi6MM3bhCUXSfn2+a2jzYegXPiy2A3EzJS1kzvxws/sgyqvOCs+nRBi3SGfHV
u1FYm4wmEqLfJ/qXY5Pf2HSUxhMN1jXMexQxzzdRnIRu0vJYsjcBpd68cWI2qI9hYJmS5O7RBMhT
Ro4QX9V/s34cC+crV/VDIxbjWEZgz/l733ebFaNF4YM++A5vVPXPW0331aSF2yZSWUOveRDlpzMJ
DeriGdX0zdr0ydAuL3Qvawj0TtTBCOMSeuRUpF5IysRE03TUFdWy7nmMWcg2IoBiOUfizZtPx+p8
TbyVjAwOwNdMg+PSo8jjYNY8qKy4biJNKYprbKW/OgeSpSSGTKi8iC1iP1K3uC4h2fY4LQU9Hv61
jobWyb8acmMcoRMWZRPppxf2AoLE5fESKVWi0A0YM3T+1T9Z8PkUCaYx1s6nzkLFpKZuehCyA918
MzT3IZ00GE/jUz6Z/YK7HpYhRYRf7s5VnyfpMJelDXYAOJy9Ueb3LsfYiU0fpByBVuKU+UeRPHLp
v7EH2dhJ5PHudXQoet2dQOIgXoOIMcTfGctaE7JalTwVt/jidhGVBkH3+sIa1aFGcsWqKKn4NkMw
ocqQRxRkHxIXgDNaOTcxDq12hT6EWEsYnq6g0ZVoXcA3jqKBRG0pPNS8iWJpTgTMSJilgKACsP2X
t+jBTchNiv6FM2uOc0tZ2es/NFy4BYnB+oy1xrGZnxLz1irQlZnERXBj/p2cSCLcAPvziPFKrll0
yNbwPCNK1iQ5iSdW6UYbchQKg9CTQZHjOpTYyzVtnANq99LYaX1gCZu24satxeq0Yf6ioU+dPpMd
TuI9Les3wqHWvl8W1UfUlbACZYkhetW1NRpWM9rI1lFuMbtxZpi5GxoivywD/313oRwLrkxuhrws
MsnGky7IhkXhvXE+92vFZYnaEV0FAUQbe7i8p17Hm61WUlTu70LsFxlH0mI36hFrxQK0aB4x2xJO
WzWzzndnGSCSw0yznpjDciGp0+QQ+I7mMwVgharCBCzTAPvD0/0Q4+R1VwQQuIc9PXGZ1juGbp19
Xdjj/Ic/kaaIm5YV7/ULlSbGRBwdEbh24DGsamKvCppnkwaswhtQKbPydG6zirokuRI2az52UKja
LOqgKoUrF1sof2/E5g8cqBl4e/9G8v+rQ5L5fnCqGA0a24huXE1CsmADsa7xdszhDTexP4JKyVVq
jY9Wh90BgzIGOSpXK+a/D9duH+4qEBmjaok1UQ7+BoGudj7ywmSjFMbY9W6tPkz28L7cQmxpbeGz
rXf7HNuVxqy6mgxGQ6o5ILP8ZGmZ633ukZ9kuFAyjQcyLRkYYhSHBC2HyjYIyHQ6QAgQNOWsT0B8
XefpIAy3ZTwZwgVagZEJXXcMJNAregsNyC1sxbvs6XmRWaLygJcKtvqAHUodEuaTRO8PWHyqC6gT
0tSPMXpJJhtlb0bR79gQsXtBrjyo8r3Rv9pgEqVzVv4+VnbU6mu613gT2c1fCtSG4WOfvk6C4+XF
+e2wGbcQGpzq9+wNmrKELEynpjKNdTMPoUo48JCEtuxG1M5Q3M/41y0IHhQijmHn4PEI4k+dMSkg
LVZZBbm+fogpaC4i/8/o69qKl9uwWUa32vN9HNXO+Nkqxx2U1zBF9sznzKxUNE69y9stI9YXzmqW
X+VhRIcLLIhR3CkVknVMRf9QIyBZiZNxJYzlqJkigeYBbMekgcrAfG4jX6TZXgsK1Ek9YBURoo8G
IhsU9DczdzxxHhZn2Jj9tk539qw9VyNT6QshwgBPhY/4sja3fcp/tc8MP66W0rlscyEVpEE9fwIN
e4AWi5HM7qx/UVALtxgMby7F4VskCwi8kwPQQXfhI7uBmqrvnprJJOIOeyM3fumQgIFDyJd07Boj
3c5Y19j5THfQ3/BrASRbjYRyQYNMhpeb+canOnWSJuB0LxFaaoytKbm0IpNtKc2m7qXl10ekT1D1
llYwh3SRg1dDrWhraohkwwAD6HvWx3EjBW0RF/OgHjWMDqRUqgTYTcxMmRtjfOGMF6y0b6F967+r
iNutTp/xkxqNDVytQq5bperQdSZ0u4FyMCooW7fwTCVXovvc6LitzCmQmnT3jyEH92VIOSou1xTh
NEwJYVLqL19oQXgvL5GBTfmQFROGBQpP+EY97C4QmFPDpM5Kc57vZANnG8+SiUTLyjoa+J1gBG/d
g5th5CsXT9SgQkL/mawd+UEHRTqE+mG2BgE/j6TcifxxBhxJCkVVedcq2I7KTP/EaAsnVf/AIRkw
QR5fq2B3v92HvFmpWXbNQCggTcTOW3WLaXFoUhBNa8WKbwxtnsQfvaHCjb2JJwPt6hnf4aUvpj+z
JFOLOxqywf3R5RgyRoRfwyAq0evGFabYgAKfWkjWrEPGshOAdIyLjJDNHqS6Vvfm4VYTtDi8XEWC
TeuktjyyC/KaPJBw9gXAXKqzo4nVyTVAEcceSB7VBx0yAMNPRGkmi1deSx4z544FWXzBYd/5Kl12
gJe98A5evL5yD5+8zUPpA3fx3SmlGnMNSeU2FYSwqEKnAUb2W4r+U0In8e52HYD9M6aG90Z9jsc5
o0aWk3FrfFSF3HO+ekeR0Vvpn8v2aQWakoa1MweJzLoQ0AMyJs+408NLe9GhOkHGxpR3JtxRMnyw
CUZcQAn876zqHkLpY346mr2X7ENDPUndNLgVXIqkY9Cp6VKspjqwRVxPHhJpOZbSYpiwpwlxu60Z
vYWUQnw+di4QKw/ZaC0f7wXMqgd8r7UQCW3g3fJBOVbZMw+Tte8rm6wk38I+78lJwoXVWS9olNBu
5LyhTDs6/5qjhWEVC0XnD4C+ZpxPDPuhZK9IWKtP4aj77fVV10GFJ4EX/5g2T0h4+AuDIRtHb8r/
3GJomR8KXjGRPWKbY/9VJ0cMgs/VTy3kGBI6S1k5zuqJj62NWfDnhKmqdYXzrfuW5Tb0HQqRJ4vm
7Ck1LPl9mLbzorqb+zUn19CznCAjOR0PPXjdsHiOBFEp2KrdehSRKx5KkHm8sJPF2cD9gXhTkaJH
mDbqlzMkOxQM3orth36JtM4T1nWQswsZC+cBWc9Lgwk56nhSf7Z3IXXnJDVcz70vZXDCDAYE3JDq
Tq8J1mZfqnN1WzkZzNnivYGDT98TjORnOwyqzvObkn357s3fi0WiHBdG9WXG0SlBisag5VL5H3Y+
w5f4rKAgQ0ngRg2YF5uAU5ni1zlZbRsFalUPZ6lixf941EoqZKZ2ChOguRYRGJ+aiXBCgGIBRZyl
E3jeQxwwMdP5toOYGuIRulr9zgoWILNqBKIMj5Qi5c3V7uh5pw2VVrzbbgvUvBrhGIgeyCbf6D8U
rr6K9RcW9ajVXHny0HmZUZ6S52yI2npfBiI3qn3Rj4M8RnfLBimZZGZ4h/j4h9IilvY/eZ8UAfQo
dd1Mo3Z0ty6yPl6/f4PkovrI3ADQoqvO/5uNCWbXWGSI2IPt4ZvYDRtoZmoQ0vdFB0pytphbc5AJ
OX1KUcICOYaLDpBbYeh8Stv8GqqY0F4LkB6Pi71bcq/yO5DDEV8tdW/9RirW2Eqi99bCMm1sG0Cd
XLqsxx7oo+Oc+DksyhAKCz5pB9+wB8MFyNc4dzynXDJVm7NbsMn/qFP0qCH+SgZ/fwaj920n+WO+
I1bARka20GqJBeVu/SbpOopDdD8f57qYlVydmw/FtMc8m2aSV3wdRm6dIv7LYqrQEYXRAEobgtB8
0b/E3PGhYuP9g3faU76BPf6hqk/R33hf27LvciOgB7IuErTGA7lTJcFlVMbk6mPaA0DknG3cFZjC
KGegm/UEm9Gk9fL6XN8+bkZCVaR9WFWcfy7LF5h6dZDjtIR94lIjew2xjZE2Dp3+B/gfvZ6FcAl4
ylQhmiAhnzPXlRVxGxntKS6HAaNHbDJ5nCB0SGUlCqCMXmLh8q9JgIobadqrHkU4vF2KZz2NuhGg
5LdbvMBG3EC+LdNiE982jlOivAZXb9z2t+zm9CCPEOpToTJR0BwyUJ1LgDf2A75hGFn+UjdDmvk/
H2Oac8f7EG0UJH8hE+2keMwxT3VpT6XQG3vIC10b5LKraSYc0LIEUIH62sdRGpGF97LJecBDOpca
1NzHGTTsSfoCIGo5y4gy7IEkHA6b2P6E+YeVGSCDfGM7pRKfrazC6HIRvxi4yPS1yccbFyro7lx2
vFXUVSzFGfQju4JOk68r6CeJhgH2LACyPx0gV4rXOM74b9Ln7YBPPRH5q0Y8Poe3LvjgZY//Evb7
wfTN+79NXO0lk2/inABhsXNnNjncxanSEmN6ny2x51v2nBKd4ELzxXSMnfCGeh5pRs2YKcQ30wWa
dpBYgcaM2ryWMBJ/3sSbolU4Wyqu0TN+wR1RPYlQCs7fF6vm1Dbh5E685oOrb7cPVk4r6UOvTk+6
5b7hnabmcY6hybWjjO3zlAwogWwyRtwQetXbFN0tZtEYdcTvj1dpurBF6Qmg95n8Qwxm5jsmxEoU
3mXzLgDB+ElpupJmlipmd0qI46pjKYlAJeSLPuPbKEpN1dVrGf8ca9uXMTd+PR5RGAcQj4jszDYp
tUYfCr6O57qUa+7/XBYLfFRVn94T7yYMEbsXpQa7y2p3oFq3W+tOFntzdFY31hnA4Rr2j4RTEvOT
nQBdqOk9bvQE0MHzDwBQv+lVl8UA0bTaay8easqIP8gPTLWjxlTwXvbmPu/LzvI/kUeThZ8vYPwL
oh+pb46HUV2Nu4LeMyDPurFd5wFjeN0Hviu6qgTn3e6gqPdXDOhEXFQJFedVOpx5+ZL+KLHtUrxJ
E1qOzcg1/6SBurg3eJPyGI6IGevZhdNMEdn7Uf9EWXd1kNpgcMyQwzyTzfNFdkYTfcQ+Rz2sTMv3
TGD1EbDWzhnE36xd2wlvlb9qY9K8LsJlkfNUDSxEmpQhNjSH6MMXKPY57+WfcldCcSBaNrLJRchx
zlA7/quyw6qOGEMB2XNfM4IgIsGh/Jgh4JOPyClQW7Pbmmp/8Wm0sByfdnQ+I96+R7g1ELeh2yso
xlo0WZXwd4yRUkgWu0UlZ5tcR+dD1J+1/SUgbmjvoMS0BausCTdPw/oS0JHsMTfZkeqz1p4vCLx9
cLqlDQK7ZWhHhgGvnTT6Pw975Jy3fBPFHhdVNCKO7miypSvqvn9FEuOvbfdHFctjjO/+k6n5HVa2
ej1zyQKO88f9ZoKTXbY3nEbxyk5ElvHseMEQO3+HUWgrNiZ+AUXkmGpYngryoxq1Yijs0cGDMXqF
5qBcITObJiWIDFOBdUJwKdfkOyP6hAmJsEzEQzQAmahkJ8thYv7UXwNb47Z4YanCyCbTaj9DCeXI
clXAeK8kYUZxx2SjqpuQK0D1lcyQ/+amsuTpKRZy09CNc5J2Vodl60nnOySPoPS79Z0xwq9AyhE1
wMupxLrFjnQvITocH3KhrfHukYv+ciF2nEqxMIqi4fIT5QSlA06DxJwtz3W+uwedo0b8BtOk2uAp
mfD5tjDOp87c5xa0YQxwzIUBloJm/UxC4e5DQ1MEkB/B8OX6BriFKLVWIWp0QMZRVS3+qWtehx8G
FovGsJDAq7ZT9ReFX97MqW2SNo4L0gnSg373tq4JZ5lhOlBO+5s83ziIYIt4+vQRqMap+026s65P
W0g0qmJxrBhJdQZ3wM/7yga8sJlUDHxOpg6kbJB7VTbRlX5U6nCSsXn0i+ZHNWp3UKeCrO0tS5Gm
Afs66bs6+wLzwvYO05UBeCu/UU5atY/PBMDGlKrrQ7VHUZa5jenEBdhhqCufx21Oo/qwvlokjaIR
T1ZLXw2EU5yJsKeHBK+NPaBkja/9HDpSR66xRR3x+3B+e8vKxZi56yDpF8eurX7ZALck0WK4zdaq
3T12LHsIQdxAvSNJ8Y8uQ/sGYve1pE8QjVIHLAIHtdTQLxqweJJZFyCjjcjTp73dOs1wJyQOkrpv
SMfQxDHPcw7YGCt0W/greDKq54zzz02F6QNVpEaF4T36K6WvRVbfj9Y1XqLmkZ/M99/OcSTLN9qK
SZh3LrmbVFJL6l9YvsFd4wHa4Awo4fGuCQuNQUJPWV8Kx0sBfZDsqmk10gWev1fdNUcmwrFHQiiM
EN5YLYK5pKDR5EJGDyvGEjL+ebJm7eqj+Aj4bKy5dyanv+zBJ7Ue4MXBAbZDNpHisiz9/7ZacYtL
RC42x7WJMGdD0dWBK7pnzIhgt34qNTRxxI92tJllLm1uL/S7Y0LN7wiYIKAL7j5rHNZZAUq5B60a
8ZVdk0Z7rXh++m3wgKG9zdaFnCXyyUKqZ+OOmFVPuG1v7I+q5WUD8qOAe/ZtrZ9JkmS8v0xvHRaj
xOSiO+UM8imPpc1ECIaiW5TftUxfaJs3hiuKIXVKSLhs1S6rIOnogQV51WV85kjrH6SFtyQcVAI4
9G0un1P/qt+XyV1ioCgh0x4feEJw9MtHAPzA98s9F1sdtRG3qpd4tWWQdIGQnRxhftVBC/SIGiLd
3kE1K3UqWPhGM7kN/1GnlZzG8ZeuH/6zZQZIXKmFSDmdpAzgXljNaa541KsGO78F55Qaluip/FOT
0azjauZQKxvVtWGPiWRo2iWrMVDLTaq9UFvup1NGJULaDmNpsCsjZiACJnILnSh33y2KqOFreWkV
MlStQvz5neuvxByZK3KE6EPEbBbCBI/Uz4V+79nNximsypvo6fyrkURTBhTuFL9AjIjBtdF+ObTc
BuBUY+aOXYClDHD1O7pz//Qt7cV9c/rh8aV1dMqD2WLzx8l1qE8903rxrTn3crvQowYFPELJSNSH
5px3Pz+Rsg+v+wDLzWS991RT/qY5vvUftozSBJt6bQoNfyIz4NHbo9+uSX0f590iRhB6WltK1sT2
UdJhRXUABQS3pg9rkKMuOepJe/qiQZW9RatUX/MVDJ0NC1Q+ldp98YI1tZLJfURrGTo5DkaOHUFO
MkWje9fTOanXbWM47v/+9QiQ5Mfym+VWAQAupojgJUEucm0fTvmu90qPZFwAWeeffrbFpPEUn7lR
cMrjtWOi32QcVwtNpOqG3hTkCTA8ou6BatAyScU/192NFXiPLaU4yXTaL3WrPfYsoNAg47kdWTpy
/cL4Rp5CINynUAFer1AWW2/OC/zU43MOBlwEfK89zsh6XMlyLCdfVp7/j5dr3y0mYeSaXGemN1Dp
gHvSM/mXRhbEmy0SmuCm3wHZMfakeJ2o+dKFLi/jwEPQoHeiHPq8anFpWefnXEvyOYogVvCpxohV
gwZZt1vgyJB/OnD/DV4WtuUgGDHClmdmM82l4UDmWaARhdsQGTcn4cmQn5NBp8MhviZG1rBz+E0P
05XC/X1Suj2R5WNyRm1G5GEP4SkfUaaPBt5bxxH0KWgdjk4bVp+G7UgsTnXD/nel43bTweY+7TO9
2ZiIrB19tbvS9l6xNJBATS5CnBeHt4h8khqEU6r/vjkDiv5QCrj8iywI62Jvj1MdPvQkvOGIuoOM
CG+T7DJQv7wSPdOpOhew0LKSFCK0Aqpf9puu9nNb9lWn8Q5Hf1lNDHVwGXS+2sEDSGtLjS/AowMp
urGHCv/G4/kFKLvpTCcMfcUDXOWYiXBb6EuOVfttqTL4GjigQSYyQ8B/mUc6VMT9WmWAsjb2czRb
nJ3eMoJfcB7rP2dEy2U9MPyJoEjlKWA5VPS/iNAFf13gLAeMGc8K6NjkcW1k/A9+lJals4YSUMxU
JzVmzrj/BuEsi6wwu6Pf+GKbbWUDzRH6+ohWanPcabXQ13C0UOFaDT9fPcv29PO1EKxfodkGg3dt
4QRNxsxm+WBShg4JtJ3FP9oAixCcJwyEnQCzkxgcfwcVCaJq6mLVL5XOyqQ20E0z5JsxIA0Jhadb
Bihk1vLDn1emY62a1bKSpP4p10xzilVASmcXSYxEZHz3UHoxRytwJkRr6F5Do9+VakkFHYHpJKuh
Q9N5Z/IBIlbwdrfnIEPUCIanhopGWmmflf2PLa2PqQJTZjJLOHo1aMjRbQAZI8nkc8HVgONOzPWM
nrzSxS+TDIoTbHMWLUZJaCkOuMqBBYctmN/Fdp6efW7sGqpg/NYK8uioyCau+qcYXKS9K+xy8Ezn
J6mEXkVybDsTpN6H/qfKE8vh/b9IH3kgzArqDOyJYw+vopS1xi59tEvQ149cCHINIiEIxO2FQeON
IgOaQY/Ar1mEA1jfPMg2MJM6F0P16DvbwoxVeIVOn8Xh/7ly3FeihLJ6QWIXkNxfqyqKlM+fB0Aw
KsaM95zqquHx4ho+5K93udnvdrLOUxuBR0NApER9Qt1/41V9Z0HgngrZrmfRvlxzf1IgQ8EKuq/C
5FN0P3C2X6rVl5EoSzEkmYHlijpMELIkv/1ysbgQVK2JxiSGdoR6gG5bTaF4Jv6xRTFTayCbtrw/
BK/6r/gCHUwjoh3VAolGMNeynkh3bHgy9/0LUO/pvdYuWSp4t0e38acWQL6PKzqvRiME8/1B9Mdx
ofpPqDVMRD3r9pOpCL4sbAtJJDx5VLg8D6nHGkCEJLvmxEnXjl6yJcoAQ8432e95T2lFjMnVMwoB
Jl4xBKCtVT8ax811lkPYwE9YQwYZxASGs3Emmdgnqc0ur0fG6Odt0LFEuspTGwmzVt+UkS7Y/tek
8qwj9nElgUFzxCG4zkMYckfg/4AVRmbspvOK7rVlxS1ltgj+wvyjUc+BPs0xGNTdtMfJLYN9uopr
duCH3rz1uGCCncshJRn7+QqDLo7QW+jQfddDKRKtzke0n77bf3VNP7cg0KyW4DUsXDRck+fPR8NZ
wG9Uwylh3wzu9azuKjFKF9dvtA/ycbHpu1+iDJlq1CKPdCHFvIZtiDDucfM5uasKOwEJpZxqZhXK
XInw1FTyVyBJErbiBVxd1dNUqxFSnivrwbKNkhM1vR9E3DQyzrUlAXFwzk4LKM+UIt0gRC5MTQQ4
t9kXJ4TGs2/Rcu1CeHCqEJ0RQZV5MhGXPhOTrV1qtOBOyRuSFY8UBLl2u2kIjbv5BbPL8xn+8ic4
fI7xRARrM36QrQz7j14RQUUluGW4Xmpr3bQNmp3PIigCvW8GSu3T4qubwuReIiMI1rmoCLOFbZJd
tkmgkjPQKijogs6Ziqf0YCrx1BPhBPBSR3WcFiUCbZ811MZPPOwEHyIEP1nyOn02gXXdXnJhT34I
7rRAfag58dJ/E9/RqnYMqTAbLGuZynZ0MC8L7w9I5l8hHFetHncYmrXoOE135dssx7glFQ3PVAMs
Lmyct6x3RoByqDd5mNTNI8Anz5iA/SyhBCcHpH7lIVZCe4t/jSJVWKPiFdPplv85smEjHRTPQhYB
4K9f071DocmnwA6a4NG8R+yhpDUg7IOQS6F9VADZaZJz7oRRhHsCJA8+ffSRzLuR+VOX37yk0Yea
eugFPvgAQQ2LV9ACe/zd23jKgcopdVKtQQkXIen2xaebYXoJy/m3LaBsEtTpEEEg92P1kVZh1DXk
+1AkvBct7QmtRrVbQBlq/O8bx09l+Bq+38dGbpv2GsR+O/XYhjXw/ex3sRlrX1W4Vs9e7cMGb51L
u0szC8Ed2H0W9hs/Orr5f0GWQ2RGXo8nQJ0Lg/i5Jeu5hslbUeG6/ghX+W+ByPus6ezaS+OWI5DL
gC8x6lAt79tTT4IICOWcTj9tRYWlI8KL/Vp4p1hJALdDBNuAuxm475Q6Rl0OLl7FeSwsR9A7P5Yw
guxmOiNXkuURgk5SlhvT+vQ3rPn6TACjMTMdZpIZgJ89QdYCJY0lhSuM0N9u/fU1Dq654fsw/eAm
bQdPz2qi23ctWLc9vvOQVenZzaHpbZvtNdFr3PcG1XG4rvpKLt8qwnDxNLPg+TQ6mPot6IxUQQ+q
Twzcu2QCu/k6X/b5e30JAu9208ayCqWKfMJcWyk3GgdbamNcC7LjmkKY8dxAO+fYLJSrQCRFJdlB
2hu6ZiCr3/1Qbg9kudG46gbV8Byz5xk9MKiMe3VXHhuupHVZ6w5G7DzdwpQyu14KM4f2dnq9KXC7
xx0KuROtZUcUB8uDfPCzWN+Da6MT5NTq4kPuvbS7hY/QcTpzfBfdh2s0/HBZ5/0W2zbAY1vK5ko3
xls6hLKZRdfbZo0ZGbawDopB7QmmwDJ638cwaaGP6WUW3/vwmTdPVDnBwxwF8wKMbIlUivBLYoef
sEGKR7Btf9JDihdLzVeorVL/pc2hvvLHMAH6hMxuBREb46vYFYwyUA5MnG9wHPULPeWaO+zIz71T
9ZhVSlmouXCPWLtU+3blxmjAYFauuQNPLsU5eKdO2R/dl1AQrJKcmOMaARRbzwarUZt85CgvsEhH
d3Dt6TnJdIqNjFkWymvx03HHyfXPkgYFtLIF5jenAB3BT3mrZXlnMX0AkLKa1C1oYjQt2Gmq6gRl
Gn0AbOrkt9PtDXh6e8x9N6ATm7Na1CJWnTGZPvbeFJ31o13Ih7RHNdNV3cxzoKIhEFzEm1OK26jb
9rs/RW00jldcuLwiBSIV533vKVuMoIno/KatFZtvjcZ2NQmo/u7dwQgS2XQZOBe87MzUibXnAv9v
N7fKxtnlzOs+RBi0dxikVbwwqRDv/kwiMVSrzR3W8oB7JGoDhi9/c+CQxVFPHmFGVwFUEUtszamf
X2lK8etxkJIW2urUsDedCoePdwdHFdpVuhncbfN7rvWbEeYKX4tkizDgNt2Hn0ReakftfOSZJQbU
6Oslg5BkTVzS5vYI6UVCZXIQJK2wuzYckEEkY44fcmho8dh09+7QAaPboZuIzFdNyc5Hejvljx3Y
a5dsRRxo25rYHaF0DZ/6ugyOHVtLIk6AF9UEvvJI9qSRPo2NpFcNtU5WIYTK9yDnknYxFekduVUY
hAN7XB91w+nnd4iICvcWJ+Z8UnpXb+HZNDscZWEyzusLOF0AWkTVxOfA5hxjy4ooxZg7szFDlNxz
Yog41VlYPH1cMqquJ8p53RnNbfxXpb0/BJWjTsrsFhRx0LA3ZuEj5TKcaRTIJ/LbeEChkMSPMZck
/l9YfKX7l3XCoUWBYoFYIGNwR3SBf99rMBpmCjNC4xNJM833Z3IOa6Q65iZG6JU85Sbk7ZH4SN3U
PVhGbB/yXenpY+17jIOlN1zntPorP+emdep6VN+p6vitDO7mWb5+Tce4SVV45BQ8Dh0ZYOEIN/Lv
Es4b+MASPVgwlf8qW/PfiniZHwvutmr2OUxXaTef//4SlbgEwEbEb46VQvs1XusaQonixNjImL5j
Z3w4W65+AfZmWLGGS2a0A5KfZAsFlh3141NT2RSEL29dvUEnz7FhygaUgcEeCHESN+vXcTRnEyjQ
8okHpAWyziRos15IVcQvDU8vST2DBWCnWnZw9p7yWrEILu0N2rSkcFg6bBBha/p3DEFS9FBWaWiM
mdJ4vLqhSSytOT5TDMuZBF/lgKsL7+DQ5Q3cZEZ80EpSjC8DYFBRD1GnWxN2LO0BnkI6ojAw2Yed
na3t+XPUXY5PK+wDaRj2YXcJedzofUHwr7GAI2UE5hhn5zxHQdL4zuvDVF/gBfU24hM7erl65y7D
vEeZ7zHTi/KmSQh7ZRnCO4g9O+SSe8IGIt6NdjoEdK6Mt9AgDWVUkLNUodC2Z+1o1E5YnTfWhKuS
vFFr5xSxApa6JF5QCY/uiju3C21KzRqeAz1V4lK/GnhxyfjIyAkD18mAA+S5JmlOe3NEPU1tqxSD
phnxU5YXRHUvsJo5rsfkVvUegVsXp7pu1sXK7tp8EWX70pu2nokGWlWVAlJJ+TBUXYILLsKWhA7I
NSjLVYqSnEDv2Q0LJXPtj1UspLQGtnKFuFaVLoIgOicuEqce3NB9dw/zxysnqDToDueRbFtZsfd8
OKyt/WvSWiIxgkKEMKN2jecl14OuszsePAsL1/yKch+7d7bBnQrvH6N7O8yhhDi4V52GcZ1AF7yZ
J0AvFffUIL4NCZkCnVait726a1128QUtxYtI11I32Jqg7i33TIsCLE6RdvHBeqnvulLDyiPPB4RF
+uAzA8BP/G5up3sToqOtOm40pmIYoFUH3+k/mXWwCd1ZKJpq/7dLwuS5jJFrrA6ekk2blHeedk5u
gfXxLePcEOFe7+cgBxnkBtiBLUGqS4ifWLTyL1bGMuvx2DC+Pw4XrvrMyF7mmo8WKAIBPbxZUy21
QhicvRl05zBPO0ypHaD+BScTlMFWwmPk6F806fHkesOmXrRCaoOekDPvJGHUHKnlov4DQgVoZ1MP
kejV/OExnMpJD5cp6g5lCKWxhRidKJwDuO1pAwZVjNXb9euHlCnSjbSPfx7E6/BcuvBQrms133dA
gR3V9/r8UV1b4NyzHWIkJf8776M7caT7iVPk5Vx2q8d1R5bVrex2WI4NPdzf77b/KdKI4ckdahf9
Dk4uH3rdtKBGlUWxNVVjhN4sM4k31ofu16DOSFCjXk/OGjLGQsM8gQ4imxm1mKKoyZb5/KOecyVb
WTEsKHbjCYEzQPPXN9yTFob0E7cfEkNoVfbUXyDGwAk/srUQfm4URwdzIQ40p9LiV80dwEKB9V08
h9/wzo9GMfXchk6jNyVCyBUEH6bwUXP9JDNtdzBdAJpBNKegMTywlAuqqIexQyMdHmIJlcASrrys
10X1+hHbTlXIJ+4jVl45rxC92WD68WD5GeTpWtb61UrWAU2cFJZfrcAXcAxDlDmmDcMNBItQ/kqw
rlJzHWE0l+6CfpQzSCClkwxpXIe89lHFdN0JW5MZ933M2kl+1zooGmRMiZ8mNd4/pCYq8OTiiWHZ
GVwEpBKMFRBDEGbrpQKJkcMirAEA5HJulvuQWQYpHu4EBdToKsA7Q8AeWZWM/Sv0nVWpMzqnDZeS
/bGkjhYDPiqURMuNCV8G4H0hvScO6/qhgcOgKHcM+BA8FD22TOkT6YNMWDEuLv/f5FpeLS4cp/yp
nrn/5gBqYfAXsgsuypYxOBcI/QmxFYcXSu4Hqq460uPurwa76FY3DhzHguIHwwvdar2/QEpPq3yL
7uHWUU+sqxjdbcfCX5fhxOnAeTe7P+eah+AE/GV+fFFNH/MchRKpR9Uu9FYHBu/GTk6+vd7/+LgF
RpCnxEfBMXEZ1OZg30cIfXi74fOMg5foSmSONmesRmmiTTH5KXpCS5C09ed2umN5gr+bdkSDPhXG
q522n6bjXmP5uZAmkX492LrtkvufoayIKALpvrMtGb7nq2Hq3X/6q24a97H164LjbOb7R6UiwC7+
zQssXEEr0Wd2wv9Dvt2mr7V5a/RGlPulHtF++NFrmxv5WIrrXMF0HXCsTNwO2uYmdUnUq9rEWTVV
shGwuoByyaA+wBi3swPw4iJRnsJ8T3s2SUCLkvIgxjMesYdomRyDCSZ5vTc/ITGjImgaOwx8xEa4
5bjAP6sSnYimDxrgGm5hNSW1nNkPfvv9HiieENCFbYKna19duv17LQi+Y5phFqHytzvXRidAB2+d
a7SI9frROFzElaJZxD33++PssMfgRsUd+GLFMjLTuXliKDo2sBf9r7GUO5Nz94bjsyjjJgJaw0UY
r0505W4ZtGB/3G3LL4NuEbuT5N0ry30EAdkc9h3ES8daA90nAdyPxJugxl1VWeG1+frglQ+Od2sd
fTOOrKYyR7yrc7vhBtz/VBhkrDbNXVxharT6j8lx85WGTLDjnbSSV0/aPMZujr0pH10tag1rMokF
jkKHHnZMS93H1UksM1dg9hFqasUT9XoXONVL+6UseFE6wheZYmrhuilvruGDZrLgpCuGTswZg/ZM
8ACFZeTZAtRq4NK4tjLBv0N2cPMlJAUcT6OM5pOOAkG5NH9oqOs/N+EYnZwWKabPsYp71jt5ElYe
E+8Im2SPjfDYjM5W+6TjuEyb0TaqS3lWmAiGZeE1mmrikZmsq/nidJO+l0ckFjDSAwqSeHqEmXfi
1bgYzMcHy2E8yI6OigX7/1UR++H+YKwiz9KXUjv/qb0FL/Gw1Dd+fEzhYBj8qJ8+WQlXov7ZvzFJ
Acq9ScFxvso9uy9rVnbQyxTn4p1Z/zU1/XuDwXE932gydgiJ1g3rgjmvlS07X/74bHxg3ca0rzSA
03wEnOQD97iKtN6HRVM/m3UuWVA1lIJfYgQQmOuVk3wQtssnmqX2a6Vf5UE36ih0JEK4W2rThYYa
RHy1outBEt5BbqyoJQ5BHPuFhK1IMlpPD5WV0j2f6Rjgvn7p73dpzVauyFw50ZPvJzV2s2JkPbaK
JP321a+nr6J1+FbQbqyjEQaU9V01yO0o3a92VznrleUvf7ltrbA+OL9wMhIZtldbz/st7um0413E
/9Nr+jO9EeWQw8vHyFZQ3Uz1HOWwokD7YbFUBKWXWyRKmF1znbQgYUJSLou9VJm3U19lDuw4S78k
T/Kd0e0YgWp+PFjce0EyAjCBaSgLDvIYdgRjqN9KT6mQEVj8sgfhnSxjSQu79aPDZoo+DVIZEmYt
QxUknS3DbpX60hSRugEYLXH7w5xhMOBHl/XjiOGTdVKL7omiLRBv3J5ukm4RYfgrBfRwDaaP3Wzc
IZ6q5soSkVxFGUqo3/2C+7YkxQjG9uAM5wvfnnteRiyzQQwdUehyfyramQ124jULSsdOfWGgsrld
LcPWcubZmngP3YrJvMokdcjcGU2m+IxO0x5u8P1J1/kbq8D9SeKMot/MvF9IFd3osgfZ/fsgKtCE
FFV0ny94PsxdpxF1zUoeZyd1AOEnhHX+HrmW7G5SHcl7/cG8OAq51K1JcHc7kY9/rpRNiarY8835
3EITWBTX0IS0eSEbLdLwjfm/CF2WtlgU6T9O6YvLJl9fdPGBrT6WaCO2JHLA1Gl6h0bHM0Z52zRe
c+42y2Yceh9p+stxb6LccbNk3KWHKDNWWfsRJElqHbafoveDy85VPOFZiFnnY61nIVIq1cMmwRK1
O/XQWw/n4h6eqDIyhlQzQFdU+QNLqeirE+jVdbZf0RJI0cR9c7MYgtDUJen05Zdn/9VEvedFSlmC
dzSbOHmx71i3KbRlKHemaAIZMzBCnE37wZpzeVv2Lfg09K9PVfRg1S0oj4i5RLjujBLBQCaUfqAC
Z1bOZfvSmZ3zry+boJ6J+S11y0+lQwUMQG+R9/yL9/5LP55Ndph+UiI2cpgMJVrHhiKwYT0FylyU
tCx+Uu1C5UiFldgPiUoWFUlJUGEFXJMCqpR+3iAhhmOsRfkJ+e6zCa4/821P2g8DyMx3XJe2a7Xs
LbP3jWywT0BSXeTdtURyvvelB2mt3uW4HHtsmLdfoXumUV8J1KcPm0ABQ5S3CQ+FJoxNz4YkFwSD
gja+cYTszHggDdbW8gqLmUEoZkEcua6ASR0YN3lAlSn2jfyn5MLFGskhA1yRjwLfirQ79xa8I9WO
BrT9R/d/0Cn3BdWSy3fMeABR09e73L/Vw9S+i5ennhZ90BTi8nP6DwgdgryYerqFWRG7k1z2nzgm
26anSw4o77ufZzC9yIu0BZxu0/xjmmLEZxQ7LSH8VmQI9i+ZlFbCqILXY+8weSajJ5+kKhzCSR3A
/eWbC1d6P88IMsjVDAsMWrbZI/f76jvUtLzso07wXJyV8Fas3gc43JvzZmwd5ht9w1+nasYsoQeY
Y7WH5nUjrlSeiiQAW7yuCGGSRQak02RgvQ2Yf8P0PllPbU9+S0db2PDjq7DqmROyJSyFBpzBzkF3
0knLfgzU08IhqYBwuPR4RlXw0KMo1dhPTrpfdV1wQnFFgnNOFtJN1r9yWwceLBc5e0W927MqG2KW
d2iLxogT35HS98hlY95TtdyXWNLHiCq46Zm0IYEyER4WS6g0zpkp8K9q6K4RBcVnet0Pg7v1a6Cr
BxMAFajrKAKeRGITffBK07wVgJvwWN5s5XIxI+CGXTM3CLIG9lY7eHTnYJWXYz09C/2+mgMlJc68
KQhzZxpmxd21Rf2GPpCj4gDMIiiDMONAaN+PCSMF0Jcf09aJayqsvvUFpYv7AxHUwqNKAxInVuZ5
aNpG1+6dYHyalNzAO553NX/614wGwOTyo9Hp6Pfom7g0iuGlRhdaHQ7IcyRGFOUKrRf7tVhVKRmb
MRKE6z7mxthn10l0QW84EBNyzDJmhpXqtLKAKki8EeJfDGUZ9J7Bd8o4/veeNrxCXYtudLWPRp6Z
owcYQf86DeMfmdV3BkVcFVNA8E8U3y9s4qNI0drF2v2dGyuwiwUufWwj97NOkmxKWSNsETbUonLS
POWd/aEqBrxWf4pIu0DO9vgqgkMV4DhgOqOoeFACJ4Ok1pvcMq1HsDiPMot3iVnPUquc+OxcS+KX
L63rNdOLxdZH3ViQZGcELUtFk4FgTtnLEqnv5Tr5Om5X7dEbkmuHvxfl6ABDgMrYkC7q8+G7Tpco
W6OTLagfzrvBkTSxQfN7U2SalHNH70YFSZrUhEDfPOnhV5KQ4nbIPQaO7oY4oRHn3CjYjaoL9PPI
Ob7RLOtm/NPUum9dG74kQjDm8JYqBVHyDDEZLYBnL0s6fczplgDkP/T/FsiUguGnGbJLd5c+pAIi
WZgCzCN4geyhUuV78b/BNjwmeKBnBQJU12ttnu4M9IpRYCyK7cEoBlVsfpIgIGcqhiLaM9v44p4W
qwIIxkAOzObe1ruz1+Vc2002nMy1w3DE+aZdEXqC2M7qmydslFyCgCF3AxEMKlx6vyvTcL7zg+v8
3kjC3n3vuudH/tbFUdmOWv+pnZBD5N66DxdbujiLPdg75RTLosQhvZdUhK3V5uzuZ2E4JjVrNsWA
SPz0UX1i8TGr4Nrx9mlsOeNbgyvuSnoJinrrT1qfpcj/hAh0oyX6zHaCMqIw5zxK8Xr9uKDtYMOe
LwCZIaPROSeKzvxQJJb1IbkzdTo68cYob0PcWjEXWTTa6m1jB0m7yDLE+vegwFPGAl57ajObc+qP
nZxuMXz0dQARoso4XEA7gdQ/xuUloWEQNGjX3W1wgIaLMVvf8d3px1EY61wUUbINhsv4uuV4nuHw
kTLPmvPV/8Oq4wp7h+BDKUTgYuktPFWjliTCElae+hlucF68EohFcQLPZKrbtbymNuD9GoHoa81D
Xj28L4IPo2z0RxTFzyjPy6Iij9RHxSyBca/KPAWm5l52/1yF0ZOes4Ezvx8pe/7ajgSyjPjfy6M/
TQxwQDONv74wmpsRtqoU6Ga9lS73ABLbPc1udagoVVN7z1Rom4PqRYbEMu163385o36dLFoCJ3Th
oaK4z8qWBydYLiaC68HtjKVr6RxyATsSH/AOUsEuPiTT/wYrZbGETtOT/bPhF5hT4GFXpiudkGfi
q+u5ZmSy74PSEYQUept44rpaHoD3IWGC+4CotqJMPlJGbxsHg7XZ3VkAguc/jESZju5VM6TNsIp9
hHfpMRpZpht4BM8ljnvmMlasmuP0cbFQFmXaqqa/ojEI+wZmCP5W+DC33Pkb2hTKJ1H0LjhaXzVM
QjAxWdHKAJoOGOZtygi8yK9BuRqLI1w39w9n1/IBkjkK+ISeLVec/88IbsS7B5JNj7CpaDCfNIgx
q3iPCCXmgIaun87PK6ZZ4CRrVAXbrre4eA5yg9jN27n5NL0pdZ0uoKEBtrDUW3lTFWmaypG50oVq
+COLpahY3rYEf5DcP2REpWT+KuWPVHTBSHPSxk//DTrxa2y5JVTVPsZQAXNHOev8kDmPF4yeq9Om
hTskeyYWW5yonfw9p6ZHt1E6j5KqsExThH/5k+q9s6/OJZ7/6WJKy0bRY82ZfzJHed9WvZVlvb0w
EOlBsc4J7NMMC0fk4jjPdAiXbPzWEZ2DhnNYQfjLnu1Ga+wdvpM+nrwXSmPcyDAa7OL//v750w/g
PtpiKDZPJilpB3flNG0NUJSfBjXR4q7LXragixLjlKKNwP71p/U1nzjb2OeSkLZ0O6WwgdkdAxaJ
bh3W2Y6+VjDrFdJluts0sN8QSOoGnEnqQVsa93Y0rFHFEnp4tJJ/1sHjr+6NXMxUMPtjmWOQtoyz
INkmHyZpbo+ifWLsHa026vk4wqp0pKl/RS/odqtttP5ZS1RhyJbt5+22k9YGgRXawd0Rrk0471pp
LGoxtMNwjCAnNcY5wA+Ak9nNKhLh/RBCoqkuhheK2mG9Q9icv05qV/iwkUgO9pLRnF0H517jEz3W
2OSBEPCeZHus6nltPCc/yVWmg6ZtQ5Ta9hKosC3742/07MAm9YXRgx3z/hx4xgaQfPaz2xGLvm51
4MdUGyNz69vmGkTNfQQpf453YdmLyWnIxNy1Ymw6SDk/yHhdOuQQnPJ3wW/MEpU+uXxnakI85vTb
+QDXmSswbdqqVgJcrlL7IiLo7zIJV9207jUja+0XQNrXlLqc8fZALfrEm64bzLZdi6w9iCSnlJTU
ucgBJYoz7K87bO8v6q2vISLQ0Lk1zORzq9uic/jCZyc7uhzLIx9Nv8HrDeSY7z73AF0OJzoFG2EU
/5T/RpsiaVAsObAyfrEXiBOBUSnRyzn89vmwVPx85BAcwTY6uAx8UczatuZQxAsXYUdviLZQcqk+
pSDh6VoWt2l55KoxkMAkDfXDOSDWb3MW0U7UQkq8okS9P+R/atQyTIfRuicEXig6faxp7Ar703U9
ZnjFW8VkyacebHcymuNepV5rrC7UYEzqe8G4Hgzm96pNhbvb9ePiVnhVRshWq9i0wxxkLWCqXRnF
JyR9Eb7Y8demsjMmvOkc3pmFeRfjq6K0tFaX++iUY8O+DjkB5RUes8dsucWEv2WrpztoDaNsd8Nn
veJSp9310J1cApB0rqXx9x9lhFTABAG3F8ATGBvFVXEyHhn8JkjCwlpP47XPMgWqt35eG9R5cQbG
Aco0SC2mduw86FL/OT3axJZmd5GdxlVNSd4lkty3Kx2or7ofi+a3rVsHHpgocoVNcZErByXku9zf
q7r+q1X7MN8kOhlvCQHK6mHD45w4kKB66p+IwLIUnpnUUUeGGxTXiNNxRFXi/adzPDFX5KHU94Vg
H+l0c9mkyYHXozbtrIFnNQZ/L6cL5iXMVmTL/KG8wIBJ7zQzn+xwk8S9Zo0S44zlrRCTqDvAJRbj
3DNuSX/rJ8+eHOtZxfZ9C3TgfrHpeoBIu2mbGzIPmSL3s+SukxJ/1FcSHjm/qi08I+VTFvU7543s
rilBM2fj77ecQ7HV6+8EKeB5KnX8hJlRNgo8zsLSqpWdnLH2GfAznpGB/We3ifEdsXUZCS2xePnM
PUkDvddMv5TkWaAzbN53yFh9u2Wn0FOTuzH67quxWvHqCYtBpAPcCjEtxq5/Caq9pwAuGQRoyBPz
9FADAMYK1CNM6ugcK4lmCLwfQQ4tLGRN968UblCvrQYo/isnMDglurC9NO3Fcb5x8JZcXq71K9vW
AhDh92AMtVponfSOyFYHnES9wUzXwcgms1as1F7Bbgf+gPx0GLSil7Ze1oPSVSzRzpaRDVnGLNRa
H02/3ojzqxdaswVjmdj7eGNBfIMwVlxMMoAIVnUQ9+4m55RldR2nT3kC62AxrXCjasMG0oF7bFM8
TUnFK/3HNs1bNpT9tF+NcXG0IRDBEM1l0loQJl1OADB9eAxfaXZQWh4wsC2ZXHh4R6lCgcw89Gx4
6hA95rZcOZb4NBjcCmC+54zUmmFskjWJ4SYgEiBVvVyThntJR9neaL+kCP/cyv5CCbKy/mPCDr+4
R+q7kma08oFV7l4SoqsPaC52YXJkM1QRHYKYl/f0uG/q/vyWlLif9CKfe5qsTCsCu9JEx5aCthNB
T13ObhhDpMP+dZf970D67hWPiMMiul1KKja8nrq8seHgEX/mVOJLma8wtW3019NWw6bQFyXxswpo
ogs4eGbvX0SHJeQ6LGUxtkB4z5FgxvjFJhjbSniltojgx5PuJTYrUQENBsy/OXSHlu7+zLyf4gVm
2MuZphBqP52qF/nXZaHA5HDtJ3HFKzia8WrfJCpN1nh365t48LoWZKGEZu/Urj78rf69MIwaeeps
61h7yWpyBAarX4TRSmUxGfJ/EsjmCzjf32f4u79NTr1lrAJjQq8DUR3dKQ+a+6KZnOEY6EVSTPdr
23rp0Lhq63fyzUzNmAjnajPYckPHjKSdxHA017FWcSUDmUAfGdmASYQgN0uNUl7uEb6tUYoewfH/
DHxyR2rWExJ2JX9ceZ+rz/SNX6U42PS64jIAcg02SQdm0rjrcB/c788PSBriZnJD0upfHXwFu6eP
idSXEPIOGMozOYl36AwzFzy+goFYQXzT65JVH+OtXqNhi5EQqKPFu3J2LLNhTtsgmtmuAWNUy+cF
9tLk0Jly1q7GHti7FMOZOVVH17oVykPScv/LGQ+8L7Q6z0oC3Gj8m01xO/R/pFUG8HefasXrz6fY
y6AzsFLST2bbAeYXXyXPvnsYd/79xnIOYee9EIgrjWV8aQQWs2YbUyKnCOqAJu/SeEjJpSSmk9N6
FExmkV3zKHTYxC8j9rabjuLhIU0K3F3Dya86KT+clYP10GfWEm7mh1+NMkBBsbbXwRfUEQlRrizK
5W+r/Mo0SqZpB7wYUrNoE9gCyqDcnVhkN5AbZ4eZKcW629zolwiCz/VWdnVjFDmZB4BSOwczqAn8
aD2WxXyhSU2myYvDJqCar3iyHGEfJSKKTtcnIWy9ajahHqIInNWXedCePJubKPkcpGg2BViBe+tF
NzAzNS6Hh+dYHkVv6shyjuIIgQCZv13cVJITFq98dJC18z/uXgvx3xAyIklE6SG7Atxaau/+jLCl
BRHetoRijgj5q6dltUqwbwM4Y6b/Stg3eflh65Vg/rs2rT00IeBlRB6Djs3h1RQ+xxEWzVY5npcP
H/fNb6QfsA+hhiddxCO4iZTH1mDJde0rUukG6WXgZrymc9l7PCxR8vQF1Z0As0WfQukEeWEfdEGg
dh9FnP9ZOYeHxbcW55ulZkaK5l0PZ3AgS/VPnZbeDONRx1NvxF7d4Uvvm66/Oz92LqXDzEcPdnZj
x8qwtyuUHF3PUSIbgwYmBz3NudO68UytIcDU45QWEwsrExSZiLo5SjqgOYzgdXD1KlrllLp3MY25
w4v8j+WR3nWui4TNtiPyUQgFVOlOi1SxT1yZWVjBuGoBF7x3RATcViZGqCFy5ZuSCKL7o5Eppodf
FoQpXPyU7gd6zGgTLc8HmT19vC6l1t4ddTI5RUO17OZkjdBWh40MaRnYT0JfSRZJ0xPELaMdgkEB
nytLrAtfkZjJho2gYDPrJMo5ixSq9mkgxGsxFFKtDfelXR2j5MJb9DTNhE7LQ73Cr0mAJ9rQPsE3
zHpZQLc5xkXy5YreaTs1L77lEaTl51WfmsdPYsdXrCI8T/FGk7WrMlqDOZV0jxuGvV/9YfByHwLC
d2pT2uodPESaKahO1nP7aRlRjgeiEAQCZzeIQeK2DHpiJjcvBk+atpPuVGGXgucMA3t7zw5vl3il
ND3g/gC06/p68Vq9T/eJbbSQLCHUrVkUVGhc+X4BkDI06eTwBHfvArq41HvNZe8yG+YC4uYQHUhE
TjlFhlzJdcfv5mccp6fLBTqJFxlklJtG+N8PgQnKV9mJmeUf5W72Oq5Nqc5WrK3cPv921whn9nqQ
d4Bmgb1q+eJz8hSDQP78qVMWG5RNqF9EalleOHKTG8G/hgTLoEBRAgbkEfzZrEQKOq55ajnQiIW5
6+lTVMHXwY5uQMtD2KWcjokoVO1tOXa5hSdhiaeYm25ticaoBLn8K/j5RNDR+C+qDQ6d+l5s3Rhz
9JmayMS/bsslZyOLOi/F3CD8pyOpdtjxPFfRG7VGDXMI+1EpbaezNQDKOG1duw0bKlQjgCnnIEQA
pRsPLcXlu01lhBomyUxCVli6Louiir9t1iZk+j2EccAMJkroX0kme/bnzbmGNX4bwi07Vrm+jV2s
0Fjfg5hC59dHzX1x48aCdAM+MwGqM+eElF6y6DDSFE0NDXNhn/zYp/Bj8xkO9RdQrzokgfWH9Lkt
XREA/668ZeTW4cyJWUJpfeuqS7RuIqHM3osFWZ3Fk1MZPu3tXgUQGO8V7aMm4q59w6sl46S+djC2
pIvY85mrl70kPh7t/frH9hyc0obdrAFdU4O6Zz92LWuygdc6nkhcHJAh/qzVy92xXwEWWkvu6DTC
RkpX54qqDkMkKdV0+7yawdmaa83XMgLK4HmbGrePSFj9BpTWdiKKDu0OPi/uMrJJNSBy7sz1VdIx
FxktEJYvO4A+JbGEYK4nTW9SOLMsoJxDL6G60Cxp7yrkUSY9D8YI1KQ2e/06eUYjzafRYBmBZnXB
R2sfUTtu3wp2+Du5cpRlZTJiAdSkn6m+C1Waru//Y2H7ACp80m3Ln7UfnqEXOErrbY1XEUoEEP7S
qQDuQ/uZPwO59qtfJMLs96eULQ4z2PP3ToQLrhuXCBPJmeI5I8Ih1N6ppeqDTaHqC3tfJ+2AstA7
Bdn+EEywVYlKVC1juHLE+KNvX+28NoKKuIB3FNWX9b1fMtZ61Y+HUbOO7LbFo0cAkpfzIpbHpzXa
kYwpkzSMfLFfJgRE27GBh2oV+pk/2cDEOKav7SZrFOBVIr9JkxDYZEyWaRDMITvzTOq3j/LbJdq0
wWsUFY0KbLi/zyoqKxteL3UUBW9AzuSxeAHU6xOjXgpR/czGcX0sKVAiV8eHDcVGtawN8oVg3Tnc
kb9zCy6ilnRhv6fg8KCKyS69eCMBPZupYHbpRpHVBVJmZbMfPdwpX9w51ejIpnbJDNyLTj669nHc
uPxjed5+VaGsT+lZKCTOAuMpSnK5NgoAqZ6mf2pQQ5lD4h6D1XKdQ2BH+/ZxZO4pDDyDNhqcY7/M
+rdejh8Si+W+i5YNsLlXqUS/L+56T7fo5Ioa65LgS2Kho8j9McEzpm27yiWpkuyJPJb7+ZvB7Sn+
sJpxUyFrJjNma4lq/mfXufHSUK+bg2R46xtnTChVf21Hg783cwyTTFIPf6McWKN7JVbo4nRYJWZD
lpHj21+FEKtVl5EZy5b0sibl7nnZ6gAwYkRFTjHQYxun6B6CgUEoHaf6RuFG1NaL3aHROVdncBBd
03XWsG+gzjkKcJJnIA2d7xuE2ez4XiS7yNvrzJFm4vomFcvAUK1wTPjyW0bdMXmnnxZMgzIEezO/
ItNYW476HwnGtov0+CekCkVn7Jlu5t30M5F59jKmk32peYhzg7SXCHFkItNfGrgVkXMClaxM5kWQ
Gfzbzs4kj3AgQZ9cqgW9P+SytqdaUWYT/3XfAyutU8RP18MO8JfJJQ1GCdQfB8ah5aijxs1eCjCL
lYur9qZ5lvgfqmKdK/l82cSSg4CH/cSCdOaB2mcOSR9NIWwvVGgUwncXEIqceDnVeVU7MIXAf/h0
pjI+Hy+MkO5cIqXP108LrlBGfv3ZbYTyQSESTe9v0z5HX3aX5VhZ9wrMn+2d75WiYRfng+qJXDK1
gi9vfexU24S28bA8ur8xTNtvCQDLy4Zx8G3xfdRnd70kd/a/qwOfy8Br0B3JboNcDRDhjurGA+tx
BhTWglC3JB0fqIwk6FFkz9zdaL5UOS3HZtpikrDEscV8eqAhw0RQnTRuErvqsPJCiuuEuyX80Ual
FINA3nA78ksMny95BmEIzoX0eqrC2tBPTYLVjYBoTH3kvC+jkiCv7Sy60Ne6Af3IvxH8pbNe6ExQ
Dh6jAP2igkeFmRZc3Q5HYFTsmqFKM2Dnu3vFbuGU76ihlGpP/N5aV7ZnWdksJK2DLFb8MUYkfcmQ
7rOMoijajWp2vqUOETSyajWDq9UzqkcxbTqZnGGb3EljqHaLDZvS52/vnc1i2zD8egVIc7KfiKyV
V/X6bEkyUbLXhTRdibtZzw7m2Zt5RPHrGFsGGP/FY0EBY51s9i3TjYBWy8ebSPy6BxCbslwpbS7S
6ZyQU6SinT+tDyVbk1enJ8ulwrRVqG2xUUqWBVS97u3bQN9RXVm5otP7BmmskTHYeyH8nYBKj4vj
RX9Qu+FpLR8AXYgV1lME9QJ7Mv1IepXxXR5IId10aivkeBnYyt1CRqe4I4AE1VHDKONhy0CVXtlx
pxAIb6XeJ8e3m/2f2iB/L/9LY26UspA+ntX+wupARRqLo3dFXv0JBaYqhL5DKgnjxidAbM8r0qol
UWobAMG56w7Y5hnN97y3forAj0OZNHeu2UWiAXoHSL2qLtym2WHAWSQMJ3uem6IExprgiVGq3OJ/
T6AEF4WPtheFwX8a5hnh5PQmHvYbQ4XO/3eUNVOWW7txmYCaTXOkFMCp6SAiUCiA3OONEiDUWQRt
yJ4CGPkBnUC5pCQGzeb28cU6wQQnoYV+hknAfyL0/E8EpymgbGbn25+l5BQiTJaZAgsKZPW2GtLe
ctmYIy5/24Tz2K6TGs9oSkoVjz5HnBjE64b4Kv65ABitrLtiOj3akM7FFHNNPU0atgkCfrQWSBhD
R8B045pMmzoyfmoUGBtRKjJRRvfCl4I1yqYw0NA9Avxta4E7zWSqsbxthrQo+EqOf+ZxJHWF+mRo
O960V8ntua+WVgWIZjaoGtyq8Z26O0zU28IQbqAuOZ6F6xraHbsgSEFYzZNh+RxKcC8XfD0+lwr+
rjsDUnS0swKYlDO+NGJa+cjVAcMTigly3xyvqvjS+yG/muKC9lONVmBqwIJslLN57yJkRmv4fkr9
6pTskjWkvtKGCIk3ZTbaiIE52PA64FjI6pZlSyPtUDtdk3VWJuTSJF6j8IDFAXU8NNKlflDCTn5x
rc/zDENboY4UIXirQ4Eiyy3xykgT9dnQbzwO8Cl+Ss3cVRSAgK8Wgb/JcRXEfJvO5fKOwcvm5k1u
+eK2GzuMfAMB2w03JgQTJ7S2jTv1gAprJkIG2O1F2lD5inaJYFZv4bCmjTcQ4hhUcFUqFIrKLUiZ
z4KPLpCIM7qz2BeVZ7Im0MdhiVo+tUrnwwkmP8TK06LT4wmt379KkWz9+RXv6AzbKWS9D40+inHF
rPEoeDCWuDYpnd5PJmJxhfciCQVMwKX/u4rkkDfsQLBS0zFr8RfygGDqQVN01Rl2yR3tE36n6XPS
TLdRvlWak1EKJysRem78Aqi5o73/lYR4TYTRPylYvjuFyjCnQbrIweSlEfMa2/45vvUiHw3HbTZW
lMZdhIXh2B6fceueujIBmSe7raWCi2ABoVkWlR1jov0FdPxPHnrHxMAD7p8HAVn10+jfkO28mWfT
qIuEmW/SSxcWA4UnK9KXvgDVwPTI11sUXkPNSZbySkYTyOHy39LY2OxrABm31FiveDla5oMr/92h
3n1VDui73hD+ifTzRYpK1UD76ytmDjG7LLPvAelb5l9A3XAlr1i5LYzrfbTU+iek4kAJY9M86u1a
kI5osQ0vETZaH2MLOr0IAESJ2s1+UnCDOmQz/yW1hD5PlRUVvYAUtJisW/5PeG4q6pQ+5Yf3M/7A
JabWNaVlt0XbF3limMdgrqMrRVpWRUs4QXQCb7gQHz1g4yKqOmb6/Ajm+z903jOUG8YvCOCDeyRe
NRYbQSCb2dfPmXl24nIfjtsZND7B3nLEZmWD467+pRPOzfpgUznIAU9ZNChjH6DB9XSSMdotgVk3
wohcez8fIZZr8bmimubbeO8uhVyRaOM+GpXCjZ8um2Kloa7JDbiVjLMHsKRUfc6wiBk5NPJcvZQA
5UMoB4+jkE70PrCWoQkcOM7T4N909lfNk8ldvJ9Ot1u4BXN6DHe66uTX4781NKlumzZJn5aiICNZ
dgAcDhhkl3gcnb9wF14jsDp5Q+A96Ko195yRk+bQ41nr/XmBt35fblD5qMMnAmx+bwS68NnpMYds
EQDvVqdz7BxUliS/bg0kBllkzjNNyEvz+91jnZzhpflSxuGPOm+OjypsOnf0AP08VCMxVpTr344b
UDL9rAAmPtau/6tTLxJnLEpy3nh39U/s4LOe81kRhhhY2KnfyXJ2szs24bnMQ3n6PmcGfuH+75ll
myZypITdjNRAeJO9u+BZRe+jlOcZJEkD1tDpwyokAmgAPnJdHOpzMGJBm3qpw1YJtuzMvXwZ74re
4XXCiEZiC0VcCbpZyO/K0R9PyDP+yqO1W3F/htSiM3X0N7NkgdctgqWNiyzP5BEgP0fvl4+xsNLK
EBXpxSg/9k7AvnMR21M0RiXMUlJcxP/e/IjtGLSTEvKiCV9EMxSp6YeBFdZIkOcpQxN3noz8cyZ1
dMIpij/3MHaAn053Y87HoYOJFJEAawMk8Jp21J5WFEm6vAywYy9B7JUtY5qfLkeyaHp14yVxuT/X
gRvpsTbcLhHRuF3VZa7DmkgBt7g7oauwBau7+76q4LkUr4ZX9RJ4lRpHoBvf3g1e07eC8BcZgBkZ
8MasNpmEKQYhiIKSyOP8VGE5mrz9R3cSlUOGPTOD7+rLdUZ39GDwGbvlZz9BVBTkVciF8EIJkwic
bNruK/cZ9N+cnDr/7u/MpcJlGlIuMqnM6B4dVusELeCyX+TiHJO7Y9zVA6AeA17kmPYQDYLAbeVk
scChfcvIzNMxScyBZeTawoANwXQxdg19oe8TKpK3cV+T6+iza9bRyPayuygft2QA532u3sQ+35Ek
8Y94lEk6E0t5jqDtzPsom6rWzExHbs1C1g4DeXYph5A0jTHCf3Y5EryFdJJ/1dafCXkI5JwgDvDN
niLmS292MlKDqszsEqyXRQQdO77ADxjQGnxXcRcXi8O9v5KaEfcYwL0LlX9k3LcqSMdBrmuBrKjG
1EQ+rCXcC5AHwgCLYFD52GyT0WcweI1TEaFWCPPVN1sStkhh6k49SKxI3/777IfvwPdT/GcS1dM6
ffERehTAQJ/zyDxlZ1CSFG/jqws0nWrOEm8OSUAEsWmQs6rGMVojJgTCgM40mW1v45xHJN6NaZdo
7u/ZkkTlWYauhaPg0lgDcwbE0PJ5UlMhIhWTEvkKX5MVhNOgs1w+OGBZ6faAFyKJ1PN9fPlhuVk8
hSKlBXU8KwnrH+co80+xZhUIMQnFCKduq8ov5epYg6FisTQGZgaJGuJSgM+uWKuY4IJQKQ+GhJtn
EZUEwYu9Aqp5OfkkV7ssX+q2NtzvtgJtxK8PHeRDFYyFeZrR0QJeN3mbGxtTJ3sLNL7kNDDFgTaK
3CaCw6EasAp+UcLpzpG4jlVtsqleD7u40SEp+KhQGZsuIH+QNInRZ9gok6EsGbS0F8FxpJAslTvh
JeqfxVg1YcL/XBgDRCzV0KF6fPY7TuGUVwnQEZV9CY8mfqvjIXsusR8sTP2hZkkHBsOEDDkVoZ1m
xtMoYVqSF3gTgwG14/QE+f9+1MHvdfhUSFAHWl2LbPoLqpkmcFSaHjfPcZ4sY50E49UCQ0LQK6BJ
uFLT8+7EaLFp6Tdvz87zNJsUeaEE22hZe0QSh+QNl28ZqYqYXFxd70yN+giU++RBw/VTeCEAW5ej
yg57q+LdJx8q3/K281wH8Xe7dl6594cc0OG0kOrWKi7EuGJj60zuL6FEgcx8SsnQjXyvXdC8sUoh
xLCVt9KMDu1uYsOlGzbB6GPeVWXBFVqFX9dFVNnfG7B9gXux+5bHPU7wfs4te96kUtlWrXmfCrQN
qlDK2YvOw2hHEBNoG+HM3DJr1n0zfHlrfUEeELDIA69Hij7l1nh7zyTysxZOOMOelRiJc3Qh6CRu
C8I04xQSoJ2HMna2QJjoCGVTP2ohWZAvJ7xFwg==
`pragma protect end_protected
