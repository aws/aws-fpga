`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
GErs8ILExhBbCwX2uMtuwOkOb/SvW4mHAPRISHydsEk7daklbQ1GMILCp9CuCU/GCLPJmWjlJl4B
XdUftho0KoU8GZ2QriiLURYsNFAtRB08HwbdnVtTHwM72NLVNOtDse+7Why4btoOmpSPdqHUbU07
NSru9umQ6IplsrJ2Vr8eLUOT8C8nDxAiHKqccnCPAZfN4iodCRgVR+r2tnzsqi+Q22bIRJ22JGAa
dXdW4XR9EOxMKMOt01tll3KmYUy52+F/Fjj4lOkdKQpFdwd5rTuwSI82bbsrCeOa0EmtvepJUF95
IdQEmHcV1TakIHi9hQUgRbX7uYQeuKixhj6Tbw==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
2oIQt5Srb9KAM2lvH7HD3DgRuP5Kpd3fCd8AS69Hbz/x2hyZmu5T3wALmxP2zY91l6Tp/pyejFMe
Tco7eAOYpydfPJwD8bTRXiCKuuMWB2dUX9u44POaPwS16tjAQlKiUS0SwpFbQNZpSzqI3opka5mX
IPBklwN3xenMEylnWqI=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
al0u0pE2FNme6rtQwj0WAl3u2rL2cc/2j9ny4aThgG54kkeUqjevHGBLDhkeQDxqCebEeKc+cdrI
yFiirk6CkEJcKaJInJ57eI5m3qll9qrBov6p0lKjHnf9DZNrkizYOuQVsxATrwWVQvEGH1F0liQn
RvLObivCZqkdlDn6l7Y=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3488)
`pragma protect data_block
lqwE2e5xCmPtX+LKHsYt6FfVSJO6exJgmgGL0ozeMP7pG3658PPAufemfqJdkJTNKSg1ryqDaBzL
+wd2YdVOwIvi3UdXNZqnHeE3/BI+ci+KU+vKa4tNOyT8EZZ5MLunYOhww8rUSrdOOGk/dDTx2FS0
wiIcBBvQI46JjRDARNf5Z4whgxaGN1AC6dZChQa1W1ptIVIs9JbdiNbsXPVGPhLaT2YAxongw75s
mJsuSWptA2XnK0RUx+8GOmtgOUmhYxQua5kbFHI/XHFzj/+l+R4U6oXKOOoX60r5Y9Uy4mZep112
yfGpTyAte9CU8vf8oUaa29nGDaAQUxhFz9QTusme8LEPeKIHOOE6P9tQ/rl2QVUKgaODpS58Ieoo
Q+lWtqfTf+peK+ue/HPHT6EAf2Y3ORRR79uYWjJ2/+GNiOGESxJ/yKRubNBxBdTc+jTa0Xc0q3Sr
arVLBOaN9D7MmnoAE3maB4jW1v97Lw5pCRh5Llx55qVlK+ySzEjY99eFY+dITT+GorCDc4C0AUl+
qr9ACk0f5f4lNXPhklsV1PG86+0HErPzX5+mooY2nkUGpMwUdb3Wuoywxv6/wlJdIrpeWsI7sK4o
UaAiXaut4ojYggbkjQBva6uRLnnyuEh3H/4a1NPeZG7+t5Zf40X35NMs6D1Ox2cpoctWelHf+9uF
uCcaXIP0KLOBZu6Ciz5gJyAJX7GOlLdKoRkaY7LxjhZVKh7E33xnhUDba947hkKFvGFXF9lQUDPQ
1ElQcf2I/NI4fXOT6uSm8x6m7AEOHmJaY+OncY/DsjCzpZyWZGpecGaSQPhErPptcu5Lh5HUXwQO
OFIIREJaAWrCP7xMRZGbI109NBqvviEp6AAkVZ8bTW768m9FWoClmIeP3kurNUUFETLywyXxHjcz
ZYDHlEWGtKTHEAk3dwDQb6SSk+3Oejna/5CNpAZI/9pLU36s0Gslg0r+ApDuSParxWEwXaglOMCV
zbqyJJZJTJNwRSZ2wlt1Lrin0H0Z3OpLvreawtnCeWIFyb0jPRh9eJYiFlNou/zdDjSW7Ax4V3mY
SU8wnyXvV/WhiYO9Cz+o75dtGCv1Je/oUPJeWpuYg2xvre/FR0ayDQQQCPOdt2Krbspd3kSXuMT9
PiO3Fd7wa+pyuYudGW0iSEhpZh3ableLPYdfxDItI8vtHMO/pTFTwy9Opf5uN1mf9IstmBO0nNT7
+wtWq3IL9XvURIGnsPiqYb4nddh0imIwOkIeBhXJqARoMlguPCTbJux9uuw6lMPezcO09TD+f9pO
IuPAkj8WU1bKo9GoTaOxIWqkj30xg9x0rrVZ4OGMU0GiO9HbcOBW4IPKK0NwKVPfwSvyIXzmO+M9
x9uvMk0LTcIxlsAnmOAJyXDu42VQe8scLVCRT/xJmoy9+kz4H6G6tnP3TUBwtNziB/j41tzbek6D
RUsQ8K+Ax/qsQsCMzd9DIGIdWXKvA+TFfwjyWH+TZ0TuA1WkWSR2/Nyl2eP31X4T8k3C3Vjvs3Ro
6wwE82xG3LeaqAew4To3s3qs303HFaNlkQpIsKmZ1DDfzT/dzWWxzyzwD30eeVjGXxdZqSti4t48
VnijZNRuQgl9rP5rZudbkIvXAibJ6InBj1LLz3RMhheUocKdWJyDVtNsCQwQ+oS1G4LvSTYTeNce
NAqPRaKPwtCGxqC3WRSe/6y+Fni+ZQPH2HAwyVyD40xpjsJJH30ZWrQlDEcChNaQXXljVGJ9LIat
yMr34cHkUILs3d5OPK9tukb6ZS01nO5fEAfBYA9k6Z7zQvIfCcJxkwmaGdqteXN6M7KAjghKsVbL
NMxdTLBU2Ouy8rQvLqC6mHSF+fK5wGHAkYyCueMHmeOH8RlDsNebUascVJPvQE3tmcZV6pbtwAJj
CbnmWoOANzogXNw1B7C2Jj8TiVGGbfZ9LEfqvwulxhVJV6wARO5mgPwgvazLwXmjmAHixxPrgKyr
2ulTzoAoVzKKqJ65immGK8+KppdBudIbz5vPVSz541WH+tiCN/+vrmdt8E9LTOiok93Qj6T3moMO
0x9uErvUrXNL1dsZeIpybx3G3AeUBh10NUqZGC4+pnMrKpgouu+4NFh8GGZU9KIKEibHSpJ+8n2K
AzWkzTCResqlB2rZUE1+q+Ngcj/5o5Mkq7F9WE+OzXv/SO3Gn1f2j2Ntx4VA+9sLE15Gqsgc1/G7
wpaz09qfPe5fgh+7gKN8uSRl7b8h2KgMwkqT1dwoLvz9W0yDDnLq2/fPLTC2DE4cfBUo/Fh8O6lH
FvYLLmoPlAxAA59Omb1UuYF0S5VeOdX2lTu/AvDtevFphiPC3k7PmgwYK7gJQrkL5E4gXqPbocah
OCNNolw/J+uOYkxv3VkC8KF+h/+ox3Ca7L0lXMAG2ZdCHEgXPdH53LEIQh4dDeBRyUpC4uBjK8YP
UlEmfhOLnTz0WStpVGRO72B+Fmcm7V9ZzegIU6X0ElChTuj2xNLPqu7SRnFEr+KJV/R0CY+0wCUc
2cUb9PAvWTuT3eFhGG9F+l/or+Hv42F+mBIuK9vdn0w/3AkCS5OTdT15HgfWNTh4d/xtEsqItvhn
vwgo1/MhBuZlkjAqBVSTw3dgPCmbLSgW2NcHMVurpzXHJnN9Il4mzSnaxk18+0ergRqttxvNegci
C+BTJ4aNQO/IboVg8yDbeDfH4D3lMAJBCGPiYAV6K1V2RI8y8EPBPev+FpA7D/BtxhLiV1B/RMLM
V8G9KInMMuNcNLNtKqRMYQQcpTNH7eaVS5q08aiuxDj32qW1l8y1P9vRkr258k0ayDWIoMLoJq17
eHBMBZ+0t6SV28Pr1W4NNSFwdw8VFRAPGfMd15ckJMUm1audg2m/6NFaloIPIfD350az54ODyQZR
AYzJyiYNpvzQNCWJrFF7TksMj5nUlJ2FOwYt6wWyYQZBeO4ZPmJh1zgcfuldogTZ7gIfILmw2DhL
gBozhLxdQRvGga8PwUwv5TyxlH1bOnqH2ztEpWKf76p+ykU9f9aOjzRVOL02xOykGlv1LFvZn1Jh
r+i2ZOt5npJ6vDNXDrh4ti4RMbKZKvsODs72EhxTtgvvKxSqaEhjzGu50ZF6L9Lue/11nN+b20Ec
zluGqATGIs/2hz97ZjChjBhto4M0duhabYPHwvCADOdeHa8E4eg0zuCDZlsHSGAh+dyjzO015EHq
N98lQSDLW4+ViZDLTQNu6iH2ErX6MzZB5N0GeDx5HrvpgHIhBbTqqfYQAHfhxUFpDCQjPQ+nfKc8
3+r9sM/az0CDozYcaQ4lh+vnn7dq1+J1zpYLUw2RTAbdJOrRfAWM6SgwmUUz8X4dqZ5mhXNLRbe4
44jV7W4kj8K0Q1cHiF82Yo28GOz8qHsPH7SwtY21Mqa1H6FgVT/Tbkh03aqLQ6yEHyfs9pd+qAHj
DRGOBV3twHA8x4gRshek8WGNQAiZ3LyZ5lb5omLlSKmevsPYWlvReOPkMf2yD4LHSqctf7WLYhJX
Jb8nfzKOiFlUNECIIzG8fl1PWqdNLJrctseqHsLu13Tzn4aRp837uBUw0Aoxut5os05aTTKaCK2H
5OInlOuEK0WK3z+IpzgRWtKLN8Hd4Wr4RITZiMY+62GkeIktH958n/jHWALuOx8OfuBDxuGFxNd3
wd+BpJe9BG6Ls5A5cVfs28GvQu5ubT/1/in2MF+imoS3PXT70CtfJenTU6q+pLIv9O4GbCXQOSdK
K+JK2CH7dTY0UYKn3oLKOmp4XQsctsxE1Umr8cmyDFW0kuaGM0Ke2G1oqfizM1u60Tn5f26HOwTD
eNUDMRxfTgEuBU0akDLPLhGz3aHp7X+fSInVS6VaIHia/16ZbaoU9/jGdGiS/JRes3HSM3GIC7mn
0gsMDgibOZEtqMyAKSs7NYaPz0+oOIvpBCLOxcIR43FPDZ8pkO4gG8GknBuK+nGnhmrzxYq/riXc
uv4NCWBre/vW9h3Zr9+rXnDzCTlweUcJeDBNSdzC74YELooHQqyJ3iwJt+T5B++MF9CgfK6GrN+D
eiCLdlAvZkUVglUZDO1fGk9BZqs4Yv981GdLkOf2NsBTTzijA82+Y9VDO8pjPJLNV47IeE/3apQp
ZqGvKfeBNgEICiy0V85gyGykkHpQnXcRsXoagjDazNCeLRLrYXM4IodF/6bfCFrSH/4ROCRCrj+H
E2xOsbvrDt6UQKuiTDihhqfsVRRCjVpK8F9f7EUvkzs7VZK4tffXMdX2fRHnprLW4bw59ZJzT6Kx
m93Q9tDw2cIyJo3OwdbQNi0Xg+xbT0ajHmTN6M+jLTYQhK+6RXxlc0Jr5QvZCtjPDz1EhFMTW35m
fplqfHqkq3otSf0sVYB9znETpSYz9/WdkjTMQq2rgqwbyai9KDUYWki2DLWF0EaC6JtJs4XHxf4R
IvfMcOkvhMT0yrMZVSe+PjiUbGThJI3wZFdlVOEEjlxp92a3VTlmYbjNu849t2jqExFIUE1x1qDd
IoOCj9P6JITEbPnZ8rcnqrecy2qrmstFXms9LtZQHitarQPkRP7N3uxQ67narZRFbjTFrIo81gwp
r5suSpLq/1lXrLi/3KRvV3t+424nvkpxVm38OxCgSfFjznx0e4u0neuUwKddUIB95/3AWiDQqkYF
8E2/DSvpQOClxQQ=
`pragma protect end_protected
