`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect begin_commonblock
`pragma protect control error_handling="delegated"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa", key_block
i+3dgAUks2H1hU1158fXl4oiKzbtv6tz4rthDoeCcMonjb8uSn+iW2G/LEIJrldhmorAsBEGA/GA
gaHOjSNpCfvJAA1X6KfsI2MpBG0q31EKgzTgfWBHsb7fIrIJg4rxlFNvBfzeTTWzYO0EfRSD5LD9
YOytyPp/kotaAVNE3MXibwG030DcIFA2o0cMul4ZLq4QDdDCKn+Y24XYtAepQ+qI+c+C8Tyc8sRm
MyMQR1+4kFWVqOvI+2+v3PU4Py+wpBL6pseqv5Iqo6jlGBtEzC/CuZVmqHKeJkBbgP3xHsBKOiv4
TR45g76Zfa0cnySsRkj7vjjN5dNUirGB8p3Piw==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect end_toolblock="PQaX4YQU4IutH6lSFlpUbq3q9N7830smuaxsrv3CyYY="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 5824)
`pragma protect data_block
XwrUN/Mgx5w7sL6gObL1gZXmU3MIiVD2KLFBVcLyi8WIbZp2akNT+sJLB4zXmrU/8o3WrTh46Iio
B+MQxsaJwcfW2McVhKAfNbylTjzn2TAorvR8oh9v6N1h/gb7f8kmVTLD6l3IB+GXxLXG06LbWd4X
4JzJSbXXmgKSHmptymgkXDVnDBb1LqkrXd2VP/jzSXMga2itoKoDhpb6l9h8qGhLeqe7TKZ2Ogfa
EEvdD6j31f0fKmt/uV56hRWey6wQboCXjv8Z867AC4N/r5EQe2Z9j9nBKOawPxxvww/aJCZxmKR0
qg9oYQF4aa5X758PfSbAZ/w8SHxVvn10dubSaymMNbhbdD5MpiygVluxAdzuybpFlmqQHKo5WtTU
RghTpO8v0grqxhPIUqtW8DQ+0dmspEmsvhyoPA1AEiv6YEm3MIdTNmX56WwF1AgVJMYYqRCWZ7xq
mv/5jmvqMxuFMEsqL4hMgutvh0UyFceOwOLT6WC3mTPwnTNXjOGLp6GYwF78QKNsjab3r65fhyEX
POmO/YSWXk6qDFwcIgYLnVCjV9T5IJpnIXMQy0FkV7DHCbvG1453qm/GFCHh0ie38oyu8xORMAaa
UpMEkESi93h6tIz/DctJAbjvbFlzIigQxirNsG4gDQGVb2FGAtMVBCRArfIkzrGZPqEDPXNQOUpT
+Y657BzHlURGmgEI2z1TNMxYLodHV5jCitD58Cume84u2tRD6LqzAd5W816l/dGSlXj75X8yuyhY
9WSdixUb5lAoqm/iiCCGVi4e/4CtQqyWXRyOOgjU3B02JfLohno0z9SdnMjxa1DqZWTeivQNNAMG
7FRIco/9gFpmQg3THn29JIXPoabQAszMgIvORX10Vdla0c+dYugxq925Vu6zd0n7KLyluPIX3trp
+n6rm5HWpUATI4dnx+/EPKpK9p+6kvlSMoL6Oj9mqZL4prMQAsA9fbPXRCTF4M3fXOgFbXTgA0Uc
oWvBlHUaZoe3KDH4zwUyjxvRiRGvjvqHYBBhpwIe5+YprtcK6vP1Gbk67gkuLAgDRlgrPTTly7Vz
djTM5wmg4++urIl3HuTdL6nxS/QqJYUGJOwk4qKNmCGlhvAkQ3+GDDymRudj7mxJU5W3tRSpm05c
0Q8e5v8MKC/26aJ4Ru5UM8hxLez5V+PebUV4zAmylJ5yJhA0it1tUs6sxYwqY9RXPkL0sFiib8wn
WnQbY2oJsmdwUM8TVS4HJpwIbwuDb6SjNB7HlhgANqX0l6BWbe+PkT2Am0r8gVlNWwIj+kpzPnXO
EC/PnFG1hTVn4alCwvqSpkoVTX//DEkWtAT1jlQ/qmHq9dInA0ld2J5PYVWO66ye9DSdfkoZcWSC
BitDY0DyHPQdMLQWhGL4UvDmE6OXBztnKmhtXEd2cYudCUKhPCqSiWs6ZlP8MhtcIMlsZ/1NKG8q
GbUkVzICh54Gwcrw3nGQ4jc/pB8VsVCMgtFuZhYvuiHnIswPO6j/eneo554h4eAEKClr8GBsKb57
XL7o/KmW1MhELXuBn7EKZLhFIK2U1yjifKxLV25taklO8YoNAIwk7Kl6MqJ/wh8Jb2QZuLxFqGMM
McksT/jqv8Y90C5gK9FA8vcoBM1Ss5rC/L6N33BqMYmbAajjHt3E7ZMtBWoU2yC7QIUbCeseWhd+
gKCXu+jmGD4QNaM1F8I3TfDRIMGnxUSc1oCt1Jw5FKxt6WR96UGuPSKINVxnoywSZY31pYpuYwV9
3KuEg/AsLbELD1lNYVHXGT56w+vPYM42LD7KK3hIx4R3T/FcjwOaD+vHNlUv/N64ydRVcPeivA2j
+Wiv1QVm/Gp/dxCLg6fCHZ0w88z7OytCvMzPL7/wsDumuIral+N9ov1JfwhK2IDf2GQ12zcuLA8m
z7BvFlxgz7mj+nxFVGG0qhpGOYEAMHQrz0Tmj88E13gFKxGZ5ZUwD5QZOBh/ZzKEa3Zg0mzteUwd
SYq/2h90V0IfCdOI2cU8Gdn6M0Mg9Lgkk87dUmtTdDJlpVhfliws3mooXPfr0zh8vELrU466qrye
a/ki1eknnCnfu5uLDlPhWi2SiJ4rSImwgTw3+3zwl14wv9BZuLcSddeZqrGTVPOuu1Y3R3b9TvMI
1OEeWp+UvQDVr98M928Shx+qqCy1wEllhIC4lbjSa6KFOq1nXisYioDNSvCYjR/eWforuKRU5IEt
o6kUTK9DCL0G0LfL2CvZwfQy17pEe/pGepmn7PiHrnCxd6rPgvcelbDkIsg0lnlpRatDg0vEqTSW
Qba5QzHDcTVVSVVfHwt3ZFShSxHwpBXy4Cm9SGsLbNGgXf5BBIX8zR+dJ+DGSpn3IwI0GX24Bzj5
DwnIxHF6ygwbwnA1ZPGzNuv7jZDHE4paDhm15UAb0qnseIAYCqv1mPQvCbJ2Rb5rbhzRUeELauwl
VqEyx8CulexjWarz5lZ1dcN3XgOg8A3q+0sj0vFxecOobDsq9o46mnaXb3hNfjPbobaATu36ioH5
AwprUk1Sgj6a/gVi0uWXQ0POI+otkSFwYr0FDjhoHe8KvdKsrF/hShbMKplVpBV4uYTa95PY4SBr
rOzzhyBJosvE6LK+Sh81/bo7eV+XzkfuEGOBgl0tPrnuZmAmqQeH4qwlIQOy60a/1RxVosgYY4fv
vZ2zZ8uOdB7SvrPlm0eCnKIofPZheehtfePs7C2nDDTk7zzuY8x3iCa1H8/pXoASt8lZ+SQx+pN1
j+H1Mn/uu6ViXjgQRF3YTBtdHT+yPI58vQ55KJIFeEr+oAnwqOm1MxU4iF897sfA4vPO/HtbjFLG
17GTlO2X3sKz1jqajTx1zLmt8LGJoem21H977ttmFJdVywxsB8uetSm9AwnFyIO5jEPNSdat42G8
cbUjlOv7PFllgV/BC0iDl5Ijf4/KAT2/LUqQRIBno30+B+vBO2PRu+R1nAd9EYPOfedz4NIqMKzI
NnybFJ6m2AffVn9+AIkeBct9Qulnm+cCDnWTiGqCD4kPMW7ouhgLD2qyY9IdOP55n/hWFfitmCyT
8WjADVPGaL+X95o5ZMiv/p+M5t0dM1IYAUfNdGyX985nd336puKL0kcnVWokeMQUEr9V3eweYzxe
xgwicsm8CbM+tsFyGVk/59kMZOY3cHuh+gpve8AzpW4sXI9jby01ANPVpPUHtmLE4tGWEm5zoOnM
ZDGsYTECdKocYxhzygHa7BDnmsN7i39tELpN2M5ARbA6cBSW+gXtiLOEp3ViOVGkA3goLVnq6kpO
pAmdlYPCya1cceC9UGMMw9gynnnGrP5L33tvIYNehIth9sSYgoVhlHI43ExUcJysyN5zlDS7cWAy
iY9EoXKcoOSs9ot51of7svSDu5NAx5nwRvkwG6Eg/z2NykLPBVeG5emDuoOYxxFLZ/JL0Dnv2KsA
R7lWfubpxdFCGP4t7Z2cwgzjb9Fb6CEgMVld3BmNVCnT7tFHDhVPJI6sENom0NPEDj0vt4NM/BDw
+t2Ifds4KODqWAr3urqfaP+uznkrZxs4cLW49i4oE13y5yn8b9B8FwF1W6+dYQpTYLgMlJEGxLhj
wTa3jQvN474/SzfTy6S1brfGZhH9dgWVoQacKI5O9WnkmIn3LOgb3xUJ7QThY9BVgBJTmj62SWS6
1GdWWUFwqn5r5fkGnrupEH4jXcrk1hhpUm0yvmQbzj7C/JvOEN+G0ysvB6hLKdsBfpxPx8XDtQKx
YjoqzWJIKgA2QS47i+9t4jNG0cfbypY7DGbtaQ/8o7zDYCgiG6WIDcbsptMs0ReqzseojouEbTtY
t0DIRj4t63/G8+jR05XdIDK2voXiMd4wdCH7+yI5GcSKy6z2O3yEDRRlBNg5lCNG4YVrv7GM4tyK
3qplebmIlhcRc2XSvc/FYkD6ZLOitcXorcExLsJALKYPM9E0xtCZ60FZbQe+dOn9jeQ4NXFop3Z6
B4PHNc7e21d2wBQcG06Ys6p59mbcPPQl4sjhs6L2X8hJeEzmh08OjS9RDx3mCgeIg7hoPOQPhYDC
JWc3sbvQL05zPV3RIDrOZFKXP8nA/VdcS3VfISM9kR0TCxRpPR42gZChUjXVWslLlkoik/21oN8g
HK6k6wLb/3fq6x6B4Wfmjxhqdc+XCSVYnakGi4F+F+vd+quV2IpJtDjfpq18M4JoMdOvr8+VzEr0
VRbGAg0bcKpEP6kvIFPQ5jr8Ts3NCAH90Hwefo66hN4bjRCfzsRCbJzmWyGMqt+hfsyNbvG7g0H9
F/wHEnbhN4CAz4Sv1W2aC5Pv7gG2PUxEDTTS3i/uIlBS87v0vvcSbgSn8JIHMZSARCEO000oUKpL
i1CxTIrPeOe6lbj0Mk8hkCl4Pjgqt+3/7Pb/sGDm6U4QaZ7h92SCBiOk6uhqI8qTBtyCaDiY38CQ
BD8PTBee0xwWIi1zE/gjvKBSXSG4r+YPja8BgRB25twNm1I+9HC4hzVXeo2JDGlXCNtGhtPzRa/y
z3XPcsqwnmkk17J66/Neq6yLTpnj0/vzTj41UYFluGw9Rk4vgrXe+T/j7hQSGxtGYzgC0QU3XmwL
lsKUSMXW5LyC5u+SdzdS9Xm0kpbmwA3uv8/cUebpwmVa3uEWAoMR2mC/HmEm/YM8mD+GlGZESsdk
Mz1chs/d2NwhLp1vEpMIKjJhv/uLFf9LB2dQ2i/1u0R8b7k3D/s+DLPp7qcWyH6dnHLV1UXBQAxD
TRGMWeYlJ8cBeVWRpaodL0b8YvHgyU2Ir+Xm6jbsYjOhFLqaFDvWkWCpkw1X0fO07c6xPEXeBKQs
KZ7d0ruEMYr5JeYUunMFkswZw35FhM4Y0M5ZhvEGLmiA9dw0YGWAlM65yLA9SKzBagYEUxHoMVyT
8XKPN6I++KkfwbAMye79cJR+LbPN+Jkl8//gGC5paIq3q4zsLAU1fNl7SaQxr4/vzIbdjuTjXX53
ytLKNfWA52TqlMzeQ2y37Zd78LRSdUuBOD/tZPhpI4EomJZizte/8RSqAw847Fft1DTqQG2l3w+s
F65A/XkmrzF6PugD5SVo5MmKUP9xs4Lz8R+qFBuEhYWgNFnO3w2teO0NsvMz3Xxm2AdBGbZIKYPS
1SAHP2Pxj1ONGi1q+c+E2nlJku1ZFUH6ljqErXxyMpdboNr369rLKCwr0VaK7HGsslVIpkrfpslg
vJjbL0zflEQNfDiv7TPTvVAQtCCyxN7O2IIRsiegHmelbeKd6YwTA6suptVrT5FSzT5LFNXUNOJ8
WY54q3jeD6EgIGXYJd0R6GKhoiTmQva5FbheGyb9V6056EMe2zI3wUZcY772SR0K43yjWjmDHllH
8HE7VRGmSFez117PtlSfCBdkTFsXdUWSzd0AOHSqWruos8UfZ9alVz7kj7aOIxwaVL1kBnxZ9AoT
j+NOV9o5nmFYceTToy3BhgjjPWV2qZjn+dklRVOvqoTeempblYkduYvV3bZ39fSMDE+glQvx6Imn
zhhbp4zVqJp1Huflr8y+ll2MUXNnX4LPe2coE/ARDEavNOVRtrtSh6Iu8Rvl2yIkW0GI2OTdhnld
xKgkvmzFhVL+jSuyWTIa7FHat50uikiyUUW9DClOfgQGTQ5Yf0J+8ucOOdGBP97S3LPuB61ubJtA
SPTPSLJ9Rk4Bvodxr0429iT/+Xk441mZYaBbDluke3vrIjyArPUD1aDVMymq3Q214mq3D8BaK9u1
hk7PKgMsyq4TyjAVxgCMXlB+1bbPLNWKIKn0j8avHAOGgSf2mvcscZBE40ZKTUTwM0HUjw6agMNG
QnjZIMEQnLEuqvNKZePj9mQknSfcy1RxD//Z+WekVZy9g6XBevGixCVgGNP7WV3JEtIMNGxl59mX
UmglDReAgiE0ob7finvC/6BXRzTRa92HeLPDpId1MLcT3Rh5H3CBq4F6yXsL6HaaoYOHk9cRVKyO
YT4PFx8Zx/bPdYWzJNY1Ij7U5obQXrOuAb9lMx35Tfm6hXuwTtxSAwuUR7pUffiOT7/pL4jUQEPJ
S+ARWUj6iEoCGPYDtUVu9d7oDoZpop6Qba0boj2QLDMKe1DfC0MMdQNfU9mw84/ZjaQP/rtlCRAw
dmy95qBcw4pNR20MVT2YTQvjPnCIs/GkxDrMKWd+JA1ogkzxXrg9PXg69tFz5uf39lLxq4UMzYO7
QJe8glFKLGxCFSNGThz1t9Zp0ZStq9d2L9Mm04g/tROH6DgXCDNbmRUPs+j3uk50UcH9zmciYYoK
KBJ+gQCB/1XkFKCCSVn3qBydo6FVT8+4nBTEmCj53dUt0kLqjgDXZsLEJBmAuX7IZ6gOXFVZ01Uo
lfsNnwuLyN6VAWh6hH+mVwQa6D3Bwg6wJH1IZpk+kisfruN8GzJNFqa7SOhi3u7H655YisWgui2k
Slg50khwN1M7WrJ+Wcjq/zpLQd3ytKqbdexIVPsFjh1Q9xD0y/Tu1jRMIxK2qZ2An3arIRwqgzt4
/sAgjh9EL5P2l0QUVp1lu3C184w0KDMDOq8gjF73i2ryZZtegOVr2s8s0gCxITlnKO9D/SSb0eCa
LZMS4+oTqWfmTiq9m1GJsHEgFpn3qAZz+sYfKRVmYaHHlKUOtXpLUnQ6ILoqdbUo7vmD1tiJWovH
zwFEP/O/7obPc7/aUYw6h07e+vP5jmmqjqiU21gFEwqr62AXUFVqZK0I4mzMxJVQuMX8qkSKnGaN
6t944W4cOLai3yJYVKiYAMRTlN6hbW4OIvaYw9zDoH5gw53EgrfZQnK6Tex+4BoUNU3gj/vmPtm0
g/89sDcg6io4ijgDh8RX1o29V4n74yyg4OO7JATJYd+vZsWUFHg5VN/ukZstihtQdqlddF7f0/3Q
caXZ95VjxlbEXVI2LaRs9wRrq0TOrQIn290DsemYgR8sqWB9yxddyQgHLjMyZRo+7liKDxQNJCX1
eRy3uJfamaZ8r1kVu79n1PQY0ZV4Km3DAZHh1jafb8FGc13OLrj2pIuSv9313TqH4rbOz2b9dvyb
5vpJBfi5096MsOFT7c+o8vzCiBJ/qWyR5S8eQESeY6dl+nAZUQtAxTBtaQ4SCmjQf9F/cOTKsPTH
N+iVD6tQILH7xFLFoJiwtdCrhhamohEFjShKZNvPdMNCyStxBd4RfNjSfwtMZurcoOirniA8zR1C
PG7aRGmqRbqBP8PeOfiPE6scpQmxJReJk1dwmd7XlKYI9AC1yB+i6nkxOtRF1VcLzl3FFz4qf4He
SMWxQH55IeGwtBkstJgoWDfsK96MDgwrhgPFGmdm4vsy9hTQWjTfq6pr59YsbWrhO/YaRhpHmrPC
aCczoGZXHZeem2xQKq1wNGLdobnlLmM6fVtMn682P6pZb8SsaMdEZOsiaBZ6I077+IPrFsvjCguL
sEzJTy/J1nK4PXsHthZ9pjSsi8E9fbC/Y8Mn+o3Ov/AJ14DNn3tzXCN6FEhBcNNuUB30qoUqzzSP
KDwQBEeCjzdWH/pFwaX5NQp6Vaz1pWfSIxYa5jARUimKLiUJILB2Dp+nxujQOESwbm6lM3W3zBdj
+Mf6j8xKsf6r5YH2asV1/+cIZICTXhZPjZfg/KQf8ek3zyUylUgZbeDe3wpybAL0jyUbwIDuKHly
hMhWLzSsShPdX+0aNRpA3PSdipsxIEeGx767+BkKpLBldeq4XNZCpKdM+V/Bbvrgf3dz9pIDopre
HLR1Lq6PX2LU+sws01A4Jrwopb1StbkTWzCLGICQhfL1LXtptlHCOuZByVoigVL0pu20j/hD0RRG
wPsekGprnLXpPQ==
`pragma protect end_protected
