// Amazon FPGA Hardware Development Kit
//
// Copyright 2016 Amazon.com, Inc. or its affiliates. All Rights Reserved.
//
// Licensed under the Amazon Software License (the "License"). You may not use
// this file except in compliance with the License. A copy of the License is
// located at
//
//    http://aws.amazon.com/asl/
//
// or in the "license" file accompanying this file. This file is distributed on
// an "AS IS" BASIS, WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, express or
// implied. See the License for the specific language governing permissions and
// limitations under the License.

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
W+XbysqGumNHsFaMf76Au8ipaY/L4WBO512D2/lZLRWBlyvP8HAKLwhI8Dc2EfEv3a3dlkxLrgMu
JzqDNziSFZ+w/tu1gngL6iADS8EmclEkeq1XWnhLVQ0ukFxtw6yN7R5sqbsY1Re6N4os2n17faWO
ozX5GOmNaBuAUX+hDyV51YYQQg5vxTpHhpvOWVzbQQEuPVFirymdvb1lj04IymiOQ1lYP23J4kCG
5eDUGP8FvSDvQftO1HRj7WHeLmfaZ7/0khFPgXidHj+5J2fwYglZNXMwbYXH28B8JA4k6O9rWZs3
RcHOEfQ+J4SSH7vSo5KmEAOvTvOcVROkmGry7w==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
3hxj12Hh5/A5i1Z2Vg4oGoif4hGU/feuFX2flxD7eVtA1DcK8PN2Shh+Leo+qRNph7XbK+ehxcG8
I5YpobqGcBBV6VwdlrHLjRYdf67IwXIuZHTWmF18TTllj4pD1BDoNPusCKFvWQaqdvnN5EI4QT+7
1k2z/bEc4JQk5dmS3yU=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
frkGFRSC9T0+37Y8m8Rr8enz6q0Gi+Ws2YHaO3IXy9ahsZvPH+dkheqU2nah3LYsHtmsO3CcUBkd
CzSxLgmNhsuAvt1/bU9vVvgC3bvTIYSYQ3AeGxv+tREoQtdtcck6cH13Ap5QKGZPPQ3qNH0Fmm5X
jgqFo33FGjZTtgocgvw=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3056)
`pragma protect data_block
xfKsdUQXS768aflth20JOW51LQCeSef/w5iezXIAOznFgs7nsrIOd0+UbdrYC0hv8iZy75bcGUTN
8BLW6azkxvjayhjeTjOM3j3oB7yu48g9M45izkvDwQfK5DGJ+WvF/+5Dr8uhFo/Bw9r0lbuQwUAA
N5CX3hcivJlwoRw2UHHoVdcv6XuunsnkLvVYh23qgHjTWHfZdCTKS776CTyAxLfUGNND3Y3erTit
LdnE2XuXmMJ+Mtee493/L8JnpmrRbKgNdNR1FVTCZOhgKqAAiIy9iBYLPftqsxRXIQ3yp7E9jse8
2qeudKmw2aNLk+fAfjQw03a4oj80l0rP05i0+xfBVITGAlFH3hbsMEoWRSql9e4cQyAZ/IRMShGR
HssiHz05nJS0pYMk2PHVOtNGqdq/MJYfCDMHQpMqCT6BJo2IY5JcS04p6IcBeij5s6K+7IklQqbG
0nAf6mSCOyvVtciTAlRD9+al8tyqdZkhgxvgn/NS//mUJDGTppnAGf0cLFyHEzdnPbXUKWV/oy3m
GZ847xhYq6kSM4q6Ulbu82D9hDpidKhHnkSveSaEHBgJbLJQ9BJwPoAvwDg5LmKxhvUSOxPWwUXT
5J18oOZxU8bXgdSvOlPhmmPQyJwQtSjs0IORgdCxuGE9V1bHnXHjxQ+b9t1fSkb1gDj/uTzSwrRE
qD+OAbGBH2B0JQwgxizstdUbQj73+SFtElgjl5vAQOr/YRUDzVrGA6yRMWifNBvMHiNIkvRUotVs
8sdgVd3b2fKXtYQ4T8Ud+8i8Uu5/z3jJ82IsNA3mIxoNPDhz7rVXRO0xF0RCa0kgBSMeTNtATg58
BjlasTPPqc3vhDj2l6kQfmWgEyBa6mzJ+9lIz+L7FTQNL+B/ceepiBCxoZjIDnk5l8wGrOY21kQO
P3+a1M1w9fM7HPegS9/cIETxNS0xzSeBW5QROlE+sxDUpxwW7tW4UxqyfH6okpr4ayhgd2LKrMXu
6DR/10WHuFDij1NJeDETahWq5G397IZemZrOvhenYxh2aJoearV13h1dgcf2THtRAki+tXNBRO05
Ldi5xzwy40j556UtINM6ABM+rPJ0loEtoEllkQ/mHKPbfhRGud2Yccqt7b+GKH4NJEM2FwGO+/BR
G3GQTb1YYbX9rHiVt4X4UNbK8FoW6fUu/nWgYhDsLxOPUJ2sFxe5S/8NbhdtArn8h8IM4wC/8R9N
XyFzp27QlBA3Lal4SIbi2LPDalcGeU/wYyCznHBTbAgB0AXWnysYaVAANBL3BsdOWFRlztsK8TZc
yEYY+DSHLIHEbxsvFLMya8H7s135XOj3nKs5+dZT18lh8tgLt1D2KlPCZq+MvBZQWW2GTv8WZuET
U8iXY0mr9vi/U1WdIcGck11iXnMhHY2jdQsJ7eJn1/DA18actH7gf/kHyIdYtjr59grYwMuRNrXF
/QrY1EbBVo1RhqQjqTCv7MicKRFGN4inNIxC0erBeqfjnmqBuNw2T8QNC8HJObQkohjnXVCQd3qc
X3lcmV4itESvi4vmWKhuiozXn3VUgbO8wAwe/kilfXgUhCXMDcGv8pgqqH9sVxx1AkuJZA+wuXkq
PgAjxfBVo146qn5utdaXzGLY7rkF8TPmCEzoBuZa9tdzVaCLQPkkhCKDsRZ/82FudJW1oZI4wj78
aVuG7wM+6vFNelQ/TFQQO+s4uf0zcuahYzB2LPijKDT1horpsR+fiRF4PM5QRsEERvozfcTNQKZp
AC97AqPcDJo4TawLKZ3IOKJ6GZR480umstf0Io4ibXKPj2DRSnRopQZZdzrLzBA+Sy+Wlu3Ay9/J
7Cgc0haahwssQhkcVMJMrdoKZUoKahDvj4yDab9Q5EYfA5r/m6oWMKs/pqQvZM5d3o1vMqphO9MB
rTwY9PKqAmnFTRUImxBzS/Z19NT3ETc0/sMwQnftJEMIXYCQ20lxb56AKE9+y0CEYyGXqITr9DVn
KgBxRCmCh6nhpXWZaNImoYuq2OPWc5NbUX13z4nQjU4hifAO5G7DOADbEU06epeUHT0sbawNyKFh
PSeydpmsMgAJmSePP57bbKBuUaKtb5723/74ua0IeQbwQqAPcmvqrZ4HG4uNX4c5/F+e++YZ3Xxn
BX/44crcxS38jCHM6L4D++btAuJtdPrTOZdRTH/L+uHWJFa1TKVsKn+htosG41WmiSnpKWuNqzFk
D2JhmEIL9TuEd29f4H6olst5H0s2jk16V5KgJ5Xuu/BYosyHb/K/HHSg7F7fU5SSej5CB4u3DJa9
oZvpAj0IQnQgxEdjcgM+yNI6FnFgjam6XRcwqMtKtfkvlloVvZQGvBOZqOFXXIkGv5AghS15R9UB
QtaI04ZL8RG4FIDJN9BjrjiAAgd5iWcIwrKUmtzkGMl5O6HF5TCb0YeURrWmXAK5pFXyEMgqnxwN
A1uI7uRqD4/TymnF/kSc1hVlULTYUnPbjdPdHxIBeeuVFROIqqVrnKjnzcAMjbS9GZXcgD8igjwE
JQ5h/jjgLol1wUwW15fUXanlu0VNW07P0r7TZ6uzv13SMxWo3ll6mdgOgiavG0XI7gsmVnRqQAed
Zm3x/RBW4smfFUiTahb/uiUSGMxSfIBBanImLZpgTDGkzuwZ9SttuyYLEeXPhwe8x/B8TFjStnDU
EeKCbiDGu8MW/zbL5M58vrSrHpFwAFJyF4zaDNtipbG7IGlszBU5bPLWZxPMAk7qPpu3N3HY3d/1
Jz/U9Xhg+6vq8VXu6SddrA3D7XpnnWCcUBb4XoJOEW4ClyiWtW5Gv3dv/5mVGp4fwGuP7fvRzHN9
FCi83VLza4fOdNDgI4jBsBXs8TTtSPwh8+3emKcDQk8YC3XLgS6ke3peUvsb9t+LWZt1uBkj2D2E
h7Hx8L+Os6Rvk1RDRY4TtjP5uiksWk1ICHpSzNG+ZgMIkO3RMx6wtjZleOf801cXjMHPVMkZq2cM
erPYTyMWc0Q4Os/69ReW7QxgUA+aXpjSnItEA027qpJ6EjAlLyyU+ard22nHj3TYv0EkZNcKZCIc
rCCh+QCtQPJSIazxjSX2pJ+aoxFfYCep+rqp336KbE3Xv7ZJkpASzZmIv9u8iJdSlZlxji48LT3Z
sE1H/iApmU+q9ZkPR7seBHWfVyCQqPMADnJDmuTN9GK1zcdWISvBb68P3NRM4XaAa8JZmCnc7ltz
r4U9oZBfVRU9JVji3oUN3eCWNSIQCOJ62s+fKG8ofstGgY83eusrozG2TEeMrQVVcBKvlVEhBGGZ
ibczLGMhnCBFYq5CQ7+Uo4wDlf+dHd9yiXGjo3azJ+BmYQDISgBhnjS6LYJE8pyaiL7GYboONpAf
S2XBwaML8IZ7FRYwCjQICS/ILfSCFhQyeIqI5UeuW24y0K7mEZ6avWiRGvMN0G/rQJ4VZFcZV6Ut
AdWJgVWoRYjEOXRbF7d/NnaC331dfSDROvk+/zXxGL1wWaBYPf39Lku2kDoitHnDfFDkL8ovv+Ry
6SYTalTLr0CgFsRFoCsnYooivKOZI3AsH33MOTR4pAM5vdPxmcr3SMaVqxJYlo+uaOEpgeT9wKd2
wM5K9PD3xUMSb0m7EiSwMKKUjTXaA+GI81iKcGTt398N17Z5ozYXFkPo9aRP++SMY2S4SAbhrtVb
3ZgVrN0pmbcpIXuJgf1Blxq3+gNR0bwAaDPusKFMCilz87ZuqN6IdyITNEFW0HiItF98scl3JD/x
hIar72hNAJA/iznpXvhbSPoqjM8vOwK3aLxEk4i67j9HTSjcvtTW47J2odvH+4/onmvyLXc19WO3
Xsmn20ODVycgNsLKXvFCaw2q85nphgmnKLYl/A/fhoz8i0qQFyR8R5S49FryULysYDSWjoHf3VYP
hvAJj1KZuCJKKmgwEmkm5lsabxSo6xPQ/LYo5Z+MQ9CkM2IhJDjzh5LiNFkxJESnYm8Q/C+JmqIX
bCTt/+TxDM9AC3wnWxOP1hT9YMUNtzzkRMeI+ViXajwaQVgGpSIxMtC9GSUrkASiIyGBECwpDWBi
b+Sd5w1Fhlom4zlkNszNK/DDJzdtyImMA3T0Qqq7CMlhZeQ=
`pragma protect end_protected
