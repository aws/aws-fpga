`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
VinOjXosxguCsieiJThfB0sdwrT1r57IKyBJoAARC+Y+uxlV8Pgzx+ofB8wDmF/1n1xBkx/z7XVC
z7JGY5USQ/VxfUH8jHa7dN1/C/Kw/eiCiZccpE4C76baH2vHgKNhJQ7EP4haMceWDfRQShCIFz8b
87xmu+7QPyLKhUdUc5OPD3MMOqz9V2CTi/Bk4mxQJX9FmjQ3s/eCAcuT/Fp9TDS9TDmVELuOvH97
RNzL2MFuN8IEwY9vWGVOUCq5XoF6C+ofnMW12Vs8JHrRmzTEM1Kh3eDvjGItSnrtwZW8q6lYL6z5
pIgv9U/ws1KaxkNNH2f92gOLT3Dq5kTFPoz1Ag==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
OUXxFpdp0TsQzcYLYuIG1uDRsmDo2gMg0hgScrMajevo1s1Q4LMpnL+TLwEhf9YAIF/VgwmnWFtd
3yri8BglFiChUMy5JPlBOAx5ZoSSkdD/SwATjzmd80k1BZOoWOhErDVhpjnyGncxSLkkcTxq7X/+
ey8KYe56ukAnqQYIJ8Y=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
KOx51JA7nL5TCbCuXVwtODgu3urrIz+KuIqWgvK8sTp+k9a+twhxydRkvGT7gjQtXBkIUqaYXtI2
+571Ywy+0ibdSZSTm4l/qxgj9v4mFECfnsmWmXIXs6YwLW1jy+4pOHn6rcqM/1onIs2AwPeWFyaC
pwJi/Ss2FkjVeHvt3yw=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4208)
`pragma protect data_block
CvmrZC0BhJRXMF0IgxlypXTvCr2ZrGFVC64PiF+JEaVg0AsWHAfpe8Fc1FH58qZP+6K4WQT/TH9P
aIMwvCCwT2RYN2Wc+fSntcwIIQocvFJ9wEWRTJ6rlL6yZEb0KGH/Gd6s5e8mGRlIg7/YySQCAA8p
0jjoh+nRutYz4B6Djjcxx4fpV1HpR+2JobWpOXJ4z0pUbvx6yu9zgAsmTcBvHSqRhYuk/CBY1IT3
9aKkYghvWJGNR9AqMlBRpawROxjpc7iyLVpaaVCwImmaSfu6E7LH05pOb+CbxjiXcDbXJ2uiXL5V
jwCTGbPqL8oGb3Yk3O9hO0PtjtK1kEyWzVoNfYht1S+EBwZS3zfjCR6ropmuaffteE3jPHyDmWEk
Mruppim2e3nyTlyr7ypoTW6C3m+974zKOT9eLY0nF2O0p6YuIUduy9g9gtbgxRDNGdVhDQWxvnAr
U+dShdUNSx5vmFBb5soHU3KIdcH/pae7378rGfa6VqT4dHvUvaU3lrfJD0URxWOdhL1vJs35N1Rq
Uwx1+YU6vCm+9q70IYvx8QksW+vVuInRdTTzUf79h8QaSIdRmxVlTdAe5qX7ApUUCC/Giy5cRqbD
YjKhz65pIl20qVfN44kILYLxLpFcmIbfMgHGv5fxxbIw69xl/LqRNbuy98ytd+HrqRYQ6ET6v1jU
OVKqI3r8oMJFtE0UYw7E5VKRE6wrwPbGWzxEdEvJTcwJYK21cQBsQgPYJW3QLEncctvQLBOSqAA/
IZ0C3kQs9Q8Hc+BeqXKWVRZ6vfJnpf5DV/b1yHN1jUOiqBQEGkMP0WargwykinOC2uRsvv18krpF
rEgi9awWW/dJP4utov9f2P8ddEzRT9XY9vIYnRAX9RPksWWEzRb4sGknPQYpDYR3qf01kpJwv3lF
izxr9JdQjTSDEwXPV6LOkkz1xqk7+jyODdAdiSnQLSroU60tzf154XUaRR6hp6uqztX70q2e3FX1
U6IywfBsJPpw875T1XTqYrCad+j9a4SBURjaofgx/nYggeEiQKlrISpHDAoN1SD0O0tLIxnxV0cw
WbX5+MsXwzhU15uwQ38Bl+vMWO8vKaWDT/r/Rs56fp7Xu6Mluzn94mDlIXftlpxvdYslpkOZWpMC
1emhrEQQutJ4VGKWYIX0EAH/CTAaZeInfXOGAR3iBp3t9+wz5aq/xSkw+iueubwtdjs5ErV3sGfZ
lXuC/O74iZfVMgcupvHpV2IDrZZ9EULPPQR96HPwOjTSZtBpZsVpVWAiThKGJPsgxC7vChb6tknH
7mNfYsGQocHCnUBMiVPIkITA7/Os/KxFLxKBsuFQ1o+lBCahFZJ97wAeaVs83l7/R8YZ3fMeFhaS
UHpM2UiczEC/+lMrRQXqkcAfCVQrILUOxjHCa79u6VZVN63KhYltaM93TZoNGfDbS3WAEB2D3DaT
xqvSs+AQgQVd3WwczWuSKATyJ61CZiAj8u/3IGY3k8bkBkXdMQ4ApgAtmBJfLJiKfpI/kdIJRXYC
VVuuhxLP6Tferw8hyA+CIwFaO1dYdWCmfYJ6wT7/aJ4TQ2yvwUq4dAlJy/Z9Bo3MnAEBatjXGA7s
MNV7tbFoIyXIslJI+Z/ynpH9JmbFMSTOL7n2ywJYb4VQCklPrrqBvcN/zuniNrrbmTI/jnOPC+k8
b1+IGJSutNp1s5YbQrriPz+BH3ZLLcZTMqpaTmOqhVnlzbK46LGbnDcLVxFRPHdjIZPUdUmfxWLq
iHUs+hYCqImLsnSPtwXtxeOGAKd5uarpnyLmOJpfg0REd8WEQvu41sz/0J6L+8QaLfK42jdZr47P
a2I27aoTlGiw+9zrbvfyJYsvfZclrXvgaxfdmimgBBwTnMIq/oMZBpUoSHmmEwC34OZ8ohgVdbkG
bSFk800ys7P0Dn0QoC9K5m+CZAgMHfF3snz+9cf3azrmdUon9FcJH18syvwXuTjaQaFPkyYYC+Il
SPE9PXW7lqudk/kJK8dXJAyDxJBViSjTiwKm3+m0Qtbz8Bnf4a4x5kmhUl2yI8CyH5AkeT6M46qO
aKxnzDr66syOT42pGqSc6l/Ur97znvKEaKz9LD7sHICl3od79Aogm4CaxHsHfe3BZN3V6YtiNb0l
DkQ1n0cZYFdn3cwJef4IL0Mu+MJ/ael1Oz+4uPqNmpApPBf+VRYe19+FW5qWfG2v758C/6V8f2UU
vPM+6x8Z1Pl912zTyYjQCjMSVac/8cDN9LUQIpoe/OA1RCasKa1M6nwFjoWF7qSIP+MlHWhAbxPb
YDSPXqEPprckMXmyloB7wG1RibJtqL22M/Tt0Cuo+UjUqowSZ6DlsaZuIJRuaRv35XHGsULHWG7V
vMESAmfY8xl1x1bAgMtPFBsONWQQXUS3an9gWzah3WpiOls3dPW0iaKT8VZIicDOQEAJDJ+MFDx4
O/Vr0Qro5B8iBcP35vCGq5eQ14s0TSFP8VHUHvx+CefO/abO2fNSb+8OQaIEsOnFoBX/wt4roNfQ
gJrSfXvVwmPOQxYpVNKya5gBpfBrKSlVJ1DU5qx//4UnQLSm2u74AbNwwPZBCsJi7KDZBaXt5tSo
QwBjCRp04IXHsKxmhFFdOJ/4d/tgFylP/tM6fjXIyyFd9fv8UgkYlssxkkoOLp0OYJKC50cY4LgV
KQc9h8sRzX9TM0xeNsIEdlXZUaxxoxHxKSgcCGn7X6xnnYKmgstBVK6vkYJfoNpewTEJo5tA+ZfZ
BII91tQBpx2/GjVWMiW5kJW2a9TbDBmRsqnOcC66lMPaIWh3Ez72pbaONK8FYa80r+vzr3AxR9Rj
+Y570NKOx5lB+tgCsmIWMYhUSHpezgpxJMMJ+6rO1HpRx5PT+WAVu4JT/EQqch8ciaWq54P3a6hF
utyEdCIHvYeJVBUVpX1Z7PhAvsVjblG5hSgFBEQ8cxDlO9MR1algN9dNUu8ZoS5cb4TVR5yWMGyi
DwzD+v2uxjUSC6vb8z/MoLY1WfEHK9L/pf5L6z+inEe1e/Kr9jr5BtG9surO3rx6lUnMNhEgOS7Q
0Wfu3u9z36kPa2om8PRY3AWOcJJOFpHb0HSZq3cZv/sxA+d9IhUzHeB+U5N96mEiPwC9Ur6p9/rR
Jy6eAlmFG5SZvBKKDjR36KKKKlpHijMgOPZ4bz3jqm1qt7NdyMAlj6GM83yu3FfyTI9QDOixQa8a
3zpQQq8JqqFjkqfqlIDl8YIBcRtpIi5+nEWSmOOhGXMfUMKHhRtfAp8s16560HzCBlCjPehnYoTc
YcRFVVlS9/jT/mWADn7MkxTv2bCVeR+nfKBgigQaWQv3f8OUfi0+RvVF+9K3bKH4WyYWI2F1ljXT
nL011VR0rqZcttsLgZQ0uhvHAExJUrbBIb/81I24OWMyaCAhwZHzb8PK1TAAejz6acbJnWzPxNDB
levoKUBeMNdhLJXLU+gqXMQF1O0IGSRBc9p+rIEM9OtEUWKsIANkMyu2d+X5FQVwMtAn6borzLil
ZCAr90Q5Lg3hP66vhjly5tCuiOD3zfUqm9aGoCCQtdy4B4XnRpO+rLIvw0ATS7p2530AR9rdoFhF
x/tsnW6u/0qB+Gyuk/7vivD9WnY2OxzkWhrwOiUbO2kT+3hxhXv/GIOZpYj1twkQAmKckdVpd6Fh
tl8cNIsJeY85osuevFy/nY8sjK1ZnRiAlb/zjHqusXuoOduG2QzvqdGuJ5tLfYJ3mbKkD6A05k2k
mRnsd3gtwQ/oyzhdT+6jZrPZy76JH52UEbyMc7J9HFI8kITuXzxt+8T/HIJaxjUSDdKxJLYL8mal
NP9bW6NCeCpx7cnF3swVmEovOqKGzfKL0Vvh7TVp6Me7ehKs49yGP+LdwmDHLpi0GxEf0hW86OJr
0piYIRSqIXKZpJHT6UC55vikLu5gyBREHSeQJxhXeoD0XD0uc/TzeqmQwqg6T4VIXkHQb5pgps91
wCckTLaKK/MEp4/2Y0sBMcThpnN5wRjo4LVxEQHofG4mm/ZJPLX/3WwF4OJ8A6oGqTBIZ0oflXfC
/xuskNqQJtXIafo++i0J+5+6ulgjQM1oL6QA1l/pUeyf0zyatrEqRi8Pzplgcl5BpgssbHsHFDEW
LZfLCxl63QnU5XaliTpUW2j10g7K248infXLgOK/Vv5zlq565NlVbmu5e0Pr8D3ETwVp9CPdRJah
5IQzxHQtoJ1iOfKk+VBvcrX3zln1RYbFI6Q1JKz5HlSHBpWwi6s8ZzQVVIzm+vUYY5pvFcsgRRro
kyZtWY/wI6GoQyeNPFPMq/ErytdIJgF7BFGLCTsDRRCSuOqFDXnpfyC3MuUNEidrY4zMK49AR+UK
S/i7zlBSmOQV9sk3yRIpIp6sVd5bAo3fYgTr3fkL60SV4/zFjEOW1yGQAnAWlbbUj+YhihqRcRxy
Nh0uhCxq1KvnALbQHskpuLd6h7vaMa2/4OwrSe2FvBs8ACbfwWSV76Am+6pYkSuIwsqn3FPF56b0
GIv8RBIF0duBgC4NEXouurVPnbhvtG9SYDWfkjCgUUG5u59J/gNgs1xK/PV3PTyVnGnwtcX6M03W
fh49Fp0zeiuLkaGASLXn8+Q7W+phlAbSL61GlJLOU80qk1DJwh+0h+WNnw3BbB7mogEiV61KOnhG
bOjrO9lUw8S7WRqscUHcc6poOTx3Gt3DHNh9NBhKsyn0n7M3cYanxLmUUiSlZ57LeHomwwfx+WtO
d47zqC7oW6etBsc22l2xO7NgyF9VQkEbF7p88zKq+1lcTLP6pkEN/e71CldHqlKxKLDKxQo7e8P9
97ZPxYPNN1+9kEPi5YUitZOCsRkPVcbwJBC+pbicg73J3YVsdFTTbZR80912n8aqBx9OeL4LNYLN
J0Zff41vtu/jqPkRR73dHAk/L+lzP7qfiuOHZY0qa+7c9iBqL+v31pMZfA5KxzoAplVoVsdiQ/wa
XhjMzuRUGMDn5NztdNDgAYwhQsRCwdTawTXHUXLgJz7F6mbEhOARsqb/FNktXaxwcLQhktBYjZOc
WDk6xxUsc0iGqpZ8mZdiuKwDT9RTo3HagZRmjKaOC5iwjSAt4rDUAyBzmGkx2I+qYFw9HsWSp64q
yzNS+hoh7uw6EERvDLRAXSHcJMOgHbOjd+Iourr1mKrPdOp3wEjgM48zb5D+pV8f8LPgua+fDWHY
N6PgeQmBQfFhdQpY5mgYNuAVybv3fqaMGpTEhRqlj13gt8PYbgHxmDmOE8Di9CSnDMffK4tB95/h
1lJR5cKAyI2DOFi1ZSGYMdLBcVA5LNKOBAILvv03mGROtr+1EEDFBmzaOLouXatK5UHXVvsYLmZN
5KOKSa81cediVSPCMCFt9zyQgiH5BS2SbWOepimoveF1jE0L9yGCxAiDLFgU/RtThCNgGey9QqWt
iaDs3tiJ4AgKwIePvjFaY2lSdQ9a2N0hs/Gc2SNoLqbnHVekfSO6GPfWRaiEQAAb5m4MSW0ok7oa
Y0AiK84u+L5q/4pij3N/N3gFen9zukv9ueHU+vyn8p7BoG5ZCEt4lG2pq0QissFho7sJqQxOhxnb
FZvyRkYJevfEvO40JCKaO+ETyDFN4wWwMFxJuT4FWSSk6MH/YtYI5hd9cjlXGMM=
`pragma protect end_protected
