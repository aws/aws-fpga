`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Kp0sj6pDYgXSzHJN01MWXiLc7uDajZBjf/VL7/+F8yEF0Mzp25UQWo2jOMKj76IEZvtqTfWOiVNC
lVaKYxW3VlURLxRXzgjzW8EIIQB2TL2T73xfEcAKN1qjzWfbAEOcueyLfEpIlgyxKHdAR9+QdCRZ
4jiJTZG8g+tbGygj3Zm4UyL2b9ckMBzNdXrAVoLf5i1CjAsfhyjnXpBJsRMRuRfU1C85Hvdof2cF
5uL+uk8qu4GmxCpKXPDs5POw+rOxRJkc9QoOdLWI2R2c0uFX7n+xiNIhHa7iBC+B2llzm8r1xTPu
v+/cpuk4PD0ljzjaNGirDGCZoFOTHEKcqtMapA==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
EJs0d7fFJ5Ng9c6gyu6QnRolhQfqQWrdc3ACWsu2Hlpo6qxYFZifhSfRs7NKDJSh+bqs8Pq+uCvT
sm22IS5qvZtT3ELAmp8DJpQK5l/sa+oM9HE119aaDhzFM5BW05M1g4WeYLk3ubzIhTqZpUD8Qi5E
NuslnKJ7NY6GMSsM5Qo=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
LnyU4mnRwW26rg3CNs6B2G/N68CM5vvXk8S+XHZstdXsrQQFBxTNXw9hInbBDTzRDJqzUU0q2E4c
k65OT6ncYFRSun1sy4h2PD7G/RqjSI7UGRm1brTmBJsNEE1WmZxdvEM1JMo343LyV71Asny4xThS
Yt7RwJbrZlvbRivOxl0=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 40544)
`pragma protect data_block
RGAjRyS095ViT068p2N5bM8OflUCZim77IB6BIwwHAxic8ASewYQ99fwtwwBHvs7G5OCVMHaGSqp
OzkB8gok0IhTqgIwufH7mMqj4PAoKOHr1pcX13k0h0glwnHPvI/xS2jluYWEUyWn1O8BNIwBUl07
JGPLyAbKKBN3E40Rk9em61NnO36n/Xl2sFmaCV4U/UShRi8eQpsEMtNJ/8cBf7ygM1Z64M9ndEv8
XCTHahDXLbxgQTaxMsBVqnZZJ/f4LEy4xACqLh5pcCHdnuvR6Uvd8rrg6lR3vYBcyvmBFtCyzZpJ
DMPH1GHPiTmhGEIgI2CuGm2rwXI73T8LgAfOp9rO9bmXSwm7vI45i6wOvUn2p/pA+6QbUQJ1PbCD
Fw6JQN4uzHg2RZG4Dl1Rb11T4x8Hs9DmB20gvYqABBes2zZAmrAgi3EyaM2QkG/vx0x0asAMdhWt
/bg177W3DIqRf0ZQvKOxMSAEkGim4AWdQU3hSwPVcWkRJPoKr/4c5+dSwBfO73SeUlYDU7GOb7Ka
NkEkzrtc9U9bIBKL7uIpIbu1aofcV98OMFBPtX3EsAab/S4NBAu70TUDB0fa5vLt/EkNhw66IBP7
N7J1gXsEw94HLdtwhouJZf2JoMt5JRHkQ6OdyPQ5VFXgWE4Hs6pZR4UOs7rrhmqaEU0ga23HqJ5r
IP1qpaH49kHO7nlPTBB308us9+tpUkV8M/2c9Xrg3qOT8ygY78JUnnkAuE7fdg9Gy3v+QIWaFNBi
EU53OfBQAnWe2r5a1zlAYFibTto73dKpwTHoFBMp8plEGASYhZq9W62x3GbLj6XTq3QLO6utMHr7
lSIkmbsjZYuTjUb/MVNmt1BEkYgb7GKd2suGojQGveXaNQY5czj+xpmwFZqYNGzv15Ah7JHFqyJu
MkZR3J/sgXrCbhyVLgaDYdkJze2TYcRhY+Dw0Hu2TI3xMA7VIFkzaffUvUwJiWQYTtvWjFMDagLh
KVwZ5wGZnVItOraExWAs15maiBQn3boUUc566BveP+HOQM+hhtvDs2ALpbD/8o/XEVbwkHjfcGjK
QGSTMia82FcOYmPuQ9uHCir9Z2MW6Pc47j5YTMswCkC7oCtnwVXgMoSjzopL7yTR3EXs1xDdU+Bg
37L3iQuThSjzbKqh1v1LvV8LlBCqhClq5C8JcQQ3rqmZNBm1d7JvWJCaDN4Oy60K2QEkE9GcB3kR
4JKDQo/Zh4l2h3xmozZQs0hVZrLpf6Ul4hBAFN7AP1vChMuTOOpyLT3hrTdfcv8kYHV17RaFNTko
g00w0BV/u6E60+l4NCW0ZxzWk0KzQiPmetxm42YFc2O56z8N0tQj+9/ysr6Ox1AxVRGEM3rX6jLO
5bc2qCEjIBm2Tx85nwfEpyu5f0cr/ZKrcz1pS28RmVnUeMSOMFPu2JgVfA7Nw6r8imo9YJfioHTp
VdGBednVPdPWlTCzMzIJ8s2HTGQdS4QU6pkvG7O7R60ToapcaJJ8JMaKvVqwGxjAJcLHJOWRckug
KXam2ni/5DFPepacjedRoCzRYWOXAYHY7scIZXHp0AwZV3EeqDlBQXj8JTiPIxMxSshHUMRfKzvh
NLmRh5F7hCQHx2bztOgtSh5sW6MHmZVI2Xh7dh07Lp3QLZCaS0hICs/HMa7aXnV4zgqiSTWWZiKF
IElGIAF8k0EyIa2oZNVEK0JiHn8TR7lSXAPdKhGQOAVobBFsptUJLpRBu5kRFdSCJQEdiafcFACS
/AzcYL+251kB3BzU/xR4QKrs9it2bUNOm5HLmdRLlcn8hdBpwdEP/AGek4cg1wC1lRigsIC0mfvG
/P/57dNjEwLRlvJW1SkvgC2EveYCfZ5W4Dc98+3+Wm/hiFCNolnbhD+SYNlNS+dXYaFI3d13vqAK
Fbq097ANLpyJOiPc1mdeJBjaGM6mY09LVFRFdky43rbK8pIRf43DjXOHA6NtPYXfoKHwH0ins84F
8OMlbp3Koizi8VPx6U2o6secHUGhpi+mkgUyCd4ZO6X7ROG+sMRFlSlcri/haRA5SuazDUwj/4zc
TuLUjVjRrw179yRbmrNEr7XACcDOm1LT/96jbf1INSIOhWAtxhXoS93VvHeCR2yGFPQSJdBVriRM
RhMDTpb+9NxZq4gh++tQsBgomQzZs7PkfVhdeB9TdzrdtS51mqBmWH+xX1dwIiunGERsn7QqQvmP
ErcS6mfztAKEcKZagV4CtVPRMoIjjmsGlZGPvOfEwYpzTpkk5ckUPE7VGRZaGbBeO6K/Cm7CpZwD
hk+Jj8BzuMW0lvTwGklB2yOeXAZl46jt5TEURABRp/k2KDA/82TaUvm0GzZODioIwpAFefboqgZQ
B7KbQKAMZvgbNfC5yMNeNV2Qyezu+kW4jDPgU88tLrikEyBtJNFVd5QhDfYsmkXkA3Dqy50nhtoO
+1EKO6dOd6Qxi4EmEFhINBFij9zWJfX2xvOGrMiSUXdJYI2Ak/3GNOzlLpdPgKFkEC0ra+GAOL0u
i+8tI0IGe85aBhLh+x0QJ8EnQx1ut/1li6cy4yJFJxQYeZKjoNechmYB/hPWrXZatf4ylNS5c0/G
xoqoJ7AAGlsSBMEVGmXLiFk0DJT7ThBQy1YszI8Ot/tKvaqc5DsbtCCOeaMi7Fk0nh0Hes/9p5gG
tNRFBJFOAxFmFXAxtiRkvnSwoJyZFAdfa3Yki3JkSmng+xU+LmLhOIdLgrhrBWNWcQPlacpl/vZp
M0kxAKGnYqdQK9RdfxzAb7V/X4QXXOk8c6gpyFmV6pATPauBCzWFOy/NVTY0N69Dlo/r44O90f6z
wZQjN9Loa8JhrtEkml8sHFOTKBNvKbAel0gp93mdStGtWEmgqC5u/zFx3J/kmpNUUMuIZg1dRpMx
fRbHkaFeezsnkA0TN7mGYfQwtIx4VY5RqZtUWkTsPkI9vLLP6bWUW8nYSTqo1FYnKK7Kgck5+mrz
pr10Y05fg1p+PhhvQ8mtopGgfBrgqgT4zHvxi/sRSWXBcUqai8H7heQL5qJ4ofm/FtN1HiYOm60/
E6V2wltzYiiAzjkD04BPD4rnLMKdCA2rFKKqfL7rDmmY2xnGT27aTAIL45VvzQ6YSARkGet949pQ
oHAXS9tqfIeydrnQIK3TLSINsOwZI6s/vBxjp9EHU17eODgKcuhTS/IYcE3WgPhK9xX1I4AK0pnV
CF/M2KM2bIE6elI4eB2qoXSEMuRS+MTO0E/tdWs6c5ixOlsAggaVGdPk1imRAg7lOjBGVkhR/cY5
lgfjaoXQbS+S7Kp6ggPQbEMURYFXQJ7tqTC6dT3Bmfpd3I+yQHEPUw9Xo4h/Qai0jquMT16JAUMb
xeqtEN8edZY9wrmFKAf8rULzSLA6gdxXHmO0tGsdTFzFQsYqPEltsEQGjMR9WMoyIlqRCO9AtsEx
YEs3L9aKKU0riHes6wpZcWuEW4slXA14U5Xj5uUeJqscbazmkmphlyCZUtwbWM+Iv13VQd4wLJsp
gAlwkHf7pX7qaFDgXaurDo5TMvaCmNq53yaw82813O5urRcf98sF20pY5j/srkWI0PospQaDQ7UY
dyEqUnsHCUgX5Q6ge1Z+/vWDCtUNnWAp4cJl+k6a+RViHLrlU7XE92WbLnJ2O8xsYm+rxxbtKXUq
tuD9KQjEeifO7MeNwSsSiS7yJn7W5JzSA5+nAqaq44zU4fLIdfmEqcWHk0Joz4xkYFeODgOS76tc
cctnt3cETuBEDQeGQT6aUfrWMxOAE1haOeuoOFrzikF7GYUR1/jjnB7SQAJqxIcB7Y6RJ2jq3NE0
bpQufoZ8ID+MSqb6GALlztw8BrH2BH7TQcmRoHILXA8yCMNvLeCF1fbKbsTFngbGywYjke1PtG/q
GjiHIXI9Ta5+3pb5XqTQU/kwhikF3Pd17goilPl/xSNCypbpt8/qaejiJkMR23jAKsaFujsPdi+A
eboQ6V0uImtOuhrOgGuidBfZBCRtE7YfUpVCkEHlJgwgZvsbm+FpzexNnoDfKDGDcDqDsV4WVxaH
0SaXzSv5ENNi4ojqhN/zfmBZIPvtNUbVTZPUow0ds0+3qAI1aKa+nenmnVHFlzS4MY7g7ojyro0M
haiedumn7hTHG9e+l6saEmcJHIsxIM5BaZdsBqUTdK2/6eEUVeZTFlmnrxhRZRZ78qHF5UmWU6N6
Q0ZMK0Z8BbW5GvOdU8uqYXdOl09MoGkxoMpiUWtz+Ii4xUqKo+ZmtWMBDxidAYGVH1pJ/d9+ugPr
E9/0nbW/7nfRnz3L4YdqoSmeezWdqEWFLUWaULawj4u/CsqCiL8+MZNGmLhPKSJnWHXHFEzGKRDn
7vbfKNe2LKo4hBZTRYpketGNCa6FP3QmpSYSsN6qTgtrX3M3WNz0fQl7apSlfjdZ74eqbinrqJtA
09DTrkeqAj3MeCs4p+ceVdKFJ4X55r14mV+wGv42PamMFxaHeWmXxCuh1akA+GbUB5+q/qUxyxSD
X9zfeOzwxI3TjwcAZMoLfbg71ToKgvfbrJ4h0S/bmDsqGX8UnTBAssnjYlne4ayyXsNYlDlwqYT9
yTJUbxcfffE2qJ+bGs6xu9KEomCxflwfIZISHVZAOS2gfoOI7vY3k5u632vOrO8K3I6dK0XcioM9
smx3Vyj66MHMEcWocl+/+9bgpI5qymud6kpGpx9y62E/sKuAr6o/lwsHVgnNjdVESCccQE8ZGqAy
k4oGbRk23dtVlba83N/7vN292oHjA929h8EJjT6f8EMusa2osMO8WtIZw9nQ/tbfvaWZmXU6/O4X
Qg5Zdm/cVsl8fGDat4GSwYKFwoqrIcGG1Z6bh8Gm0S21300GR7B3KRR5OkeXp/VcYUo60BFvK9Vm
jcET8Dd0zo1meO+5+7hbLhHYwoG8uH6eQPg1zeW46jGNPUCXWvka83HCLiWtdTBJHsZvwQHgEfcj
g53MDVqIHbmRswWZRUIVBYGMjYy/FW2MxGBb0n/8pPJBvugeogAo3ylNJ0y1XxOZadvI0tDRKJDX
KiXPvCIeMwtIslKpDdBPft2zemq8SJ+ShV4pLfQZS9V6qaaBDkmm9r1dUmgh6yddVp8ZimZRRJJo
LaJ+ASTBuxwBbuLlxuG0MGjDBtHd8z4w/xUzNBOEoIfsPjwfG8q3esxL/f8OPY1Udkyi5Gj1A2Pz
8wXYcBu4bFHv22igQy89i1Y3igIXBqKNnx7CAXuwP9OOMF/SbRPXbaXABPIqRYDXm0wyIfVp2sk3
OQyEZItXNhK+rphpno4OgBV2O14ncnMSqgMHIlpKBeaAGdsdAG9R46N8DL+N1/MaymSfTXvr/aLB
XoQFn+Ka/0A28KjGi4h9G7/HiZF5d403dEtpjEbuh9EwEGN5cFioQ6YcPY8ecumMkk489F8yvup1
8wVBbqhTd6aH044FtZCqWEIxzTNLDMQ/qOxjrF84H/s2hUh5/D/OJWWQ9gCAuCBMCOoFN089tGlj
tUHJOfetSRtof20i6cNDWJZ/1BO9xSJZkCdoWdJxrf3ZAgv3qbxoNY4BwcL881Ox/k+4121gFAEE
6c9djw4yaqSQ+P6RyI595tk5RN7fSkM5oGZyfOR8H1y+D3fQnWQiN3fPMVvhSXhl8JIwt5VrVlm+
BANqPLDMTJ2v4+RYdw0nTAgX1Swx8rcbdy4LdIpT/LAuXxNGAiKNqjS/Jvf6ZeRod4/eHhPx07OD
Q7mHezarurtmZrYbWpQWAf+XovT7kOrMSqmtSlaW1FgsFKMc337dt7WvX/IyUEq47dAIrGEAA4/W
Vn59Yw4WU9Cl5jnQsToLxZK6iF/qCdAc4SA+cYWE1UYfY+um0RiSeyarDpY/JxCbirK/o/vqkfl7
9C4TJ22iwkxB6wEMa48Pj0zVVTrB8ASX0Fqzp+UTQfEhp/L2alcfm+2OkNRfNGKKN2XWQv/1Jcet
XS9jrVK0gfcY2/7xfhSdoZyGb5qkJAy+n6zLD0pggBq7bG9+rYW2tauVWDONZq41fjdSouNHoPIU
GAVyZ0dtEiA4wcIBx5P5H9SuzXvAom9b8Em89VwLS7CM/zMHjBdJL5pQgA4bht53O1C9UoTWDh4V
3ratDeFMSy9ll+pIttZiCXBBlp3cZshe4j6QuOM4v0QMJQglJh3g/IadmgRvaaKfI4QfE9shnVle
VMZMIeCPol+n7eRXWzUz1MkiRKH5G4fMRXG0OKhArthWi2n5biDjhUwi+8+9CoYccIf+HtW29ajB
NNELPWyzYhhO3JIwq0YQ3suicaoYqNxyFYpXK5uml4QEvnHa2ZcGX0VKzXvy/Ml1yot09GX9LxcL
jZO9i++EZY6RuCIGcbZpg0UuyADj/E6Uxb7wthwF7pVQ6Rd5Dq/t9kdasiECmnSmNLtCU0+G2hzj
dO3PqRoyGhnfwrR8nv70lsSkmd/2E3mR/9Jq8CfWbBStuFoWghvc/l3Xvy/htD+6ZNEtwIpATovv
DA0oKkRs2AM1UD53dhBolKxp2oTYjCYUq6iNtF0awqyYPTDVdSR5ur9GUUG1FMoWr7wu8Y+ed1SO
C3d9oiff+4KKAMQzU3ccbTGNPE1lSADPN6eWYKeEaRts5Wq0ZkdUJM1vGMgC4e9uTK1DkxJl4lqM
gQqO69Hd6Zrzx24p7E9QB9AAlVMhFCZSvZgd8uLwmvRy4QOXmkPjDgATr9p4NalbxD82WIj4j0UH
bPmbUsa0fGEQHLTQzGKpUrd+e3meSzB81hAkTH/r/03Gb/ENnvA1XZqCySTylX6zfreHbx47Xg7k
j3nt6rYRuARjdEjZxQpn/qOy0fs9lpKZszdDPd3qMOs+bgikklDiQeoCOhxEeU4VcTRGDgOPva5o
EdWctGPoS+373ShcRI06OCZIoS1zTfnayI3j7xzMvOprsyNZwyMNhUfKC3hvreSlL5P5xG+jZy+a
OUMXGuvnhJ0pZe89/IPf85HtX0xoa5u/JqKoinEx/hbPLyCI6/xOueNuHYlMPYkBMx+MdQqQxVyk
xDghzLB9RFx8idx1FKEAZjtPOCKbPpZyBOZyg8CknzPk81yKqBis3xYqrzO8xXd/O4Ho4NqV5O32
TeOsDrVr+ZRAED4KF6FsWjvmTQG7wPyv1UouhJmpIn+Fy4hArN8XdjtjUoE9wkrpu5+R9GxJU38t
TGQPqHNHtBh+aUcnaNYxUsbZy3AOf7xRxKTzeFCtU//xgs8KQqtq57UZbNVhm4JlL4LZ2VnruCSv
L3KSvgzg1tZh8Znn8Jh6c3c7Kdk5G0HuMY9o8I4GPiPm+f6elSQE35Xsw+0HDCz7Lj5SvQLDOz6u
Q0FYBTQJqovSvTa4+YKdZ2tS8sQhGpsgJO82keSdFi2iPeHydBqQVGPnVID5mPOH19MGT2pw5mM7
2Bce/W4fJoVQ/hzN/6gui6qQDpLw9aJQ+4ynbQMBgVMVqyK1Sk0aT/QYiWP037E32JofLiWOFiFw
Ze9NjkJKNkn8yCUbUQbCd7jRwoL+OFnYx0vqRKghtrwYlHHHtMgI3cV/VUXwXv83J78uwBbJr8HN
WLRg5VF5CtOe973Nvfnd9KgOuNXKJkaeMHsXLhb+qVO3sj7/qnVYZcasxSjItnbnfiQgTvYBPNrr
fumsnZ1oHhYRixxviRcSXa7Damm95kDCWIBBF/wyEMeDuF/gHQMlJi/mv3ftczVrKVdIGTtYVSGz
Ylyynf+DVmQ3MZukvayZ8ZKbKtUAHfN6JnGIyCqwAmap7Bk6KQAId8ThwvIkMHXMzzGVUA3os7Ee
JfADm14uyeaOdgfqc30qR22v2wbb7MgRVFrKDtpMD6bs9iQJpjGD8NGsLyrXIv7gru+ZADFyicoa
kSBia8STJtsZKAbBdQswZogw383zQ2ac8qESD3nB7woBGlWl4IX8/LH1emh6apZF5ER89eIoSbfU
h1pgA9dSSnToY09Nt2/tcn7DoLfydFYqxleDZlyb5CxR1SSrly8fnUm7HEMSSqmG9OBLuQoQL/1a
K/4Op/Bl/MqUvaaOsWunW8SbcnBg9K8D5Pp3ig/Ts5N3KMbJCXTx33jnER36TzIWOcxPCncm9+o9
K8ccfkTYXRcDbMbUgFcALiTnBDhX/NGipp2W7tD+7ZXOyRpmIiJ5dcynyKe+uD3/+kLHzN3B6d3M
D2ZXB82q1ZjLQujsrmaXI0a9JX9n5Nff0CYDGbVDpXkrkdX69LQmdxIpF/rbP5Bcf5wPp6QqCOfb
4P421jbPh3kwbebcb1AYIaIxreEri0ffkdnFXl8xNx5SsIJJqmkq5XegRF6RPj0oIOEb0h1dZCTq
8pkpRZZHZQyg+sGdMadV3j4iy85ScuqHOU6mA1Kg0/QNrL3E3QFJxsB3JwMDdR3N01c2THPmjoJt
zWC/ljlgJNGjjgpiLypUIgp1kKUx66ytNCyZa/li8xGvE9ua5kivzeYF3FavfnV5cCPmQZZBewMA
sXrMsshi0PiZrf056j2+2Ykzms3PCJ8XQX46CQYog2P61RQH8rPzNw3ipx2gjp0sXj0zedvUZznw
55PWctyn3s7WXxz53IIgLN9wKtygnpeGYTxzb8AC4XzKskCLSmseWs9E1IHUThBLrlI8KZFJTuti
ejg+sNEyXzuZKoVbxicf870w+GhhIUVQTESgyZ/02e9XZOqylStA3kaH9QvxfDU4LdvqTe6D/Qkx
wSAJzN1FkNKgVvXJnDHe4ikGSY5oATFqxnSjRhBzNg8JE9Z9ZMTo+cAUJrgTtYrgJQ3JSQehZaLi
f7IM7wof7VH8EePZr8NsOgi8JTma3Ty9VK7u/zSXOTA9cwK8hQ2Wni7wiZHsK1CP/CTC6x7WPNOB
SCPDJVtvzclvUL5yCNXQQK1R72vaOSocgsS2YDddYNsKFU+nyNdqA82VriAnkX1DvOxZAoELASR7
FIj49rT7N33QSkKOY7jt4HRiFp3xBNg4ShZ9Bd3abvYv4U446DKrZ7+FJ0YurUFjXjXY1/Z63CZg
akYg3AiMS4ocYSPBq2suNM+vMtQOea/bjM+pDOXdb3x1CQeAXHKzeS3mavl1AePECPd2gek53K3V
2j0y9LBXmASpuuEzAfM0ZuzkD3Bw0oshQRc0M63+pXmLQa9oPc4/2gcSdEMTq1jvDiv5Ep+FFEHU
fJ4nVlBoYvbBrNAVRNoekpBH+PCOtw6wtVPx5aXdBS/NOB0eQaOxmBjwi+VpanaBes1LmM+nYUCA
70eDg3pRnbGGEqu2ip5/hCuNtDHzkLa4RtnFDU/3NFbk2BbwrpaHJFAX6xGFLOPJN5wN/KLvXf8z
XYOOwbc1ChMzd08npPmMQe2UI/X+7sSVZmU0HQWfocBTqV+ycja/gVDEnSf0mng4T6KlQ0gnstF+
bk6ptnaoqv8oYOhco4AgDrx9XR4JxiS+lUfizRieJOVi/S/AOqRpSHkpi48uYHnsi+xFR9Z0d2Hv
BE2zSEaWGDHriYUWQOSxQjwobY/Kux0WoUp7HKU+HxzcQiyZq2IFDHDbDn0agXh1Lz24awOqdZ4c
MFnDJ2XjJU0oNjRonE6/+yomFbFI1Hp99iQmmIYtUGXBaOx2J8yWLywbGUFAF4OX38t4shM+PNYS
Nmwa2fYqkm1ZmOClqDViyw3fELT4GSiVd+zSGIrXw++d9w8kmm/iB7H00GyWKip0Z3TRbBWKgYCo
+Hbr/sMa+2USZz7yXadJ12zSIPk5r3lvNtvjz5Wj/ejvzyRtWOALv1D6IU9G097tvyEHKJVb5rDW
l1VFeixffMQ2ajP5sM5Sd+7dbqQZTcFT0+VeVQsMSkpSgXsOIl7bir7kUAi8gHO93p/KXFW1VW8D
luZZTScgrBpbYudku/XFCc3BmJaXI7RWtvyrVICZHm9L1/7pWFrG41FxJLWcRcVE7O4wVIGubRpM
+Cy7PkQU47oUNN4Pt04DK9AZsE6hkV2Vurj3ix88VGel/enx1AeACPhfkuAVvs0YwzvnXnXDhgHL
Y4hDIduXUO5wtJTOl/qYCtGdKN2YV+DCFhukjb/q+Zs5sgIQckefU2ISo6IDwqL49XMKD+/4Tn30
zYCZAM7Mp4c67X7fJk023uNhlPRU9xW3e/JGIv4i5ktQvDuVTUi9BuEVOed5yzZUAqnVQWwb/CBD
TaRL1rqt4gkdMSr7DyfXkfRDjozFe/wdA527FXN2BZuqet68b39jufpMXR0Gy/WbUWwx49oPTAoM
Zsub3oMOCb+jjWO2nNxekYUjxsfFGAsllU1C94Mo5xH0DsJL+4AWnJ/bIkkjrY5oe/Zodwxq0gJ2
wsTzUmlKQT2tBrUeqhJBrSen9Eqszagp4Tp6FByfNjXJnrkm2McMNJ+m4YT6cHPVjKQCDU6Odi+4
HaOAmIosGwEc01jndIAOXqI/ZUOV2clzbVw0dUaeiOdfur0fM74K031DfPRKEqrfd6FDzEXi6vb3
K29jHmdkZN8cONT3D2gI1ZhVeynlXOw1B3uZf4n2An6jl/YL52oXRO3mScPf5vvPOvE4qVr3fmya
VPP7fjYGSMHIfTtw3kBAmd1/SFrLHB+tZJlrBUzHFxwrHh6bdY7b80ULiQzCcaPYhe/WY4ljj3Et
LadcwaX2Ii/vpu78wFUWi5HXvGp20qwB+Hd90TG4Gna4i1xjrSiHGXU1/AsuIi7uL9tlJTTyigm5
fklaivuPBf8vEbJ+nF678sAm6sfc078jV9GKZL5UgdLUaIVinLas2+7GbJ79GrREUwo1pPFPagfq
d3cb+NIiVEvjtdQKRpFCGSyGciVoZaII/wiJawAFS4K+oNTcVUgTg4vfUZQ6S0hb53BlfJVmCkk3
Qplu/KLp61wmo0vd4g6YedDUjcMMSSiK+lEJTbeRy/8vr/CoePkgO909bOMAKEsAQflC4UnKKIX1
jTm7ieCRTEac0IMg3sStHeLwfbFxkq1BV4pYna2LLD1cjH8n8q26Cx59hqfBCbS35mm5hWmgag2X
wN5l6UFBL1tETOjcPqf0tYHACIjgAc9AjYuXi8Xyac3NjK5gGtLJhuMHZFEE4Zv7cD0vkw7UK6jA
UfMsF82p+EcfHFp4JkMibA5ARNKOwVK0FfUEfR77SWl+m54eiuFlta4ADPxsvIcR7OV4ZvWmdAfz
UOskHcTUlUMaxQExZ/WdkYcdlOzqpouc63EB/1TWdHXJc4C/at1QOUW00l+xPLn9F1xlDvOFvhQQ
g4X3QNktrfJXuOPiS3GDWXjVXU9odozYLJJ3Bi1PhOewHPbvK0fpo1SFUkiVil52S86KxGaciei7
dtRHO/ihi/AuYrQQParXiWW7oDceD7KFSWDVuDozEU0dOTdTzwNkPPhdAr+zhoqHdZIFRt3a+d86
bbQaDQSJD+mo5X+pzTqgyYaBXUDrhboDtdHOE4XA4QELEhCW2IOYXvZ78YlpjhqkUchONIO2NzZO
lIck52pUvxQKbaFt7hDNnbcV0c3RyicEmnmb24m/zco4KJKw5fvn/p+L3w+9AEltVWCoHlDWy7B1
GtY6miS/vb4YzHk5BRSMIZwvn5jsSz4LsN5YgZoOktAP6C6Lh6HfVYgL9CCh9B6EI3P9qEppfvT0
mEF+bMdj/380XauRHYnN+4ps2LaK3U/8QbuzPDAiER/XUIhasDzk/lYEEwdPrucN1wiALl0gaUM6
CVdUuDCUyUqnhDWTmOQ8fj3bE7VPHwWlglHwhiGEohHVdBhPyuHucI/mcSbO8W4NLw6y2RO+5EiZ
WJoz83CqchVTvnygvRp06IX4G3nQ7WfFV4wmB3a5vo82mYtKLaffMoh48ObSaJdGYWO287BIsP5y
BQTJgTc2shHG/hMuPLLK/AVn9KwcmvSY63LC5+QVLTVbF4lDtbbnK4+nXHamWKM1f1I4hD7ZTqHg
nk3aSuu70ibALnDFNOv13C2sFeDTGEgd3hBiZj4f6eqo2t9AsBkcmS0KpFMVlmvlkV+i6LSFJwIP
vpLlcV9NlHajOx+O9NFVhCEnrEo2ctFIuNQMce0ZvIsT834ncGENDwSOw9EGxcVn+lDiq3gA4Ra6
Mv5crOM5/Ve2/v4xnDLRagoelGhPzZn54b55yiOVoAqhfeyRPB9uJX0jpnfvBbR5fnenqUhWfpoT
zj3EioZGFvbXOyz6nND7tBUhEfhFHncyGJnyFjgZsB87ml1zTxYh2lt9mqhKP4pZXpIfsUxoBJmV
Sl9D5kWuKEAaq38XdYODpj2PLscHlYJTWst1gkSFudofE/pkrT4MHXOSEBC+rqHJlfCIWP2JY21E
z+i3fVJkEQdRbBXLmvaevHb6EnrEjyt+j1sfZAdniqQtZHZijhhFgdF5KvrOWAdlWUCLc3ooewgg
K0ef5AGvRc2s7JdP138e/2vHL1AtPGt+Ra1+2wf4j8+W0KzUqBLmLCv/HwzPLVHn3Pvj4N2TSMqe
C/N1ugbJ2M/I14GTvt0+JBac3SuNIHWDOGUFyRVZ6YSdcaVx+bAdbG5V3qza/v6Mt+m74vEM8XRN
VYMBVL/hJ7EqxJEc+AxoWagHyVGhGEWngSxUBCe9++Eymt8oqfquuj0/X7SRVSeVyRVZYyaA0PNs
Uk7VV3HeNB3siiIwwpTUh65HkZF6yhx0J4zABbwMiqpb2CnQqg1sZDKjwaxvlIrUe8V54WZrmYlT
H1aoG/pSskvMqo8+hP9G13AI4M6DCVhlROFBceTAZnJj31c5MGgW4InnfLA+RngmuJyV0uIt+Lf/
LhFSpy8n6OPjZjKk13ga9miEoAGH9h3m6mL6iD9ilcXVfooEBVXQQm+fhIaR/ZMBxvpdEiFhhGUG
uj5j72eIpj77AvEFI9Tk6OrPRCKZ2dUjrk1FW/GCRg6TYZJ8P9H6I4NTGj9yJh6AXNJITA+aI34x
H9MAzKs1cNcRhBvh1JkHydNyxjEXaUFTpl1T38D4dJCotl4IUbgRTMivEhp7dnwCoJp6c4RD3KLS
NPbF7WysvJ9k4vQhCZcaNlCjgAJ3734Nc1N+aOL48hCzsNFk0uLnOuEPazgjSR1aEssOzlXAh6Gk
Qx1jZhCN1t3ChLgzrI8z9Yr3JQsa9MDM8p3iw+QaMiVf8YjA1MADHMayeO/FAA2oubPZTpxGrCtJ
qUHmuU4M9kk28nhT1sOOZaGp5Jk4gs6yYwvIT5VoOFpulIImxpI1lqszjDTXSf+wcpj+foX2DKoL
XZSo+P3fzt5XG21oJrDmpZYPBZVeIvbfiClAjIcFhQa544ZnKSl95BMMthjFBoz8JTkkxYDaAz6/
HB5dZzCBJV72EHVcDLerY21itCMLO5gy+y0CGc4Ewm7m2MBzS06tnHlbTsJ/NNlAs3U9QEQQ4HS0
pLCKCCMyS20FfWyBxM5pq9l30Uyn95UunmkTDgZBCAILA1SFHQ22mcQPK0We4VCYaCk8iWr/BucB
JvNjIwEkFebp4HJgBP9J1pWLetjEbv/RR/tjpCJ6+3kXwskUQAGOrUjub0IJiItOe8FPD20fhVjR
3ZYebAntctu3DdaLo3hi8wF4NDob5u1Qm8nHDiTNzTunslpieiqa3y6yf31Tp2JSv+ZVW+HyoUTh
RETf9+LuApn9YvvPVk2spcXQ9dOMHt/XwLpmMW1xVl2D/XrC4XNMeFI3zedS9tvCklAjIuVIeApA
eHs3lPIfteGQxiD3TXtbPR3VyW4/Vq8DWJAGMqryAl6kyT76kgywape+wc4O7oCDBcnOEGOHKc0D
MdMgb249KhkyLYwyC8NBvJTJ7jpzw6O/0BwtuZBfnohtk1Z/pxuFBWw0lsGdZO1EY2DGMU9w+29v
jQ8Xn+e6MrblWobR2QXiJ2wp2t08LMM++kK88ETPjd7a7FhiH9EXdwkxYi0q6bEAQB+ddHwxCaVB
Vhl2KgpI7WTcD0+0+ITepE9Zr07r+ElE3FKdWbusF/Wnmkxi4Iu/aqutPYGw6vKF7RcFbUkpHm2i
iOkoqq9WKHxjAtQR2WEODOql9XzxsMv0LUBW9KRE/AaNZq9EjuHBIZ33j4LRouE4VURvk4+C+WVE
KbtcfrJw9RPo4vaL9m3UuOkStEsn5VHKnDzCZFNwzI2yfgvycgv8YIKqQDWsMYThjTuE7PpTkw+n
T+huNIh3ftnJSeamlf0tkzWJiKmM5jG6naiXoGZKCGLVHm/RDa4/KseNSqSn/1X+bozQwfPmpVps
myogjKyYoqwun+B0HfCmuRdIAPd4Y4M8rmeSsiaVnT1P7Xd16iD9SbIdDYYdUstaTOgUfCXWKZdl
/PWCvZ7KDtBJ+7L9jbYkQLB4QRl1uUr7MIfnTq3QyRMi/uIdKShDSXWX99Y5AgttQzo8AB2xnKmV
tqtRjlP0kV2X6qqaujk9QHv8jPlwecFSaoxyKdL/CbMQZIxqFB0Gct+IeEwpTEo0V3Z3GgFeAxQq
nhQ0TSJpTCVhS4kZe5nI4FkreMGn2v/S+wneVveNWYLNnzTCqnl5mwgvN/cAkJ7MX1dY3pVnREgh
h+eq6Vz6TupTcAWw07LcBt9yDZQHQGIB8aG5Ogm178wXE4Smkxh2L2bZrquz9JEDS9cph1xgPriO
8xsIZYdgwERioalX6tHZk8BXPALLbqosD5ULUC+6gZlAXDpOIrmiIjORByzWDdez3ftjdkaf2wNy
Cy1Wx2QTCMDYREwDQeSan2UU3QsOIcKdwljvl4w3qba2LB+7HVuYVq445h5wAMzzHbcODzN6rjmk
J2B2SbxRtqZlEAiz83EC4RPBBZZUyiI5Cbg/haek9izHdpEkzEKW+gw4zUXaH+eBaEcs9xEhQOPl
Dc103FO22U5fd5vHdz1ZvNK3f8FMwsYAya8KLh/IcOeWGO+DTRNRksSQFCsFFX6cj/xnUAElI/Nq
5apJ0VEhXymqLCgCfa71+Pj2+mSGqQhEXxl9gE5Sb8dvjLFbLnpQxfgdgq0jygscYfspGuPNjcdc
pavcTiq9lko+ecgNrSCfjtOb4lVFe7KrZyDl3GfDxHfNDKNQP3qLkFJbSliRTafQbMQI4MrRZyDc
VPyAmqBIQunEUSt0u2JMiyIMZTDZcDCWEuHF9ciGYdeV9ctNMvTruZ1mVRrsX7WKumEb7ctd/yJt
cqXPoRtr1qlRk7rmA/5+WCV+Qzr/c60lIhx3hqj+XBTCLDRwPfazAnWuAms75ek/tvK1wxT3sOf4
Mc+r08PLS5PYNYFdJ3T+1rlPMFXCVDUHq5M11nNh2/geCBXTMr6Ag6oLO0AxbaliTe0K1epbEdEc
yI8xfTguGj9ioy2JpVdE7qTq8/20zS3fl4ImdGfTeSHtIt+oK1MWhVfYREyKmf18TDyFyYYju9R0
lyOqX9Hlo6SfZ6EShRnFW3IbPzog7OzI41mdmmPMWQtvR6nqmY0CNrAirImB0UvKte5GWz0IomKc
X/0yvvg0pJS7oj1Rvz8qKmTvB4L1s4/hraE9rwQCC1C9yBML6RyjZpkI7txcGDufAQ3bLkP779Gg
xDSoh2TOBtwfeG7YZxzmKjU8eJdywcwq9jbdYwgMKqBWfYYhle+5aQHG4bnyhdmZBPXy2KKiKbnh
MalTQ1Q14y+f8h/wNLUPo9ms8p0VFMaMwlzCfYfITq54/jaaxJ2OG4pqmnXTyBTw8c0xqYgXM1hF
Ur7KZKFqDyyQobcm46bkvIJqiGrP3KEuNk2Svndg9fc8O+vhOgNQWYKx6yF4PLCvwfSanABnhGy9
UBI7DbOviLRiPXyD9amuYRvZdk2/6ST0y4KS1oCnGBYznUrimgapdBZilbCvq91ZQl32gBD5Flke
hl+sunrSMNBKzI2PL1skRuUN0nyVdqHslchg6QraR44IwUby90GBlGCiPKTkJ11fWHl4R4EElR2C
MTtYsVBy9XRhNU8UvF1Wf9JNlnH0Bo/qTUSnjDzwUqnGhUeVua90K+O7nytrRyjT35p610Z7WwHy
BKX8R4KsUNVj3R8F2kDdDfaSQGOI8JT2G+p4lNEGzktzbKYMgBu96uf2tRdDwmeBzpG/cMuESOV8
OrDZPWq5cYVg9YOpBUsRa6C1cHS3wOqRtU81xrH9jt4ujPHYQ07ek1eOOWf21SxnglACOMigF9kG
NVD1VgQMCWolnT479kz85JEdURwghkpjY6+XZkzbgpGJZpG0rv6sE8bq30/EWLNGszAUVKJdi2+f
+ZSnMNqRrlGOHTC7LtXQPPEs/7sJLnQpnGh+ITFwTAFiRQf2XO8zo3HB5/6ajVPZ+CxR8ImtDFf6
UvPILAqaWRdKmYBjIMUdQuhhuQdC7zSDAXxlA2hwhpMU/Do1TEWrCiAJQjFs/qE4e2t5Xv9gsnTT
gpSuEdyfJwAtuXx7rdcNvYvGguNjXSpWFp9VX/iAsa5T+RQMDgHlDc8R536ir5SP0Fm9crrjQ/1u
2Vv9P+XdgDtZyZVThGsPA/fKS+vZunZT5OwIYcm6SXRSk6+k6+unQmAEb3aKZ4CEPMp29/Ws4Vpu
apjMqVra8/agpRZyFHA0OppT9/GQAKQ6XSh12qdFyNWofth1aHhKpHY/Ljm8Gdk//g5DauJEbl0h
NhIqmCuuo4qa/YCF15Iid1U39CEr8IBGu20T+d2bjAIXabFmLh0+qSdJakfwbc5+JJCeiDHnC7DI
wEI+AzLElH8vbg95vAgzdB+AHu5iLKBse2CvGW0asdFWjSlfxDIn3/exGwA9yPCtvtdaua8cvxhq
ouaMNj4q3xRSqI4y6Vj+x3JIQUxM8FHaL0vdHnFqVD4xl9AQtZx739GDwkw6V9Ph6WPpSOSdgUXf
o8A9zouILH2MCMzXFlhfJf54nL7eojyYRxzNDE+7NGA69SqelBX/dRP6J3NLV+AACsDYdKl+0U+g
x3aOujPpAT+9PBMIZob9i2vK423p4AFp1zG+xOJo8iCKhJzwLQfq+hS+9fQnRJIvtPdbhpTeK7Us
q2hPF9pkkSWDiYZthxAf7O9aoQ1OrZTw5fclCvFqtVdOWmtpUlB3GJ2QC1q+T1hdxa1Bklr2s0mG
RydnuiMoUMeeNgsAZKj/sSutPc1UhPIINFx/Th0S5QqiWdr92SJkSSqDky0WV19rR3UQ0qju/YB8
VzX/tJNJmPUHZRCR8syAr8EYHMj5NleOln7jrh9qyI68ZoBGpgidMWLQlwm9V/YltaoaL1OlyGUS
W3j1/X0SF7x9aXA8J2Lc2vMt9SRca7sbsA4yEPuqNieC/8leo7PRPFPUSPM4do71rm3GJ8vaEO8Y
Ei90ayo5lJ+XtCW+lxGp72tsXxIXOEefI4zL7mZuZEowFVyq57fmx67vntvVj5KsuBA9c7rfPy34
VJbj7n+141cKol7C7yhhAlWQd+lxNthtT5n6JC5yWRmwSa/8MpKoM4xp77unUHEi6EtK+Pa3Ewvf
TjY72+bSH95Z4pAvkmfOxxRIxeYdieLD598fQT+mFhh1jgLIPV7tq2a4cJiFxuQNPehhKpZIDwTQ
zIRH1N/LvtGT7E9GDBkrWWJjaeRU+TfI1e1DsUFTC6JlIKKJZ4KIvbvxBvhyfaA2g6QGwK0TtGoW
WuOScehRFaChFhHoZt1KhfsoLxY5PFfli4YgUyWZ6BY9PPTRhv/DgU7IdHHpnwKWWuoxLdAUpVV+
CUjugdoN4v8ZLPV9k3RqV5uZYhrLuO5oJUC7zl4pKDAQJliPMWvuJllaKiDbErgqLk8gRdeJRIrx
BmDM5kbOQpvP0mN381QlwzaGy/5CDJ3nS7erRWJ23ny3UiiwBZINdIfm04sCnkYn7C0hhCExJrQe
oSE/D6NZIE81ro45CZuLXwpZ7Q86a9tvC45qN4P9i5hI3XFaYtZZGkB5Pii4k/M9mC0XnfVOKRM4
Xu79WLo6hoK4drPSbJj1B1k8Yi6wXghldjPNO3vTJsHQ1gzCtY86Jl2gRLP5R5lZ0B3DAUOrAHJH
Ozk3TBa/YS0s1pSgdGvZZrgfvix+p2xfypwSxSeniU9SR5x7qVk+hFMDLtTGajV/JqN/IeippY4p
/8TUOQeG48rkmYodxHiGQE9FbNajR8okYQGdcQEUSHcygM0PZBe+anIPW0gOcpd0HAt7BZQd7wc0
+/2BWTWbTuJtxntARSKzqGYlj2FawkyVtJsMfz4sLLyzm3JJEmk8H2ybG7iIUIqJ+aINpOOa8lIh
YOq2ShCGrAE5R90xoEEGtXvs45tiE9gK+jFClGjvJlXDdyyEZshNluJkx+BKHZfxe4KEWD5ZhvaE
jfNI3772bgfOq7g2HXNutJ+UvcIX9ZE/P3jSPCiF1AtXZLXNlC5ph5KbWQPHh3YQ4WmoCpmjNZia
4YY69CEH6Em0GVvC1AgEC0vQom2l2/iLr1+h7JC88pxDkDEbtwcTMUYkH6P/Kp5r0sm5Pip8uqad
OPm2rZS4x1lDh0yQZKEaMTstDPpDMGUUkQmlJNo7jutvvUWSUQfOv69v6cUOD8LiLrcvYsOLwjMF
4xJnP/iNxeJMAA0kQPIDqUhBvCCvDB8R3rjGL1k5k22Qcveve8WQPE1Ul/w7uho9R+KOpDOt9K7h
vfWTfgjFer72GMCotoBoYTvr2g7ejR+rTe3MNhVL4PgM9nR71Vs5eVk/Uw40tsFgN9xAKCiPKh6Z
W8ONrhjSoB6z2+D/8GqbtGj6iDt/pzwUMH+eMUeZiRXA3evLH3HUHBmaNGuFDX0TqQvB/xj8UT3Q
Y+NF26C+9+3n2BsAeeKUITKM73VnRhgASAGzDQ8jqLfKqipBcJUOK0AbrAs/Fs1wDh+SxUvySOrP
ThS01TlicSwFNCfDx7rhcOEIPnzlNxErjNmUk2is5W+ZU96uEfevy3DbZMhQ9A0WRCI1Hlmo26K4
Djt59zEHw8l3Bv+5d3cQx8uzAPtDVkoi8boin8QnN7PUCe3E7qdBdMOfpTfq6m/b4XbzS23Dq8v1
jBucbyabwT6/s4l1Tz/Jjyv1tD4Oel0ncu5s2BvGgCi96P5/mm75QbroES//chGSu8cQk508HijN
UxdsoyPXaMsPPzViDhlnszRx7HkTZuo9QUI6QUv9R/kFsPwhdsD+Dra3r1qDyqMYPSkJla5JCTk0
pwu6f0DBPF42kDGgcAksgmgRtgwPYcrRtJ7glSBCSHYG4ypuH8gXcxZnsZgfa/WFKkjEc7f5g6bA
okyltdtro8wPXwtbt75SFuEH35ixRqggtpWd1tWJeUVk553zrBWtN5jn9mivOzIwyIj5k1CjYzBp
gKeaxiZVQGi6HhrLYajWt4KSlPvNEF9OBWd/Ag1D3+dV4HmR4MA9Wmze8vkGu1xSmYWowW2PJzXk
1XN6tuIg4nVrVkaui6qawdurtPFHVenuFUYVBzqlyuQmk17aUxp+3txoVPY/CrU53QH7yw+5jd8a
o0bOZgWtCEfbb2W717b6rH4u3zmehlf6OACOgLRmVksqQbMk0TQ8CChU1qUYYdeyxiLeL5Pm48hn
SSpKoeiTvFMvAmYIDldqrKF/p0bcYjW13PTYVXwLCbkLkJoprVfpJevGrf+8yommpq0W4SpImOTl
wZCT7vtnBjDkO+RUasx2S4u1Nk0jBc9EVEIj57Pq4h6kWmYmndDhyeD6RQjaUAp7UUa8NzrLuuyn
6AOelVfoZevjE6LbuN2G+P43rqlTx5tCbNOLVuM6M/FrphUGjDL0AB/uIw8al0fK++sexkwSW37h
Xgvkk9D4IRnrmfz8+inw4n8pN4lkCmYrigH1eiGH6EJ2ibPRRC0gPvWsQI8vrFc8SIiqVbk23wnN
0Ku0DivQsIvUsg7RpsD85xUVzkXbs8hFAwdO3+B3wkEnL3+bHihche0TX7yXe9MsB0yUBjajfgwo
pVLaNzKpoT1X0ybdF8XBIwQHHfDNX0KiA07u8nYR6iwjVY0NwigcyjzVXJOrDu+IE5eq/jRLUj8W
HdupVvC4HqUY03V7DUinf9YJwIJbKe8dksP/9YnxlvFiU15wyNND2aLcngUmvS0L4+WTWUAtbhtN
b75Pr3ML6LlVsj5K9iCjTaE5vxBnRHnC1HlCXJ+RUK+W4VXEI/ihHZUeTcuhpnYsbXj6EuPhOPGz
ObzJIjnEPIQ249LN0hg6XT6OdTeznDOxw16ey0RAGhh7CVlwy055kFY3zlmsiDsG7V2mEGs8HlzJ
ILJ/viLADCOtq0IXgdTZZ0HD10b4SiiNQCxyjACmbXIKJyupBS3xxeRkHSGyFt2dOyltn1MJcfB8
zUR/sckC9BvxW4NmtbSWHD95v49ncO62/c1nD7ZeKvezxlSeYvm//88b2n6LDfe//CY6MbHY/VSj
2QZMHl4uE4QxxWjeiVh15MlH0PYht6+ex2g9ZNGdsS7Di2W/FfSmAlwyTPcXJ6/u3QT5Belvj5mC
/idbeeAJM+oBNXXU+PatOhUaijx6L0qSuH8JSYW/UH+TlzlY6iAN7D5+Hfz3U9ZIzwYI36qEqLqs
PRV0vlkgs3vS8MweZKss4Vm5QTQRyZWEA1OV78LSUpLRLSHDH/ZBWx75+j7AvKIXhk3XwZy/w0ph
rHobWixIhBmLshDNtq29S6pmjQy3JjCMNRJLFfBeN3esEu0KcZgbEdOTBCaeQ4aZwjN5CSkcdf8B
5YCQ1sLLzUubxd0poHKpqra1rDNLK+fopjCFD28U9SQ2vqL7MZEBl7eI2iXt7l5EotQ/vQvJMt0F
hB2ku2a36OyoDGOxXd+YSkdO5a9vz9umrbp0zyr9WdUQBeBoSYNnNzeU7c3NBg83taFdnmFDdncD
Qv09jKGYXKnC87MnNhM9eohUM1cCf8Op11IlfLEGlVADvRBAaeZ5p1TVVtXvmCsg3QklAslbvxZb
y1Ax0vRGU7igT0rvBOZK+SK1fe+EqcgUTdd74DE8duw8psteWPc5aIQFbgOackQCMBU0QPALqE1l
LZCBGHdDQYJzRPS4HWQE4PSDlWIOu961ybxs4KaH6UUOOw7U2+fuEu1QC8eqHdfOB4eJzA/Dl2zQ
13TXP9ZiajGtr7MvOpjn6rPVuNfL09OQugeNwb+Qcv6V5f3NtHM2+pUu9e7X8diH1Ko+L07zOGaD
PbNKylboE7hNiBAnU5Wb5ZR1NW/D91/vyimnlFyTy1UI+o6vot/0L2iXC1JkgmgUtoLRPppZL/qf
KW5UiBY1pEU08j8g5RT81e6DVwyx1KRmbTDhHMAxJK/Pr/jSeAv4f1VMqIFMixhEwjsJxm0vr8pc
OF1YOZG0ze2Y2nUtwwpMZF9PNw2Wfc4oun2REUrsuLBf79+DaFklw3vgtyC8bAKxV1BqgDXRYfx6
82btdeHCJlFsJnGFkhvihu4Bd3qGVCm9Zl5L1h4zKAlulW17tlNNStJnYjYB+zEdBhWImOm0el9i
fj5HTACX6NiYtc0lFfzUdc9Z/bw+hI1gB0w3TzQn6i3jRnTMaz85BNeX1osAAbSpU1nIAledyt/j
4XYIwJFM4J8gX+BMuk4/hiYjpf5VD1A07zCCQf/zLaVFRxApT3WMWrHEBKWdQkuR7h6RBwrSvXZG
R0sdoCDv6UMaGCsjjdAjAGSU/nxQnWRfu7ZZsCPn9nb2XQD9jPy/21+V/iKHEMKvDCbP959vKz0G
BqE6kNHCZtDJada+WLxYK2EfVznXOxZtJDN0Jn/U2/vZnCHEn44Frc6zYp09z+3JIM5X/Up8bz+h
BCC1xSKqs8w0IDV95vxvmJMVr9+SF2RvuboJUAqfB9VVVeD4Ya0WIsYN6EqeI3tMscLV5/V4Gjmm
S2QNZOp+WwAiKdRLo3v4ECyvL27cjVkTCwn+tVQD9kmrq1v8Fy+hSHBhkYJ6T9cppajE4J+kSray
debvH8oQMSF2A0K1RIbBR57WHo75cmCyJnUqp2sPQHFv15ZFZWdb4NB0aPP12ZS1P5CWDsSLI/Fz
exhMr4LPu9/+mr5K5SX+z1F8uF2w/glJ9yD8zP8/J/ckrHlxENQE9dCyhIiL1KCIjdWIRDzIXOff
rrCgLc6U7wn9DGWM6oG8Lw8wIX5cjOrJUwpfLkqEVF2l1IiZevBgFvlOgw0/mNaMJqk5HhLBxfFy
4A0E8wyJ4QKhbVDdaoYD9rSHsv8yGCmBJnYAzkcUx/NiJ7AT5gKecwcGrH9nbw5smN2D9NObfvnj
DG0iBncEhcmJX4BXFP+9a7vni2LKFJXUCjCJzd/9/kz6045H7sJSbOA/EwqcMTqR24xk45bbwExM
Ajq1WT/ltinn/1NbKKoK2CAW4HZdT2K3Y6FU8wCF4xK7/fzpHRMvnpzaxIqT98rrEzbXXUoYrL/N
1GqXtfj3i1gq5MxXXHtWCuGR5UcSUd69W4JRvybW8l5ZAqAW2RWV+Cf2CKyd1lgUQZ8WJoiIEP61
0UaUT6MzkMcS0jDwFPXlMtPW7cJwNecmEFw11ygWjv3qD6slsg//aaECy9PFT/waQBbS6ZiB6pEG
UCbdrWVPpuI8j+4Kgu4LfzeGFr0gOQ25XBvgRZf+R+aHKoVWgaRXO/clzFbhLmOIra2rZqyguYw6
VEQXRWkRZaMbi0Kiqd8SskKPv7nDfBkbbMkyzaOcSyw2S9B3rNYEOQcxog3wrHbH9aa6N9xewwrG
MAVV+RYQAZ25adfKfR/kvCQ3Ih7mNUz7Bpyy8gGX2QBcaz2nz1MbAnzow0TejWOGxw7dgwUtC/VN
lj5NuoJ5nkBXK6slcIUxqwTJBjjKMyqJEKXmXZyKgndg6v8vM25sc5YvSmi7de4ZF5K7g/loo4GU
GGvV7eLuMNXjEVJ/CvGOg8KDvzdljVQhyLNAbbzs2OEOWfk7EVQ/rQdBZzSym65rDPga5DmvjQDo
+KM9Mm7og9z1RYfCzAVi2HY8vj/IkqbSl9/IU3mSsZSvDEr+QA2TH6vZZ6pyxlljcZDIgG6OhDp3
t+ausG5g971jXVnJTIV9enOf0DasgRruP0kVZUtKH7zZAxDmCeBVOc6WzmQOL59TrzzfaEGqIxTB
B4oIK2+pcy6jAckpjxZ/f/OqNZLXcjjv5wDcvXfRTKIVSIykYHwELTFW9Sed/xGL9XUzdRoT4cEW
eqW49zDxYijuqqSeLXyR8DEIefl5WG8a4ku52qCv3wrVN/ugDsWTAqj4FZvRWAWPEoQC33I7vLLl
hPOfv6SWFKq8SUeZlq/4+pL4hpRgm8B7dH4zGMGrM+rIVyh6/WWK9NLtSlOXr6UnOoiOB2Th73EB
Dg342kBj41rknzwIIZACshH9NXr+4Pt4neE8Xjy1J2Zly+XPOuLpU85JD8QgFtE9evbRJKQsPGMZ
yV0rKSh49Xwgg3OfeCmzFVw17AF11xq0Ernqx+Hojtoyt/QO6EhpLy643AOlpiVCERPXvepcK9mo
aB5D3sDyOTkpeScNhRtuh/iUK7V6cdpWID/rR1nxwEMoBJG2D/IGEXlwSAQGuZ+tm9jqyxTLkF1w
LTnwhd6zPGiHjEyVvJzQzvB/9eC6k5RZh/uTGVUdDuC//qwaVaqdEg9oKIysaAN7CqdwmMAv/tj+
IS23BAzmTVMkBndiHpL8moTJhuloU/Mgi+m6R3ec/aXubMiLDmTkwtaOP+WKEbQ8lpvut6V+95Z1
jFXfvix9tV4XEnQCNJjrgeLLfOfjzAD14QBqgDha5hhjxn/UKi2mk1w5UcEOTM+GpVG2s4+AV9/y
NhiObaN8aJx6gE9CIO42IbqzFjsomz5UC9syaLH7CWYpvUjo2KT9DKhCqpI1vKAnqDzjQFcKIvck
wxKrYDAJTbmrrd9ZsoG/hFSeokSsj4JZ3QI4cKcel4Sm0eOpzcCNWDTZvpxdY+Bgoc7kGYkcdu9+
x9PDMztcwHMepaPGVMX9SrCR6x16ynGucD7Ejh8GxUwKnzOYLiGme2mRQSs7JGjcZI6ENkdZcsfz
Wh+T2ZsOopbG+ztWSbeViuisbZdXYOUvA7yV2XplyOGa0xVSZCNZQg4sJATTYC0OG/50bYePdIMz
RPuIJ21s9X8ECrvWv/wX4QnaD65dpXpqncaZcOT1+1l5bgrPoVnlsiJMP5Nm10ysPTGZFXBit+qY
3Ehbs3Y0ewDqTvzLpghBODopHVvjUSWEtLgHQHFK8exkagEQnaXAgTUhpK/hZyV9UJlp1wHExygt
AU38UqWtBYNSjffOlkGjdrA6Ts0ZnX9Xr2a0fNPUB+sU0OJUC4xy3Cw90QT+bWSnAhdmwNblwZCa
FESMStnHkItT3/Ev/EqR9XbNrIaSp7xxLcc3pvEMgslv8QopUSmNBBWon6LbqKhxeYNQgkseoq7Y
W9ucIn5a9hyiQEALDIFQtxEd4O9lHhxl+a+pJMhPp7wvLojWWFY37f92oiiDjuFp9/IfvVkp1PPh
IxuSSttAFD0Y1ZMscwsy1RmNtHG9OFdKSJeg2uKr5+EqXoX06E6knxwxdw8rO1SEHPa+J+Xr/KCP
4SB+MTuEaSt19+MMPIR/G+8iYDOWvkX0H4/UJvHrugCBrva6XFu2+DLqyAw71s7qLzC59mJEnqM5
QRvNOwZEL3NHxqWQvx86/thhiAcjoINR+l/Wnt4QRfPRUMG8vGl6AWC4gd4A0XfBepm5aMM/xoFZ
01LdvIAZLet17czdcr3yzYRzBrxOXevDiguVTlj8uvNI2zFMjdZW6gAGHmAS7eYyHscVzCDyQM9X
Vy4gUzWkK/z7GkwcTet/Q0pm8XK9CPJMYGJUv254d6zPua9cr7pgnC1Xm0t22/o+dg+K59/pu+SC
F33kHZ2M3HQk1iNDa7p0XyGFw/9q5tH6I1CQKoolxvQqtyXVpWPVBDVhTY5pFOK90qQJY41zcjG6
4qSQXWFl4Guj1wx+GuAxJgYYTyv61toCZ8YVCbWvckrDnnais/iBWHAW3vWWk+WlBkIkI6IUs7aG
Hem8g3pxvszL8ttjmV8mRnVuOD0mDVE/QpNmbAT6AKEDL9RCeBmWi6A7cybfsK7q52ou7AGTZHWi
BuSp1tTGvJLAA4x0YpogR8bSKnRhelTyH9rhXO50irtnVAL2WwNQXJZW8xrQo2vmwR/QvUkP0205
BYrO4Nd+yt4UGBeks7R0iGex3nKBBH3bFmNBYp9rVdN6J+6Q2T8f2Tw0/USxlnpYjouxW+OCV3sQ
HwuX7cl56M4pLOHjsimm1yeUjEkEGQcM1I43+ew+WJgkoN12P4nyfpn9StklTvr5k/lml/rywSC/
+MyzZejFG6pUKJl41kJ07loGBfwcRHlLtl2wFGZIx1iZQa1zvRXyFlj8Ml+pgr/s2nA/v+eBi+E/
DycPamdSzxPfdupSO2r5hmfejlevEL1GmXybe5enG7+cfidtl9rlu/d2X+b+VYELMibk5H+uVmmv
Kcx0uR/EJLnG1rGRNzkkqxb+B39NHXD4OpZ0pLU11/Q/ODJVZ2lFy4M6FEa+M+Xzq6ljEKIEkpGH
59ZMzRtDDgbYg5oxq8Ijtw0WzkM7gIwIu2Cp80WmPlqgIAj1xzuJEHNv/eG2rBdpZ8wHxSoEI4Sn
BdCV4AdsiDGZaQsl4cqhlvvqjcbKLNsIXB2YPR1uybVeom/GkM0OoFMH5trvSUFBv9grvL1Nt4Oz
bZdFcBxH6gPJlfXvbRgd+Pclky8d/0rv+Wxqk4Oo2UVE+sJJo2GUMacZkgIDOEWx7NAHHJHCcd7E
Z3nYCJ67ewIsOD+ZdcC0VAhHlHa3ZpzdaxVnauehDCB2xLT5YK6ff699M8R+sezNkM3iJeJ/UyAE
R5/trLbp4mATqbp3riSvauq7KERdnz6NkufFKHRqmmQ4uh5WYtdKYLqrkWZtz6RCIPhQUlQn1aWY
8qja9KtehAv/1aXg08svrVwg5jjzYnbBQdguCeB2LsKiN/hUvEtuvIU/EGdmB67K7+ovk9+XNQ62
jX2hfg5dDCQd+3S2wRFez4yOFi5sMH9Ybk9DnIvUD8m7uGfGASJGSA/mwajeHwqZVEb3WUfIlzcS
r6ggB/HZhd2kfROmjmm24la5YqBNELBF58QKoqTqFiU7mUALjuEoQNNBIbuBM3kZhObptxlBjZl7
cV7AU5/OW2ICcrhSyAVw9WfFoNSrRUwdR7NTEzP9QB7AkQwvXX4fWGnCBw2bzBp86TvQlxxUxfFF
X8aUznEc7S2GEk9vEJPKc3rjN9NpHHpsZjN/XxIopZs4gDZ0+gg18yLg7S6HynlvS3GjQpK1FnSf
fqMrP0nah+2myaJElNrzatE2063/f+JE0AovrLLDtc4heB4qwzSYpwNydDEI4y/qFnclZ3Syxu6N
0Wn85HaxMvCdNp2AJAWjvBpSaNvvdjygBurOUO/eRiAhJgLuhIzLGbxtJ4rW+JatMdAkvMdfDdbr
YumLxusEJ6Jcb+4Ey11rPJ2T7FNO4xTGA6fMr9VH87r4u1JPxYKkpgu1WwhK3qbli/ljhYd4Bju7
C8FKj4EGAZqrWlheTYp6cTwYuIGyS/CQtsO2a4sdJ+Ue0FWnPvdJUxDG7+dtIJOwh0NtQPpBZk+Y
RHZ1yvhsU4bImQICqJB7Eq7aDScFGD1Upc2F8OMkslEuVl2p0JX6SmTFrqf865ABGJu/LlAySpPI
5X7U5BMuEz9skBYFSwKlixm+Rcx6WdCRQh9IeAXodu3nS7bhhgmje24NcrtvZwSSBnroFH4iuNfR
MMQsw6woYt/aJQwAEnAXC3rrUUysNS3zfjF8Ssi/2St6uWgzLuchSCeE+21tImz61KWF/nhYsKkK
dqsCzHk8lYzdLP2Omuj6w5UnaF3FpQ/EnslDkTctDeg9shKZ21EVI964u/yLGq4jycRrtZ9GzBJu
OeSW1YLkamoMHv6BhHzz69RokIgKcj4WUa1EVTmB/FsMjnASYh6Xy1hPwxCR1Iy7efV2dq6rmvrQ
hzfCgs37bGezB54I3BVFN039sK3UFFQLQIG4jO/Gb4Fu4iL0dxu6kT0tBuKBxQdHjiKq584vz1I5
MKtMl7vaRZoYt1AbPvmN6ueW1jY/NtSmNn6w/w+paYWaRS4UHiJ7EWtLEe4JWrdU86+EtnJ5JQFw
ieZsNHHY+H1KXsHj1d63yTxV9mvsgnq3r6WeF/DWzIRNaBJrb4NPtFd5UuqbxuA/f7AJ5rOhqKUV
za6jD7d92FDuRtdw04YHwtYQx3ujLYw9rzuHmbPboWnmj29Fjfvm2qFQaILzB09PNv7sIyozRXaF
ia8tPHXJDQQNTOdYhQtIKpLyTLJ1L/CAi5l6rY2tiBurlWkWjJ6e+Ulfxccavu1jCYuD9bo+31t5
YXMy/ux10y1d2KjIahevPU/Y+qC+6eYDeMHca5uA4pTF6F/OT/NqEI0UdAMija2kyjW82agDWlNL
BO1DKVU7d7sX6+fbUi2lZ7zI7TbshUYmCuA1dAuVqMajDN+S1KO9WJv+r4v7LgkofI5O/NL7maw1
eMAiSaXiArKF8k1sZCVJH2oL3Sqd17jxJDwDJc0v7N73dWzb/lpCvL5yjBchh+iTRxcSID+au7iN
ChQ6Dw6149jBorrPHXCZAyw95IirLy/nre3d418vB/F/1+Ajp0zJkUNwOsG40AZJgcCb7xnjsO2Y
RnwHMYHTuP5EyjZ4xZHBHX7Q1KNuVKEuUCxwSpefmi4CutKGLj88kndoxzfMVE+E10sK64T+Zxb7
IeIwPF8kwMCMt6Sgb/vcPGZbKG40ysE6hbmgCSgLkSvMQpRkhrUZxgCCc+/Sqj+er/f8fzu0YO3D
1I8zFGxisk5hY9EXFH68F9+3WrfdqaQ2q6lui0f8saQX2PIBzWJ+zYWVXmIWf0vE9AJmmEqYVHyt
qU5DzmVxz86jYpSjnbPQvQ/+xdHyuuU9JI/snprNKmcBnBi2b6tsgscgsYP8xaZjXPzb/Coxt75U
gNxFXiFexDad0PmRFiPrIcKsSJuYUJVe0TUzZ32W0jxEdht5zn8L71c++SDHvgerO1kNrEAJdEHe
HLtTA7R9DLvDUrNijrIsjL+f5kna5N5bkEiH9rkNGYfhCiR5QRoXvLs1PFBOEmLAv18wWFA7go4o
0j06aj10IQGeNdXtVF5ShRQOWdH6ghED46cWUZ4VwyIy7wSl3sWbxpuGKvlJwC8mRKjzuLaWBhDq
4KSzQ8eqEfS7acsi/we4qImSBrARqZTwjPCt2xe5R5sVdiVPr1lTobn9GCGGEpAJ6bCeMd3zbm1/
U+O8GRAB9zTiBydmoB7D7MXHomWLjhdSNXba6KEVwKoGnDodTzeQQ72d+45Qb46Blt1KX8WOFZEI
pnp1xRavRm7FazQPGOtDpl0g6CW+SG9kH/10XiyUApZzf0Iz8B9Sftzqj0H0mb8Fc8lFjj7JvEtp
LIrWrhwbqdyW+4GZFlb1Pkq66f5Wv5+QccVh6bNLFh8+8UTFESNS8xXhaKwoI33/0GH3iJ1VfDrm
Z6DFV6offni/Y0SlmGyOhAc5iKUHmE5R3n7DFv0vMzksivQkxk6XtB5aFlzM5tLn2xrwtIKmruph
qsWYeoM64FWwGAZvPe4L361+fO+F56iCkcjjsLpvZIlTrbsGNPP1FQi7SJp88NUaGokCcoPAUsPN
aYKGA8uhWqMaHXg7evTqH3oXu5iTsbInlHFZ24aOVzR7nHLCdYKpjpIARSBk1SZRuDwIgE+ti7qa
0I7U8XSzurytykWpv4lWMu5XtNOR+d4+A65eDJIDu9Aq6PuSywNwVuOU0pnHzf2DlmFLYuIhXaQt
SXGRRhb2fksCdn4VQGgBopSvAkm1VgmpOilfLGETmjrV5RcvFdpJ4y5v49WAl0sjR4DD/Mm2l3mH
7RsrTxTxoB66noUuYcg/5JxrU+HiNIVJZvngeJSk4fnTuCIhC2o+6CAFxRymYdEpZXGjLs/tzYAw
OwxiXXyYxOCH0HJoZk525bAPHoSH7KO7r6jAiJO1967Jvu+Q3sUxAoAtVgnv4iB8wYNq643JzLsb
DG6kft3Rv0seZzhdvhvgs56WMdDFZ65iaCM7ygx1Lv6E4SG/48nSIftiJ6g8zdpsfHrBJaZ6g/GL
LY6Wnt6stZfxfydokBwdRov49ytSpzTQC9e7+18hf4a64VkOXivOtiYXpU2woONlKbjqoBZXEnKb
0R5RZXm+V/quHV8X8Q59xHXkKHynULo25/g/EBZiiy80ew7JUCFenIOlM4S0hNQBW2bIOkr8SqKw
+v+WiA95p3CrJYtW0OQvo6VjZh6lqeKwkwbHqAl3eTItvAcA8thpqTQ+bms8yz9dy/t5XGRJ3AJF
rRJtHdN/pguQM2ZvOdgFlOAX+j5FN47rW00hrM0o2wtBse55Bg0wMQAg1mJECbepWDvlb+ut+1gW
Mjrl0wYCfUhSqHxRYFNXUGRK/JTI+4qLrwvkdXjqR+U1CxHthAGDEa9oIWml+7LXWzwptKdrh09q
Gx2z5RtbLupNske0z1F6iDjEDcN7wfcE4aP/lPt6DghSmzPwy0i7czIRVPxp/GEzpeQ7c1IF39zP
WhXj0jbKIr7UWdFaBAQfIPh5Dblkr6l/hvqvUICfqgHEpGcEtI1P5Scn/DqrUiKODPJLFYKoMUEn
vbvrRAMNKkse5T0jQ/0ih/WOzLUlFcazSAP2PNrSERVO8dr4AT1Tw0rvTsgjqQqzAOd3XNIKmAl8
oRs0shubb//W92T2GC/K/sUu9PvYoBMIcuLknl3/pOQqQQjMnVtSwBWOEzSE681H6tGhhBwUgUat
4TIGw82Iqa/UfyhbRAFuQwO7KHQeGKdKcV1LR7ClIaQHY35pfJmKc+NTYPf9qteiRfruVS0LgZfX
TxRKKDM2wGx+4ckeo08qFZighl+rLPM83sQkvLevjaUJIdiXQYfsGW2eOppPPxjb2txnxbH7MX3y
SWOm1Rge+Z2Zql9NEzxYYu1PSX1FoQQuWKoY8r3TMqCJJ2aokypw1DIdS1H8CdP0HPTMZUpRDWVM
zKwMJMxHJs6uRGGOZaC0kP2TytCDedPjBPCgdt9Up14KJQAKGiDAUdkQisGPpfHHgttPb5wAqCit
LuKQYFfWpvK8EpDB4/Z5Z3/BNdQfkTMGB9nsDJUyGF6ZxgFwj1Wiv38jN8to3DxUyfR96lS0fF7f
SYLWj7U0rDPs7rps95F+AS+5A9+eBE37cNpApOIC2hqiuhLyc3oMko0SwyNFXn9qk6fQlxes7eSX
Yp7LpIDCDz6EmbOV46dbi0k9WRhNhnxlWGlP0yZYZ7gnXkNESdz5f6tGtf0jLWTg77JcWyjySL8L
D+xV+cCNYb4x3j6CHbJ91GfK65JR5USCTCaMFkrtaff65dkXt0dfpNWZYN45U3rmCeM2wFCX69LO
u/imxAb/DQH4OLGw3dLN3E+nlIOwKikC7hyssfUsDYzmkp3AeB9HLrGYwoj8g64WdhzCBgNmHfoT
6plCbHy3G1UuB9cqfFvoioT/Dic7i70k0xqYUkXmSOiWbdZjpNNZliyrSdzXDl7nd2YNJuVcw3RD
MqmRt/ccDLzvKAQugxtzLLpAqwW+tLhJua92JhhJ8ou40yXEftS9NFkG3x1dKRiP0/nJCexBKSJM
ydpoS9+uCve3tslh7KJyCosUxTb8XQNYlYFdxGTBGG3bBbfbT32UJdC/vyR+pTcWic9V2XD8yO5f
ZaeRdgxnBoVSUOOX0o2V8K/vJhVGVkPigEibX/meDXD16mNTaMbmxhkY6y1BXVkA78TPsQjeNbuW
OLh8OcRO2XV2vcwDD9kxiFg6NC6zdWbETpGEfEbng802YVdYTkDqB4ApAqAsZCpACta/hsGBywiv
urN2yW+0NQ4dihTG76qJ0giVM10aQ9NAmdH/zi6xm1+sM9TbuIfMlO2H7CS489caBns+6ceJo4rz
aC/i+V4Yk134rzUX+imMObxARKgJ5lqRfgtSLqFZ89nE+TSMBNlJXLL/yswB2VRIIeBEmk5NjLsE
2rdw82TmgeaZJmDZ9OxaNUXz0dZjModYwi4dYjKDgYT16opBNoiLWVpYYXBsGj8jJkf0agDfuu9q
q1cUliVQEZ/67PUE/yOJqKOCKicmJWCm9KwGzhIaFjolx/b8SBlrW403QS4TAstOLD3E27O9zAJe
XXuKtfNDic6kxnABzpk11PkcX0RtS6rnQMAop+Li62HiFim6a097BWY8Fd1UOHJY4kBaagtEAQMO
U7ln/BzSfSrFSVGK2yG0o4KrtDOB1Q2Voo9t1Z0xRcKEld3fNB1P2QuFuA44z7GQCog4crizK5+/
Epu9OYSK459MO1v98Ho6+9fLxz/Ido+UNt9RaIaCMYitxSog6uZNzxz55zKoYk5czYdY/pi7rE88
PH+5AborDIH/6lFzlrX1HpsGzHvWP+vhnvFx1BlA/sdv9CtV+EzGMxGaP/92xDEQjqc4xLcfT79Z
01VJKwzu0EpnF7LF2OctXn8CStcquOOc1LDCNM8W1yp9d0H9NYFGDbRqI2AE5xOViE5AMxRasp0T
nlElYkYzLw4djQ2IzlBbefhKJO40ZUfJoIjVAhmk3R6o+rwQPyRv+ije+faNFT2sS3hCOOYb05f/
+ZXxAwLTYlzISjFGrUOPfeU8jMVAer66cql3FTSvlZkRGnlsFsFz1q7pFBGoPELLDTH0Yp1m5mDk
nauhCgMUp0+D9andTdfQnpCBi52eBZwLf7hhYkC7tzXgYeKKMJRWlfIZtLz32oD9+V3SbJRaXVHa
Aa/xyqMJkRvN7l3sXV1Ns/Nne8hK0lKQOJm6+ZjekKmJ6UFG7IX23P34bgAHRGPbG9YVk5LInqcP
4szmN8J2K1i6yRwwoR3MbGQoruj2dddgNa4GUm7JeYM+Ch+/BRQa9GQ8DwGT3nRVqqJpmHO4rrTj
GdcYLkAAPy+7JJ/AMTe9bfMgCDNwY0fHgBTYxjSdIztfWAVI6d3vx1ssDzxaYyCFMORK1xAJmPOu
4JIOVngFoBlpUqrEXRex5Eb2vYfUX146vEo28E/Zy8gLtQojhsSnzcOB3xzdvRuR4ZhD/KPYROR6
jhVOAGE+9D9auh+cbNGz5A7CVPVe8uOJdT/I7/6rd5bB4RZt09xh4FiwrbhMM5Pu+v+18jHcZg8H
HTNHa+I7K8uYNHEQ4ZcSOFamaeHi3JKLLmskgkQ229PR8dKhdpBITrG353cC2f+wlDOiPXVkHeIW
WbLTwDIFaZySRitrTMlfQYht7VWIJIeMkCdqo/FSQ8k83bDuFXWrnnYuD624RtfJBTg3zDdRH8jc
bxUFDe29VuwjfYxGxDix93TwqDU5wSwepxvTrL159/tCXnhwVadB6ymiqbXrH+B8aTNWD9qIgWsg
E0NA2rlQHzUohsSFgyUrogI/HewjbCa46mkzeUEfc8AFaaAdzIn36FeY3H18abw98wkQ3du7kw21
zrl3fg4wfBD3PFFQy4Cvv1YrhnUqS83PmJq78LNYPA+2NkzsChhNe/msl9dv7FkMugMBpuQYaR25
K6fo2YiD4JWKl9sZUDrpDpMKKc1GtEnk7fMPuqM+zvoBZUdINUR5B3vuypfEUxAp5E/wjNSYyMPB
xvuC8kjvrdjH1trvYNjXw5neae9WjUu36ktbLvqyNrEy1tA0Eblmp/6lxysj20w+5wKVD08plY9m
h0ZQFmMRgUhRLe5Re4x8OMP3ui/ncxXBIzUd8w7iL9KeW7n5aqVTdF03cLTsn+kOdXP151iNZ4bz
3iKIQ4cw5lbAeHnEg82AqTKMoBYJ9gfppyjzZvPcfW0RUHc8249CIc5qCMnmzSf1/xwT/XjS5Q3p
YWQ7O3Zq4758VxCh9KD4f7JtdjpPTUYfUBI1cyoKuWl9h7xVFDdvYuxR+zrfPe9LIznFAMyd/d+a
Ze63wNlcdKbiF6Vj0/CKC58cqXSgNcN69DShLNucBAgO0r2Myr9yZBL7bYWgUhbx515QZUTCbbJF
pDNIVkW6p85fwBTDuVt49uVRUl7Q8ygU2YxXqbdOasKqm8bPU5gk9yktacTZWcqbnsrqQ52DVFhq
3gNGMLnXF53ClfpMFMBkqu4RzEhN6b5K6oneNEput/YYRi8X7mnf7DAp40XblG1FQCXDcySG/vUk
cMuA/ejNNmYHUm5JEL4Sy6HDx9yOZblbCUSYu6lIw0tL9UUEL3hUrD99tYOfMQxYoeFOMsZFPVMD
qXy3S27Y0Sq+NVmjHsZLMfoZD50SS+VhZdkyjZ2ZRjfzKWnmAvB3CxswqSvwu/w030E04YrTEB3T
uiLogKNvu2eBcf4jPhSwBXAJHpLeGFwAEOfRuoK4gbNSX/kVc06TJ1S3EvNSjkeClBD2xW8IHW1Y
vtcZQ/hHoy6lXg1u0eKng0h5/hDlrbdcC3vJbxE+QZbmo2kjOhz1sId8Nf6RpomgchyyyOYS/4zn
sFj/BTuTqzEfvappypcGCKXUQ1bX63aqMtZsyMbd7+AHcTDpxDFxV98VJGwxAAFaiRyOlVOvPg1F
lAqg44RSLupEmXMYDpWV1vRCe8dKZeUXDqf7zcX1lTZygnYqkRismwqRXk1xKUUMt9Bz3apY1c5W
LHx7V8bBEPoSMy/GiR6v9s1fWypLFLb7eMuj0zAwKsVahQmIkuzKObmcLKq/tfnjs8b/QBwlq74e
chmIzzMwHotCftS1SVpropupg2WG8LBieopYU7eDQhsiiXzt3PHTKnHQ2K2EoshsNRK4ScED8o3e
NqsCONZPhsI6gDSRfWw+qcknyyfXmwq8sD8z8jbs/YIXRQak19gmCS4w3k3MWVO1URs+COJ+y4Lp
yruAya71WwyiiaGhI1rXort+OQOWw+tPcEdb6unGFfdsnJlBQhAFHk3WgHKr08MxfK64T+R6JVHt
Jh55pwCuermMKrG5HixhTvSMzYT5BCc5xix11EN0HtahMyKigcBKP3oIQttYvcwFT04uaVYuuNB+
KNM4dtE0yiDyXdh4ddsIyMlHytc5AITkTaQes/3nUVvQBTAitCkbslfGv6E91KXB7zvhP04df11C
SQQlzzqpGVIy5dmMiB2pspCuG31lc/KAsF9YTrTcp+CYV+4Sx6XTfP3xOSs0TPMMNIV5p7aG9dup
1U+WnVVI1lL+i3V8bndhF6e1xgNC5PVRIkmeXmpe+mneU+K9OSpI4aKDpR/A73dgyj5ZL+JCEyxD
njuwVKTL+5G4YWMZ9yN+Hfknin+AWjnVxSNb/2MjFBv20FybIgKzUfaiUC634K50PyPP16wOvk2N
31LG4qhLH6TG52ayTa64Rz1rmHm6w0/eUHnG4RXt9JUyiV4BKByw4xcFiAGN+vW37XS11v73yi8E
lWQqdYxq4Qdb6piKNe978h3ACNz9dpLlRgqusEF08BNDMw5u5TYoz1BlDF26SqYgnWfvgyzYAOA+
NL/10Jhq+qD+PVcb4ldaCmQ/EthQEwdaTZiXGrxSYHXIGdDG1iG4liDy0IRtENt/qS5TRGOpi/O2
SHoIF7XK6SYm+5Cso5YVAckCD20+6LFNiY2cNP4nXrc5d4aOomU5YqplFScC+gX2Nyn1NsQxtgqq
IxWkI2dmoQKD2BHSQO6FuLPt6IWDQB16/l8XzdwgMuNpkWcM24Lf8KpXSmOPDDuDELgP4E/RmE19
wEQPllH8KXfmESjED7bI5ddlvTpWUm97RD4mvCF0ZoA/9ao56JjsJ2MqNqJQ6vKswPf/eOR9B+lq
osaZKU7nDRqF5LuGWwHp1L4b0UpSat2SO0NT5segK2eddBIeT8EckWX5N2LE95mQ4k9sO+2pxCzN
bt6RjnaM6hG7EAUYhoB85KgOZX6rP6xpJYlZ6OEIkl2vN+5pscn+wnsIa+TzsrLdrI9yz5X4zcFA
OyYHdC2nAStIHDQvG2BTTwmoz3w2jBnULO/92csh8fVQF0xjrE4VKCJmovR4PYJUQxLO7x+Yvehn
XiOjs9ew0NCPXvaNe+CiSuqj9ZOr8YJ0cEArFPwgFNo71DFFcBqK/IwePpZJyQKI9qRwN9qDh6Ow
qrKBYfce0KhtsyktDH1fD/3AvQzNI2OuU93QKWyRol5V3yWCDnJWDZRQAmyYmZL9ez1Zgmtl0+l4
lWn9nx6vn4rIgz8164lee/SVZVisCXnZCimzmlWCGjkrFt9OmnT3LESRpadZtDrffQq1O2Ecc2Ct
oh8h+fUH3ZaXDkVP9LyoUgamgB3B2LZsvrq6tmoO23TzgktW7SFVvPQd85sge4eIKqpWQ/4M4epB
KTAs+a6ssJtK2oCU7bwYxztVvO1RfODw2KVqDsPueP1zZDdaRjhaW6pGeaWcQTv1zu8rbY0U7GJK
95Ixe2l6BeODbs1dDTK9bAdrkZD6EgT576/mRPGbfK5v0MYCQ2IZTJ/JKFIfLLX9Pm6ARy8wyPTC
INsYmpW7ONmHUYzhVgfVMSuugdE1DioteCmtz5bD9Q1p3iuKtrt8WmA5AKN+Ft784I5VWsBRQ22o
LS9Ky5AXSWvPzWpnCsH2BvzBpjUXIoDmBY0A/ipWXsBzxqPC7QaoRF3pVXHjrBtZJWoBUl0IN3Zm
Z/+RD1eXcvrOtHHjRpTy0DcOIuOgXuCd+hdVf/tplfvySdRcPhGxnleU7uDQHuwd/hx64lfvuPwH
ZO1KlAe7soDXDAlFLD9yW/2LvproHUHPx09oyRKeR19hjKM5XBLOho9+HSzYbS6LUruGs5xxsZbY
O+RF3T58lEis8j+23orEbMygZ78QwYB+Ggl6fMsHfloacgKimkeZN9osQ9em9mw5EE5kU3E+KCWt
CT5pKUJMHdBhwsPExH+7owklGzrNEwo82AeTtZevHTAhEsXIZEjHnimKfnt8I/HRyCUDTnkDBrVM
6n6sbUiLK3LICZHiLOV/t9hCC1fzXdijrar7ddmXYsCDjTGlCS+L8IudxuSlN//6k4SdyAaVje5p
TvLsxT60kUqSY47if6Zu2A7gACoSQAc9l5hjnjEHg5j9TVG/wHBvaQk31YQI+8Oclyn3QxlxLzRs
NUmee+Sh+tEr0bA4hZtWeeV2WHbrAhWVA54MWTY0331CNYeCsnNgszy1DFVtNVH3CZrPHdNtTm4K
Xm/AY8P95ucn9gLgo/c5tRJOvjoau9DmU5b0f1f/EFe+I3EV3Seaborqi3xUzESattqLytvl5Ocd
VX1nYckEFNdhylbIcEUvnSipJQlpGP72aY8sEFAzbD+7la+/nOM0D80X68okHikPnNH/MNs5TpVb
I/vyjgKJD8Bu7IYtqgJtvhSwrd0ep/CIsnUamPFc/7uoZpGGRz43LBglddX0b0SL5oYKrj2ti/uQ
kfc8JTzEcTYEqazm4rsA+XAlssh8EcD1NeZoBZ7Ntk3dFHS5zEOOMIbpNNio56H8Gt1tvW+SgE/p
Qkk155V8AL6318sKlY8+NvdpHjVL1EZqyvueOy7XMF2VNkRfbq0xiW8URdY/GcRagy6OpD1t3Na0
X4WiR7QIKNb/VRgScg8sN0kQX2B1lqpuj5BQOTAWAujLXMuM9RV1DVfNsMm/GCDFof2SlYRPL61s
OyP/JrVRP4nyjvwqVCaBy2SwHe2Lpg61k6n5Xb5CcrOZL0JcbQA7AX7BQlBNZMvD/AO9FK0AyvMY
I+cSZVtfXDcDGaPvf+DA438NsspU3uu0oTNmJMhvlkHMMNeM4tzR0XOpuEC9lfP98y7Mw+P22CeE
sCzYZekiOZnNymXeU6ek0QJY/IIfsvCEtj7BTN+Oh65l4W1x5bdiqS2NA2xpp4kiuZH3BRklQFHH
JhjY+/ZGCrcSFgqWOQ2LUCIhaW8weMlX79BEhLQu6TxMzZAIkAJDex87/Ra6y4PROQqf6VXqhWnN
PkV30hbvbTUuGI3zlmuW9//7acAgq7YoekkhBM3ZQ+OhT7IQ4fDQRs1VQb6O16kfiDv5sk67wfay
86WyfJ8wQ3xNezReLBlorefPtNidJAKILle88XIQ5Gxsk19ipEp5k4nvzb+mra09xvzDkCrBZP6a
rMnteohr9qo3GwVGd1VLldlkAMJHxB+1O+xA0b5Zj4XJeR6G8iXGCOhoiiZi3Qt33qgp0NHXOtkr
XmIyTqXnLICzpV3rA0YmTqvqt4yB8DeMsvK68zuas8p6HokVxMv6FyP7LGSjpwezMP6/XnWTiIkW
0zdb4KU+pvnkjAggbQ7HbUvGLyJGx8KCwOQfUg/Jb51EGckJYYI9UAqKCqL1W6BCz3AgvQGvwHVO
SXNc9HJZg3Cv2vTbGhZTzQtGOXR4MlDSuY9iZkLvL7Q5onnjPlaHeGNujoMVRPwI468uY0ESDuCc
vUkmEcBtP8Mh94se5M7NPJXSxfYqa1HL90+yiQWbT9ICMRQmiRhW7KP5ZPUrnpoNWfVXBSFFFocn
qYpM9mgFruCH+NfZCgwEECZD82aC7aE8AfCOObi0O39iMLYUFQYvRmn7mWN9f1QzOfwQwvRtsBwb
BLt2+QqxCTgVHIXU6tdD/1qdgtNl8YaMoDcDdj6gxPlSUTIpaPcQROlny59dXXqcJBIx2iASJ0O3
Ufv+FSYuu2XM972jYXsxA1DDaFZ4SOeBz6tgT8qrFyEKRSzRmDAv9UwhDg9JyDqzeEBL2D1QWZuz
p3uyzrxHYAbizka/6qjR4kGYXsBLRWkBUeIMBfLOYv8YXv5tHvQXZKV//5pj3q9OwNWdm41dbsav
fvOEsxz8Gzfv5+zWZTR6IZxEGUOy6GOZjmo1n+myDPRaOEaIoJhpoZwmrMITjdx47EsVLDk0YpId
Btfb9tL+kMj+ChRERF7i3h6UWPPumI0u9VDRpTSTgCqCjlzjZVUZ6gFzN3UCF265v84wPrC8w06F
8/CnhHTghyym42comsH/A8h4IIaq4CWaGpgxJlQtXiy8QZ+3AGZuYuvZ50Iys3+Qoz7pHxj+0Isu
+4W48WOlP5Ll8m8S2DnS9KXgOYYiRRuaxiD6hZn3irDHANfNpxhRqPtul4JOYrD0XsloXWhUhVlw
2KO1ZjEFrd4TcSb7PlyNIgPiwvjVKA23cmL/crxDRp5wVU1WBjfXl595NZftgEzihcuPiMsKv54g
65O8VLzdwAbF4PMwcMZ9Pye1PSFBUrKidb/bM2e51ZOlqpyhTzxlIQIMOSrKTN8EAmBmXE3Ab6Qa
Z/V5n7g1sSNWEkGVkjM1YAm/ds3ck7DLi4jZQpwPmuG05gOjicXiEBYfcQG1kZptDBpa1aU2Ndc3
sm0X5fBnhKEdOY8zhXFdUJXLVrnaRi9lATP4PoW6SDG8ESdGgM2taQM/k7cFG7pVX3dnczFIwKy1
+vhedfCEL36IFPnUN29niVoHJfkCIU16tybvTtyGigE+lrmRBnkanvv4LcXC0f2k6TVLwTt9/7Ko
fsNHr9s7bNFBVUwR8Ql1GbetnMgScMmGlHkErLKaWfCEtbrlJub3kodlOlGFYoOGlcjIUQhhjMTm
Ocsihb1Q17QFJ9rRu267ReF6qMhOE/OMDYPLpity+4FgoAINiXv4y4g4g4ONQtVmwIFnOqhsv1Km
l9bzEs17b7giEsdi5p0ELQrlfPdfcUuHgq7p31Dv9xe2VSXDob5yZ0NTxi/7hgPJGnZDZgR/hfaY
zGfuotkLXOKSJ2kVtjVoTpCIiAR8TT5GJ2n1m8EUj15uIY1XAMtwHJz6c9zh5lNfOnRx0Y88u87y
lRnzehHQIGgp3NkYKas7X45fRevxrSeTpBE0Kbiw7/S8e/D6DD8OYJMJEsS4b2Y3w+GKN0G4THBz
evVVLjria9P5OWLWiFnabI5AOKKyXwqw0Z9/zLHnRTm2qCE3Id7jJjbCTY68eoWy8YiDdyHuR66J
2qBhA/hAtBZ08P7d25QuZggA7Yk6lfhlMC3ESzo49BNUwFS48i5rzYCZQLyGHSyKSE6IpC/uRVSE
QmJa8YUP2RBP4JVShr0IPW/BIX2qnL6b6hjQsr9gumReY4O+F1cfOpsObCMbaMZgfaCXAEcWBq7c
nbL7rJiXRCm2WfBeahx+6Gt/Eo/QYahloSzwrw4ST68DK27f596SbnDLjRZnhbFw5bFAukwledo+
LExWZJP7qfOSujuXoBesHe84UNjz8qdoPSOET5vHzWu+JOwm4uXX6KEqzEyyBcHN8/MorVPkFSfM
ltHXrPH2MFQAW+3wuoeNukigqrL9FzaEfkcK2ZQ+151epRdDqb0q7g3AQK+fxPG01YbqLPv4salf
cHwB48wPJhhhQUDIcyrwPloPrhs50R14QM7PqQGIlhk31t+QZEXlRERaI9mvkUKz860u0E72ICCB
KnyuVqM6PNFUwSixGqsyzYCZWJAPBotDMiEM3w5LPI1pPKInc1uMourw7XGtRoyglQ8hI40k6pST
kaKP34sqRh89nanePrgj5EU7zAC+VF1MgIJv3ZUXtoab1GCJ3b7Q3xQecSanVtFZesjj04CWcoFe
LMd8+0s2fbq+Xa/g7XqUsde8d/dWXFEgpCbhQEK99E45T9MVZWLkuCxw5pJMB37J9eWS0KW/cDfB
lxU9D5gsXDxaHIP4Znz0Kt5S4Yf0PXTrvHhx7VvO/4E47PENWGsSFV8NKUKf4N8NMlLB1O/JzNPA
gsFUNSVJ2lvvAgKp56GJFzbPOEgr2gwuXJyNlf8Prv/1mBpMmK8TqcF8Nd+B9iNGNE0GdUN5PEHr
WCWY+2mvryh+/nXHzaMGwMb6gcgX21TPAl1P44c0EPNBKP+rABadqOcb67LjqB1cU6Vdtay2Z/wb
qVOh1/FxmPeV67QF/fOy6emC2xz/QjVzqFFGq8m878C5kuag9aNTNIxLESCeG3sDqjyGlFLpm/cl
FXriouDAwKC62k3YLSWGbqyFtf675VBrElRJBtXUOd5OxE6vFBUQVFQD7r9mGEXj7xZBHgej7fM9
X7BBqb/8442/q2i7cyiAzTHMPscmfZ49zRYf6t/3zTBKLYlvfOqgbRq5i70Huw8wHuyJFCvAWxZ7
4ql38qQJv1lY63VdPXJrDWBGcpDDXYMW3XYAMFfdj4btxiD+qwfcilL4ev3aQkMth5Ia6md5GBVH
BW0OFZ4iuscMGELQchs0LjxpXQqheZL2QJGm7L+mwdOG2xALQ6YhhJcWmjcTIbi0qgutXhiDP6iY
bxOtV/tNGo4M1TTyKsugEc6jToQxtmgs3tEMJtbNdnVV0zLfjOpb0dL5PC5eK6sc1tRG1qg+KKSy
8MyRVy0rCKbVf0dJY3rKNJOhl0jX3S8thFRK52kweyT2ez7/H45Ampj+4DAL4+LLjc09d6/BQUsT
QKCHnGmtz3PA0Sa18qw6AJ8hIiWbKIa25aTERNj8xcVCEyhFkQJTP7CQI40xhP5uZ1dN0HBhskqb
FzZjbBMPrNtvcBJB63Qvy5o2id6wtXRFw/KBJwgcpKVs8JS8uZ81pbpNU9QWlQK/s0loEBZfpopG
30V0cYcfc195NyVl4Dfo3JfcOCIBlHTP5uEJs/hhehF4QJ1J8eCzhpVfce0DDSiNHVtQK32APzre
HPScTvFbUUnuXjk0FHMin9el3Jl0COdLG+aYPbmBHdHWAY3LuQEA6jse2ZhwFEiHlWsf3mJJ9r9h
seG/hK3Juss+HGeIHzClVMtDAubhceVIN42POmyn5sOaf1cZ5j/XeACxKhcjjUyAeWygltpXZPIn
AfHNIJra4zKNd5QMmUl7c299sqOdI8NXCzV795lOldtVTAO+aLJRpwPKFBXKdGTywLxc6Hss/dmc
0fsEIog41sGgjVa9yscNzL+ckRWOyRIzlJmShhJ3M0g0XJP1akNatLZJg5xNn8AyPDbyoilWhZ+m
XfxSYCRPfk/9ORcIJVZUBqOAi9BRXLeP20wHiNIzK5OIp/VE6TC1KJjdQu9yF8Hc3TXgmwx6hNSi
Mzv/xtNWI5WEJPUjlulIY7609xCSGxuJF5K9o6ha/ZJSK8ReO35I84bz+newfif7dia5fnZRYmNw
P8emBOXl3C/85iaEq1ugo4e+uur6L5zfqMbLQfS3r6wgrO/sdWoi01eAfTmkVGqtQ4X4ebKx/fXm
wszk1gy5fBjMmCRtrqZd7+aF/+PmYTf6Rwsj5APdl7JmGsnqmwUKErRpmEtmC+DJjFF920sy5N/R
2cXfm/OElsrS3y3V/j4a2Ysro4vjOmSiL6RQCJ4oHawvXgnphBepI9N1OUZg8mQWVzY0LaDoHldx
QjvaIPQ+NkmrZzRrKaZRIBq0obmqGzWHLEU+c4bX5t6YgFFumX2fFX/8irl5WoCiOjpbRCvs7o1I
WegQEJ2X+YpbIIAl8oGgfiRwfZRrOv9MI2WdqIw3TYe9vXj34Lekmi+OGyNB1W9USDfyEMWiOmGz
minLU/7yDOxSB+otHoLc4mIfOxxOIGGOpJTClr4MjHLgfoQhPYFeVv6XjIZ1L5ZlCZlV0lFw+D9j
nehlIZsv0ys2LnR6Ki6AuaX6CBEyD1E71PmzuzF9nn2QL6oLLJli6kXrAIj0X/la1ap90/sFdRyj
+fDRz8iD/vHM9oIKwNgBjfHsMTnfonrttAOv7QyDfMn8ZnI+/lVtMZJ4CA8c/8cgBo2ZCe7fFc52
bPrSaDkKGUXo75thkAI8VNQAdUu5OFD7+VCpCq31mV5s9ZV+JeVqLxNmsm0r1v8w/9Di3bW1wCGx
oEYrAveTX8HNK5K41MRLRijTGKzj0YfO0vU04gMhGWYthMItm5yiUwjbLh/0ot7t97B5e6CLCz9B
l39QQk8+wOXkexAq3HJriNBzNWfjYb3bTi/9pM97FXyUbsbSsznIRm7W9iw753vDkDh9jTJxxre2
DyRBxDTjtGSey1SyZ8Sja1U/w2eCUZp8g/j3nrl2oCrq600YjwiyuqXgg6TRmpJVHFqCFMzt0WP+
sxxrgSzpYEVn5eNYs1w6CET5PyRhMZileCVNSGKkF8EdiWPhzCbFllwqSJVUzPf4hsJmbX0pw0+f
R7oCx1MfLaVxt2ZXjYgses8tUUp/I8k2jLkwrHCSR+/VuCC9ZYFxKQbaLkpNcEacb7gjRJvA3BIc
5wVTguG2ut7k/oEF/tCRqvzpz+3pBEPqOu32aK/jtQcK+lblu/Hy+LvDk6KHja/gwttY0n5fUY2b
MLCw9Ly9ayFZGD8Ts3Hg6tXU7wmQ8pjlgenIIh9GV+Z0VdaRoj3iHxlmk4Z0LuDOImMkFaevVvpu
wukylMDT1St2aNjZ9a+oB46nWKIx+gAQ6VWMREr0pxLCQYbwpPnktSxU8O/VxODklIBS/DFwsHlS
1BbH/vGB6R/iNkcCY1N/ps0NKuEyEmle5hC3OqAcXIlPE43Ut7wyYdaMfQfdz1fowfUkybOTc+tC
oqyu1F1ftShjeJIr2IIQdwQ6967OzWUp+DxJMN4sUqWystVYCC18uvyjDb3iKIHnGJrMJ6xI5Gl2
3wh8+sDhDAywekcbzdnqYCQXwhacRXU4Ghot5Axv/2iKt/3BasPvVBcOkjz9LmgIGHqMO5NvBtJO
aBPmXVfmRx/qkHA4CG2m4H2XRnT4R6Gu/k/lqv7W27cK1rEbvD5SFdDt8sztzJQXgpWKMqetlRcM
I+cH8kQcr/0GMuJ/DB7wuggVSDVFUh5eiHJFQiTLsYwpg1HaGKDq3mprjY1Fa/XI9Us02AbIvzG6
8QKs/YzBQa5GDS1/A2vQiQp6yOzF/6mSD45kC6+JA2Tv0gBmX2xrNKPshGGYVVTpfH9GGXPIEbRf
/txCpF3WHjNexm4pRwkXs7Fa+NPX8TDnOjjx7rZ9BVyiN1q9vVcF7hSC9e42SZ/jsRXMkDScMcc8
/l+MoVuGGYFt7HjUOvgtvmHOZMgorgILKUp4pqiPuISBVGqiuCKW/56o2Q7ct2pp2y0ecv/NrBC6
IP/tcjMGEMHIuxrqy4bUZi/TNKxmslNTjq7TuRh+3WLaNcIqTAx+ysQRj0YMFe40WC0nHgDn0BEr
CXK3NSraCMkamSLxl7LQE+yoryQMz+nG9in0LlzpKBXhYM6XbwSVrqnJRMUxVEo+3IBlD+eM0iaV
QM2pdXPbfLar/WUY21CB8qvbqBjgUkCUNx0tstWEHtD/cRHJFAQeQTUIZ/2OF4Leu01DXQw+8N9C
RtBo4Ee4uhCrrtj21K4uNnSIuygCSek7n4zE+EuQMLUjWPMJtsvmTAuPxeyJhWlgx6cAXxV5hRkc
rZSmJWfg+gtQcKbz75ZRKTKCLx5p+j4sbunAZ04fe5I6wNigQrlCJR+ijkidZtRFaxbaloWTnH7r
nEW6EBFB1EXMXsXjLZaoRCPq1NQXJpErK+4gWaVS7Ja7Hys4pMeH3E33P0zux7wYUWlOCJvkI4Th
YNWQ9uL/tX30LCSB09EhqZRJDdHZ4V+L97JNO6Bo3nlSeTMBGL1RkXz8qI3hlRVnVG011nGuCT2z
s8zjubexhsAcY+Ls+lNfiyD+8oTbzOKTvmnpowc7Wo37+Jnmke3cX8Ik6Id1q1yDKUCxiJlHfm/e
RarLtgNmfal1dMPfX5U5mXuTxvNVSGLObbXyxCVcQqj02KPfc0cCq9g08/sfkN0fbFgphFvs1cen
aXEbNpCG+l5XSv7NNF/jfbn1FC0BkVNNo1ytZOGCQFiBqwoB9s/CzEPtDeXEFiMHo0FpnOeeQuQY
9GcV+AvbR4Dji0qILkpytzRULl8tPWdiud8qEMp6Tq9FS03QtHSi1YNCvxyqg7NLiBQXAgybcO9w
pvhdz16MViiegiTSNRedGREId4FXToXajMkbHoz33ClKcsNVdqJMI/Bp8i+W75UelF3Iatdp32ba
I6f6eMVONI/71DNXWB+Y41eL/IJKa4UwNiQh8vhwpBdX81HvOD9bwHdPuJXPa0USoGzXO/1JNJ7V
ulhgdDMrcKBYvDkidA0qJVhRTxbg572tJI6dX7YxrOF9TQFKBw9RYOTULO8/ikjhjtX4Hm8Vti2/
jbtRsSALM1hmmdGVnRf8Itu4E98SyzQaB80U1trhACAtXTm61bxMiToe0ADH0RNASVKHZ6WASY3/
NP4jTBxdFYL9ja2a3Gjb2liIy5Don01S2jJ1POthJwml5hj5gZA+Y7hLZhOdaoeQ/d9rEeNxIjsb
rzm6bbg1nIraYsMSqlbU+d4FfFz6FHrEwsf9N+5I3JzeN1Xos/mRCmCJHtR3zroBFMjeD9WD+gHV
2cXjsYzUu5+kjtrTRqiT/u3bF/6hKGwaFYaEjBF+nZr80K3n47jwa6KxcZwzA666AZ0wl1KfeNIV
DcK717Ntx5skpVJouzOableHA7D75AuLDo8LyifSiU7QxxVxvXFqqnmTgEHFWlktO38gCUZX321M
l4hRuN/288uNUqnZAk4umplbvIka1lkNy8PM5K6eJV5l8ahvaSUtpNx+gkSR6NyuhqrprdVv645a
xku+mD7on/mXyxbRZXOgYtZwaZqHooK4romZ886m2Tpq+s1MpyzYMXYMd3U+/qHp3JV9GtNKWlV+
e4qfdFissuhgFO+MUwYczdb84yWat9iol8cX7hjbTnvZCmfcgUlc7dVIH3UCtNWOnZKHf0pO9yN8
UxK6VK4UIfiP2dIOYr9pVGmQ8OqP4ZABD4mDljg5gFGZM3rTioPAbOXUjhZBzfD2c+3XCoUkjlT7
CfkBliKlECPxdZ4rc50wHWuRqhj33me0ad9Lkn99gNu3gHQynGEBp8kXmWUVZUUIaOzuqq1PyCk+
UeeBAzkdLGcJAjv6akAyXy8m2fjrJp6NMZwQ7CkOcXRjIvL7MsZJvuHSvhgg1mVqPJpd6LZ/Baaz
hByTMTXIlVsu5XNyIGIHDxWZRu2VHuf7smF4ehDUSg01L667UZMVoga70MWMh+ph765ajkCWHMAy
nM9anxHJjUWpnIpor16U/HUlct+HP65KRIvN1dzd7gaZLLJUDqbxvDppuMcDO+ce+QTqzIezjwHw
SvIt+01yAoCfYYn6S9TsmkRH8B5OK412e7E6nyfxCvKU0CATGoCtBaobSvcHIeXp1NKZdXG6VcQ/
jvXKTFEWCQb/AGed9fbcjNpEWY5jUZZhDKmivFXXH51qhRUU0064kpfBX9RsKwvhlYL4i1ugD7wH
ct2/FwVSlLgo/RS8ChYVcsXMh8+8KsGtYRx/Mca/jIIuiPwLbzoa5T1thCWMrqQADywMxWm3nlfa
4NVsf/kJz5op3Bp95rT/7vvhrnoOxZiTz/v02MX71iDTYnF9yhnAPfkAoxC46+0kmjnYiuXCe8LM
tVHvXGbyiTXy+0llzZnjTrZfak2ZYipz4xhDy7EwbYW8ro8MghSoB/M9oPHz1ZSp+SR9jsdiPHed
odft8mFiRRHMSe7q7hP2sVPJVwsUmlAuDIOWx8+GA5P1xOAnx9MgiLCydYqHEqVK7I5RVB+mvYng
dAT9N8NkmIb7lF10U4lYz+/vi782usVwGof2kqOO5l5Y9XX/ezuHb7Jec5ZL08PjnViYahYYA6q1
h/2sEvkskir9OEPmPSM7WwrQukzKWfnVMa8dJUmQAINg2Wu+06eCgUfYjUpaBNzaRDZ1xVwwFnnL
LxNvT03NLJJdilUZfaNeOrljTm6DRzseFN01M+6d0sXawySjSLd56amo+hoct7HnEUr9L4j0S6/M
mkhOyFFR0kGgAYpRPRgTqDAmyscae0zp36hnjuy6pw/WHM1KqWgYngcr9ZSM3S4r6GQ3g2GxwgQc
aNiMNZT4spWRdoBQ/hXME0QWLEEhsA69Sga6XrATExSopdG1ynTy12k0p3D08CWEhXvedaFHbu5u
h1dtZRou2O1m2cVBuOKUrfSyv6Jg2AoOenrNHRCDelC9FEM1mdro+dZOE3KN0bi+biDaDNHcbBAK
Xwon1OMTMOv4rCDhG0bIm6piq/RPv03467ereL5h1hsqed+yDoIu7ma0dTDXDHxYzYVdmdVnB4p5
dhNdaC3KU75YcxdFs5AwCiFbvdhxWVeJzxrhO51v1Q7Z7LWQPktYP2ATnH8S9Ra3hDl41hLeUySz
rZVrcJ5/CyFJEmtlo+pVZ1hkKTmJbzcWBf5rTVoPBxelwY3+6Awsq4aA16fHGx2iUV4lOhQ4qX7K
9eEZzGxl9PKuj/oZP38+SnqGhigPrN0uGfmomgyA58EVj6pclXDYrrvCPl6kmjXqQM9Ry3v4v4Dv
1uRdUNCNkDreXsUAj9TyNPOH4q/3LYtn0dbcywxG0np6HhVBH16YCDzt5y8OTR2ZIDnf1o9j0Kig
uYk3rjoVhOCX+nbXNOyzZkdMNONyAYsYpP+PGQMlcyP8a/2RXVtY5edtRjMGNjxcGxhDZ8Ysuz1m
cEr91vMRBVDGcyS7XfueSZv0RI9wz5esOOPxla+kkbRGzxJZqAcjFDTbeoi1mB6MT+oKX7gkaI4w
N88L1IGSupKeTVRHWzd40tU7GIocNmFVtljgBMMePzcuWjkgsL3+T7oCykumY2Akynm22/vEzfMd
e6Bc4d+bo/hM7g1sntMjqE/64eV0WoHSErVUaKBbNyX7L+23Tk2UpymLnxEnwmD8sNhZ/N6re9YP
MKEpWXp3Hn8YFKZ2vLKz6A6FcbbVz3yCZO1InQurSFa0r/MtM0T3K1iSg1RDR5nmnl5JiZ9irKFF
QSbaAEVPCEaHMkvbIyH6Ha3GWCEvi6OStAnUn4rMXXVoE4tynddFk+VagshrxiAX8FznirJvKqc+
0Axh7KuIBdK6QXbmlL7E9UjpcwWVHkkhkbRaIPabz7FHlLoLQOKSpy6aSDcoIG7Uxm6+WjIesqig
qyhXyjzCM6TWITLCVNhqr078YQ7vPvgUFoWPRtWa34L23Hhk84w+z2Vwe/kmRddlvVaWqD+nrinM
UV2B3kDgGQnzJxbN4Vno4J0rifOVDsJB/fuzzufLW8cKkPjd2Ax6c2dCHZaC32/5Cnk8FEKs05sp
hyzOusHIAzW3QXbhVcdpQE2bfGoQXbCWWOYro/J4fr5UoMm3ocz/gkwGiHgsdRpbTRY9vDp76ujC
HRpL37PPLTcYBJPAiKo/fBrqI8RGQaGBqki1ok7f/3CnmKkpdPXSSaBBBVd4DNGt9pF5PkCNoBDJ
O2dsz0YfdIEQquwLQaEG3Oiz5ubGlIrDiSrZ2u6A5ZBFmh7arfKnMV4leU7dToz2hmB9FKitO8Ll
Wve44G14CnLtP3DaPodLnaeF4EDNOx+1SyxPLfPfDDzuDCTOtPHbSkcDVZgjUHf5I02N0d4XQYyq
ntqAlUuBx1qIG35JS2+Y6vdhQYR4i2v6ESTUtShG/zNz8JLI9blmRa81ACDIkezJHK2/P8H2bDtM
JTe+e52AhTBSz07OeEZsIoK7PaawW8y0WMbbStp9yMusDzyuFfh4XLdR+JMslt3Kjzd+/jAWYem+
7lRTkIJ8E/ZMRF1I66/OhxZKOfUHEJUI7J5qZQAJkOLej/3fXgAW7d9qND6HaZU+VPjFtZgoCpzo
byt5rvst7krUTSTpBP/oc1MNY3QAeXXEPKLJPN8MkAlRZWuUTxRZd8d/b1GFt+sMC23nK/ViP3+W
EA1r6aHqcslM2t69G36OeuPm79lAFNNCsZwZUfRsj0ULbXhdZknQHhqgJzeH4SdKhkgiUAh+OBWv
5/ILL8dV05ax5aXjAfCuaRm40cHdHQ0AYx/0c/Y+Wpil5cdFGeehLYasgBsKe0yfX4RrOrCb1J1s
WW2wzFurZWLscre+i/1GstESZ9AJ+rm36MInSRH7h7+0+Fhozav9C9CZB9f1beq9F0i2c0pILr9D
XkestgF4OoOR1P0manh6caWwfJ9/HZtgEEmrWDfioBskKD0BN3vGhNU/381PkRZ3uVcphRyN2s5H
VZjgbpapaXW+hIFj4uO0i+HjjNXxhe2NfJrcTLs85UYnXWpsH0jqH/JmUgvr5C1HgettBbLv9yvW
zWg+4dzZzO7Vhz2K9BwisV7PcN7u4hSKUQ20PyKJY2YnSWJ/wkGGpnnnPI6114HOKZcSUmOioo83
V7hEWnUOczbEycue1z5a/pnOGhTO9Ya7vzgNfttoIQuYQa3TJNpA5z7FUpvzHMlwP5B0tlAn+wIq
NVvpjvwYDDk85Bb2cl1l1CnPRKZwWn6rzCUR1swBwUe7ucrx/wzZqPbrcjPapT+mBoxpzkUzHA6e
fXEEQBd6sN7+Ci3e4KHWQgBRbQqovJSiGTF+4F8ykNsAWN4TuKueIHpEngdsdUI0Cs11nCUPTYie
qW0ebgAw4Agen7avVe4Nm0YKEtbalCeFrmjNHvhuaTFxUhixsDHT7XY8htKMeXp8mxbBwsSsPGrO
KA9HwdJqR9fzRY6JloIm4hetF0K29kuKpCcYlwODyLo2DTaoVejWF8uhMtWj4Pk2wKVRgLpk79SF
KLdw+7gL6g1BQB3yXoowQuyqvCHTupQcjoBZT0Z88vm0wEH4+t+E+3fav57+S6jlRMGjwFt0m/bI
9gttbj1BUMHv2iiXfGLKXCafFR/ipRVh6JluRPBYtQT6LB5vWA3ApndrjutBB+I/eg8Oji9YD8U/
JyEYjwzfrzu8J36cJQSMt8VApCE6iQYK+r54jxdy4WbgXkKs6ig7OaforNRLvJywiockjpaBbNTT
Q4cNoiJtZVL1J7S5PiVRpXdbpg4xOtzHImPALgrzMO0o/ZV9yLbIsywfHP75LwrxOzSlSnxDgQsR
jL3fpora5gWGTQfbX2WQDkQ8KJD7DDEDrPXRRlevPT88TU5kkQnhNlbhF2ZJczRop9Bl1+6lH6XA
Bbabv7reNHpo+Q/o7BL5q/8Z0/NBZuLBEX3awcb6bPPnA/46g6ZTWFDj2eU1iBJDQbE09mC6GCqF
VdQCGuVbdDU39JEb1ksB5K692eI5nHmFvQBylKGNKsGLJ/iidhTSmSoiBm36WSXmBGQCviq+0JuU
VpKkivrA0aflOlN6vKhSDtgOoe8yRHn4tYM0KfHmAwH52GysdTLKftOlyT62RkAh6PGvJQxbEpn9
AEspFh/ulP92a4jWvOgBzhOuPJPyfgFzngscyGW9Qr40UPs/lgYzM3DPGqR5PdRs8n5cPI0ljkrQ
vcbDfuDLGcRp+SwVM6bEH1Bef6Z3BVB3TIAnZc/H5QD56sUDqTuYLrNIyy2+sCjbF/VJqgv759o4
wkUZGvrc/C8SYN0sA0r0lIlR7WzOVqLPSLBeetwOK1WFYitQQ9IRAp6YpAdFgRr9NU01J2v9Whoa
fFkF6PqUhO4y52DNbKxAoesdg038BIsVgKZn4KMbOrSa3OVBchzgjqOVuJbMdckNrS1noilo/ZVY
GhF1mpLpQ4038L2y78GNyZb3a31cDd+BHB4OZfsr0GXx5gELN9JTSx90kjyjnBM/XzgaC0zWH0xs
xv6BQPK0T9BknlyjaMzXG4U0r03Cp1a0Vwofo1VvhEzIN5aJd9swso1b+wRrIIPTiKXWBXD/p275
jDQRPbIbE3VapQZ55hlB+eLr8fD5OM43qG5DRqQs5uCFmP/QbQMVejk39KofDdV8S1nDWVb2K3eS
gDCvVvqIL55rb/p00QHaj0aCAeDcq3HQEgKMHxwJxKsce7tKCMcJOA2vHKghH861MYgGsg0dqJ7P
Yi9efCvErQPYSkHU7nMotUruWTACWngYF+nv8noZ0ezSMHc3HDQ1lcfpzgwq5vQW/U0mXd+rkR3w
xe6zXaKNFoQiz8YbM6mFQN5Vp8uC1+pcdGsrivN5AawmoO/6OVnIAqw7n0xekvFY1acSAP6bZhFz
0Z+0TRLVdmSBUVFiPGCDb9WXD9oBSrxOv59UMVrSq9I2nDQL9zSZi4CIateNevgE58LCS0mBWSiT
nmfBTotXtdbOEv6KKVqdHCwa4zB17+MLhl7yJGFQa3e+cWz3IeGzneG2ladCzZ3KArLoTpNtmG1N
twsP97Bo0dOf+wwQzdbAPz+zlA8f7kw2kbWfdbF0OqKPc3p7W7cTKcDx0I4RdyLC6yjYYNvrmOZZ
vY8393kDxB+fkEe3zKq7Duuic11AnvIIYcQF4eRLzUgyTKQm2RT80WJLgUhrhKkxgdjt9c2HmuLd
GL6h0M5sXpFV2Hx8BW67/bjJko0xJYYBedvgGysvzgz+Tmih/974Ggkjf7fEVFM8V61tHr3qrAyj
lVXmAs5VfLcG9Nu+oARumrA36woBUDsd2RV+i8PA93D9YSC3raNhAwZQ6ZyhvybzlSjnbOFZ2H/w
wCpYnHjVluFvOFuzzL3JO08zn2eznTQ+ijqn0MUyar037NgrMLFOG/j0tnT5QhqIwKr3oMciXpgk
oYLPLBoq2LNumcluFoy3iV9wUKewgz8ftiqyu5sj21qPLeX5z8w3lbWVEctTYMC7SkoSkzlmcW26
wktrzXNjAlvKcsd7tGoFd2SK3taXW0juOw2mYldLXZB08AbuAsx2XxgWI403KeaMfh6XPxuN4yjZ
XLmEiIvNGkfZPrXrsS91eBHl2O0Oj8CELwfpkBHTc8mkmKb+65GkI6MjcxPLKrDFbv7ht5QuTYb+
FWqsYVto8SK+ahDeA9WQ4zgSVnwTV4/xLdjBcwtEVE/awMaJr4cXhlhLo2FvbJOSx3qPuK7XK/VY
+DQqFDOMv6R+LUVBCvhEZJ4O9mzI2N/6u4aTcjOLFOPVL6AsEDk/7zBDVzz1XemDpu64+mDHd/f6
hDrypJimnVUruPRaVHo1yCqyqBPJpX/lbIdp2gjv7DgqNLdRBYdXKRgk6N9GE8Rq8NhaY1B/kepc
aq4sPSAo7zsSHMx0BERz+7nmlE65xqSbEzy04QMSaggpLPi6KMAXjW9amdgUwTzqy7b/zqWFv3QK
TydZ/Vfrj4xJlb2EVUCkLX7qkfiXQ5PbKVTmORADfsWXdTVbSkNPjrEDfHP/XqPp3scuhyghaDYP
+rKJ4N9KgAKsAvKKqZ4BV58xc/nXGOlu4hSy/9ckOCOlp7Q7Jh4DqBSH98KZeMzrJcILgHCBGk1g
V3JPmScBBxluJqRL+/FeNBf03JMu8GET9az5F7w470+e+SHDt5AJ3Gwt5r3xWKrLwFVZWuFG0VOg
GrPResAJW/N7i7wFi4nbBDMzDjjC0Qbob5ElKAn5zYFG10ukyO34WkznKOKEbT3QB0U8mgAuqNpw
fWcP9nO6p0sps9DIvfV0GDkiqlJK5RGPRaFx5NLzb6bzeWTW6nvGGoJdd20DFuikSKTQii7P3VFK
THm1EX7RWLbAQuAKui6b8xd57MXTX2+Kd42knOaFjI+TgKERGlAjtFmQNWtIDjXSZbL4sXK5XTyr
2ovbiK3f5w0sJdTWOXbdRsGxsIC+xeS4nayyCrq79rGyJaQKrgN1wSIII5FBsT8QxCPY8LpuDpBS
MYh1v2hr98JK/Z3+eWNy7+fhrPFZeJyLlJU+S+Ly8v4uWbhUsd5FgP7UaCLRjmM4sh12Tl2Kj7Qe
BGeE/J1tOFfBzEIBiSXyJx6tlsSDMJ34S5146z+vP02SsTOK1rNXld6e+rZeMxVpwlqrZy3TC8+c
p9DQhSzuDdZph1+uLnFeVlZOt7PVSIw5lzgWLjSIWJQoTgl/sgfPwO7XZv0hS55mVMjTeIE6cI1L
pFOT0saqm4ML9JgrV7DI/DQF6QJfflJ4WflxkBcSraaVmI31bVgEtuXXJS8o/YPUkyCrjR3j2oAN
WYuS7uoEfRN2lZTFDEMVguTZ6yztxdcTA4GW9ArZkPmXtyW0/wAE0dylCUsTL5yQ2wAb9qECKgY/
0n0PJlOzsNrMV8A3rxYzwGRccNx3QUWTOFZolFIn5XUu2hjEA3eSdoxLZKRt5R5vEupz9zYe+Enb
OyqC1i9QTtqZYFuC57xflMkBHf0a5ImYnwCUwRiJvaNE5TvaQrP37UHJMHfmV5yByRA+xfaybqmz
APNGgKk2OvdPHkrGFYjFN0xlPqqvbmQJAVGFKa4tHrsEzFEOJVE+DXHRxAOdQO9ETuUZJft/sF6Z
qggpSQIiitRVG1yEpvOCy1LDy18t57sYnE+38okM3zx5K0mqvNoiOPmJrbwZ5cUXQMpvmeommrlg
eRaW/SKOqsHjMPUyy8isjMyRQ20uKFx1Bnfbwt/DlHbmXJ8IQtZdyp/sxaOoeT+zk1s/O2caCcf7
0ml13K4J+KnETDoywihvFPhG9FLrnOrLfonhzU3a5V0ajT8UDx4dd7mH9B2FepKTcw4ju5w+pgUE
w9vpdVa4mgz1PKSvZB4lGS+GxKwZPvsO+onvWviKyTm2eH7+c0E+gqvXzRmZFuPUp3ew3SdHZMbk
C7VC2bzAuK3IiXM/nVRi234IzZC/7mwNTVxSWaRrx+LpfFM75DC9KoP5mrsZ1UMUIIn97/kvNjQ7
1PPRCYQwD9WKk2b1+c2BPLhexQbqV9u3GmE1fsUpn1ATqtIPY1Vv9GWiUeCB/93+znkSdZ14SJzM
OC2fdrujDpp3EXNpB+lDx+idyLDLefSZ99z5QLMIWyixp6E/v0GfPCaLaEFlgJgCH/aEqI3XHF28
gmsdWKnrCHwk3H5cgQ21fre/qSS2TKTTjSOCxozJsJMdR3zG1iaEq4276rpvgCGCv8jcQz/KxWzC
nMCWsu1qbUHYU8j/aYOoVA6Vh3Eu5WXZRWinaewwskHPpK2IM5V/Hkc0es3Ld8sphQAXokgfgtT2
QUteHOF5IjiAO/BS7x5h+Ti0XZoaTS/zWTj8IrQBQV8wfFONW/X/bJmEk473ucMCav7AAbny4nRY
ZLi3VATbMUZOjgwODY0cW/vZxeFv3HFNjn6POp9hjxOA5W8RYcRSNqOP9xkusBno/hgMwkcGDO6B
sxH9IT45+rntUei1qgKxluzxBt23CXgvt27RTqsLovWxcdpE4IcuaHA1sSz1GsGJhAm1FzXYvDDW
2JORoKULFDnNcWJ1LUntteATVg75V49f4cvleXhTPyIZzdnAOuTP+9giDUReduzw8Bdmzp20FrnN
tb5du8HYj2+czq72L2lQW34Gi0iMkismF9/ityOIu9hSMXl55RAyAO4QOhSMUt4jQkybnw3XAgLO
oTDU0YtLJ4wGgNOImNIzRc/17xIP0bG5FyBLLmQLNC4iMU18afvATMvXrKQawMhvfoRIv+3NYkBQ
No2INld12dr2dJgUcEm5heybvsZxsATrK4cqKa79t258WiqfbTCkBur13gLadFfj0kWes4j/ieEV
Kg+5BrWP33QxHcwr9rdgL+PkbK/0IMtNd5K+MSimmdPX87gpbfRtrAOf9QATGS9PZ1+fpBjmzHwv
hH5Th+w1nzQEs2j+HjKdK/J/yZCL8YUsLtVlGct+8jtblk9tdpmgFG4DKm7ThihNAsdANpd5I9zz
D3adYde9cvRd1itXE0mwvLIQEP+3QO87siZwiv2gVDiY2WXWKbjGqLgKHCUbUk9NIxJL6BgJD1py
8563O0gNybKyuGd8/MA2lbw+26LcdPPHz4aoJjZt6fDXwH7JuIWJ+NfkjGKZMzhAfRpZsJgP02Oh
Chg/KCnUSXODclGJhUZB7Zs08D8kug1xSctDmK6fmaq4jy0oEkW/ObK1W73GLslM1K657f8z4MXs
KQQcRLVTcXCsydS3sD0pBMUAnDUgvVqfXI45Xi90oDK1DMAnmcUQnZwpkMTNpsfmtTOt69gTkF4H
exep80zQMe9E89WGux27PBq7cqKkGObmRulQFzTs7WZDsKjCNYo2B8ObzErMaAD+/gT8Xr5twQVC
XraYUyXnAsiaoFFt8/T5ksRBjO0P11J8y+fqHb1gQ79SilpeV3K7iVDdYVDn3vVtzdkZ++MJPFnL
NY+MLyEq+C0GPBmkf6DuwKhG1nDyqLvxz0spJ/tyKpG5f/aXsdPTHXP4Jp+mJyrtgX+K4PnlQVON
HmJjtKwrU/Rfm6dPhE3ryu66mcLDp0UFzC5Emhf3A3ukHWsDKCGZSNgRFgikifqtQ4AQOkeHExAB
TThTlhRakV0/UyFq79eqZaeAYmFY5Oq6tZYNyGOiB8DiHH+Vec+f7wd/O6lJIyxxWfZ+JJLv4iLh
tfXJ0nM4ibm9jLnSucI2KWlEFRhrvBBadL+LwtvT+0nu8m/MI4jrRctbxXuJOWBvMZHL+XO05JSW
/1P/8Ckp5a2JigihEeUFGcZBgPTzrYN3P3FWtGsJOQbo+K/k4G5Gj039Ph5RdC6YC0Jjmk/1jTwl
ibLBZpJdWT1s2nAlkM9kgWKNbVdwY1W2JQEa1+m1KCG7meUyWQu2jUKFSSj+HF+VF8NamTm0XVT7
bZf5gNv01u8GWYX04W5I6TeRshMVHzTjYqti4rbpUajdLuTGWr4h4Xa59JLyZU3IeE+yH2ou78QE
XFlMUsCMXS71PnYtJSxP8PY=
`pragma protect end_protected
