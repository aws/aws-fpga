`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
jGbs86dhR5KLiaI7GiptLiIURpVI3WIsx3//e4aTJfl7imiG5ElT863FdswOLsZgVz4/ML6l9pPQ
H+8Pnx7yKSePu+Vn+4wvhUl41MXeNebeaYJltA4VoaQis02OI3c3BzUI8YPT/nTcpd7a5XssEL4a
fjhBaZuMk0gnvV6aPPtR9CPHjYUAUlKIpyqMGdXi33bHv+Py6BZ24GakeiGfyKuIUrh9XgfaHIEg
Dil/gF0J8b6H9WPN1pj0JxYo+RkXWed1hhGJ6OLdbZSpLMMyQR1u9d+apwl+DFIdGPE0lc1I+wOM
y0Q+0oQQqsiwhTjz8f+fJM6ETtx8KnMVdcZaIw==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
ficMnnwN6ihlHYkat9z4MEVDLSS5mJ8A81PALop4kwxUEMvZINdzxHfdSOWnFOywkkgESftlix0Z
toznBYxBQVMaGsn5/09NhaPa7WyC/+aEeP/wRTAOAEfSRn7egToioDoB/gQTDuTC0Sbw2eggA4qz
9khERpOBCk1/fQQNk58=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
SdVRLg+xBmEkxzbBuDgrnNrKuQpZAZHzS1xIu4yr6vgWjeJ32IwZd4tqSbVsNjrrG/0fDjW7TgVr
xV8xnOX6P+WtmGnAx/kr7Pxc/egHIjAZB8CrK1Q/0ForOX5GuMWdXFTK23UO3Fz6IwWfJLUpIBf2
LyOdydrtFp5mI1oktpw=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3056)
`pragma protect data_block
sKLmjHG3AkdH2+GiFYGCD6XqNK0Khwd6C4WGdeBqdLuKhMIKOs17Fs+gjMeAxczYKhZvjAN2WuYs
v12vXmHlzJmZkp2mRU9UlKkNAU5SQ2U+5UPcaALTMFAXtl8POJkE4HU0q/L+XDAum4rUjgAfNxvD
L1CySZVPIdLNz7gxluzjc78dF0FT2gU4hmfNpCPVKcgnUALX06Mx9wdmlpPLMl43Hj6wN4CuarMF
xtuo0WHQeLTdOKX1w7TcM8HOePJ5pyfm28OEUE4EwDcWaODYlqd7iD21ljNM5TTjfDCnQ7wbnqDU
u9dPbS96wGkEYx2S6FCsjhexqBYz6j32OZWWbDp4dTNW0tBLJTU37e1baYMw+nYiHzdKTdjABCuE
KYpdy878eWPFbFG1bB/BJP0XCOY2HOOchoDlIy7/DspvK9qrwihVokIIk4i+BpgcuDTzU1NFDW2T
3Fg64bYDhmORVd5TDkcM2GIHdsvHS+xp5YKZAM3cxZLf3QG0rgpqp9eF8pmspksfv4SVAUC7HTfl
YdhWCBTI/V78radzkfVBVAp4c8fOnpjsNKO/gw4t/2co9EyJ0SulsY/yHyYQ8a0D2Ue5zZ4YGvZe
ed2PmMiOPURaw9vTrYDpzi+5YjfxjJifJye8ie0zfkYjtkHU7+uZ3gbv1JixKt0P9eQT9gcrppcs
MsjSyr6MyvDacoUqeKYgNQt+4pO/CKxLlgZIscAKKFXmBxeJoKqU/SVWTU/XnRWvqNoF3nFJmvGJ
AQPjPm+IUO2by2EJ0D/YJ3Sg+oM2bOws2lpvnah5h1Avh+9jv+6ochMNeXKeRuGqZQuGoHAMKlE/
M/PbqhQiM5J5hKGdxJmCtMBOl/88ODcT7KLmyavsIFMfVGHMyvdkHu6c4XtS+NxznpJQHVDS8iX7
Ack2CjP7cChZ/zc+A8VZes/f0AJdFDwJkxuYLFxQVBy2sIxCfS9QzB+wmok7sn5L6XHBKXyOSOCZ
AICAW5ES9pwCuPtZLIE5uuHdYSrOBcml1tNEcY5u92ty9cLrWG8g/E/VbA/Cbb1yifWesFGqYwCW
l8+uh+bC0U4UUV+HLKt85kI+Pg/J6v+QZsCrggvSk/jua+4brEWp+/V613NYfXlxH6xqKTSLOAfK
MsXM7KLVQMLndxp/CC3Dk+T3UlkOIFWSyEQSEvexU0t+bWxuuWPmmgiBQdQ/3mhZbUR0F6IlWM+c
8t5mSCghjKwmxwskVWAzFhAqfSqbRfNkTthAgq6Cgq1EIIEkd7dkuZbleFQpdFKdrDBk5CFfE32a
cOfyvdskYuVfT6RkNpnoiy3K3Fex89XXrS2x66ZFYb9pNAMatKkGdwy/CP38sipUDe/zOQFzFkIq
x31EujHaRl0jgtwRCncO7wR14WXelNPxogGwu+sKX9Y30BeREHZKilxLHoY531G9TUAUQm6kt2/Z
n4d8LuGnIQon3sqGVznKJWmkBgHQ2hZbgWi9gc81vOIzDQIhn/ORoHx+/bjTYrbgTPz5/HSbajdw
8FB12lKRbU3W9Gesg/a6tOGqiBlYfA1P/n1mw501QaTgczg0K0BKNl7IamZJnTV2Z9GlZ65ONiVQ
QT2ePRzDciqWf4WBAfiXbggmulMYLgi7404QX1cqawpq1GJMH87D6xcsoCBRVt03u0gGzufqBN8p
SIzo9hiyxVcEcziJdmLiXWJZj5lH9Vg016KHOdcJVrYimsSaB9WhSzmiTnhjp549Ds/KfR0j1lM+
jcmK3fnNa00wixo6TAQYG1V9aYwtiM9fHXICQ97lM35kGQc/i+/3AgBBgnuEo/0rvR0jbVpp6NQk
xDOvMIhikP5cxL6AEnz+aBTrf4SSrd/x6xhKXqPqxTcZ4M6WDC7uloBpjnYvW0oJ0gSJFWPth4G1
raDO5iop051H34FVTi1EZqPNR35L3imslnt4z6wmGozUopPN+uI2sF20yuSzdxmpRT4cvrVh/M1m
NPwTIH4N+xJGvWPf39MRdxZuRWcbH4A1u9XDJmJyK3RZ52Qe3lGeoB/UuOtfWOnCmK69LYI6/hZk
bbH1PyN+Ja3bIpyta15GexYvBbNJuHMsx/7/Ds5qein5ynuiCVOHqjlwdxgAr9311Um3m+Lkqez5
7x6kpMm8YUJ7H8Yatz3gY7xtPSRxst+jdBk1xLbaZB3lM/e7NAHUdut84/Ory9ZepD+0ccvh1VuX
Y56BPzqlNDTM46KDSEASm4mlfFNADvcG1F93Cc+AwP6Gtz1RcGIOrzzjILgpVo6Y+iI5poQGRMGp
hgeETLiiQ/ds7mW1K46+pruDjbzL09g1d1vwzw39HBiloP7nYG0j6hB3PfntwyJ57VZuNa2xbmNv
vUhdZFsFN+TBN75Uf8W2JctdPsY/xhZ2YDgpFD3DsKtZncyTrZ1L+tnnEFOruHe/iuuiKlrZvJN4
uL9UwpLz8+he23JJAaIciH8qHKy6AJhqrLHIulB0TrIImr/32V3/r5XVmSZ3QLC3fK8qkNsYGIGZ
K95wtaEAQUfriVuSxCfJMnLhFigDEen4OGcHdacp2Co2R6IjpABu/ceLQA72eYQejrCoCrKA6AB5
ZWE8MVK7Gjp91dWcfaoZYDfbp8rXXRehuncZldxYl17YXrzNuz74NPquZo65OrtUNY2orfJVDyC1
sgFiiEw5VMGDdXs7Adm0eJtSFJ/9KUpfQFklz//zkZfF0U3jvkhWNr8GDASLgy3HXaIgAZl1EVOS
rcRVQ8w5LuJ8Ecka3yQQTeVSgUhrsd82Za4QsNP3IB4zkfx8SEH2C7zhq7yrefXEtGszDT6K9+t7
Q6KI542ohTqer92iqR1glS1BQaIjkjXaDDYmKBbyEVVvoKgqAeg1ZOo66LPoJZmHqBsax34SZQMY
l/ojb4f+Goa49vZF70qFqSO2FbTlF6fD1TNm1O8Ub51GhJgAcHS0v23f2spoysNf3YYHYopOXHFv
EeOYMo8gmwdOByjIhN6zMPx47I0LLzySaRDwDj0w9e1mlpAXC6AvkerPSWNTQ0I3/E2KmPY3RDYL
ZkFks3aaa1Ve75gAfPgyGTgUC9H+gAnRvDuHx97Oeq3NN00hFnxogqNCteWqVfLR6WCcjKQI32bl
Otz0zWhNqUEhsCLuGVhj/pJx+PfOWuQdlRmJZfLB/EywE9G+Z15ajQYXUolWS9huvmN33r1UJMnR
UBNO1CHw0BjKDUXz23URrB6rwjGQ4Ql+iXvRg19ef0r8Ks8FtGUCT2IF41KiBYAwfiDQw4VTLzPD
nQ/hZwjgT7ui4bcMLxpYgLdT3Vfn5dWN6021mIC3x5SiVSd0RaPTyj5j7hMAAucyU56ggejQyQcg
OkAU72e+RU80dwsjXXhzN0ROJQLQGpeZuWoL89nFQXEQVN20IO/cX2tVmv1bLC6Nkoa1Q0kmYu7T
F1+3ZnrKzOl/HgXBTlEhEoRZhhHdvpWCKIifhBqAZWiwzTFZkpN6ECoOoIrwMt6qZA0G0dGoZZEo
aR2AQoDlF5ivk72pf6CfgSOis+WxAI09KvTUtJbk9ZICUZTS9KcbH7bDSGqtxu52968xHHn80fVT
aXMsfUGkETvNOnHd0pIb3+MjR/t8ispEa1pyAR1tb8NsabkqjvbggkjJ66EYzf0W7MtzDWid0FD6
9WpFY7K1MrzAxQmxFmst47EInXjPbZyOL0JmXUaMcLpF7a2F2yscqvbAvGjXtumC6VCXk2zGRX94
BqOfsabxXXlnNlvXweNPOigroWMokoR0aBRUVKFgYenqExMRZhXgWM4pPJwlX2Zm4tChokbJSqOu
UWHpsiGsDM1mc+VnzEaZXQmYmhzr5+NuwZNwh9Pzvlvbvg2iIa/huWmIr8YPOdH5cCPHHoYFRazs
eIpFN2/k+hJQedG03rv2NKWLiOxhyyXq/itwpLEeW7Nt1pMbIS8hANBXtYnmZNFrxznwVlqhGfzA
smlyiU9xpTCD3mCna9IUKy3o7WhaIkbjPqr/w/EyDo8r7T1b0m8PJw/id4V+tne78uFLm2XjTLAn
BguqWEAjpS2C2irbqB0sLnszEOmFP0rJlBFryZ/zZSbvv0I=
`pragma protect end_protected
