`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2024.1"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2023_11", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
SVkk6URD82soGZT+m6xKtGRFtjAs4ypYIvFDCW5NGCp5XXhZPyV59y955ou9ASUe8qPjNGCIxCtr
mrhpU8WZC64m9Yy3IImOVzA+6tl6yF7l3FPSAmE5y6MLrZnodsd4OGhUcFKMY/0BQAgIxiUHE2Ac
5w9sEeiEh17IrC68Mvp1VsfIq5r95mobsTbxBIM+dFwDVySf4Ar23mJK+kcfiXYa5kxZqn/A1B6T
06UYZH3xJmLEEahjj+6PZzRPVXdsvagZBD02iDHH/0X6Kbei4uuxWnTGp4zXHGiYCnooSHkibItK
zmNmy/i2Hr+LPTJOmZM5CT1g9WcvubJT8TjlZw==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
g/MV9ed799jOraouFB6YlSCfrMw+JOs7MtYh1m9LuWWOWpM3KHPndmuhMMJ2qcRiIGv5rQxSVj8P
0lSsUhf83GG/qWN2DzJXjFutfVtbGiMj3z4zVUbHxbteJPqokJk/6kM27H/V5qgZ4oEc1M9vPFSR
97wb9K6b7Nn0+e0KrEQ=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
BWnqz0tknhalamI98gmYQfscbBPGKpwlCHrW7z+3z41TBzPeb2wV0tFlD5YqmLty4ztgMh3c1s6w
tPMCnoEWSWPWOKyOXFEwYs+N5ajW6/M6pTDJZUMa6PlqTitgAn900tHSC+iZYe21qYqXWeb0Ns+l
LU7NovcHo3/Sr2QOKfY=

`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
mnNdsw1fT10Y0rKThqhnzB24ez8eXYMhvW8Zrh+fs14XRit1IssziNkk/YUNw9DgRToJ4NPhx0sa
b6PTIv9VlQ==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 80784)
`pragma protect data_block
HL6re6oHRl0qa7m433gJlKZ051TduvFai/hQlpBCpLE1NMujxd7btKI3yrjEb/ei9dei13HFKiL+
ahJEF1jONZ010GgR96NLDCsL28n70s1wH1h0LEUh5i7nqumGbPTlT+/6nEEImQUmKKVjzrCdodmw
GePPaY3lF3LyIBYE40vdjk93FPniIufK6kiwVtVupQJBWh2+2Y/mTNiWIL0XAWGM5vOqcPj55LWK
vmyKy89qPsGrvYdS1PgS6CbfmGfO5SY442O6MpgYkTQUZo/knJIfuPJmIP5GYJZyD0cbaPX5Xt21
hWl/jnssNrtREP/D30paH+n4jrpg43nt7PIiuM3+f73Lf/zVWoP89OgM/kGY1YHDFnGzZ6B0bbaw
k+9SOvyGU+rV6lhYuMV3FnyxGfM6eMPjkbDaHVzlCgT6Cy22LBUWv+BwrHJqVoexhOSclWLFKcdC
vvK4wXr4eZRab5KfOUJJn1TedQGdjA9GGQDvgNXLBLn2nlLXGMLDPjhvSOKGhGzptJj2ork6DSGq
GOaHUOUrB8pciWGj66RqMSc0PSbvSIJxosbRGn/Rb99V7Zhn3nOXGRNsCm89rcKNcgzfnLM5wTr6
Jb/lhpYMKMbmSalPsWNURhSGacjx0gFDC9DOeCCoudhsrqJyFz1VJTxH6pn7VX6AxwMtsR/XHpNv
7s3JT2w2rDqDEss9AWDX5YHDs78EG4xvF+9KIdBMKGSPGGj4TxZkh1Qs5+mV3mdTKvXPc92sJ25a
HZt4j9iqF2VhfupZtSkQ1rBRiSE3h/eCVh8/1m966c9P/sec3hPIszq0vpvLjnz5UHaBt18IXrR2
5Gkrog/kuRHFvE58wMgqzcPsbVxftbDg99DNZPULUdm0+gDd8lQvnVHUG6W2waHs8FUl6oqfTARY
mfp6ycHdHM3vU5s5lpUU0S7eTn661HatM8tx8W2nQxfZXRkdmQeoOuR1UZMNjGoxQv7KsM3X1j84
GWSRPdUOVoCnCXgDoXQ186m5qq/JrBxl0olrSKFiWQqY1batKpDB0REv7dYs7JAISFQ7mxb6doxV
1sKFCW7sMbZerJp1mGymtGF3SQuRqtIFJ2KQsZHya3ug5GM2C9ysixzcMCxZYV1GhjcVIVlR1ldc
SHVP68uGUUfWL6iO0EELI3TtGWXJLSo7cNBubO7JCFLWCpLRA6U1QBhE5YPXOG1NAl0YplPsqzK9
HxDgLL+XT25AjT8EQB7sNU5mHH53YrbI+PCZq0uaEzxsnfZldLUETUGeMrezUEpobkbsseKW2hoj
vFRzbQrKMVR6+btRnTN2NQV1iBW8+b4EuS/rQsFOsEanOBVB6xOpTo6iKKhs8UHPdewF5X8R5/s5
xeS8iE00LXRXqXxWQqGyfnEZsTrlgebuFshz/R15cI6m5iJdv21cxAi8wsK1MV0KPIUyORpSHBlx
wIO46nIKZT26gZoUZh2BqAleDxO/Rt14ISRVHCE4MjMcbNXMxbw/fEwZG1h8DjUluSYDbMV77j+2
k/BB6Wp4ZZfe0VKslv8zYSRuL+7rKMwsWJCMNMnwzd71ZAcXtwyqMqHJIHF6CZhAJ+5DNNe9s/5M
jSvu7yNseRXfwaqqLl5R6BKhXc/DrAfrAqjs3GE16xmkMld3LJx5JST13FGBCxVYddgpQOIP8FND
tPes5oT8YNHZXl9HQwpoF9kU9hzJY6v0oaWOEHUSVBn/XpBUhESrm/KuF1V6tibGTj0nOi+UJ7gr
49ptpbkTY+SdgBQUzAlXt4v5acjsucVfK2fS/YxMvfSQlV3kyPE0Z4sNAi3u4FFcVHiU7IGAxZ2t
ABnAgLCvFATomf5E0ntQkQd9Ypye69dM8ilNzc0YRIlMwJDYm2wMsx97uCfvyBHWRA/df0MUuYl6
VpsMI2Rlvy2z2NFZbncplag34Y2++03Gmm92Yq3fGS+WLqadEmXcLh3ndigj2jrwTQrhtFyRi0dF
lGVT1SZrW2pvanqcaEKqeHczQ5uAg7JaEACDhFFIk8vdFMJv7qv9Pn6Lzi7laZ8tBWqb8aZHC+kT
AOc0DE7hKUFYJSMps5cYF18DsbcAM1H1Qfg3H0tcJMsPXHxGcN6+IgMt+RU2NQQWoID/NOuFr3+L
zKXgXGMEDSKZKTRA49i/UntpeMU3sVoFzg1pPCawmZEc1P1kyDooskScXz8aYxMv2aVm5/uEksvI
O4ISHyF3Wu6YsHZb412rAy9PzEIjcaB2v67953nR0qlWUNtNlF2Z86k2v6YYiTVx7Omu1yis14Zo
ySB8b682viFtBEBzemZX2j6vM13F1KuzO7QPAZkwteuZyv1gKyDmC7mh+SzJo/uR2jAENRYnfn0j
qxI3U2DGiLlDeT+rRI+e0s+9y+Vc2E6AN6xhO8X0+GObJ9Xx1Agc6WJN8chNBPmYWlyt49VZUh+e
daO5ZxZyZWsOLZ+c+AKSzcbsa2PLJr0HRS+8cRLS64lnFBhYmaMdQKbv6Jl0ebdo5vNPwrZB62cG
iVFl8A/zv9hQTFHEc/roB4a30LYdFPbYZ6g6yBZXU7b2xwDevfgBJkuqvFf8sNmKPiGaMxeI2uIU
922qgcvXoRu6yA2L2379fNdRzG9hpOhYSC3rHWaWI9VEcdOkrdwqCZfD2R7MzGvC90o5dhZz2c4t
Opeph5lBsqljsf6uUeM35nGlfzLahwwe4bHlYF5Sx0c3CVrpsUgiJqVDEnIrq19j8NrrUaBXxo1A
hZwfhPoTRkQVHwgUT+3hYR6ZxmyzraXjIafxAb73b1ElNxFxC0SYLhR/eqMPVMhjj93G7xXiz86D
pay4SQKe5w00OtnxQkNnNIi0hkT6ecKUaXru7DDQp6H/ehS9ZKR1DDjMuMvLoAbQtn9dN8v8xA0F
mIN6RLeIyaER72ds0wZVMJrdZQxkMqCt2B7IR52h9Vy3NqjuuMsrOrH0pCU5LvJMX7AMrNeglieJ
o5H3Hj0e85SEXaHeaj6HZE8JsIUAFh4OGlG0+QaLYLN99xU4TTf6m4wwZFSZ1Mm7cT7B9AXcC+LM
CMpJT6T2oIFYBpY4Xlu7ik1sq/uzCibAt+QbOg99SrMdzQwFNYPCjY8wWgHLtCFTxxfsDthVEgED
jzHtwo/Y9HfUQPonk92Fbr9TTk/mYhLspSpgGJ2FucfdJ7cSAzVoMmg5guuugOGoBV2r+9XWorRW
DHzVWEPywPodw+bmNMVVd1JpV0vnWpWd1JUSi7DzydI6DpRYEtClZsRdZ4ZmmXoCQ9cUvXW3R7Bv
zLnkUpoixqX7/C4xcD42iDmCd3kp80IYyfG5L7FHYwpO4Okha/rE4HonpnZnda7jPKrdDA1nqp+F
4PJpAPmMm7eQumN7jYs1yZq3TajgN0tl0R5I4IKxZCRFc9StHOWR1fheCOeBP+9HA3tNowdK2Zn4
WDK4onV8ZaRDdnXipCGZpw+cn4DYfTuDb5fsfI//iR63tGc/TF2CYNKggDlgiMH8/nRSOaTynhHo
IKIi5ETwVNTVFEHFeymIed6Mj1brUfgpizZ2srU0Nu1cV2Hli/HSn62emPiMwXPOuggaz6Ssv6We
Y2MDvlzqILJrWdsvC1MApQaG2YG+eAP4s4WiSMuOL4truyQQOYpFdiG/acW06tTRPkQKos6HWu//
7fI5d1zGOjN1/LOvXUVPoLEFuiB4zTWfSMOzFtn22fGcc4LeN3nSfu0bctATRfll7Qt5FiqdDkJw
Y1mPg6Bn59SkI+pqY9tZJ9a4sjuOwtmwwChAc+/29bfpYNb8VhaMaHU9fnKJnu4+HjKyrm2fbJDU
in2xMsTGxA/AXNZoHLPXapUs1L5NVDy7KZxaPAvs7cugTupGCFGCgDVGQjEXX/L7A60ANrE7jDCk
O0rn1u/qqGGvpWryIgxgsSE0SDNcQ2ZqMHu1OzrQLGO3PMLjwfTvW2H+ZEoey+Exb4HpXtBMneAF
8Zz+QZ1UixP6Tkpvo3JpnIVTPbPSUbjh2hR7Wp4OI2Ev5kZPFU7wsgNXd1T/O7En/onkE5yjNGoh
2PZ8WQjLM9woqwlErZSrY1uxLtgTDcic7GakgGDW0DlSvgKioKYjZxhzLhp22r5ofUrDM2UZqPKR
cz2TqJI2qIZwbcDLXhIdaIZJTy7PEcLuvc3+GdWEN6PtwwY5+GtHlPnwiJcOY3143hwpCICgsto4
Q5HTOBVCdt0tQOPTGy3q3ibxnt1oinZz7+bm1j4Rz4LeceR3wSqwiGWNMx6tIlvu6TvMQQBsURmd
l6HJb89z7jVfbO43bbrianYT+giubqbn5bF9lXXv/CkDr/SQWsRgBHOz9hOYM6P+1adj5Od25cxW
SgO+CqUCSgJOU3oQ+XLkPTk8hPCSfGHVSYhopaWhVbdKmfC6jDx9XJrxNh/QOSbuPSJX3tIb2TtI
cegNYM3d/rsJg8FHyV2U9h48/+e8Z33cxyNCNOwtatd9oLFV+bwac/sW7p7wOjhhgUpxUjGc6s6E
Z5qSuEupcvwUYofhtTfpZ2Xg9ZUxINem38g60qyC43qIBz7K+m05I7WC6wXQN8eQRhL0R+uPeQ/k
yCm9WkIE2eeO+gyco0vJsy5L8Y8+HawtU35MBq3qTDThETQRiTbYlSmW8hxoOFSk6XCOqoy4vU2s
i9Ft9aRPg608O4vOOrUxU2RX9BI1lbIxnFs4j3LsqhMFcjsIecxCmkQ6JWfqCQ0AhpF+8P4hCWLb
f/lIukY++pBE9eDu6MCbWIM6fkeSJ1Jt9xlR6CoJL7DKK8EHgLLkBQ/D7iXQiCR5KgUKzDL1Su5w
Z0IZUvelBV9mwTA2/OYm3JyajB1gBvZvTo+JFkF8jGnuzKGfiGZpwQMMjuFoP9BidGLsTWl0Nw2w
WAtes+7oD2oyXyVaKZOYKK5F5H5+8Aruc0vajqbZI/z1mQm2e0W7Thse9AQb3LSfJQWxBMHSU3R4
THoglrz0OL8cMeC0I0nWCZqjFPQbofuo+szoVHqoGQq3djrkm/YTK3rQ5kRcwFVZlFIB4hAMjIPW
ch8ravJVcW6FAgl3qQNdBMEXl1ZiBfVL2/tCpuHUPyW9sdIV3TY2ebT1zKzR3hvnBCr8Y6ru07jP
IVU46bkiGs1uyvbFIbAosIgbxywsvP6d+/JALd0/BW057be507NKHOOM/b9C/aE6amayOegAd86p
uD44X9aYx857TvIuhQUb62MN851P9Qow3mBfnjQKlZNOM7t5Qo5iKSj+vNW9STAM88SqfHeKm2yk
3++5NlCAM+Vy9ekZWCKofnDTVC4r1Mh/NFVhaYx5etGFhKSPq8yd5uGDxCeAF12WGJsEw1bEwQQh
83ewFalHgBOdKSIsifN9oK4y0WIPbVYXILdJ7ExyXr22j8md2hcrvLnrsvDvHpIL7EiX2vnEQ0+w
1RKzWaEphYZ2LJJWCa0eLoc7HLUgJCFUSK19CpuYZn2Wr2mVcK1Vw7NzgOqls74icRPwVrcptFFk
XkuPJnmnfDDTNbGUy4xjag7V84z5ykc5EUn5aCFyLDX3E7qYNNphDCtzJgtKsKs2t7JRdriBxb5y
g+L5qsmrd+sUyR0whPppKeJRP1dBm+DwXfdLOc+dCMCUAjrcXZowBJZQmyO6yF0jXUzooV7ZXT6k
SPMYjaKO4UCVAfSJptbKvX7kQM1McryvVJ1g3wcpI6r73sNc0YSRsZKqppv7BoEp1zu4zHjyGppH
n8iT4BsYNqLoK5ij3m4RHXJ7UgtuDVOJ2rH2EaULVXebkCv6hfofk7ZVCH1Ncwji8Ah0T8nY3pPl
UKR0SHuxs/ejGiPtHapIhbtcRS7BdQeskWKgTpTDBg0ioguYHS7UZCjjxIzRjDLNayaOXfzwUDRR
a2GsQyyEbk5esyi31ju4qeSJJFYvS/N5fDW9b8zFXBfJ+QKYghlwth5e/qnGaOVSya7wOu1JUZU3
MWq7jnR/K8RmJ8zLa6P/6F+6grJCEuA21J2H2iSfB/sOpv7B5MHK2ujDS+F22sp9f+tN4afE53Ym
IyIko1O6RC3VS/+/q4POToCR/s3pY501UsIU2c/3bKHCfayp6ct0cKF9l9A31S/PScctqGrGgDCZ
UOd0JOsdZ+vUj5LbAn8yGsIWaTxaqvG/vNgbouSO+aGj/GQEG99uctLN25W+NsAj0jbEI5j/D/mh
i8DTN4mCmARpSvEOTc8Rc/GIhaDXGuD7EwpyjSFFfsTzi8+msHdpw+M3y0J+6/satU3YXEhqSoHI
uNfeE+MmWy65RVQamcZOyMGj6lVywNhNHCk5pDNtUXzrIX+rN83Iw8FVvF5XK+U9hRFTUrH5L3Us
Y1Q3HP4oqc4FsJgUoifVRYe6xm56+rIQuIvVx15bBnEWV/eU6ilwQJCpwgecOnjaEKdeniipNv+I
cTd/T/m22LyLLkkMVlBOU0OSLDCteVyAwC+GUsSzQVmSoqF8TmCTT9j2xphVEFQd/wIWr2A4yEh8
gapuookTzXv9xW9osh+cN/mqs2zmYI/3LvXyhJV62mURqeN/ZEAUebTzoAqS5WxRmBIr0N0o2AL9
Y4E3ITulJnY1rnmYimR0ucO4SxyhXftaM9NsMPLxFSIv9aPrt7W0WP4RcmhjexQRjJ38TQ5f2/t5
quMLW2bRlEBjPAVWjWMmcRKqFhYQrSNVKZYeSqJSIJgFyn0A5htntNZ4SKAgKoHlnwhOjZpjNXFs
hgizKHvvdNgdn88RgkYCE44YhiTORJpqUqmRlZ7mQf5kDSZKZoVMOQoBxN7nezVaJEaR5A20P+bV
U8ZnEvOsxN+pVq0A7Y5p2MByObZsfJvSqzVGKZye/k61CV5GARSNSyjET3glj/rzOm5YEs3ptFoh
usJxR6zqdSIH+mRSpaIF8A5rcE9VRJ4qYbBPaUFUVYRkrnNssnTqOSvEAhVVXivwgEUzR5dqRZjD
9NprF+0bmQUEv8J7zv5VdGW8AyJ0mG4SmrXBc4FxVFUwt+bcI9LAxLWrEwJKYDMXvVqfPcq3Y3Bh
CpkSzNFYYbdF0mwjxlAGJRpR/KuNH5FgowUX8ua5Ho0wQXdHOGDHK8zQRLrOu101DLs5wBw93MS3
S8qRGcKZtzDuh0d52iRrjuKM+Bg+zbFnTlqjoxUYQs/eZOaRHRLOBzYHyP+22l4S/F60z5UAwnq+
pRM4kmfdYWlNn3Gxpsq/71pN9FyLKwLzFT4CINpp30L8psBqXNn+JjTq/PCj/OF694qID4RoFpuk
gUK9vZhT6+lDOhZkDRSwynuQ/TDpw4jGSQqd/iOvk2yKN+60XKRRYke0TXAg4ql0BvXeLQpeJy12
1R+3el/Vf/i/pDGF7L2cgLixka1N2y022g6XjskGaLFc8jrOBjXwtQIGBc7NNLj8xhg+ODHoia6u
qL9t8Rsdmlb7ATGFPk1GUcXme2+A8XxPmZ/6MV/qDZAt75YkQmM5Cf9XFZUy9AsJ1CB20SNWd8WW
9mVH1kht4LLSGyIf0sMV6B6feP540n1ORCJ9pAukcv/6RvyYu3IK3jPwf2cyZx4S1bH4ssyv5Lto
atsI9UG1FP+n84yhwMo/aaG41qtA51/dOo7CqUEEwR4CHJBK8f2HsEf3XvX37Qc5hDHWHkRd6tl1
mcSc0k1O1YshStQmkiiR3CAJD4y8ScRBGgWsKRx8zIjfJu4YBAeC/YbyPbt1UiutgrlUI154+eoo
XItFropxChcGG6q6dJ6UeKoFz0MDmGJEHIsfAVpnJ6Hp+CG+oWn8E1KN+o9W3JGLdvw6cqS99gW0
oaLYEkZtKd+R7Rix/LzH7Gszomju/q9mDyEVevm27tATmI21Tnb/FOtGLXjyFuwkZE0rlOxxsny9
XgFu0jsYr9nFgNhll8CkzBhUsn2XLsah9cERYHvXTdys2IERRF6ur9sw4Nbemq4UtQeT4NcjYhPQ
16XUGiJ7Iu1fQJaU46jZxRcLoPLgpJMOP4tkD+msvNFKNLhBvd80In7lAfeN9ZBjABJ6iLxRVvgz
NmqmeR2ppUnWCPdZdYxz9iKLPfZrQLxFjmi/46Lfw7EVeoc16IFh+uIXUiowE1njHOQVPVYlDY5S
JHutoJwHbgN6MouAZIDAL/Kry6WWORfq41VhLClVKo9a4TIoOLTcsI/XFSQeUgIteaA1yHti1Afr
+2dvVwfhej5559YhQEPvs+Hl3lChtTONoCbVlzqy2cZVf/c7qgsHx3l3mLvscqQiaSJLpZM7Zgil
no553BgGKfW4URi3uwopClBXNcQgWqUZgoZaodGDymN66A0NyI6oafWNzj3XJepeXs9u+9XlCDdT
a4nlwGGc1Jyu/muhSbuNnhvWFxeBsQWGq06Mc5WjDabyLiU3sFXWWS0n1pAmdjxtkKjT+ynwlNgD
UN/DPOhTfsgJTY6EkBoB0le9kYHETVH55VdeW9n01w5lUpp4I6+SbJjliqQZie3LBT5mTS1vKpV5
+qH9flP5AWRtHPmpanixpkP2whYMa8HjpK+sTgtecToPqNLNNx0F/Un58TkRCNsf4W8ZY4EhHZcT
ZmdfWPburG36QgCwtupw/7by9Akot+kDmW8LdxpL+uHF3QJB6XyRndZIWie37Eh+6gGjJr17CAV0
tznnszdGxZBmvppv1TwiibRwKZkne/vI/0StCQi06IChU7Zyd9absGO34Silsd/Y1ihbIy+C8g5J
esnk96r7zOKmc0vrn4wsf1V6fvnrRfxYe55lin7uUyVtQturkjWvGJ3adBn9kWj+HcyMI0oSmo8e
oudY/qptYi4wchwk5u5mVCS2elWqvgY4bXq9kZ8khsmgyxaHZIAeiw3aNPsUerC43oVxrD1/dS7S
VQ7tvMoBDE5Io5NdSe8THXoauoDF2O56Ln0PuOSOpBVAG5+ijT82Rpwq8PEcv2KjdHH03i74X9DH
G8GCK31ZqxTPQWNJYgKL4gA0F897ojEoqhIirqXxGtRzx3VyxGU6NWjdOK88cYxRLhFgBDC3CZzE
NlsgROVYY15znqVqkiJyqF8kyPAkGz7Fibi6hVCU3DSV9xhlLJTh19zNPvgDTjtdZczuNUqQBu+g
srRJalMEqd0GWbcoh8lvcu/8JWGLG1NYWJQtViyUJyw8kjemF6sqQ40qdsLtV/W4gcPS3wtPLnfA
gLJsrAAEzgk1VKf3hsjr+jBeBgnMdNBTuSvLZUkAOWKl5YmRU1/VwkOnUtE7wJLvo5uDOmprMZTI
2WoqR4KXY7KA8l+Vh92uoqo0hrHU+KjABevshyx4MMmQhoFZf+4Ohjv+2s/TAuwr4iCArYncSo6r
rPLZmeWJR3lYCAMKpXCVIrQJl+6hNTcy9rh2JOUiWjivKb4OLkucbDWQBsVADg7fR9aNxmGMWspM
1uC2mRw8wjzptk4aardOgCeSnV9jk0GRLvKZHDq++JRF0GlFoZ1Uadm5sxDwuiJngrNX/HaR2f9J
wH9zrdx3tyomucSr/XfKNp+EeYPoBGe+IJbclDQFE8jrtBCXkID4LtaYZX1XD+CElxi+fNdOdlji
iVw6IwqNY3cBgvCbgqF51HTYtfffvdseJA6CbqAe8xMPfR8k1wngsrw63YtuklMOq6cKM791kxJ8
2nwDShfWuY4m2SYbkVuz4KvDSxgkV406TVe4rz23zChpD+doAwgac1YNy+ag/IkzcyZLwAfm1m9s
mY6pPmA4ADFTlvDk4W8acfEpjsp4TLKqqmjwWkVk9tcMF67EnFOcBcS8iHa/jOTvWnDRDvRpVIF6
vLSinfo+WWULG0yXX71CDJki3QF4wOaAan4dRvcw5i5E8g3Nc+CtnKJprJBWm9Mg0hXsKmxhHaD9
rotk403fAGxWTF/jqIbWaKviHgKd1VTLCksAUgtZUj9B5Rwm61ZXGZI09yS/eKFp/+Zh4c1MsLwM
cW5o8DGgd9ePc06YnMdAvIANcGZ3qe73nH5DfnVjGqciLtqLKX76XSLWYNJMB0bkFaU9sYZGN/HK
pxiUBJAdXQSSOcvaAatSU57RmPYNkAXCmIPtqDfjZCTlI1+zZ9V5ViDa4evJrymvjyHZ3+dPPi/M
PIqD2R4AFJCG6IydpySDw208uaQJRc7gmBcWsunesC4tEx3K8umLKUNBD3iLI2B9qrtQc2bremvI
mYwX2WP2Zst9n6Bz9U0obv5ilabJT9br5uPvTs6Q+32HpEGDt0PZ01LTBayWrcfJg1X7XM7jciEe
/LQNG5dMyX1YJVkafSaR5yRLP8zCGjIoNufZIlpN65NU+E1HrL+865Aq36EV768hbvzlN68T4vGG
7KExWwyrWrlrsnRVAAPf+ELGc6BBeNs19Nte8vlFObasu/Jb85ao0LSigKIUzvWNPdCsvSBah8HI
1ZF9Ra8Ff7Zwor0zAgAFBAwZ4bC5/TvQEVcVoSslp30q76/lPk7TWQC0VhMMRlUZWV98fvuVUZZA
ocgWI8muEciMIffZxo/hipVDLJyfP2WyoKQkm2oOjc7kZaVEkXyJ1J5JcwcrR7YpaDNmAg3RpKBc
aaSdtFGJ2fwAGomf9JescAuE9pl/2RDzBNZFedjoEECN6EK6z8Zx6L+Qq4/ReOs0kbbqpMpK6gqr
767T1pSEggrjiC3kpxZw/ugvbtHgPUJvL97RnXgb3qvbObaaesr/uDjqNUqMX3chd9kZOKHkP7pC
yyZX72zv801280ShriMgJjxUin+Yp+gPx0FzPTNIxS9Dh8AnuZjpQ+ilIWDxJBYy5/WCA0Zsb2RK
K+GBCLUTtShOfue09fpFxE50b4x8Lj8njU48YHhc+yQjMtZQ1P2yzMACz7ysbTLnUy4WRp4RjBeq
i0v3x7qb71B60fvFm+M9nxcVseQv35DZ7818hvjnV6E2t1QQ4KwAW80s97TOQuG/+wjOuDxm4ls8
LTZS4yr6zsbjtcki8UzrKUCWWl39jtzlrjbaYNz6Pcgj+JpulGqXtlMswFkMMbOGNHfyyQRU1E7c
0woqxB/qphcYSyDWSSWH2j/FJCBB9ru8ospiA9OCIFSmZAoBuxdLcgIIORRITN2xxH31QwzVx69J
LmCJV8bzVGvkENEFK7Xc+BNWdq5CMPh6SZCRkYTH/Ef+4iH8+zvbnNgSm+jPzdlPp0f7PehA8Dsu
dxPhsSE83lhlwU0uNWf4n3InTOeD3mizZzqCKiBW3XqWM7rgpys0sZ2HVNyBcqsFsY3gkmhWk+Lh
jztuV65yqb0FMiSUjWkY5hZdLjlgE0LtgICJ/xWnUcj7U80srQaBV0A4eNFbtq+Xpkkpu30UOREx
QrIk9GQpn1FKStjoATXA8NuoLU4P7ik5MU/wJgrkjsimTGtycy9nZ2GvTa08XP/IVHxNqO04ttP5
QgRQpeqGpu2cPzHn4yD0G4uPw6lRXmgkEvbd/+GazlIn0UfnCkqRiFTYNk5N6IX6tTsRATk3xlr4
klXXI9TX5tRhQWJtLWk+/f/bGhWhS6oG0cL9hnljplOQ6hRiZ0YV/kPq4LXj71MM/KcNWEvFYOxU
RR50Bc6cyn53tHbUvPjb23ZzIP6IUXwrZ6u2GNVt+pu/rRM/0emC+AAwTQ5dADVsNUVrS+7gJF/4
PME6NqtpMKF6l9MLA/r0wDz0ONpV4hg9gYluXrkUYlV+jXi3phGp0nBd6cMBGHeoo4dorfctPM64
HScwlXuH5CEMIlZiwjHuBRxXtxxZg7eFWBJIkkTj0wa3F01G0SfLV3KV4XUFfpQhkb88Fjuh73+d
8zXpgHjZ7bZBH5EPqN+sLzkslQ+/7dd6M7SF3hJKel3+wRX9hDoIKBlymBYPYSHNEXMpgCXqm8ZV
C+hi1ShZyEJO00eC57AtXbhQlZN8OFJfsk9p6IbFsbE0A/5U9+DclVAEwzrfFb8lI3919tFv8HWM
MQjCyn6C4s4UZwWDoe3A2GmTVYTfL+DsUKCAM5LlzwLCL/3onrJkoLeq9bv0I/EDaPAngJtYVS4d
dSMix1eEq8jb/te9y6QyW2t/0nEkvMhb8TM9GUaHIWZUDesPkLetP+roFjl/UDEBogGonBd8oPPc
aReOpmx0auwiM2ucuGYBjw284kQGXAZH3+UmPqxKmz72qdAH9vCBFaxiuQRNXmOr+KbEK1mlU9c9
p74aIn2tDPobrKmQaVfDY1dlp42gmliO29ZuomrAqO+fXs51+y0ekUyfw+QCTkoZFXZOz41/r7IY
KBiksHb83Bllfw1bNXdSHtzy4K+Lerg0QxvoksIl8wo4sJBNiEDxnxyaEoqMX+4AfFT4Eamwj5q9
vhg0y7BvoGM6SYSKLBCY+btBUdkFrW8g+zP6CrFKJ5lC9IjK4bZN2+TdJzkemiTM4t3Jgn8YGQNS
oGZM25sSo5hbldV8S4iOlcNaSOkM6j3s01HNhI3o85veSW0heX8ZCCY9i4xn5wg6xExdd6Q82kp0
IRmfjLA9GbCXQm9t0iZXUK5ZSeDvDZoG3SFXCS423MXv5DM/QJf6/JrihWVrbDI47CI44u+IP5Vq
lYGYXkR4jBFnS9kqxJuBidNfhRItwg47ppY6snImFDvFN0VP6maWzSLRZfKdV1wnX2PrYTcjRjz5
3HWnfjgWHNdslOgfsR+VCZQKPyOSocE1ybJfwnL3NSLL87OonySEh06qSJARd6K4bAxYAlipvIVe
YtPdGuZaKIuHXDebY/sZabwCchPhepD82btMYx+UlQZIR/Hf1M7csmNS6lH2oxn3m399vyjAksmL
MwC/wuZ5mITN5pYxq7KdNPUEevYSy99ykuS2FLYjglbLoOqr5WseG0jKmvpS6AeF/Ps8/T7euuRO
lx3Vq/pltI9P0CF3HEjSuuG6OQJDOunfTHIi9/dCXuHum/6d7VV89B2LzeWhrAqBNnQhss+pL3pI
/UBwLYEmLMJMOhZF/mByZjLVh25nobyKcfGMc9alJLawCXAE+qN2iBgqibk3rrYjZ5YTXgraK2Um
aS+Yyc6s+ooGHLKMhvJaI3KsKIl//XuuraFnb+cEfySMINn30fi8ZHQSW9Egt4MOez0iz0pfVGE2
5reKwWNwZ/scQSnLHAcAbKDfrPrgEkv2Y1M6zggHlyZy1FkHdm4ShCaGhA9zG4H86fYOxluRPARH
2bKfV9qsBee/Rzk+OJnlL21bLtE7IrGrzzhKxDW4HZHcLY90daZI21++XYjhbH9sZ/B003DuW/gj
bN2aQl3HLy0cbu+CV8yJBSUBVP/rVtsZcXm0xUcbPJhuJmMISVMMLACu6VrehiQouba6ltE3k/6w
rcgWXdx6O44fViZVEpHcKcqkyjt7fCYDRuJR/rhKamITNxxDZBtQXS7rKusx3r6vwWgbO7+38jeN
tqek0VOx0BwHaMub9Eyw1F4/yCbZJ9CLox7qZD/S0qvqicGDRAo6skIUweFKvnayvHPrY5yww0rl
aUjhVVpMUGcnBZL8agbzYbsBOhh7+J0k8yOay+fahsZQfZtmvuqZSxnyiRmExvWQ/qzb8cdIhUBS
JVo2WpnfZdLGaFjXn1SJwms1LMPfqVk4j1DmFsGrX1pkb132SxtjcbG89K996dRCboVDWW+qb7VO
46ajn1B/yvma48JNpy4g2KQhfwOKu4ORsi+oWFQ3vZRXMWQCbDGuOJ4cyAaXiOmONMBwX6ialpb0
SaduP8APJ/+QF/M8jsivcKKCaq4LPUlaCGZN70s8goS+u1tgAGfF9wBPSd4MKMq3fHsArA+FN3l9
QE6l7N1iwmiFhT57tzxPr6Bj+sj9zba7ZFFZNA71Py+0+uYQ+tasJb6qJCPge2Gws44I6+/IjY4V
n/V5WhDDXiAPmwF4mTs4dJaNHG4UOI6z3iuu8HsZrdkp/3sW7bo8luRx2dpCY2T4IB/tpNOfierV
TQ4yy1a+12nQV7UthjojThZfH+S6DY6nAounakjw7REy/oVfBQrXYfKd96/hqU26PWECGUjc5ofr
VrJTvqmF3KLJNAgeavkbKPRy/p3BhwOSjsCpCeRwKv//CDdPPMhGR4aTtL9qNQ9S3hJ3BJmQIrDg
PvlYezj4elvmyzNK2cQrIxnqeMrWnlyGTuLYPEZQ2y+GfI981ATCVVDQSJY2yzt2xNWdQu7zjFuH
Ve7LBqFRlyv3kpqAb17Kek564eYz0A3cIyVX4g0UI/3N3R9vfEySYmEfGePWcrIJCW/iI3lS7JHj
VTKtXWvKgGGAElcq2DnDELA3g2+URSlMqa0QKH6E4Aeqxar1LG6wnqEFQ+1eSIlwb6RhXgkrxGJr
NHsdJ2cmov98eJcXdhgCkwAGxYOw4RPZ+px4YEtMJnndY4zviDng8m4wwHzCBZ8ICDfAN59r0SDB
zF8MApdOTyQ8hTq7estUoj5fI6v09qJkEFTKIr3FSTgByCb6Z6/IfxZz7dt0c0R+MSlvlROgY55J
lEOEeRZLGaWlBeSoLQNIU/ZSYwwxVT20KLNfUTjrZb50QP3IlFGBCUtlRBDm/SHphV5/JsnOZJvj
vTrmEz7nnyklapOg2yDtXLO3+aw5TuhoFUJnsf2mNucATGOQrL2gTVUu4pw5AIwzzI3utglWkC4J
/moeDe4tg/MnnFXVBnDrgn1K43Pwu5GZdOBHPUZwSfZWvOEqjPv8fsvVjMiTG89kbR5Nw1UBI814
PnVu6qluoNylFsNyJEfCfBhuWal4r5jrNecCcV5rK80ifxzX/2ATYHmHHSTuOJJrEHFGPO+Xm6W+
FmRRaXnH30CqNom3yhdifueopaJ9HEVwvIRXHZmDtBwKViS7omtea0neYqaDYCS2X7qE0nnGzZWv
YcSnQZisaTcK3KVQz4QDlB3RS8NHpnd5SKHFlysGBfZmN3Dj6kiBq/TI5LRUwzXJWtDXW6lkO8Id
Q4Q5clECqcwqN6Ivk0Uxlf4WYgZL5owS7n7viMPOLzl6MHn6vHOM4/NeBvAqmt5h6g780gNEl4aG
I9CN140aZtzc921kf0lW/oIEC3S/WmWOPcZGulhTXeuqiEOwpiwGsKie2Xo50HJ1YlP2jsoBpGmz
e7KWTgog2cusjvmmlqwKZ8mwlUeJqiJA2jf1AvRt88O6JPbnKFonYhKPZwTW2L+4FIblfD9C7Z0P
mUy4qopOz1vNkS2NLBS6wSJT5tHEEiZTsMBfiTPFCEXE6zl82OgZwALOV8bBjYVc7NY8p0oZAQZ3
jj/xK9G4RKZ7g6dxe4fcwDomL+CPe2cLqjXHTfubPa+6iM4/5pxv2Q2RNyE9zrLl+f+9WuKkaJPK
YxNjzXT5JwlKUmP+8Z7udfSeX2CG2oc5+5gk3S8+CWk6s5Fbs16LzQ/LjxT+g7ePhX42qtUqDKpL
z1rw3jEfFmUL9sPUf11Vr2YDNb0vIvYrOGXGq2mmbkEKHPu2pDmREkQbPwUmPxGlVzKQijGA0Mrg
zyMjjUXsYXjU9po3MxliqWVu37cmJ2C6KAe4Nh4z1dalysBslyL9x3DgsIGh8ZrTYVzeZIbGOTSM
Kvc5zhF1+wGOKgoK8SFwo8/iN4/mZvZME0i4teQAAL/7JKdM+HrZ7r8GRcY2aIG46TCIIEQZ54Xi
auy5AgrA533EAlm2k+JFfLQjHnGdP9TC/kszRuJLBPsveXswsZhmq9Q4LRNXAozqhmeurnpZE3UG
+jpGnzLQIq2kD4HAOk8L964O9d/snxENy19r+q+F6g7gzWlPrP7zzmvSTxa3CuMtQQtAylrpcnIK
Ca3+rjyfCsI5oVIPlXUstRpBvLukTnQX/941/c+BIzReRUA+ivEpYjuIiUcizdovs65Mxv27XVg7
R4nP5aouenfExnWCfFj1lurdysYvmBurY2A4I1SicZUidSUnU/gQwxBiutH6Y5gqRPkPnGF3uuai
4FhC9gMEtjjkmXgz0+u2OzewtwMAwoEAM/uVu32OKnN/db0H/IgYfgqvgOt2iZdw3qAXJ45PbkHc
pQoG7dEbEPrlG8gvTpQ9ZzzvdsGv61dACmxABzKdMm/Y6pY+cuCRADxTpRh0Gu/EYb0h4XfDxepf
GkLyiNDzNEeDA5v3PBtrSGHs6sXqp3Cw6ZcAdtlgn2AmU4PG6+uO55GXkPwDpefCyos+oK6+nZJ9
Ehmp0tUl1GVAOeVkodwhx0taUe9FVxZsLxeC1dvheRP5az8XZ0qI25J3jJ+lNzZbFTx3FrL+gJAe
HNDsU5b5XQoYbfKsYugno7hbqCrk5PxMAsu6uB2vuQD3dnNMBX0JqxsraK8vB97sWeMnqidfY35h
XnZnsXISJMGbgVgJIOraGgb79gRTFGyF1TDoxfjG9Q3AS11Z/bWYwpMPKj+KIcBdV4sZGAQ77odk
4WffXBxXrjr0RpPWB8z/ahvXANBjbSS6sLoF9xIWeM6Q5Y4Ni+CiP+HOU0JTjXKCntZyz4be1itG
Wb4JMJ/hNQ87aLZ56EW5Uoe5YGLnaosOWPJHUdblcsiCUjLm17Rh7PtfCj3xsM+oOLzJSjqrIuFp
tn9lOf7wASSOLKPoDRvB97yAw/yHZbOAm2LPjTxwGKXCmXlz2aQGLB6ih5oYe1/hmnurwr1szigl
mZCLmi8Aqk0i2Bgyv42qbD/+H913YPtDd6j1jfYjgqLbPKM6JjwDJyi2zWXdqvy1q6AlmKqODNa5
wouljD0tnlcigfEuyfTtpCPGAqj8KZf9E1Kj+OPPKlu4uhyacgZyznu7rzgL2URqves+ZnkqpImH
YKNaVZgrWGRyWphnAAnomqx97bHQjRD7vjh/TgEJkzkrRtq5nG+317u6dN0JjxCcZO9wb6ZCSNLS
tM6qfl9O2dAx+vJxQrqJlz9KHcOk3Vdv3jnCycqxnmJQFiMo4tSXVfBJJOeo88+pv8uP9I9XJjLY
cbjFR8W1JNxQj5xG8/OdF9dxUwO4e0ztbV3KGXRchgjUsF+nhgEiBcGonqUvSIoN9WFNWBzaRESk
3+j2ofDaQWMXsVOth6C+guhYJLH63uqaxiVH0qNx7Pukw9E0LQPJVwhrnIqcpVe8a9NtDX5V4iZa
uj3vuseR+eTcwvjtpDrSdRgSXq0T+7eMU2LReh7kYRUr4aW6izcJsdfMps7G1d1cdIR0cM6ovbQZ
yzC9QpMHIuPIxpxsHa9OiHH1KM+auFDXU7zSLHcv2FlGWfJFplLzBV1TxpxejYoequUce+1R9l/3
8Xmr+v4IZysvUAS4zF8dCivC3V98B0x3jiGVQRMwHF0E52oSW0VMfDTSbK2cV6ATWjq75QcpljBm
ZNzv3Z2ey4TOM5KJO0puqrrUMYMfF3Dcxzc8mI76ekgKMgD2bTnoSFxnXOopg1K6KT5DYef4YAwP
ZsbAIPLwqgDFvZZVqsrTftL6whU/fvMcl/hAd7stgJIaNJoCACJ7+lVRp08TgNA67AEv7Bn+poOm
ADowBk8XpZOAxLcyiCNmP/qRo69fvP1ACN+4NqJKAtxV9Xk18zzvNv6SLw2F0By9TDou4j0ilCYw
ywtCepJaALVMztr6r8FWVa7gFVKXYdME+ZdsI61UVI+FkVgDwijAtPxRQT+2g+YF1gl9ijSMEHVv
lEMDDsNu97GtGLT2okU/tgiX0GjGOdSmWRpMRGF7LcSO+uYitDwENEqVfMtvk0UHX41aO7fw29XB
FCP6Ux94Y0SY0x64NlNf5NnheslZ2zSXKdKuhh5jDv11v/TzYWWEOkMgyDkNumEUkv4X1Gm8tfu0
93+kRRsjTJGFR/uG7Ac0OlFf73qZ9Q0EEuCIHJs7QavgyJ6QeVpqPVpG12y5GpVCdDV6i18gqIt1
r3WnBsfdkKwJmc5d4pYIsflsgsdxVuAFtKePokJUTfHq/rQ/Oy8kIYoss4zE4Gd/gf7yeCJt8idu
lrqQwvwzmvpeLjzgiicDwuJete1r9pDYZCDIW8auSiDSXJeUkHkGX0FUEYAzsewGZ/5G8IzzppU1
qndbrRkYGPGH42M+rWZ8fBeQrt1RDgelMc9NX8liSwiLpxWipueHlbnOt4BJnyaSRPvH553Xa/X3
VHi/CaZXUyfkNRpkWnT6U6eS0O5rKqyfOpPuYRVQhuJU5mu/wMA5ZLoKRJAZhWVe+V7am3KEs2Se
eSCKrsOgM0ZhE3MU+qqj6Dw2bRdKxSt+3AeaRl7Tgb//5zgXaLbOq2A0n1lldMbtjC/Wh91t2hz4
irq342cU1rsgDG5/0lXNBKJUW9dCMWBFuksx7hwHiJOv3dmwSG5iX2YSd9toax/lDFaRcowqdkYM
DQCgYHh6P13irwKH7uZM8IiZmAEzF3ntgKJ28fVco20aqQIREzs/osSjjpJRT2GMQxzgYakswe8M
gzR4ZT0xsAcOu8aXsIGYsRDaGx5Rya9Gakl6a908+Hi7kb14Sq1IrBbLT/KTPIeLIviiW+2DGd5H
uZzrt45J/agd1d0rj+AOIvUSiY4ElZ8rlGlyo2bXOl5j47+ZOif609bfXRXXB3Ifhx+HaqQHVrib
DhdsDTFqVKhJYi0tO0035V+hqpGQ+9/2bGiPAmNswtTEr6t0HaTXpgkaM0odeaC5nUgppLoQN7ux
zwsbmirHav6VUhGo1tUiUN/roMIDCeD3D3Hsl86Amug6+KbEjWNGkXxzGlz8YfatEjKoIPCVDCWA
8E/ANvkfmanR9qc2Ihb2+VE53IvnrEOeDRmHtFAyvntQMXNAf3n2cvqpoyddEYxSGOj8qE9p8Ei9
uou6F6fQOJhJWK8su4yedR7W1NuBG2S85fFCt7mS1slOVS3WreJ8IdIvyGIuiSvIRjG3h5j/LLKF
eFqYhxDVhnTZfK/0JDxyUMHm5qTmPt+f4zhFeF5uOdEwP05rY8mzMMfEkg3mluyNw6pnOoHOJL8C
/Ko5gGBOwGYCFdPuDQhawqrpq/ch1WsRBY0oi0Cml+gal8ZJ5ERtyj8qVeF1TKQvK+hk6gSS2Yfd
HbjjXXeHsY3Okhveriu1DLl6XyC4gYbrqfC2fqIu7kzIujH0n2irjH5UhTEe8a9J6iDp+9OjtDs5
D5qPsD86JiwEviXALesosg6IolzDKu7916mm7CMZ++H/lS1sJM6NxkAOW/pH3KVI2YikFwA1qzoT
0/Jt3AZlzmr3dt8n2V3A2jAP50R5YJQYbpSYJ8/p33ilh+TvIPZKSNiMquafxKt3mRkfqqSHz3Kg
aM7WUccJhhMQm0B2haSYVNCwwKEYQLAPdUHYWp7+Fjf7CWvpvOLmVtKh8WyIsIaH6KPhyq9oI6BE
mKwNMWjHEHTdYddAAKdOVLxUtlJw9P4AicfRt0yf1nxwnZYRBmjZldV3OoF66e9HC3vwtYGHJAFW
xRcP1/eLFakOqaK6pYylh1rIkW6KT9iwesY9g00sK5QoGr5tGt1BQCMTT5uoGYoc+2DsLPv/Nr30
I8JBuUhW9ErJFNlXrQv4TKA8MAfGYw9q6R8CtqsI24bUvBaqvISnoPq5blkD+BlquwmrnTMtwyeu
clU+wAWN+ShLDX4LEHOlK//aXxlr03jbUf4Y5mFOiBHvrYaNrOpssG60lWJCOc8PzhzfZRWZj5RH
BPrEOGnyJLdsaok1AyohjAnLC1PEl+k0pCH8DK1ff2+6x/rtg8x+Olj3yJTbWJoc+XVGxTJiGXII
pY6GnUcq+fek2mPskJUkz82nwXZCHdLoBOIbPnFTjoc7BpTSzAvpgPFeZtnv4A6ailArnaZYTlxc
JPVXMtgsor3lWi45qWK+GvbosEun2zpiOzgQ980FKsdI69ipjK8dC186S0ffKhJ6N/WiT/sAm7xw
pHwd0Lrd+ZuCTrNTrexjnmrsabH9pwtB6v88pgFheiS2zplBhcrve/UvvrSqudJkvJRpeWzmFF31
g+fzTUtSyFAyaQoY7ZpHuPEAF6+GrACSQLdFl8cHBK0T6hIwSJFJmvl/U4GV9cyhot3w+MGuaKT1
5C4Ngjbk9r38ndEX4sPOo6ToNFeIPM20joaO/sKYnXRfkTIYMNhhvmQgyWEedvmYZAMcUEVaoGZO
deHlLcyYelfmVtu/nqCYCNU9nPFa54SAZdN6OiEDovo9fZECu4gXvKGhqj/1eNZeefyyP7WdZObU
mK02QF8uMJjgTr35fNQBxzfvmNcIJu0RgKaNdQetNCR3txa4TIGc8PG74hdi1LadAj1TqjCZFmHd
5esiZKadr7GFT0H67yXEel0XV+kko1WROd5R5r5HDek/m+RMpTFO9hx48aQuFxN84CHxRBAVMleN
r/nPfo8VaWUNFszpZUmSYkVovuS4vrnncnbUSL24w8SVnlTt3Z2ILkFnxerX+uAPvlRK/6Rk5CJU
tCBcyT/JJrcGeFi07jx2lUgdxoXcV2E/sGxDhvXydFNQrcwfRNjr9yiN38lp1MCnpmO961w3VRTF
CRmJUFcp7yO8OwBz4eUPelBgbBqycjSjbjAqjuhcVdxOxaVFVqYzJTjzsv7KCjJ4LJV8eHhTFXri
aYiR1EAj9bJPOGmiUboSxnsqfyjRI4aL1s5wSoEsivcnG+EaWMUc+UGUgdY6Z4IOAHwNBs0udhds
8mCa/ImmUXl5QeIGgbuVr0KwvVLnEx1q/24eOZlStBkgRHi+ylT37zurK/aOF7cLC7snpnA8Qisx
RqjuwnzQVLYzEuyNc6BHFHdIoZkybuP0F5kEmxKQ4o5MWKkRkaoQKanrNiqkG5PpUgl2Xoc8Pfc7
pxsBdtYSEEiNmbihpOhbe+NFgDbRiE14BHZk9khUH1CfiXRMIaiLB3yxb/C+A1JiOIvR908x7DVW
IVxxLokXKSvSenEsOEMP9yHpJffDTpHVouwrYwjeEeq9RAPY2W1wBHgmCCujJxm8Ugf/cI1mFRuX
KiG7fbhMj6kRqgxvfiYbzlBfgXqKubmbK0W/kWAGoMSj0N83abNbvcv06vajtcKZMZgIyNsHAQAm
cb1lFknaHUMQnO/zAE/ZnYBCZkg5a3wsrfOUH4MBTqBULHxLxJGQFWtspn6elF+cvcQp6ulTz79a
NU+wq7u2F6PMLgPGe/O7WuR8sa8qx34PnoOmdXaRypA0cCvZEUtyAKmTm2Jh33LcVL/1/07yYSCh
pb+4eoxGpIxpo5nEB3Qp56J2ci4eX3cCGnTQijgQKlh4XL9jSQpk1wjkaXDJseGlnAaQBFJ1i81G
HkR4oUSo81T9MWGfN+BADrdoGlUalzeo3vJzIb1VvUBARmMJqAlt4+qMNDLEblLOVbXl1yTOOuY1
YhUuavVxASID0g1HR+2No1rAbuh53raL0+VMA+/AdtXgJZQA/lyLwDRjAsSrrO+gi7xg+yt/sfR1
cv8vFVIcJKXrEs7Q9oGLEGQaHo4hoQMlmr8ZOGrTKYoCLHTcYy8VeVfkF9kLv2EFWrx4Qla5Qq3j
CwYgknSnimCnx6Iv9NIEf/rOz1MMCVh+9v0VWg8psIi1TA+0YY0Lz9f9wnXYBgGU9yYmcw86ijSi
DfsvKjNa5fqsOzJZYuL1GC+WrD0pZlejo9PktqdppFG4TovqJY98VUc+8LeGz3roSfjO1oQ2FueS
2aQvqiUo6yI22biOa+7sGqUH4ILDF8gsHI4nW/A4H2HCxYsINaPhRB4z/1wasGFQG+jurRkVInhU
2WdK6aIlWOMrv2+EP42PvnsqEJx7JtfpMidoKmOkABy2gPNhxLlSqJLcLNJh9xjeYcu4qFBVsQkg
SHmKnJvS+/iEvyCHr2NZzuYWK0mFFA4Nomp57VNefRe+wuOPfoTysnPxfC8xiaMNI3g9DAOVcE2o
1PULptOK2ipagnFEYbnMfGs9fTV/7F32GAPXVHIgMrlR/GxATtzkr1o9iF9EHb/Zg662PORnnfw7
JSdsAHo3OmNggxugI6cmXKN8R1gDiDb0ovH3NDJM2DzJMIkBBvmIdqfkrLpkK3gbejYlYVYnJWG5
PVfY2DJWFfxIq1lKeWDPHFgQudL0TSKmjXoE6f9mG5rJ57vhaBKJiITBwFjBqAW9MICETpksc1lv
VMO+aU5DJN2qGy/CwGmQKSRKoF30amsf4iRMGzMGs+R+LR11lxtH6C7CTqQJZTn/pvjGkZZd16NO
PW69m4f9YjjHCjvyMGBDzVSaMRNCAz8Z3yG2V72ZLceKVRx9gcBKsP1UuxbHylxCB0oRqkuPr4wi
/F2aCVsZxwMceyheH+qBh7vRAsEM0ke4JN2PCE0czWrPwjQ87ExicyiAdv1bja/ESb5K9JjpDDLg
6tQckKrgoYT6X9SJZjTc9Qfd5aE09oc3fan2itl8DzH4kigZNso16K+mEvso3s/zNkhi8UG0D0gE
1qbCHgAE0lGi2cGTStEMMp+Efhm/f5rXIfT5ulf1kbYKcNIEv9JDrTj7lqjxbrnjVdoeoQQRl2+a
+jWvqOYON/4HuIjlCrdEn7dMBjiXV7JuMgFaxKsYAyfqj80NX9am5l9ieBSkFyXRMcVdpkeTUerT
Gugbtu34+6FB9jYvXmBZFkOCm+GbpDx4lqyUMcHug/nkqa8Lo5uSywDbRt//ogoBuBMu9x+MnjKs
MXUK7U5bZgZ90RiAryYqXeKiAkEAJUKezg4COu9Zi5E/Odszi02EaRBMdLM4e3LbyaTsV5Q1MxOK
flzqJctXSWXtk08uxPcYRnDYgpYQsHaJ/mNRPs7qiBNcCMdmHTq0TqBYnolK5vXvUqc+KB2BtT8k
KycpKlTopApnDbr+8UI+JrxIpjxao9GL8YVWysIW8WIzTgwmGbUYD0RdSTaXSucgc0Vvp8AsM5XC
d8s5Iorfofqeom95PeInD8peJYxtjtY4Ia/dBA8QEbLkcWkS1bq/+l42Ubvc98zbkJG/f3rshFEq
gBePXg1sfD9ZX+qp3T/kRZgsTzo+jfeMMDQJxHyFNNzXdULj86XLE5qxSSSnEwPwPMoWAlSVWbpN
ngrId3HxkHeYJOWPz0f5vWDcgz34IhN4ki8ajmpKvkNipOa1L3+FTCaVcJ4uNoTkUs1fJwLnHIJ4
IUdrlJJaYP42mDsN4MuBsV17JbTOETPHc1SexHF1LrqBG0Kuk2dYY/Ym+EDTqqeyt+9kq4VxzJYT
mX6KXjl62OZ5eLxQX4mdFqVFPEOZYenu+sT9caAWkImMr4DOa6wKHcmqmNA9t7/eQbbJh6wE7MvR
hoMGqGd3ZG38cUTLGBVvtxmTc1ftaNDeBMIfBUAO7lGXCXdnBvFFgShdQSWFO+y41vqyxlHQMpo0
LGHMvB9VuHHts3a4WWCzmiYgHQqscw4EWZnTeZOJoGOaHL3eVm3zO0mebadH91PUqbxqP5iz8Opt
Q3XxUuoRN0i1KiSU/yNMCs+jOZ6JLI+QPkJCJWite2iP3gaUKDu8Z3VXAyjJG9hmzWWQe9Lwp07A
8sxUjVET10mVXnBdDkWgZTIvOHZGoN3Mvv9Odn/jDH4BVpYymTlzJnumLYY5SMeTN8J1eCl3wLTI
UGUL6lPYQegAP8StrCQfeWIJ5T3jk3WCoWEyDx3Igjhwrwxbj05pfaR5UD+Gfp8MTMraPwGzkbYZ
H+eCyZUMMyn5wms6oPtQVdvFtGGMjtOOs8lZLN5KpV4gYniKqAuJAWVeNVomgK47axc1umSCp8FR
OXV1BI9nDOFFT+EFaPVS5on2DhmrGxrgBTdFMGUMQG4mUaJdW7ROey+gGmd13CuqMi2lBVsl2rlP
HhiyV8KtUgteDNw2CdjgJSIu+7VGZNYDpDQYjz9xAXNO6bQtDch8kGyiLsnHsChM+P3B0r2LDR8F
9rGGPa9vNMur8W3deF+mn2/4UX6G6Apdrx83gwTJ2S5mALZeKUyHFpRqu4BwMeMCzY7He6rpgRX7
oJ7cndOm37GfkaO5UVVIizTwvTcMsQoL4QS85hnltPa/CgFIvSMs+it+5i1wLT9UJMgKiIuFAGQ1
oSy3cSk6vvgOwlJrmANuKxTQZ7QadtXcVIfMgRM+sSCsg8ezJ/myxaJ0U8I16mC56mY1Bxu3l/7o
CjzWdRZmGMuRMrcbkCoFsjCI6b7V6rNuIb5fuTDUHqkKZUb69fa8PMOWN2PpAWFc7r0hvkfmN0eZ
2/UaMyC8OM0iGN0qE7k63wH51GY0Np28yRvzb0sUglAJkLZfQZml3opTGyAxwANFdrcjWtuVql/f
YFQqB3xkmzTCiLB4lhYTxCRzMALjVkOAx8boIZcSVHDUqTJWh7H8W8SqqFmIRbd2lvD38pCqrVdw
7pbFB844JGkRhqT/m360Ulwk8CeUFKle+0nFnsw/OjLXTh0/asD5UtUmeCyQ1AFs9H0PhbD69P/T
LvI+W0FPl1n7fAwc/XwMHK3EDKEYsCUAazo1cbAGZ1pOYK3G29kdoXWgU5r75voY94YxUL9pJ1dD
0AyXWoNZ00VW10w39n8IXENYhhH6FpTuixcExVkmpAdb6/J5jtHaVZBLROJ5FuDy2nGg0a3i96ko
OyJb/lzXwRRcjhwHLZzB3rJewdvlT8oZM21wp7z9yGtvPMX9Lo/5XyuGL6wYo+BDBb0x40HsXnRU
w9JejZiKcvg+kR8xMDTj0xqbgJAXuak++znCOb7HorZ8+aatw9rvcIcJrnK4nQvqGTheRQtkP6Jr
s4OReZ5mjBt7MXWoJcORnXKow+2OgBaHS49uIMDwtQFAN8ayO+XPxgjdCq919M0yanZqmp7Javv5
GaFR9BzJQVxQXX/fBrGs1MvBSScHUV14cCW5Q17PKwH5dPkvvEjSQi8ne4/LBr+e7ex8A/xt82Ix
Xur39yiS49HNkRfBnmfusELg95EPzxc86MfgCyrID7msuPbpMRaCGLqbKf3znr038D4itCidta1p
e2hD5J+6eE65P3+g6QqFd3oj4rVy7ZQbEflWvBm6EVeGihfX64V6ERD6K8TPh1iJUyTJu2DywsCo
t9KdSlm5e63MUNrC3J74IzumpAm4Lh0EkHKIURj9paRXHuY3HL2L+abGkvMz8S+jmQSuWpWty8LV
al+jpaq1W5u8+iqbGAEE/Gu0/L2M05NWj5kQSmtPTnc5ffcV2h2wdeSk82la7qWS5q9AIymcpU+h
tuwPUVLUr53hf0In7u16ZuJ8LWPCyzF8sdWKB2RAh4ySwCQE+EHLafOyxI9aeiWoTZ5Fiirtv8F0
j2Io4B9B1Ii3wHAeJr6IMydVxn7RoQ0m13oOIzUOoHJnzA58wQ0uVXuCqGh2w3/7fs3eRZvfyRR6
1MbsPwaW/m64uowdW94/LJ5P7XjS34SlTjbcpgohIgFXAlPgaMu3Zt0lODlbAkdiJzVDctnZEU3t
aV/B6qx8kwNI7of2TZYcOJWnrQr1XHQAk97o6gx0GLG+v9ulXL++LyLM3Mxg+k706Y8/hnTOMfW4
WgYXe/PgXTNfZFlP2TnTGNrOdEBM/guvmTS1FZkbpzIPeJPI/VtlMPmfGPcfkfnNaZbsFOPOsNNw
ndf2ol/GJg5DKim+UHv+LzVxUnWHdYCbXGugI36IHvurVlca2oZDyG6pf6TK27fb/FXk9GPeR6IZ
EpQt5dMSO2dfAEmSI49fqpIdGr0X6+zVpiVYoj3DWDjSecmvdBWEubUVNJikWJ0FGxS1/RX483uu
E3/ySHZ92MoYY42KTUoBxV544EoQJes4K5uqFq2lEBsgHbKCHC+M0OWzNDqqgcj6CghN0dmbqUDy
1UGqVynRPVf+wo7qzQBHmu+voiXtWuGMIKQ7611YGi6h/hBcHugEXc/IOWbvhTEdxfqJ/Vocmq1v
YGHVDww2zH8pKw/OVz/F4lbErQhSh9+vljXoCXHLRfewwLrnyEu5tnpwjT3n23tbdEJw0rPKYsPg
ytEM8nGugdEVky2dfViAG+gd09bK5H0u7fU1GMY/4+ZUxdXeSFCWFNUIjOHNENEX+nbYSAxKUM1e
RQgEWwzb/MImID50WeTaVUg3IiuttvA/LGGYjWsxmVp9nrQAOJbUP04sP25H9SMU/NZz1YJd8Ty0
MrD5dB/gkRzb2kjr5qh1wHzOB0pOe/VVnAmOz/nMmMgSZ/6QWT4GioF3oljYQY1HPqe2QTsRCddW
pbDuKSNC3VelANVEdJr/O4JUA/gbBDCMfYHFsp4N4wuWSuvDf1vSeCiFHH1dHqC8uLrA+veXdYJm
8G91Cc+I7ScBdO6z1+77CoCWXhzAFDghVCsc/hBphKhHhos6sfBuhJI/q+i8cNSjoNQYrnYitWyY
kfQVsN33XVkWYBSVEzwfV/rWSsr++uaYcaa7pnmYKM8/WXIwh/UPKUnC4AzVI6lZtKX/KJpzzQ/9
XECuJNC3KKupAGurk6Ouck4ekyBd2+IOA089E1qvgpWAb62djeYx83Gw7IGBZHoOhlhDU17cm1sW
5ZAKvfe7O6AN7urCzixUESbxNL/1ST3+0erAVF7BsXwVDs3A6G70SadFWVaouyjBQVxbqwqR8DVd
vB9ArzGmUBfzeCL30DPTcBpp5cQsg2q4oNZpdRlNo4ldNTvs/JS9hBG5MvSTTlln7V3m8HpUSkYZ
vU95Krpe2BY7LSxUpZnC/rzp0TmnZBNiU4J7IZCiuQbIp9gRMzMzvkjScMrtHJlcdQ0s2kVHvZgf
XcDuhZeWfOFjUtSoG2OxI3V763Zc7tAxmFlQzlbAVp4GbtA8jf/mPZnt871DhkAJar4zbf3maqOL
0LhHvwhgiMA88OedOciLI7SwOY/HRjLHIl7M+YXLI0ISCfIvQqKC28WAiVf9MiiknQ/ZLELzkss1
rOtVwyfHujNMmzyN7clEfQCu09PgSss0Oy/OBAn1Cb9NK3MdB9Yz0cb6xERR6af5E9TyOhFKOrwA
FMxwwY/bqXw0GEiFInSthPkHkFvshpTTZGbqvAr3UQBTi4GjHNurXKG1sOEbgHi52kX636b78NM4
gsgI5DwM41HWf3ha14w/5bApL55jL+zEtCgzQZF+BnecWSfJh0NdTGEV3/DTGZBGZWTYW5CbhDJe
h54UGGiLNHC5CYgB+HnD87TTOBcKyuHSLG036eamXEQowPA3q+BWnwdaw2YO1uZr9ZAbnZpnouQ2
asLssNB5z+rpIZ3bL7NXS35ZP9TcNzlKRwr75/DiIeX31gbR34ZCYjJWWm67QQ+2if9dbjU0C7Qq
tih9TFbhoYoAmeaeYi5CxoKjSXA3WNV58UWbcD1low9/qBrg9Il/MKiSF0rzECatYonYJXjmlH9R
PsU0rFZyTRkE1KcIMKOObWONdhAXfOhOwoweZhtMBXPbNkMPvk2XMWCLDYyibkp4jJMnL2pb9AFu
kh9TsFiLzYjGHj8NFooaQ5TnR+fHXT9fhVlWYpz/rIa00g0aqi1YhWBsgp565ZtjBVfPzuiSS56E
YW21R0R6Zj2Wo6HDrztIKa9WTX0fh1Oe6rikt3oGeyVj0uTfYPLnBxjokpqgH9g4XCnsXkSExVyp
UUahNX55oIYf4UjoY8moEB5uaIRXyFa3Uag9fjWB+0ToIUZk4CyoLq1gCi64IRT5wkK+wUNoNPWO
L3XEGO0At1G006npIx54GWIOtCk/Ufd7a/q0ntuAScIBDJ6maAwDl0yn3pqYyuiGlI2FvgYlnpvT
zKS1jaTQZ3w+O+tfBJzIZYEQNhk4hiDuG1U1leA9dGGdtFiVz2JfHPrQY9dRSZq8iLl6xltxGAQR
+rAA1NcsDC21wSlJd4htWGVjoN4pMRraWQgY8V20p/XDD/6fwP9gPumsk9XkyRoAM6SsnEjO3h/j
wObulsloRH0fad0C6tX9ePapNAAa4r6vGwiNpfsqGCr1MQaQUiR5d0s4ZxGraBM5XvANcUu+D6Ll
tocFMkMnO5zpCQJyaZoRTieKKEyoSNIl26pKCO2qH/rKAst8M+wCaIMNsgSvQOHWMjuM5e/XgijK
l7nQ1E67YUN3hOhzxQ9KLVL2Yu+a4GtSc5HQDjLBeyOeaX7Tqv+MKwvSWmYrSW6ZEdDsRVI6DgJ7
XmtVAhRbN/izr3oqCdHy/9ArTLZzcBzNEXCbaa0Ui0eJpUdVRWQHHFJcSANGJedfCxbIROYD4baC
MrTTNxwi6qdDjZ0/FWL7ujy44RFHFm3e4kb748m9mH2/Wj8+W9GalLn9WC03xtiKNTMRGseMs2Jy
yEWTaPmcyjjORKqMGQGPPaZcM4hAVQoQWbNk8QVhH+d5HFGDtXdzWHr54K/IQyGcTQxq39JSJXuy
4rL+Uc/92Og++dYtJLNMNmb7TKTKKndKtbh8oPAvBtXIHIrHqY4k61Jftb+uhOMzBTfh5hRIFq2I
mPfgwVP9+M3l7O2T6ooqYWN3mET9F++2gwsQ/rCF8xZJ6lCywxaqypfFtRrtzB2qxj7gHD++B1so
5YxXSCtlVQItPnKGoJrPp2ZhmtEtc3Gqv2VGh36nyQ5yJEmUtRfg/1T40VmsIv2zaLU7GD12opbK
O/Dml+dGzwwQmoFZ0Xp/QS3Kk/cOxsJCUXiF1LMHp4ybVtrJjIvqg3Z1XgDfQWzs7Dk8djYj2kdd
obISZzSWeYgk21yPxeR3+tYpIbmwDNFzifqBghnUd4NNVI1IwbfDWwkIPfMLYgndR5QcEhRuUqTP
rmm+6So65QK3sa/0SA58nRNkAZqTQ2WNNx/60Pdo7Ubthvqw37HqxoEfDL5fzdMDsPfNC0s0CAdN
yd0EWwbQ2Og/aEr9/kKpa8PgpvIeddFTUpfOvhcvwSGZDNRY1qtZbtVw2ikgqfdFOoooIy99rPk9
YpJ5wohTDJRN8EEOOTVXmlySGAR0hwPKf4ZksEUKwcBgrZUCF1O47uPXlJjnE6PjIdXkdXr9t36L
u/HNwh1nQdq+6TFvi67binixBcR6W35pyM3IrAajBWcIvuDQY5ubAG0zIeQm5QZDte91JkjXAlKt
wJZWBo1lQH0gpINVBjxaDiSlmYjd3LZdAnYitl0hwsDRe/lXKAhY3L7jZJrbOOfPyuHzVTLEktFD
aMXtVS7DU1lewORmJgPyDrYiuZN26nnnFsFS8AbKGz2pwpbd/JpA7JTd+6/LZsosdBwcY2CyLL7M
5bNsZLfkSGGBRRjuwjjJYvjhckHZwc1TPUW4MUSpZNOtHiwCdeZ+5fUHO1U6fJnnC0HjXyuZdmO0
B4Z8u/ljQMKC67EgXCK2cAN79IdqrIIawiAsfspPPibCnInSu2RbUd1j9rkWNTxETd43h6tISAcs
lCMUTiY8YOQSbQf7dYYmbRzfZPvbFAfwsTVjjV5vQARwXMOUsrzpHtQL2EUUUEaPUoB9LrCQPLhH
UrruxeKvTteOlZ8tttrIX9y0NExL9ZYKAABFcKKbgm1JUDGWwbgz4xyCr22AxNuE58xPIzvv3krl
ZTEMxcHGuCRswb1nXpajHlkk9DMk7o20DHE8Yaa4HYxAysJvBOFdHEyB5Yupuak9u/7RyN0Qx2H+
8D7EhSxo0HlfIMs3No3DvnD5f2HxxABJ77peE5oeNrh/BHVuvytNai9yH9O84aALfRB3mTJFvygn
lMDStkKjHd2MUPqWrBe9WxAEN4C0lIPqQeem+sOYHd2puJpMlm5VWO7LFdE9kMquMfpbgvL80tsd
d3Pfl43IaZGs8//AsUXXFDr+KJiW9/lnkIfj1Si+NcxIZZvCPwCe0GwiuGouXmrjlBwqOySzmyxH
ZeGKMF759EWx7HrufEyF3AyT0UmKAASUn9UJ5MZGh0lMtnBscOwN6JPAaol0pHP7RlgDPd1WSohx
Re0W6cnRvZ2NGUeEyiJQvFiohZ5MxLUrqz0F/X3bECwNvBeMPtE7DqCYQSSS7WhTfEre9MO8LTOz
m24T/4VnKJ1BBclWKzn8ZHV9/gZAm7Sw+GFnk9yAHjhXDX7ZsBTaYvO2wYWzgu6mjQedpHav8t2e
KPcUw59hb8cRwUP7ExLru+fbb30C5STMtlFV9PS5WVhqi92YoRpbHerplIpf98QecZgoPUnShB6O
xlPoGV2PnKM7VTsMDSQ+GzezmAtOqEMlseU7SMfjdVQg2ENwNh1SmQpeaYuMY/t8RY0i67QgoFAh
7/tifba1ai35ZVl/AgmZH9X1EYBEYwKkdUSK2sJ4kmA0HCFbZLL79mIRxZmCHHvBU4j85bW6lITS
jcMIP/ZL+ueA+2yEMDlu9z8o1PEfc/VHBI5us6UhBC8tNN5Eu3XkFwMxPY3ru13PZLRCw3t+q4mn
/rY+UrlU0zh7gi/OKNMJofYCXTXZKeSfsIkaCiAVBu8LXPTsuFnOIbMlK0H4jONP0UktyUJYTawV
tRDNCiotKBmTWI6OH5qoZe2dPmIiJNqxwR0ITCjkpv+U/jwTRMfI7AUe9fcMWGsUbPvDpDJPmdHy
4pVtlLNILaBRI4YxYi3PWgTKMIKVoRhXbP+iW7wDzl8WUX4s/nFUm1INFlGGTpdwrMRwayaUCL3K
5D9GFiRSOg3YRBijxSpiKIOveN5utt5KFIZhhQzzw4B39lMMWWof04LaKISldVQygJTZIiUTb8ju
qqrSjQTvITzXJbQhMu5UGOk+t5h9TW8RuskxBFjxAmDUsX3Vk2OEwLOFBB6qRj5gF+Zgj5l9nBlI
B0BS/HVzQUz+PCQCCwKp8TZ4NqGs0qsFdkv88UTcb8ypENFOE62VtUyvNptlWTQFCogqtV/go3U/
3s5o4sV2LxLOfk+/HQs9PrYSF+xBf3W1xCJpdIQ3nTZBe446HeTEPE1H50OHYFgfSWs0ZsZkdHVz
RLm+cIEloGmKA6VhNrWg0tusvGvyTjNWNwuhV/ku2n3i7kJvLHU2vvj4r+ck6x3JKW31axJ04LSV
EqpectGuP8Qwp/3X+9/rFXhdJ6EQgpGVs3O8BUnpI1qbZGNvAfevyvmJLlwbwFrURcQ/YK9nNycU
bJecZ54IHjQBABlj3Zlbn3DhJz118ifvQmEu2eiM95MqcSr2wqphrpWjRkfGT+lmGjREgfrRNjLB
H9HBsEvbINstpWNDDr+WmRXTnB63fmA9f+LOtZXRCbB652XnN6koV4jmJvVWIleJukAWYDTsj324
ugZG7sg5ycEmr00DQrwdFBvI1Pfxbb9MQUTOmFMW/BOREiszZMq3dZPi71akR+AsheaaYrC2VRxo
clazHomWk0Y0HTfL0KATl+f319pN0DxaHdkEF0A2pVoa21d7TCCop/lGfd+p0RhbYmSTMQTSKqnv
5tJ6xCFWn9kOAr9FuZC7WXtEkFSXZdw5cTAsYWK36aUIJLAgAKcwgxQX9kCZDcTE9mhLiZcBb1Li
vOFkbvzwcwUv+CEMk1PqXO0cn04J/xtKCeRhjBMYU67F1lodr40/85VbAf45uph/5qBzk/aptsH6
CgweXQxwEqijxw2vQ7v4YkUkmkXV9rGh1RHYTeIrtVTCBirfA+k5V1k1KGB7aoQuqWGMeC5tt/k+
y+EBSj2f3HvHvg2FoVa1r6aLe7SdM8vh8/8ZChVy+SkhHTLVbYy0AU1WDCuLoBzSivNZ5NWlyir3
txpJ1dcCca6PSR/b3WRDyqgb7nLM9GAY0NMiER0qnPEBG20zi4z08qF066bce/GZjH5G6lYrha21
lCVIT39O5QcjF3TjYZ8/Pbs9CDXywuL0a7L1yV8toFCGtpsPsOrF6QZ5tpqMJzA39subiGRz0g2J
6ECaMt5RjbWEOAHgWhryis4n+VBDXQfc6cwlZutK7gtKm8KKK9K08cxxwK/WGitfBmZ3yFobUOjV
hJuJ7elWqwvq0ZS5WC14r3R4158vYqtQiJWFPShSZvpUcq7dWxH5XW3G8zfWF3sqCggbJRqDjy8/
dfN1t6Oj0h/9idYuI4To50nJD1q6X+8aW04gR2vlTBTHxnIeOdgeRyQ6sCt+4RnUavBrjeNm16a/
9oYKhoyxJsPDL9PlhmP83SMW0ueizEmF/GIdpSC4IuNznHWDc0abbwlFkExpBtHcqUQgxqMxevHO
9NpYrdaIszd6J7SFq9EO8MJwTzf4O0+8iF0leXvvc0U3gxaDqrV+wsvUyQqociW7tJMJ/x7HAaYT
fUe9P/mfD4Gdh+1g0XzSpxxhmKUjYFL+mtWj9CGuQRh9qWMuzn5GK3Ozf7Gm4cBv5iHo15yXmfDc
WmL5Wsz2sf3mA+ix7/tuD2la3OFaq7MWNdgzNOwDp/1nDJ5FmLBRkvG5Bz3Fxoe37KF9PXfD9oY7
NWUIbos0VYpHOe5Q4eXCkVzbDtbnhUVlxNvpK43rOo4jcgide550BfnCU+miaZhCkULFtDKIBmzP
HSYDUEB79Gcih5Ivo9/ARG9FJWdAeylotMr8YtqMm2jdDVrAbOT6fcrV7B1OWo5g5d9jTXWJ0ks9
bcJFObI9lt3IuVQpGNkOG+mO3JOBQugvdDlM3RuALjJOBIU5Qe3TCVcHGgTs+qeOMs2bYOQ+VxWK
d6GMeFmCIwNyVBcANIDsBzFpGviLLwPj8GJOlU0Fb0TcDCJ5VMfaf2AM2FTz3L13KVlLwjzPQfCQ
J8yX/DD/vzdGPMz/sfbAdBC8MeM3Oct9NJiRGH7cCiyCYoyXm+7JaBIksrAGFkWdh17bx+8UqvxI
12w07DE7T/io5BY0XxKv0n55Aru1+cIxZOG+DgFwpy5fuqPj+OFX9BFQBji02fITEgtYg9X4b9s7
qN4aN9YwCMH4uMoFZm3KLvsuSoZMmPqquy5qVDKWCVtHi/Lz1mJ6xL/Qex8SJz3zxKqVY7PlkiNX
QdNEoK6bLc5tc8oy+b6sUVfyS3n2Cm5sqFhSvvLuwNumjBh3V95aw24c9HehHh4wVoCzuwZ83DxZ
Myq1qAm+9BdPHuSZmKNP+RE9OkLAgHOAopU27gPfJqyTdHDNrQJnF7HxLgAfyX2Z3R9nL3Z9KHtT
PvfK4k/+oKwicCLUHXYEuyf276Wauk1D56MtznKOmzXlj6K62IIuxUFXCnEhX0U2U3vvQlUH6oUO
oClypNMoIwEHGapCMLRaYpp0Mx8NAn0mfvYzlADYaz7dIwj6zxUUops8E7HKGUJ3j8vaTyST0/T7
yPoV2dtMA0BcePlmVXhyLb9Wxen5cBYpbRaEjZwmKS7P8pkTN27/GvuRlin4hvaEYlLONqqWuGHG
q+Zli1ijxgfCw3DacxjIGSk9rjZdfsYF0ih5sFc36IQcKIqYK/Qr56V2NWN2OGdfbHYcpiFPk0s5
tAKvI40P5iqi/uH0do1Ri11ZnPNjOZau7BkQAQLxGt7SA3cGOXdUvDaEhC+ahYSY/jOaPUr1sUYd
k6XKDInJPRVxT3PJeJHDYoGk9jIcmRgM/PCSCl/ZrccEgHaw1C0SSeZ/KS3U9y4BamDHbgsv0m5d
GAuCMq+Py9BhOzW2s7Jvb64TE1ZFVmmZE/TMOGGVtkeSt3r6J1oJwMXNdYerLcEkClQt5PXpF1ui
Z0LJJ9ApAnfmewG40RpC9+LwS0Fqtk2rUzf9yUrcZvFsXO+DLHuGf8jSjhYkq8vHfK0u3FXLKY9O
N46El4QHsa70Hv3PLOHcq1gLFpqcxWfUpTf6VseTNpL/ZuRwvuKuepRcIlT2nOyJnfkifVKsNMGd
8P+yYNqtknBvWX1PYaJFvsCNWnfIxfqkc6mEJv87vmcZDKDNUwHyNOqm7ARJIMV6c238zgLX89La
FWtcjl4R7+AXL6DGcHFZpmypimPZdfbkwUwbTFxg+NzdJn4z4TPDvYui8qX1h5O3RrWJZpPl08Zj
fqe6baAFNbb2ypXK33wEpK9uY64OQrvDop0q4sFEJdpRivTPZvQbAt3uuYzTH/Wn6ep7BWdwmi1L
j7YOIIIkFlSnQOg7GCAVHyIk/vROC9oSXpRLE8up/5N5YNgn3x82YUsi0Jl9F21ZChDG0xVU2xkO
wEietJ4AQEI9XnNSJpGghxBdNbXXk3o7TXI7R1HDJOPXHWVV5DInf8shyb2uflcyXGrw5zcKJKej
tZPCk0A+RV/tHkSVEawjt0QDHt0uMS9Dv5BFINNPpnQm6rbfcdV4zLaWteVYIcA6CETEwqfFXoxt
VimTp0sCH3h93SK96ofDBErXHDlpr0DZaqdd0eMUIDivW3H00PlOYy5wD9zKEMDNKHM0l9VVNUgh
kAM+EjVFlZk63hoJarDDD9igUxhFTYEbFRTMt1SDNOlXafnl/zEdZ5KrZR/sZmzmfSg7npPeLk8+
Jzs5THiNfceYnkJmPpbOpZBPoEV4epWdBIyg0h+ETQ2dcAWx7EKavCYWqXh7ieSzwy5Viq+eyB3w
xyK4XWc94kthblUgmd3asko/vUwzt3C9TeK78Us0tLddYCiWCnvphpbH7JKlLS7ZEVBJ6wZeOUjy
lBhhHuYviqHQVvRzfLOUyfDrx1oYIvE02kdfP/X2vRvERY5wtUY0wa5eK4VyzfgR/jM6T/UJBB31
Cc5fkYmo5i1hb1hKtmx+SqSUdx1UWQNGOcjNIJYKdUql65OzbGOWc2KlOzVo5XlcUNuzkhbvvQgl
MvtvM88zPdN+LqZ5Aw6O4t/UTGVO+6UK0UNYyQLhP5TMA1m201au2TutuVpLxJm927nKCeCbktis
FcRkCicXPbdOk7GcIikgpX/wjNimvxthdCbs2/J4nHEyGV4DENv2aqoGK2AGH2NggwjJgZAH77fm
rWlw5YgmLSKRAnAlQaKw2pYooSPDuuI5yUM1McbwhTJfHyfPLng2g7HoRFI0K1iPmofnjlflCGJV
phX4LEPHkZJCaBIk7Egp3hyx6b0RrqdBTdxMnjpCkj3we7TVmbCPRitx7u+bTiLdWEizj9xa3H/L
I4gMNCd8TLeuzioPKYFNGC1JtcO3hBSfRCa9ouLp48B0C0tY8NrL4Mf9u1n9rX3G/uFnUaTSyic5
8tvyxaNEK/tp4nh4HdVA0j7TZtSdDq0B4nVxZpkiurkUab7oo59f3SP8VUSGvTkVoGYFJQ9UdPBo
tDjUIfzNuypq0m1mOMR9D9GLvL/BOeA1PhbXRZffL1RfSnxwkbgZSvJA0DB4vDpEaQ9bIRls476r
TpLE+KymQYgsBKbZGXVHRpdf8Qcf1sAe+6jwuvhK4UVIu3+7BFtALRJtpvIjNBcX7yPyD8Xqpn7S
iHEti7e+5eF70FJpoiKTsTLDxPe7dPWXrntZx42bB0sXhloVdFvwrvUJeulvhhvyhf5ILKHhHePz
3aAZv3UjBTIi0PS55kcsVh8LH5Mqi6m/WUCIeUdJ0HrVrs4sOod0lQuzgHhrmm8NqueXOElhYPMS
dx9aAql2GasZ2anSlye/KwmdM63X+4giwQooXGzORH9bjXapX0w/V/iKAgBJwTnkqhmwZXffzDLc
E6n0YWuZsriNulakwPWnDL4A/RpKZvdmPF8YhwnaWTNp1uPQ4DSahC6Dboi/wCk7cu+X2MJZgV8e
gFwtReU7Uj5KtGYmN3/hcPJHL+a7eubp9uezUME0OZPSW+vvqvA7JrlbWSFPUH9RWj6hNC2YotiX
jYRjZRERnz9S0pmm9CLjiOGEzHQ3Q3srkqErrsLHOvBL8wyhvWBXKA4vw7k36Dquq2I9PIYMAt2J
kMgNP5lT3QxoLADySYaUClfJCjoWD7fstMBRvCuSp5t5JAU9ECQR1RyGIuJel0MA6+L8E9y5KZAH
9EEKxkUqbUc1t/LpZGz3LPkamPtXZAHzEORDmBTrNYF77rdlFh62XNddj7MYRCO7BpFnUJ0iOSRO
2lRzGeddG51MYQmHLzMZMHoKFZ5nZIhVROVV0CrCFnZGnEskI9UkQBHfNlVzBflMvitG2NJUW800
uo0FxMEiGJFuhXpDkRMJYzCXy2v7RjMwu/FsAtONJRQWHFhzvhiiLuqEUVNu4MocSl1pDV0NGU48
LSIgyVlivREqN//5M0nUgek0UWplC4AyjniB+ZtrHc8WB2LtPPHOv5Wp3uOKrfR10cLiM2nzENuV
LuBRQaA4sI+9mEVRgLuWUWQQKlL+zTfVc+Xp1eiYrl0vTR38Vaex3X7wZvCUs8GxZhdWrNHiC9gh
hFvPnUuHoEwlh+LJLtzs33rhMCh0pn+NUOt2fvz1mshF0dpMH13opo0tcDtvsRueZgnzNtqQJpZc
fUPfqCMy6CvOlrQwMaP7vDIkSQn6/b8UyYv1qOlPOavKLieiqxl9NH5ZzD4tCP1/UsRrQ7iAzfGF
fGwEYJksYBa7KZ/4UNlGju1vO89A9fP44NHM1+RmUNKMw5NWUzMQXUlmTfyzTLbuckwS/iQAQ+iO
WS0QjY3JWzBSHVwogEwPsUR05aafObniamQA0oFsQituVEMGB85GBfN0IfrN95YYzzYyM0br7iqd
y/kqQhRH+3OTsHYT3n2KVfAJkaSV0oqfrCbKKXspYe4l+UASskezJQglUEck6IX0pIOZCttpMEem
ejGhhE0TIjo24WoeaoMx3rEAKVtWlqjXJiNcYJ/3uJyUu3+W3Beeu9sBxUfRy+MgBk36/Frvuh0t
qKxGRYdySmjvlPAbyNlDceEXo+314UAsNhT5FhNN+rfXHJTUlF0KewOCPlQ47gMEYh5SrWlrtNJb
vcpL3gmhmWT88VR+wl55UaeZTRFfUGN7/kTLV4OyrdMyNgJmtn00+R5bP4bwBg/oJo6W782AGwzq
OzALQ4xwo+TrN8xnekLWpW5mlCXoBq4uehTUnJ6YmMBLgtdb906l8ShYpnXeM9mmikP6eOmNsWpT
8UGwhv9MJKUs5I8q+FQPyERFbX3V3WVBHR5D2vWiHCBd0sSZLoqHAJFe5ssRp0zXxfsjfj+n6vj4
unl4K99I14zEds4ZRY7yc0TUmm1sJRSu/uJPDz7ax1MK+eblUt/2nH66wQrFvFoatEjiYO7vsulJ
e/Bvg8gsps3A2cGadZFqxbPvyq1MvQqObIs7sF+ApfjjQtmt5wNDfbg88nviP5QKmCQOn/Z8jhX3
p05b9b20JaIi5nTD2NiZIAyh+BkM+DG+FUKdj7wf41/9ercob/LI5D/oc/wJI+6euhdzvNYTWexP
L+V4Cv0wiWnJpdqYbfTdpiRaiAz2QkXyC38BcZw59+Y9sqHVV0ysSSKdrUg1PH1xc12zAOzArIsc
kbrR7bO6e2kkpvH1c8caMgPkYGxISvBFaijDREVWErMG6IQUfsxfcJjpFDWnA/1ArIQY0tPKlv8X
6f7gEN7XSRDmYCvELD8QwHAEdaIoYj5heYXfhKViixVE1wWMAMI9TOnXvv1geGY180ltWwqzOaXA
yTYNgyXegf+oFTN9+4M8dluIr8nYkp7c/GS9GMHiPOoKUaHo1hf6ZjFIsb1zEL13H2vFhD8/Z1I5
DFs1jjBgxi60n7niY5IEOXcpO8h/VjNto5LoEAJjHyBGfLpa+WrVBDB9VksgGrygFcE+/ebUvhMm
Zc1U2amm+qy6HnfRbj52jspdLI6ELmhlyd8x2FaLxaA4Dh+g54jMeJELCgGXooZN5EQMb/xMw2KO
29F+D8B38b/WsOnIZRSXl7+MGYJpUla1ofB36mfoo94oYDJYNFTJobhPtLCDdwFnrSmi5E5Ru9ys
6R/vtAnOK8MdbGTo9guB7dZ4A6k2VGZR+0LePI47wZMlIRArZ8a7ZIEdYjvSx1CZ410LN5S+Wmq3
+GM+tlYVPjXX3g/B1fSagt8SGytRAwgZ9HKI33Bf+HB+EKzXVpsyDuoXyG52RJSZzz+XM/FP9ljc
i6644r0K6djJwR0GwlTivhSzgTTj5kpZyeXgj0gOQU4AwzuGWt7GF/dr9Cl3isNnITr/3bilV3NA
vRnN4GSyZNBihziuqQMAH4iBVwo6uU9LcYcDX/80ax4yIi6ZMEXdmsYjW4lTM+mh66Gv1VftLgWf
4n5Pz7sIq5a/wiV4kOiAeZqvObuxDVNXu5IwMnv4BKEvOwWdkkfttorspQyzpbd4cm388KxBPugL
wg0x5+HluamkW0MwG1c/w/8AIRFVLnga4u1TUUTrtrTqWg/3JhB+ra3cCRjidlH+ll5c4AwOWq7l
wca+fBUClKXS58QSQPrq8mugF2ZaBHEog/rgb4Y71nNZd0V29GxcbnYjjkFMkIe0kTGO7PVi/5vC
6UzUcC4D9oEw9N2dSpn6wZILVPEYoUUerj7EGcGFfDzIcosuyVWEHhraeC8983bvwj+YD8Lb9DcJ
bNJfUo/CxtVmVX5x9UcNbsawDEEGZasWV1n4YvvJlceiP45ywJuLiMslUE8P0O0HSkcf0L6my1C4
FOfkgVhFFzAq3iva4a1jeOpgwqMGOmDnoXPkGfC9OqazpmpYvyYuHQIrF/xcfnsWZ3EZi9SAM6zR
/CnltDHgt4KjOPiubfZHDgPWh7EwT/ZBuzJR5CWkjIHGknJt5Ha9wEd/wzOgc474FEVxMePBmGqb
HxEXjFD1T5TXmUp20itulf/aqG3W2najz9Sq2xJZhfv9HHsD4L6wOd9vJipp6U9kL3gC5gT0W+K1
K2oUP7Nlt4+N0mRAiW6vaoOvTXLx9t9N2LPnxr8R2wtaNztgGOPCrmTNyvs7/sRxgBxnWFo1Nfw8
jxb8A/4+q73M64B2wrl0Giina4U/OWHYvU9PYQBItt6sAze1EAPt6BhSzGxhC0Pt1VZjhowVBBES
DOG/Kj+Tv1PHsnFWEWkyh6vrI8GebXUViWKBPOUKsy4KyQWKQzNRFEJcHwyUT/dAG1AzKPC/KMZq
ONXl6mtl97n3j2btVhURJTwQP7J01SW01JtZz9JrOkeCCpsnHxoXoSpRhl1cgNGzkpJ8Wjxqj+dl
ljJvL4FSWLkL0Y1MQLmKfPsr/+cT9JfniMQJg9iMusXC+Qycoei2SZ3MLssGI9LbiuUNVV62fJeR
Pb54P/t1JaYA3PQYSGzr5kw3l1I8WpNgU+FFAyDRGno9aVWjTNc49uyu8er44I8nYcAmbTEXNWLv
WdGIkIA3Q6UMDg5+QsWDrj7MW4IsHxNToen2Y/chSDdx+6JhN/hDoc6GehxPlQANKW5/MYgBBNks
Prs0tAFRcGcJtVG+bRyjsln5RdZpsyOUBDPzxpmowZV71oGg652ofa3r+hK0CFp8EwL/u3YmWZTg
swBbvXksJCBBctzUARSWw4X3CxZ9bxTllgENXDPtvSwV9jV1t6JGSt1D0fMS5LfMPBmGC/HbQ50K
ZrYiMs06VhHKrZMxkgQONcIRTITpxUqqmR0hNQcz8bhFt7jjDdaoFZSiayXq3dIHiUw1KpanbmqW
QrqNaAivYTZGeqgC0ol4YAfXwJYeMdVLM08Gvd0X9geXQj64BeDMc4dhJcNZnHAQ6c0kmhmwRsH0
kqzXU6B8dbk2j6mGn+BexdVVAPBCxWauCoupCkTwI9l8UcvFIr5NIsW+5iK4Lpo6wChYEHuqOK+E
UKkVuzXcjxKBqHNjWII3t/wGme+vMEFsswzRc7aTtFRnxWUkc4eQUqZKw+I8WIidG9KcauhXKo2v
xmKNUSkOgBCuo7NOIvqIwx92MPK3Jk70wrIHF9UxifxfhebxJtiW8KbrvvCnkZ+NT5rsEyoz1ve5
4din2BqZI5/YiY84xqKMQQYLtdcHm5PSkQCa2bDPWK5gswKw/cwHODH8B93S6gC8RjjAzTMt4UHV
P4QV8Z+/QO3Tx6nHFp25tJC7Ith4wSgqSMyC4OcSCVaSMkQk3ilyUiouBSBxCglHN3gcK5kZ5bjm
ehxa9pnJG7JWAI04aLnTa37bzvnRRFDrMAqs2SQqcd4A8r0WAGwQFmv55wEdWmLSehPYht6hhcP0
CdR6brDlfU4BE1/nRlRbLFSedk4VvLFOB9UVOpxk75NoHoMo+mQe2zDZ+qfY6vtLXTEgzQy8FQqA
nw3C7m9AgJIgzgqxnvjTCMgiMbrmOluWCBEaxUXn5H1vI59ZnysFNLKS2PORAbo5R0XPmUPjSoUJ
kCn+oz1bwD1yyT2+ey2GabYOuId0Pr/bY6Z/ziI7aZHupZVy1zRonD3S/NS0GZQgPybG11w1vzKL
oJwb/KUFgK6uJa6yqv4MVCe/bGUHs2E+DiFK/BuYsl6yaaakS1T6brmVY3cuD72NXWCrJ9hc5Dk2
sNTx/uV7X2N25WyBLGMOZuZm79TgRMgFYtJwkctY+XsesKu6EZp7vXWUPaX2zBEmRUul7/4LWQYL
qBBPdTAjziE2b0JrUfqObtRH25gw1ZWazfWywuzKas+Ug5zO4Obm5WqNfxUFogO0uXIyDczQKjuz
maHZ+/jlNme2yfE+MivlBQ3SZh8k805173sN27ZCOVOnKD7s5fun4mVqCBpj5pjhLWJf4ubw9tOd
mThPbkNvWnfJb7Q3sQNYP1fJABucwyRpF9os2ad9m70/nrVmmsNUoyJP1QOfqXk3agwWfrlmCSzb
gueNeYbZVeid0WJXTfHhr097bdnM1FOUe1sd0fQtYphme9bO4t0qffErW30yhuj4jyfQDFYUwYwu
dHckIAnw0s22glENE7wDi2jT6hTkakS8MPi5qIk68i0a7hvxhOpLZJ5x4444mgwHq5CBhYvrY3r/
9hugVt/f6tbIZ4uAHnL5SZko7yPaCJzFuDuKwjpi2oNw6K2raZ8TiWB4SzKfQrH/3bYZN2+bTpgP
upfdzC9h5nERzbMTAhuJUvBnynAxkQmdSOhygVP4pzUS6iE5WcHcIV+S6T3INSPwjKoWl79PtTvK
QxjOeGmwXKKHxBY+1PLxeYTlGqc0oj0HUMioKyxExfuDVOKAvYDhY55rBrf6QcmqzGZnriTk1Ai+
VZAVcMSfARs69LApadn6iATjXhucczPeQrcZjShPhrfHPUfvj1F0upbEssjQjkYHXjOEgcmFcfsn
FIyspjqO6jQgIy/0B7yHicXseASx6q7RPLreaEVbl3sGaPYYEZk4zKv/+gNYz4B734Ch0jtrjlkR
rbKN8O3ljQ18cVWXDmgGsEyJ1QD1rjbvNWxLNXCz3i5UZhG3UJC3FovROi9QjeILepoxrxXve3WW
HA23pfEquWCFFq5a8mxyTdakvI3qrxov3BUtpAktWttRfkPcIGmR/Ys5/DibloZv+dp0N8LymYeG
cZIbCv+O5g74jiBIprWTMYoz0tpmJw4MjeqC9S4dPmrG+P1EPRDqPu0BSCADodyV8mjXIWQzcgME
/kNw44EM1Rd1NgpcmXYXcJRtsh7jZCOf4mJ+/XvRv3fzC139eaoHhs/goyiMypH/4iqPQqOmQ9yz
Tm4BHFnxqy3/T7t/QWSvyTxecwSd3AUfoRITLkgELpZK3giF5fdK5xIoqFWZ3dcpg/Mm9rlwM6nr
zhFcz8tGw/3Wpm2o5AYysNtd47yTArilPcJGtHJ2+4AO6/kBcsbYvyRXTlVAh2vUI3X+kS2MHJ5r
IPO4F8X3a7Cl4VkIkYdTnPmOsGQ+hVtYeBXZCHnW5dSWytti7RWHpY3SkH7KQjC4dJKVpmUj1ZDK
taFm2SfxZR8tl9KboLlzb+1dTx52pCa/B6D1NM2rNt36wGHanmml95eL4jFjJzoCPXPmfEkDnGZq
i+1vPv9b+wuXM6Pw2cg7QAJfNTrjWhQ3ReOxeW5Yc1FpjKg52YubwMAI5uLWfT8aHXIOctEfLz96
dE1cHzZhlB7S8uR6fUs5ISKxD4ivsAbKQUnVbAke6Tv+MsQuYCWwffVQM7N7qm2zpNKh+B3fcjdL
MenaFaiUBP0/XffX8cwSTyXfvKZ1oU0QUyno5QOrn2hbzGGtymSaME0I0x3XVuvA3zqkCuq0T0bh
ta2ZSBhNRdrkeU5Blshnba/l3aDtVHVKY3p3atAewMItT1nfyPSdeUFH/fq3sW6EG9nI1GdH4vQT
BMoY8rHShm89eeB0Dud655Ib0yaQh43jYQ7GbqwN8K043ykHSf1P4N07Y1xdOseu4JQWK3EwkNfA
WSdBagHFEpRHF74otIDF4YfNPBjULjvpx8N/jGF39HXbfbjov4nDFWhnDVL11ZDdFjRZ21r02qGT
x1UJzNfxI4VnWKdQ1DEGg9IrDT0TOxCCSNzvP3QAqFAvn2iOFkx/D0kkcbsA793ewPe+PJC5GcUa
H888KUigx6TvMqqrzHn9AMDqC/47nNUilQVeW+R+smbkDgcTYcKoiIdEE3H02Xq3xgXnjmjxcgIY
2zS2+GZBlDTtkHIvUc2egzhkIc0BnJS/6mzWKkrlmPs/w69Xtok+G8YvM2s5eE5gEKXuBwKydEKK
QrfXYVZUU48ErKSt4hsgkJabaKIZR+OTPrjaL78F/68my6mtG0n4amVhkdPPy9fpVXBe0q7RTmbW
6aR8/uc/cY4+AChQwY0EbGPU7JCET4dgQxz0QxFGMAZOyTaV8QbUdMcP2WjOe8hqn5pdCDnvPLcd
UvcsFsxLxYCa9uCgz/POOcWuxIbSkxB5XGXHAPbyoCKPNU3nPJJlIPjRMyK9etozaeIUP/qJuqmm
jwGLxngbq+anlfvr0Zl2nvjC6+p3qKmh1hq8okVtLIvlrzm+HKcYiJ+IuyWCG4EmsrWLr8cILUew
RSqqQFas/3rno6jj8X+VXxI/Xkka/824BTurxXj3yWzIp6GqZTMILX/Hyrr5XE2XdO+FLUgG7dR3
wQbPBERjvN/6D0pTAtlXADvuh2UbI6/FArbGZiC0p06PZRgmjJYreGUTSPzDAlbVCSOV6eY+Xjnl
HMHPk8aGgFUIi7apA/x7DRBJ6FwWj5IMI58u2CIdvt8oktZT15HOU2OxkrxVXdgmFLjMUMf0phnf
8tWn9wTvKRfZ3Nx2UoMwCJR1Pvpf8w/jlZkZXDSN033q+gQqsA1Dmk/KliO1ZsfZkFY4HVP615XI
lT5xeR/7sXywlxwFruPI2pgoKzbJ6D5r+4JHzinfDLGl2prX18Jx2N3Fr17Yeh9dTBSIC7hjKeUu
Bw7jEgYQ3RJOv07sF/wAH0XorqFSr+Nba/2djuiuELzVe4Advb8o4yofTrE6J5CZLRi7NAKG1SFI
8qO6GT44ph+0i86OXMafEzQZaYiBBUc6CR7zPL4hTGhUMhPV7T6aiskcz1eKwWB/RZSKLSyPw4q8
jRgHfAo8+SfQLoqIOrpqeNQGJyKC8BHvrTYIrYtAiltTzLkhmKhkIixewrbrxXCe8gU0YAEWELaN
7zOMtubrAPrsPyPEpwjDMOop4VfOK/A2ACHdSsb/TIn+RPtA2acysfdQNWVorURqClgrZqKE7TvG
u7MZ9VhBU9uLZEnUZxTbrRxebTZQ1sd3MojG9abTgyueLCD565DZd5SGcn3vXsE6yS1ksxjip6f6
kr3J2DxU0nHfpUqlOy/vYMbNPPEJGaYP/CdtS3+bB71peAZvWfP+zNz4vGB6DZx98bUwEttM4y5m
kLuKbwQ1QzGqCmm6yf0R8TLDGrcRhK/hfI732Jcsnc275k/N3R9SFHh3PdWbb0DKV4jhNPe3c/AO
bN3p4lM6eO6fYHk/zDzFhQWOZzCLupJhFWAZJ6/hrF7sauHkKR2VmmMDCp0oAsoRvS9ezuUNdYFH
q65Ro2souO/TAhnQN2+IY0l4Rb+0xakKsKxkkc3R/m57SEui6v+5EHbe+10j8YljMUeSOVnh+Z+4
9OCUOIHEnX8imseiPJRrbiVbItRSQmvzqVLYsijwQg0+W6OqJhaNY7uoDaoEZpkvx/NmjiQE/z+u
DXMFHS5swZFEOp2KgVTfKyqHB4iCJFQngN3CkbZD8CsO+ry2jGF7C3DcQOZKQz1aiVtYSugTeRC+
OlGWAfPGmRXEETvSf2NsLgVSGLSmemXsXHheEuQwMhUu7pVspNZwhmLniLb8nVTA+Weac3lC2eHl
Z8OnWwMIfn5QgnYz6Ky6IdRR7c8a3cHgoIdvKFykXW+z/vU7lkKx0F6yzhWe73+BvICTszxbsr0r
0W4G2pOdkOuKthkz7yJEkYJD1eTagWj8JNMJrb3szGs2O3X1AkR0cUp92t9fCy1VsYib4dZA19pQ
mmXcQa4Ipk4LVIDTr4VTY+vjw3Tw9nFAMwUhbINxQI+CESlffBwBSvtHq3CiXfUGm/24wtS697zh
sDpwdRSoJeGAT9xd2Sp4H+mTfndJIR+WmOrp2Zhbxl65c77ApffzoNfINf6/soWjwhKjc5Q0uM72
GDl43VIdVt6dyWlIRPI0I9Yu3pIqtV5POnK/DZHmLfsa14i281Wg7yGRSqS4kwaiNokMp4tIQtUs
gm50MTurQv5SzKOlxFf7l0uwh2G3ua89aJaP5aH0QSr+bJzjLjmiuwF4ah+33ogAhMLC90zDuySe
+KeaaH24LyG01dgPlhuOVzrF1XX9web1P3VlIDAhcmlsRmA4o7iVRsbbjvluIoEXR0euExvxWQxS
kzQk1VzV0Zi6GSZS+wGcnoSk7r+AsgzSADefLJLGX8UGD1x/OwLSTzvhbhNHcz3h/4N3D2yTdD1U
WcTmODVcNkHGkAph5StidW2ulmLKpRrL12ph9u3MIQMV/CRU+wzD6khiTdcvxio2ZNjpP7m2tsu8
cQXHk3qxRxYZAeppsGwgxsjCDvPmpMeV+rgjfk4MSY69JRN5+vsbsrIeVwyxb6kA+lUnbKnlAXq+
UlUFzCKAjKxeHxg05sqLmXMACefDmiQQTLSCxHVR/JLflg1JZjqL4pAHA5e87fUa9eXkQ1+wKtrG
TqNK2C7XQj6lC26WPEDePvvf+b90h2RGr5bblwQ+Oxy5v/9kWHmOc88kqc1EbUjcI/X+wWvXLAOf
9APVEZilyB7bzEnin0Tt67EjtMOA62WzLFaRlXIL+wCX6xLCm7s1HZDmbBvEq1tzqbVQqiDKE7z1
dMp3c5+0OT1yZytcl5DHAPxt7dlvmcNkdlNTc5zcS3pZlYcBzQ+0PQ4YeajWRFOhATnyLaav0As1
uW0B7MRCfZcCBPLOOkftngDoJaJvWih04yebb7jajz/kk9hk363oVOD6R+ipDZEF2vLGkBh3Tab6
cD0j+Z6Dyk9AC7AuAIXlBGrMo19v5AYAdmnCZCebXCmRllXoMaIxz9rzXqMOeqJzey4J+QfrjKs9
WFKmBG2NLFSy/2GhWMMJuDBKnevoxZAVr0ZtIH7ncYb1lRYTKRUaV/JT3eI65B1dgmi0BBoLF8Yc
JYZcgH15vuARM7HdP5pNs4IBo0i2Zoq8oF5pdPGr2dJ/A9O9+s2zJWdxJ5DeWUUY+67Z7E68qfC/
uOTcOkWxipx4mxCjRJmflfngsulGonPowgqGjRiuKAaXOhPlCwPLwKqN5Ex6aQPOqfx8jncGET5q
J7p2LA/EZkFHsCNS8ZszgDHhwymJaHG0bpkCQDqHAwSPWUTgT0NG/5x9e3Bs4+mDj6XEjOMZSV6B
yB4cV8uWagC6rRMV88ygNpnPrc5fq4PGaOAYI/eC7oFNC1VNuPJWDRsZET4ZAxtziTltIEYl05wL
UluiWUGQlDZFoxtr9WX6ljvtMDYRn7ink7f+bidkVZi+SxEFZmDbfjM7OwkVZT9KjWfTkwrPM0+T
/ITygWHl/Ld8e7UoHLCPlNEPkabvzPlGA2v+nIll4HFZCkfHy088FZncum/4rhewLL573mgc3x9E
Mz5o82g4bfufqFNGAqG3sqccZhlH/aAERkq61pu5ISysrvJCTqmGDN+EOGNZOZYWy32XP7lUilnY
pqHKBdcp/t/dn/tyip2fyKpE3MXxsbFF5VdWXalNjsDvpYBfKFVu8HiJKVFuAy5khpq1SfgKts2k
ESdUSh7kuOZj3wKq6yMidQUTpzjRS8sLz2bJkxj2pwkQEssYJebnmrAxcfw0kZ6ZeQraU3wbSXbZ
lorg1TzsaDM5RyAddHun4HHFy1/tGAhTiKjL+oLmB/pMir/bO+xtFq+WY/47sGZa0rSFYIOUtCmj
fqbF3CN1BN56/uIHSmJoPEtUxcboowj2bmtxYfImF4bpCLSoX8bQ5U0RdAHI9tbuqk0idvF0CMi3
phaAM0J8VnP3bXJLtNUXKb7HDhNxMkDTLQdbWts8E2Bx5zW/n2zeLOrhLucTWxchMf217txiOC5A
aiDl2t2Tz0Jf3BOg2c+kchtuk0VbFztgC8dIL0qo6z9FvgxfkIzkTa1OmuZBHubK3z9oL/XNgcLS
ofoiZ2zGZJOr5tEAbkViqc5GUneMuAylKVhYqHpkNtKfxb8ZzYK0TCaKBlSANw/LOBJde3v0ziuw
7Af6e905Recx6AKKSBHFXurDOwSjkVYKpP/HyYpdvdSY9rVmM6htrXA7zHXz7j23A9ZMFOt0RqYQ
QNH1LvgY4c4RJtDP14zox0plqb4yKHoAVdVG6+TyAAoQiKq4VgfaNS4PGLMcVr5CAcU0zDefOTjG
Vj3CAog/mFDVlwyLZzBjeEkKPUKavxONMv4hKUejieZFI08WzOV0VlBBPLimCnkO3RezSY7gFCGa
6cFWAc5nvavIpeqUFsNEio/pOM93S4PSpfilKnTwzGNnb44XL0+jv1Kp61hf4ijUWG5xwupNzGLY
hNppgJUpIy7S79lpcuO6oguYZz1urpytTEF6b8iHkAz9S+zmcZdMzKDVsvLchD44t/R1qpP+QsKX
9s9EKMFv2Nscwu7FCt5Ti20P3EZyLGwlls76mCSCS8hC2G3noIl/tZVzNT83nqDxO9SsMplaGABS
qhtqooNv9x4EI390FQ6TsWuG9d6OOmXTEDs4UV/o4g+9fYHNKnCM3AfNfwNMfnRZHcyAMXp5qQB0
b8poDiL2pV25blIAcRYJxdVYIaKg2PQXnwOOKJzsJKh8UvRwx0dEjHbD6DCZ6uPycTewNORLH1fY
deOfqVaQAv9h7lnYQCnIFWd6kGr1X+D8U5VSyTsynE7px7G+II8HHhAsQ7YiZib3/VOvdXHl//Kb
ya4fUlKg/b7UutEaZhOJXa7xKo7y9T1mbyfNV+5sLB3ExSVd6frfy1Ih/K9AZGTxu1U+GVYd8baT
oTMpO2w//OwlKTwtMs4WpvtZKTcK+H4xcunbEZJDswadePhvOmREbqk3jeNEKa+KETZug6g47aLk
XBFq2y0EtN91l46/NDU/3frNKSNfDGwDQ2uqqyhAQAUXhu00By0L0kuKnE6HiNQ3HRTYDF19LTYv
e17pzL1onqkH0t8KPnZYWOWJUHPQHhFvnX3M6iqIhkIKOT1jrBcpzMop2BcVqXBMEi/4PfH0cv89
rQxPlImAgsH7vOw/BnBbTZb1UMIB15OPaVa0RKgzcoUialNnNgZochrtK/ZIWNxebkh/T7HBCsj1
eCb0mxfixLww1PbOUKPCpOGrBLuDu6DR5WKT9W0RoeDlIPYWKEPLCOJ6/YgYnK05zQWjCFDzM19G
aV2by7FwspTB98+W+j/RSInf+l48f8icmcWLk97z5dFceZZXjQqHMoTOWeyFRuSfaRBDZ3HQS3YI
B2/Wnm4v1ng+wgEYAxknnu8zFpk86fKnkj/VgvUE7x9J5koBRI2642T21ngLg149Yp39qD/cRz9I
8YDBFXyWxSye6US/NF45KsoNqi+vEkMRNJdpArDKpMbyxZm50QEehw5m70wJdzfReWJbJKVPxQ5A
5zOg1KW9z3htXbRvUT4e2EcSPo0Y8z4XhkQmqBj1jAOI50cfRP0LodDtHfBQf0Vrc6ioAhMImhPg
5I0ga7vBM7Yhta74Naz6Mj0bhz1pueNK+XotYdVTzBiB7l4q7eZFKxrycLHwaxX9Od5+Ouc0nCbi
8Zolp5b/qA5q/EpaLtxM1lWtE+JjyHp+SZmLetiatj02WdnN1JRMaWJjSwrZR5E6GTSLyyHtWE/+
XWPrTEDuHPoCRWp1pa6A1eRYq58W2V+3696e4naAxnzz/4nqy82VvC3DkDB79wFGDmzHXAvBkUNE
sc3ehiAGVbET6ZwvJC9zXtjXoUobSpJiAL3XQv2MWtEeFPIisuAUXDsQXbfn+vV5RDncrnSn/cry
PhDMif73VNm4JXn/olGFV58YjWM+CcKx7ob42B6vgba1qsvTmb9Buq5jt8uefM+ejQw1TqH0YIUX
W4NUyP90xoMGEK6pOMytWNuaRoLROyVwjE47zVQ92LyvYJgvFL+DvaU4GU07BA96r3wZRvSDkakM
66M5XEt7sX5VwXLzyt8bCQWme5b4J0IMGAloS7+lfzmu2W6HtvPcswfw+ze6pPO2F3nJsGXafTsK
yg46NEqT2MzCCp/U+cPakD8EUNaoJQI9g9d8mn3Zw0dPHmylrkZY8disksmVc6qi2fYVm4cLc3Yc
2L2PrlaIpOO3IB+oNGzoLtiKBjV/EUH6FwccquiX3mm9alh3PvJGJFyqztpXTVcKV7meRSrdliC6
Rb/BZ2DD7DnoCpD/aynQDlsrON+AagEZ55wJcxp10oE/U1Gu8tKC1jx+7J3W5W7Smh3wtAhcQtbJ
+15QsdYKeOVvajwHMyCRUdnJmaKJYxan1TqiLZoe8jQw46DuD0YDMj1QwpYHsAfV0ENT4JnYM7PI
YHigLciw6KySL87pOcf7abiMXXoGyDH1oXViIkkx2BpB8Hrijo90WanBCbE04QOjR35K5CzQ5mnl
LklChmFcKP2PztKVDeUIegusX8lXM7vZShfjjKlNwqyQ5hu/sm9C/YSUA1PXVvGnVBSTj6cEnSfu
Rf0QBWgL94lhevxS/siTPty60LLX0pgTEiU+sfiWE666gRzzJ/o5B7s4znM1UYtTZJVXOgWsYgU+
LDmmB9C5NPKl+LtIhvI6gyqsOJWnRS9rZ/PqIPBfLqxlMM/dmdSdl1lT7PLU9FrXxSVO81MxkKjR
3o7/XUBG5DsAvDpZ+jtsgSXccsj+8jTvybtit8VhzHvJidFbnn3YuFSc2M/i1AtnIf7KEiyGP2Ga
eSspp05beeuPhKIrtmGvzQyyxQX8hvfDtlfV2lIJx3Cq4cgLjip/Efl+V9r8y7/MmdF4P0xFK9kK
FJjkPA35J+Cd4Pl0y+5D5kZqCB5hyk0CHJN7GStF7XpyUA+PtkwGyf72lyOPIoZejsRELvqazTK+
3gIvAhvZo8kR2pcDGmm7QLusKPemyRSvg/UVhHUq2lpNoXBY7IZrKbfNQ51wyNe30dCYjk7zq9wj
kMC4cCEuY1GhX0v+0zubSZPCaVuTNMEFBqEo/IYYMv1yp3TKNsSI4q7UoecpdA8ZZ1x57cT6/YWU
s5/ZWLSs9oMr5001RkVab1xELHWq/WAwnO42JRyJqZaKaIL2BW9x6iTgSAbMBvZ2kFK5Fsnk3qD3
OYFL5CuLbZGSGJqzHMS4uE0w4NV9JMjZ+qBlq5Kvtitar7MM3Hk6L01anxOx+fi6ZgulxOPFMI+e
dWL0qe5nszudGoktoWKaHdVbstXKFI1aIZ20VV+mLwguHMvfXdrJq8SgUwnRZIrmqGKBI0JuWb4f
ukKBpi9PcqUeWyvRlf3Zld/Qtd3IO51zYdQX9fmuZFgQMJSnmPtIq3zNR78zN2klFi73G7z0LTSs
Kc8NMqiB6jbbnAbRIHw/rtm29nTtFZkzYEhjLJmDY2XjMCcTug9oBFQ3w9VykyvWIM+ju+IDQw9J
PghMbUgwoupuvGK6uMHm5PkGFEE9tZVTvAaROr/ljQk01FRl+35NSCqWc0I3IrnKSO4zspWw8jgG
DBjyDqjTaAFgi5GUB6Q6ig2lF2VyIW/ZFrJNKSGsqXa/MlqRJ8ACSDbCip61LoyrHwqZsrKX1GH6
XmqqoFiDeiIK+yRpn5rM+phh3JcJ+vEB/McqBZMNP0CjSN4i049mLAKqZV6c/Gv50CncqSii7nYv
mM+sGZOpZoQdL+YJlndhAmRhHbYnFFz0RMTLK9NilfaPLCNXoyJze4es3lRtpdMKJWwamqWcIBBP
7tEbtiotFN+ehv/gf/1jO1uK5QksXYfGSOD9Xa7zx/GE0uvTWImbrYEjh4uC8x8zHp02D+zHsvrR
VRSiemBbuSv2wg7nuQpGZW6g63ATSa5+LTfGXzrjzo5nqHq1A67NDmSV6s424ZdFfw8VtqxSn0a1
DJl97Q3pLSwTUyQsv1o5BXyb/9jvOXDOxTbU9cOjJ6syP0QFJbWt4fRf9keUy7P5ziV7xsRiySyk
z1P0llIDwjE3m5FGeWKRajfv0+b2z4oL5ZHhrvqREmVi013XgGiRQ/9XaWDcdozyFfE/Awt/ibVh
GTPWk2mxYsBIAcdj47QncTATk0mnZWTe4br2PtTcsNM+XPniMAtCDM7L6IomyB3D62O+5YJaaaW9
Cc8TBDtL9VTZKk/qMPaUEd8iI9pWzTekgYXj+MQixccuAgn2vDRsgO38GxdGISZZypDInzsfCaxr
0ynydSODA7HSJQno2mzLxbcYCViKeFYQT31D17EfFSq1uQ/RXNwWWSucDU7O5Xyf8pUMDesVPhgd
YFSa8gCtrvOHdCtlAw6QcPAom5LDc34DOCLlQFRm5REtzzcMb3CSVuXkSnBSx+QobH2mH90nh+MC
MG2JtgTaiKqzEBAvLq5qUdknREl4IACHyVlWjou8NhgenBVFuQQj/FcYTmrO97P0GlGf9FnIKASa
wTnagd9dQXDaiBPjOyreMcUTMoOHeZnBcqV9W1HSDb5oIKVk116l27PPVuAE7ZH9zyIuvQY7BChv
IRUJV3yLn56TKvgpaOsTsh1uBhxN5BVqHVkTZrecUZLxaUK6mhFmv8xKJGTET/9PI9OdFopIcnz8
rYxsYW/GxgLrgSwYm84k2FSi038bCo/2kov83PTGXRcbOTTsAUyO5GwSWJUJ8uH7B7PxjJfoPEzr
tFJlj70+nPrMTnA72RNQ3XNumjL2ba/qPimUdYYBX1hRdLKGM2hEgqfiaOWxYF/r7lkrK4bn7w7j
V2/jj20wou+/wbK4M0LNRi1j40xJTgcqoubKofPQyE/VV33MBPbiGEU/Ar8WjPq5ImqmPUGBL/bm
wKzSVLwJNaxhAzLM0uHL78cMpyCbgMXsLxBUH1+gRec4Lu4jvx0qcwKdtg2q2T+jN/0OuDfR+X1z
18aBANBdyPb4rjN8GPBDawdQTqCPYlJBIZHQxAF2IT/1os1wFOeQ6Rf6Gxn8cN5zMBOBbaQdgvq1
io0RhrUcpo6/KXrrDxc1LVm4iyVHQSwTs+/MJ4mNpcXwpDhdgN0kP8dcEBQ/QwHHSQkmxT25tvnn
WqO0yKDD8494Ng0POyrL+kCV76OyKqu0kz6YEPbJdv+4l7uSUtaVoVa6Fu0sLKCr6kntp8ahDr0d
5we9fFPTuHpAKesCMjmBmgf00SIO0dxNgiafbIBhD0IyP26kA954XRAsQ3P7IrAtN5k7L8nE2eKa
mdx+t3x/ebQxSsfk9BVb2tAx2RHHoKbOs2OJtp2t1i6epZE3MR0VJxTUTa6PX2Am5WQW9WMEGw9s
+VJ4uE/qRrGjOtilhrs/w2Qv9P35CKAMI1x6lDwV6zq8gPhBNRsN5hK2nfXfWud9y5wl7ZjVJtSr
eCvleh5FGsaxl5qYgorcmMGDXqxcuJd21bs3gX/jPWw4e3nveLBD6l24e0ORby6TKiFkE3qDWnqi
XWIJhQUUcYggAUO1FYnhgkCat5Mb/AzpnfTmOcjOYSQ5d8Q1ceiBxkXSs+GSZDgK/CphVTmyMDQp
a/ePgP0GugtrrMgR7yuQPxgQjsnCkUYTAxD2sfMv9DmUfgOBwlnxJP1C0QCM148p0qYywKaTOd0J
3LAKaQKu1fZeQJkccYdBXWhDMKQiFFIEENoXR2O/QRcyPEL0o9jCB8MPT57hS84JZBtlzNVEUNiA
z95kHC9shIWAyB9MMligdluC4T+AXGAfmWB5ZjTifOLIQZHbCLrqoK/ckNh4nLiLM0vHHb1nAT1Q
fUYfp1K2M/jjsl30UHi22PpKj+VNtO2N3T68w7rQV7skUzPDgDrvRWjJdYYcOxM5SY/ftBiAKvRE
QfArYGc8PHb5CULcSBtCpISpInBO782pzVo5d94R2rzUF5wOFvJqBpAdbS0PtZZLmx8XRCHuPQsW
1BgT5huJfy4yCn98bTq+JmC/O3xx9UTo9zScMEhO9FhisWoKD4tkYgudGIeO8TlDDmhr8uvmKSOO
vdWrRukGwR5PxX3zY65tZ65YX18PbbX8fY67aOWTCXLdJZ96JUBpAnhPodZ6/wtOlXGiUFKqWRuT
0q3iv0+ppiKfDXoyb0oIic+oyS/JoPWmabJm9Evx9qTuHZT2Cxg9TDMKJAzzM4P6OhOsBZUJSnYW
aOqtdbyqg2D0DXT7UaZ5sjcrBh5H/RKeg2SIO+DGbHzKKo1yfmKG1iJtoj/YbVhexmcTreaQ67Vf
Dpb8oNmtqcO+ZIJ3F0v4QhKe/hBGXysTw9nLJyrGXB7gje9FYBnnqeknJ4OnomF1eDRIzMDrybav
fJfkWR6zqVQLaREfbjz22VVC95Go1ufEJOodB3NyEUfrnPWpf+BtwZssyyay+/UazpJjDGO3IhtN
E9rFQaFOFJx6aYkw4r+0ywRJx4yjiFJZ9EoksNH7AK0F8vEkdRwGYwrhk9XpXYvycrauor2aV1sN
XygwWQGovSV3oLzymZfoJNNc1htS4tlzKCfgNwCwXf+rYTfWhFJAYi9bnMnCkoQ0c5NBesHyZQtw
FVlLyd2G3mIEXxKzWCgLfnAww7BqGgzMqKQV8LNJu/fbQEuZ2Y1MKvd2yVjWj1nW37MUrYaqUZD7
+nYGnJGI/Ys4ppk6qxh4WAJAijJR6dSdIas9QYs0ARdd+6DvktLxctA8W0mYTReA1xQAq0bDVkwI
Q/WVaELzSAH/agd8qXnVDTD9zOtK0N7l21zzOrZImnqgHtnXr0IzvIIBQomzjvY8usLGryKAFw3D
BU6v+KdI6dupwyn+RMTrguCAFLGjnUJZPAKi3DkJIkWCJy7BM1MNCZeLNkuL3jla3Vh8lEwyBsN3
C7YUBsvMaDk0czw6viwIGsYozQpRBTtx4ZxU84eUqWgPeaxlY/lo4vAmtqewFt8JspTK7YBM4MtP
IvoeKQTfruKBRNBlq4P5GzpdLAigSQE+mzdswtrKnRR0Kz9PvXI6Jzo+ARqXpTHMZVg0X6kI49mY
e7zqEn4XLw3fh9/eqFELUhPy7K8G11S3lD9vLW+a1i3eK46+q1w3MLQX89rP/QGJYvqRJvYVXrDo
GgNFiw9H6mPvTKt62kZxxz+M1D7r9cdk+YelAOlQTKKLJIyhDB6x8Q5jt/ncRHYWe0SQZFiu32/1
YQkYHxhIGAz8QJSNEj3qIaT1eFgtc1B3LlL+1ZfghQjPbpaddksGmqzzOtZXdpnDQSWcvNGRJeWt
ymc85u4ZSDw5XEcJFk7JeCVqEkCXJO8YRaImz/3IBVCoH44vTy4JAMkKKNyq+Z2hezX1TIYRT0RO
wMfnWbgXg969qvZVLIxu04MtAE7j1K9jYfiQc05Z/EPAZ9vmp0YitQj3hm9I8PNQ3ydRsqWDdyOY
x89kEhriEkD6zZeQ0prnj7TBhNeQqan9kHI7wKlM6aM0Kc4PXHeo78/kQZ/CkwkZpL41LL7ZhWSo
UHixbOKgeiZEnwJv0I0X99HpCfXLWtJ3t81RlprVDkClzENqwvTEvVG4wYP1J6zKx7GqJr3eJlys
oXF+4GhDQgeT0LfymWKdFkPyS+db7EDlu/PaVy71x2UzzTCWOPfZDPBGEmeGn0pnhj/nEc8S5FW0
hCczRWnyjfkwNLYv5Px5KVDeRLxwpbIuuScIG9mBPYfJS5YzVRiN0feLno4jdd1KYie0kRlriEdj
G2mKIZRUmam34RpKe0QMVgXCI+kINQYcReHnXIbXvhz/JGkm032JAdusUqguznPbd13anwDMh/2d
z8SCqhaaQ1d6VSIL5X8PIqWF/+RG2EJSvCbMs1R/80P6GxBW6XaXyv1qsptNaWoDsP2t5P9wZR6e
wG0MbSBycq1di9PlsnOuZg+G05MqPxhJO9F0SQ+4USBTN2J31u5y0c8o/ShbTFkisDqUon0IwjuT
Iq7Z+sqVk4KZvB9nvUEX5gaJFuBVuiNVP2VWpeR2ZTMvC684MeGUA2gcy9+vLF6ABN9oFcnv+7Ad
d83Sap2fmb9wZwm+aLVYHs06zfuvgZcap+4o4z9+y4w19VsMb5+lNWEu7CUrONgNeXwzvbq9fX6L
9XCaRA5fQMYMkGB+XhGKuBP7qup4Ypm2kHWqcZp1zJD73xjpwQaSRS95cZ+nJiNMWI17I2WyUpJ6
MAosqcXerRCbEVhxdpvCkDOP1c6/H6rQQ8LewiuB85zG+uBBSe2QsUWIFUaA3z/FrbADhYeEcglk
xlWlOyOSj+lFOjn3P1LyPFNy1jXQ0SyPhDPhBYgRE5x+0+BWOkIwU947bhBqDgrLsLxuMKayYqyP
ZlBVxs1dzPouZaZ2jkxLN/+bqRTh1SS86+jbRHKDcgbNcYjz1kCb73OQk3r1tR6A37eOqiNhgL5a
6NTwe5zNJrxD+v5EJxTaDaZYzmemoqwZ2mdv3/piI7d2+kZ1RlozNVs4ZH69OsYnkVybvGjoczhZ
vhZohWEiOiXwxyR+yR3yS9vBl3n19B58v3Mx7hloO0OKDfdCq5L+PJER1K0l0T0jwz7hmaFjTNAc
xkKL7IPZrczW4lT6xLkve11kozaqIVGtwvCETJlcTnL0qlOI3jiatXF/amq9z4kd2QsusJ8XHuXK
k/ctK5VLAnCIabKS/HlBtcfdyCRJVv/BjvGH8vrUJvkplrnSn5+G/VN5EsmlOfE4nJKUzKzn2hWt
Fviw4C4k+xbJ/A/jE1cm9iBRvglJseAyb9fUEVzJBCRcY9Ry/4SEeONEhX7/UYk4TDIp7OfJj2eM
LROvsW+ztHcY5JR1RfAICjdCx1VfqO5MUf1BLpKgkO33/GBjOZ2JWBqxOg53j3qEsGamOifPNY3L
3Qj28k3W5CrBvOId3yzvv9JOcHeL4ZPHM4Hy1K5djiKWEgxkOrAZrY0n0gLdJz7XdQdLsTPOg9mx
qxpiK3zpR9+RjgDlr0Su4mVo5CNAqNVZkulucaDoOT1EfSJ2H2xJfpTTVRM5l7fNdlNaeUF+MWgs
slslVlRaDpjNnNMzL/+udn+Hh/xQ62nQa7ma0CsRhdf4Rn1htdLt5wA+V3DgJmZNppOR8/x/0qOi
ofeZ1OCtdcLttlbzn+gUQEnnocQ2SIZr26j2h7rRM3jt3z7iq4ZCEhRkG/RIn7DN+0eqzM/6FybJ
odSsTF3XbVg1Yoq4W2Zh3r/80GkEL3XRMl4X8YTh2rK5AY8gRhAq/KinBJCcc3qWeHzeWE5rhw3D
fc2T4FreR2fZX5xxJyBnYz5AyEhPdmCLQ+jzPxISPGJfciM6pHsiv2ABts94f11YygVifCNUxEZb
nhkhPFfVjDNwZUtmzp/iAMK7EHYoyGF/vTH2d4oGO1VywMoSMSarnItP0Yao/0Qmdv6WZHSMKNI/
736xTUJpoZabSbArS3oSDpLUgg4oz6g/whfpx3k05j4C5tklqvU+3tqfZx4lW/DrRAFGfoN5af6y
Cuw62WqOE6FLcKnaLMlXKiA5Df9KZ7byiZ9C6SQJ7LAL3LbaXrXRyCznAxoL/CPcXLko3V226YDm
zX7v/i69CB9gdLi6tobreCTI+OU/jFVHHWPA4Vab3zFpArNPDGww3g07+roCJqRhtkcex6ip+gDs
edOfpRi/q3Hom5V6ZHCmSc2z/182mnlUQrWt05dIruXgeI4JUxVHEnme4ZmQr+kQuTFsQhtq+A3T
6PAqZCzSSNuinP32iWyDIi17fIjznH8WBuhLSjH3MvExDq/q+7tptSblzRVm5IAZpDM1rzYKwALw
PmYXn77fh7wHqgYuZyzwrzXvBadzWgYDOkGS482caed6QSsu/K5Ko/1pMltVtTR03/XhTqZqicV7
OK/ATpX2ecxjJqP2VKB8doAiZUSNB+nIZL7BI3fQVOdMLsERULcGE31xCztqdX+KvLnFZz41dvKG
f3cBke250ONBTcp484hhDeFKsrpIsaz6Re8dCj6voxuWHBjAz8eptXq3e37CvV3TqJrIiP960SVr
TQ42FAQg7i2Uc2OzjAnm2z7SeFp7Cp3k45/r7RYYZ0OMqxoIZ2qkGRpBWgxdeQ/H2WlmAx8ydRBD
7w0KEeHuLJj0pqIiI0kYi5YIRavq+AA1X7fsjLwqq1Yfawf0I95DBOYk3Oz+kMLi7P67pi6uVnH/
rp8cQSZBekpGZpsWN2trm0fNmRyPxEbg+IhE13rRMP/rHE4UxZ5o39c2ZeJ228tpcF25qCTBLGlo
XpYXbt/qb6g0BVH+IjzKr8rDX3YzXojmLHgmGvtDhhkW5H7P/Ij7rqFW0p+7VEv/xyW92x+lId2Q
yhmFEeiAnVy0gZfIz+kAuPg8LoJP6PIk9c5HcrSVhAnCzeuOXjisxzggPQdtQmcuu+pds92EhxIb
mwtD9r8K1PD6OKgw9HD1HdqFBHCd1ch3VhbBq4f9SL3az33aI99Rq74c+UFsgAT6ouELkqTQmARd
yzezf70LWczpwWgce5LseA6LaHtcRf4pGd5Tc2CxTVW31wbm0Sf2YMRxkaRyBlRGZkHrpCfGag2F
G7F09EL+JhwtFmSCJmSYUPqUa0YkPNAL7fWUTL0FUcpE5h4QvwJiIrQ9FPvUYanDIG2oKPkCE6g9
D1XnsgeaJ8f77lcKkLAksX6iLycv4+bMLtvo/Qig9uhKpeHwnub25HQj4Qtcp4GBGiYnBpqJ79tG
FpaqyppehD9eGWo9j2kyeCx2ck9qWtN9PDJVBUu+keSZFmQgcnXuNsVrXbTmttsXu9o8hT7bcAHT
P0JV84GdOhTIQoW962Kx8Qdxi4L9KuzQMjSYiWYJoFIAHZeTgew2XKcV/oqjtYO+ScTi9/RtvtcB
mMfybBSCN3gMoFaQeB44/u1jRjk3cUxiaXcDxMZ8BCsNUfyfFDEL+B8GYX+BmkpEozcZ/FJrpXG4
W2gGvP7fwx2GUwvJxCaD02+s6SU39EjRty7YYV3EaPnqWEvUXXI8E0QRtrENCg24N30fN6MXH8vt
TWdIVBV2RqHbXfM5c40f44nYHczFBUV/jV7aDArrVhVVV7f89hw2ZxY8FldP5OIaqxa7TnLD6gyP
R9r87Q+8iu7RRDU/EeOMArUysUmkPRKISmQ26INaoovRK4XV8xvKsottK7gUuts3UJp7T6+Bu5jH
xeX8f9yc9cnMtacy9TgXw4pf7vF/tHZJ03oWHcRhvF9bZAm0tVAgQeamwrzxJVr7W7fM4HrmpSEf
G/d3o0elKw7sWFFTvjCw7XRMeQUUvIGdigVXDfflJMNBlY3rm6HLneDghoiMH2wkgGDkSF9PAMI+
2ydoo5DVWOALJWR0VBLLj5bMn3WtSPOUNhHaBdJgWJx1KGsHI0Kllc0XpJFNV/MV7WJrxu5Yp4m5
/AMXWqhmv2MizkcJzr+39mwq6lqHi245n+t8hZqhH6ArL5s+cmB8nChU1ZUT4A6HLjXKeWYvUnw+
CxBBdb9X+HMxHdcbKVRi5UbZRjp+hEdFDdqsncCWPKUDMgyTyokDs6j0Od7wu8Kbx7JCAFLiYCcw
8QLGR6/J6UmUwv8XZS+of18YsxsRiARe3/rDGNN40Qgv8QX2cEFMCKV5ne417N/RFyZgZWN1uJvc
l7zlz69E+cfiOUsXkesulD1dJ25DYD6I/ypCJjlxVDr+EFKVCVXohHBqfjOnEoNTk2QCzcVUrmT9
JSFUyhrLmzPahVcepsoyVSqonzbEYVL+7Fi4q3dN6n7sBklLOA1Bg6VrVfyz57RrVlXLP6KavtUM
STnz8xf9er9JcqOULYokfgMWQZbA6wd26NEhH2Mf879rBUmIfzAgatFFyGpOWVBgcw1g9Ng5tAm6
ezPWIby45yjRoltp50wyWxUYXc+0Df5IL5LsIXW5bcgqUHOiAhRbHr9Jda1Qu4KyBFs5O0Jk+pHZ
EV0+4Cy9ohn808yNYAkVTiiUHicPfoEieaMib2RDloqraHoUnwB/Zv/3mMqjEJSosW9/ENCm8/CA
zVH9wUwv05cIPEhrLHo85c4iqMiGNKR377pK4393Kvzfv6xOPT31aj0GcyrOk/hulRdVM+gQoDxJ
sa0meWhsTiR9eWIKBY7Gax6RYna+KCC8POopyIai6deFdUj80H3q4VBeX6sWPozG9486QPLDQopb
uZQkk1/IDRRhIPdw1/LRLeOvm/S87ucf0m1fMwHKrdGueQ0a01taVjrLEhCqIBfMFz2QgkxsIKk0
ZCxM3x8y66PK/UjoiyuiY/+9LkTKiwIhiO8g07YxvnzNeQfLQVp1TS1ZvinA9ucSn1AxKiZhovm7
JG7jQdNNtlygiiUxDXmBsLmAho29ELqyI2mJhY0jHP4763hJl1ImO9KErctHXdUMu12Z2z/AxVua
45ti98FGRqukmaq1b2jQ6mSNGVNiPPnUC6xxMJ8Rx+AD32MsLStg3+mGDLQFh+RbT0WRgEY00qK+
tQjokzaXHueAyCpjr5ziR6EJAIyaH0g77NX5p3NqU90vg6BtJSRd/MBAPNBsfQVOL2ve9Z1r4c9v
kzXJLgyfcg76c+Qw0pEHQ7hHnz+oSC25LmAeGnddy/esJmDfJM/+cBPF9E87vQi1qstqGt7z1O0e
8InD9g+W5dpXmtTjCzmemMTfAuoxk32AQkLjmtkKQU0P6LjAow6d8YycUNkBMKW9cdnNO3FMAH91
zQ2WeG3kYMYH8XbhKTSNMcd5fVfE8l5f1uEoO/EZkNTi0FS4dtopAIgNZxt0FuIBRJq+OAUJVgl0
XVfX54BJ52CN/AhI423c/LPNndEn7njKwhb9uNays2Y9C6u7Os9hDR9E4fOGI6/Iy881i7GPR7kc
n6BTI1kET6NnGMbohC3ouVlSecNpofaad3VEnovQHJ2ToMCL/Q4ke8G9WDZRZcAxsCQoW+Sr+bzx
OeSxtUl8nmONm3aayMBdoU2UDW7bCrQcMJtigbcP7TwxllsSAphHAkvi0hcTcLWByKr/wtnUqrwh
D551vF+usaA1OMR9WYsQgwWGzJCisQxVMgmYTbQUNTI12vypQy97kUtfozOwCsxLz2vzwGWHCbMC
iUfGEMBe1A9ENr683Cm4Jlfdd/Nrf6clM25WKJ4oiTuEQm+21WVZPpkKFfl0eoBsnKQwJzzyIGKp
y9J5HjspeH0yPBMf4gl+H27pBOy7wcXr6jJMi+WCn2TEm2MIa7+Y45W9REs2Zo3mP/U3BmAo4w43
8IXPMlZTQHOYyOK1+EW8eS7h6djxkradHwfEJxnfmDlikNc2MqQUSx+ijq5tMWTDHl8WMZUTdeht
oiBppBEipw2goT7pUxvV8ZcnZr3S5eLTs2Kqg1ANI8YHFHh/ZMA4oBUVSpMcGhS4dMbiuplbZJ8G
pKhHReWeptxm/MDgQRz8KPYA0QAS1B/4xbHGO/cVX3FtIaqb7Z8fuZM85XoGLk6e/xO8H15H91Y1
gaaR923wCllupP4l4feEkdFPdA9w2mU/TEdKiva+S+mBvcMqHMF1JpNR4HWtd8jykYBUYxN4yceo
NCEaZ1D4G5Sjqo0v3cYY+Tl3lomATQzzYz+MUKNU0MA0w9EUsmdwm+2ZY31V92StDePRNSydpEhp
3ldgSymyutjf7UJ/uRIKb0Be0d8aE2wspm/o55wIVChIwajPwQb01UBnneId4zy3oF9vMUPlqQoz
hobqwpM8V/YC+QAGwu/GDZjOjukHMfIW7j2Qv8+ixem7GCV+4yEAOh7Oqvrx0H8YZQb+w8OEOO67
GKPfNEP+SE4uXKjjJzOb0kLBfoeEXlwOmg0HZ94d7IoFydZ93sDxkTl7Zhv7zGgWfgPW1Zo3Q5W7
vdc0OtZMn9aL8GybqzsgnRZV37OExmfH4lqK4IkZlV5XpgdBCuMj6DncuvzGjK6bzIimz7/XFZTr
D0MTLhY8/niGSWbuMm8lkFPisZ1O1rPqF8Rq12L1UhcZ6j+bnIH0paVxpz0KVSjyB0zYLnOMKRFV
zFNH+7pMhTs0/36vH1UmyEl97CbsvVg/7sTjnbMxLjNBxvW2hWYwvKFiNXP6JTeExmVi0sPZcDof
E4UsM/OrMlVQJt3jijOUbEfEW/D2GgApv1bdQJqt225anGq7nCxk3jjEIXaXUSRIysXzS2znOfp2
Br+xaCcXzkm/6rUoZz3JEM+DEmkU2ykufPbum7P1XNqIrcS6h1WSDrhjRGhBRDBJdOmw60tzuDvH
c8LoC6rIxc79sYCMJ4hUGORDWxMKraPtxjfn4cVHcgoViNgEOJb5Y2jv52oD2g/d9zEu2VH7FgI/
shV1wqPmyfqT41CPOEu600DPgg3CFZkh/8awG3sbW1Y/l/uCS/EX1kcbwjQbBELfTa32Mliv1fSt
P4e6kR62Z8KOGfLnB7jh4HnS7wuO3xOGx2ySMxCJ+oqwqtL/F3yYbLOJ11ijJBRoYLfNPibb41hL
kps6+FU3bMqDseOZox1+wqZhBF4wnAA0801w+ZOl/Pq9T6FtXpJoGFdFgbfbiayhJ7avYju+8DlP
vXJ7JWSRmr+XsgFFPPEz5L4VPhc+P38cF3GgNwx54CeSvEg9IOIuOei6O3DgzGTSMkGRC6oXIwTI
LGFI3m9vRVxjIH4b3xZ93C4JnbycWaJPMifYhe9lnYfgbzme5IscsYQGlO5R7u6iqJIyvD6rnVOT
MGy+qHcB8YiqATkr2Bvcy+WoiBgq5xl4nKbIC/NGWbAGT96o+Q4i87O4fk4JRNdsPOZmAQuOwuzF
+x0gCdvpdn7XIQUmzddb1Qo30Pf04TLEMnIbQMmEm/NY3e9M/b0yPCNSVtO+FhQdixOqlYvHMHrh
Dp+QfWbfHT/vpbhne9eDt4cIasNykXgLALGzuVhrUMWK0LZcTHagYGwVow1c2Sm9zd+aJo1lsKLP
AJUqVs0OaPEqz/bOvBVtPmjYJ62GgH0VCappUr3ynCAA45LcQiS2INOrTaCnYOfI2tyDY8m7L62x
clTp2z1aGjnTWW0uraGdaHkpIWdqIhvmkRk+BDN+YjTBfpxQxYeYGmG3TalbJdXU4yyQmIQx3YaD
WHjWYfFA/nHaJfoY5OOJ5UVEC7gAWQ6YtTbwrnKqapxM9fbAWUAlA3jxSPBBnUuPOYK4B7B9ITrM
5YzCDCxlgg4Ni+rsO/w4S2d9YeG+9jrNaUGh+RBnDFmgm95wEhZSUXHA1jWgCUBKJcUHsTEKkX8b
rgXfTP8mJBQaP+xsbvlUC+zH8TFQjGg++IJyXbkU96PUl/rUUN2IJATRhv2z/CSSFZQtPTWheoBR
PwUoKugyVDEtdJTjPUNt5LtKGkkmM8PsmZDsERtm//Pwgw8jqWFC9G/E3ooDJPv6PuwasnQUH8i0
57k15GBKq0wPCd42ULZ+z1iyebUx+XMa2M9uCJU8HonuV+U18U0SGZfEXE0kPy5J6laFCjxn0Lww
sZEmLQw7ycCOO7kwT7u51B5M3vpJnTSJqkuXvysH/V1VBPzcrHt9Uho+7lCK9xGn/3qV5OmnTsnB
qkiVZ24m5lP3SAcqgrdRpID+C5mddvHlQLWgQEEm8HPpJYY57SgHaKJOb3iMcJFqR/v9DYqTR/0H
GT0m+bBjQAUW8vm7oVcwDcFF8QdDFb87QifzeigCBWLKxD1qSc+Tnco8uv61FqWpdNN/V56qWV+R
Oz7yJzZybmpdKTKqtyUhBlinzgbc8wZ73Bmm/DgdqW9HiTxQf0GNXc2s2tnhYSZrv4U+bUjDJvOZ
rOlEOM3CWuuiiLPQiHOIUse/rF+mH5wxlfKJzumFbwRLvH87Jr7LI4AjX3vHWHLjS+rYPvWZdvRd
3MTQnXfo++bsF3yqtcrHJ7lQMNCF++fo/jEI7F5BHsWw335NmyWX3fOPwWC0uzZGgc1dalIv/PS7
X2iYOYJUbI9wlacptbBKXPJZ3gsGquIhhOp4iaGZemZBLwlChQXUso1n1QmnHT1VcX/v+B/5I72J
pTPJHQ8S9V1kE8gusw6OPcTgSa1XNxRSAA+SZ4J3NbcQozkgrOBwq44b/WLD07a5fn5VHLtb6qGo
w5sUHbjGSGJM/0VdgMXa7klH+8gK6QMHOzVbxg2XP2qHBJpCf7m44LoC+8FpIBuSRa3jljVdbh6L
sWEWOpKjjnrjwsSLJoAIUUmTu+uiD84kbjIkxZ0gQXz6RKzc6JjSqZrgau47YYomK7bxnWyD9ZKD
/mj8fuFfn2H4+B7GfzqaBybco99iWbK4ZkkKjADx8GdJM48NVsZ/5+ABwzOO9NZRPywrnoPsJkuQ
WImmoR0vs8zPWKsnSeEbRocDjSG6RgybuQIBya4BdHyE/489H6pnAic1vkKoHRnAPogh5S66nm+0
X5V0Oy0LWPK62uSAR1ONrr+cxgrkFHl2HrsuF0CXtP0VmWVk+Lg7sqPiEI2wU5Xg6Ik++Bs3M4jx
vwfm7af34SDwinXVlgJkWyNgv7008oVTow33GLHrQ1yL7mfrr6u7Aqhkbzl8qJDA+me79o9u/M/v
CUv0GCxQMmx4fBBqJLXaK76VQVu1AoaL74/reXfPRHzwWzFhz6mCgXvV30WXsVgIc+ZNfYAblwaY
r+OcM1DVfPp27uj1svJL4+FEdAfumZ1Qu4yiqQl5mVMAdlTWBa6tPYdG4l4siSOwjGd745UkP31N
91dDl1EBv6qpiEYOYH4JnR6wJ4SgDahtx2/XW7DA2Kb+XVp2hF/kqeF3mDboB4nPYrgjSebQyKqn
PFZwiJJ7bfKU9wCDjLbVOCnQ1xpk4Yd1mOf3GyGqN/CdKMaHmoYtMqL8jDZkSZjPmHEIWEMIZh3c
vIgfaF0CH4KS8zMdKi9wwih1lnVBrXWHuyLKPVnfP/qFun3Y5FHVRYcHV8YMT3e4GAPKhb/eqlAY
R96+oi8Jo3hiMbCaTEDpq5wbrR7ejhgisQnHhlu7/o50OBnuZQVCcMwQKbvNxe20L1+hFlazV4Zy
VeFX1GW1w911uZZoseNsDnvUT2M/1Z4YrXIA9bQjw10ypCqydetNiBYS51QNEvv5bv9QEUYnPXj8
S3R0vjzBPGYivDglW40nVAqQ+lf1GMtxlQzLfmN5RGhzfNeUsn8GPHtQiU34xjs+9ugBX2KuPApS
8n5IOw9P/orU6e4ObPcNp+6odrG0BhjvtZ7mAwDlK/HeS5Xmcm4xgXBhrDlf0MkTX8TyPo8XzQH0
QwDC45z9baNO8FHCd9mrYdYsV5WtWUx5to7IaAlvukBHClu+A8c4FNdhTeFNWZca4XGKmG+FzfKH
Jv2EHaBd41snTpwJue9yV+StCbQ2SJCV+Nkoz8DX1dtBWL391O9cWMIt64f1z/HfmiWKsbST845q
wlhSp3UWMMJmXNCNNC4YQbrWwnsQDaG9RmFOiaGMOJ7tIW+3zyXmOYES8Jh9i46l/HH7hG4FLhKM
eieBMPhtgq6NFByATyyEetO9h22DjwquEcdcVHGZzAo9hqf3oLrFBTFA3J2oAT27iP6OpTVCkDMX
y5uWjmTfuq6J0cIn+D5m1jJu3E9OuvyM6A8Vu3M3DzHNSrmusP7I9dq/F5jDf5kfWjHWkB3kvVp3
RApqQPxkgSEDlt9XWKqdLfJtxJ0Q8vuIlKZ/Tt6dsTwpN4RtInk1LEQWlOxIMhYjgV4Q4BiFeCOx
o9pyFzQj9FstAuXmOy9Mzsun1jMsWO1Nra7Sx4WBaxK7HwuRDDodIzcwkv65FbNbcB9bu4PmtW/i
T9x0Qg5hYdMrRQf3a4Or+eACja1AFIIiBSV+ACprArAMdM3DoexNMwDb1n6NfNsrfkUfm7q71sUD
qynZLVpAPSZaqQ/sI+IxQSIKRIqhPM+TsDzkG+Tfr9FEWK+aKXVXs+zi3g4MDbpXH0hkb8EwiEVR
iRkzVXxf11+j0mTuxkJlUidiN+BJ9VkOeaYcjmNlS8oos1cuyGS9FgABXBBRaP9EV6vYb3jrgcIE
Ak52rReVpFmxTDKkF3T999yVu7Ine9j+Nx0+FLlHrjI/pWKRsdKUZV61RNMX2HHql+Z7yCOKVQWZ
yNx/DxBM2lG7ofFAMPNXusvLVqp8CiX8v5u/AAdJQS2GLXrfAVinnOOClK70+T73L5uPkN1nHBdM
3VRhMRFmEeIoaS1tD1sKmA3MGiSe4C3HJvXY0XaO/vSaXBP2+kFQr7DnZOAIAxL5CPqtfqmAaRid
NwdZLqiB3bMtTQUrkqGI5G4pZdtIlSCg1qCqyD8k+uMslHjIPePZ1tgrfFeB/yTCLR3oD9D9zZLq
r4VLUm8M75HSE3gMeuGxPfGONYqTWsTrQ7hnqA6GKg2OYX/0WG0jjr5XvVSc6+t+M4uqFYBbNfp0
mvVCIqwxO49TgpgsrYfFxrsVXJLjbcHiB+GhDoAxlbYHuOnwQe4yvItF6nfjc1BIPBe1SJsusYWZ
ivr7wAl26MLA7BBKVJTRGRVChVKhL+tET3YPAC6NOYAuGWouVAsWJd0p2JoJXQkAzi1Bo96r/T9+
ZRUIxQ7CCrYexpj3H57MTdPpW6Ymhb/bapNn6dsFlYpbfczlcLziScg8G+jwg3eltAKmVpwTw/wq
kWk3OZ+3GZ2up0ZJnkdhpKwlwov53EXfykh1k6EnfbEKnvOVXRfJDRxK0oU/gFBZSNivDPT1rm8J
bBo/Z/4XcYnuEIFM3vFGxQlGZ/yQRMsbk03mCxKkCY2HuveE3VLmMARSvJRAuR3ijUG5ygQSxQUS
KFSql2Qxb3Ar0jJNoX3fyzHVe5QbIHIcq1QEWFDO48Hqwudrpa1/GhuhPiJ4NbvM3Bbl2lQ81zlq
zjes4xtuJON26jwRYGGMkTUMMngfLm5JvLLfzZyU9lWMkNPItp8Sf2D7MhYF/zNQjrRp9G8Zu/xz
xpFZ6IN3aFktk6UTY8YZd02l7O3sGOab0rVfUHhQuLrY8Naj+5IKPLY+l/XmKddfPtfPlKq1cq0A
tuY86RtCOgGUd6DZ3Xo79wTM+hKGaJv8v5GPjVv/Y9OMCJHa+ngWCQK60Uht79ZttpSSE4HEqiL9
j5NyhiilDz736nfL47tQsRVJ67XCTvwlValnr01l1sfv8PeTh331n+C3xXEbbh0tHbzL0UKDY5kx
taC9bzzVepm0MtvuvrMrND0MVqbPk6StGQj+Dh/2oeiAcQ1xrtf7/eWc2X2yZrKnq4Xc7egg2gGu
scljh1KCLxWei7bkOWwOn+hYpnNY8NhhmIkdCbAJS9ci6++xVeF8ak47Pk5ArG/oJrgRkAzxejuB
zON/bk/K/aIxC+RiOxmM80cePpexfsfLNpcAoQhcNSGaE0ZjBRCHlUkmhSi/v8ax/DpY5bK7/50x
Ck1V8GPf7hRVr58Ds7xzNytFUh1SHKtL1qazKwGgbs9vraqEPLqC2tagEtcGExAkFk4QzlKeCRmu
VLhC4w3ATyId2zkyOZsei0+kPeGW0pIWx9LcUArr/xPwnYe/qepm2OMxE+bTnXFB37TzLESempri
1zuJl+RzpvuY5BeKtzQ1EaHbapmQIwGBUZTHsvfbMLfZIauJV7gpWrg+ghTV4YTpxb/EuGE5qK9o
LDW1LbTb1Uya2L9miYE0bphguDswr6KakymljYIGMFs4YUskN9wiZ2PxocAT98/vJnn/HFXRYTzY
j1hmDLOIuKE3zIxGAxN6vHORSqorkAG95RtuC6qPLxoQVZ3M37xrYOl5ahOgus1u0EWWfqVgFqJC
KXrZsNP7Ip5ZGNsuVBRYHwCNWpVX/A974KsR1dGP57Qw0Y1POkHIFl6iHDZwP2lfG7AW6sejxxGS
dcuX0cR3VadUzBa0verApMIOieBEdJq9WqdRJ9TBIL/Jo4K6wQT1VULhzpkVeaa9nyvX1ZS2iASO
fcjjf8vH74SmhinY/EFvzMmxFUy2sZCVkhmpVIc35kPmjnho2GBvzW+WlOCf0LPkVmjaOVrPkmRm
3yFht2FVRuGmNTZ6ldmxeREb35sga878z5UQOmufxplKCUb2H465a7gHQIn0Q0vW+gnWI/69BkmX
tQrOBcQeH+HkkPD+JefasdUAsjKHN2OvrLUbw1B1bLqyUIPcGO6Zze6h8vETYRlTr++ugTE60qFI
HcIOfqsSCWfkBV8XMHzO+EACaY6ow/UjJMhkcEf5g7Sw+f+k7gMaRLj3XH9EVRu1MISawbxUOGRq
xROaY3fkl6hUHn4iCS+xxKlFWBF6QidX4U62oxFmZItbbmNUthvPKaK8iRWkTNTZkjgAbXosThXL
8y/Ao/E8RvtUQBu8qfmm173XsMJ1wmtZTcDwv0gPl/1Q3Wileg0AcNQ2I1tiefiCLE33NpUoYpRb
Jjr02qWgAL51ihW2onFShaoWhXjYuw9YIS5D6c/wELocViC6Q0bccw1KT+j+lQt1QG4y0gaTFFS+
PAESkILonHAY9N6OR7Kb3yBosfb9PlujDooL2TSPB5r/TwcZ7UjHjtr0yHkQyXaNWYoAURuA7szC
9yJkH5ZEt6COtpqhC+xEVuLlpoPGQor24w6Zkvuv+vEuXSA2WuqlIx2yXxTVAjdC6CJ7/1aK4cUr
hXQ/kFaRIBiNYVQX3vvekhln0zegMVSOxzsbR99pT5RXldnyPJjtF1RdQh009anZrQLl8KEXYlSZ
AHikuCcUsyTrjv0cJy7cANPnWqg3EDxRrn1nheRTzD4cfmGnf2VXl2BUFkymGpi4BJO3xQ8/Uj2g
a79gHHAziQJaUi+NrelHUjMjO9CLmdKz960+rRbBCAckcygEH5Yj9KYXIVQ4VL6b9RLAiX1FufaD
MLa9RhKymdQ978EzsOm5S5HosTomLnXRXlI2ipL0hIDEfAbhnPooABvNQsXRnPWg7DONp6bildI7
gJz1iGDN0xeUjxBahg0jKsOKYRmTRwRi89zK/EjclGiA/mTs/Yvb3z7HXmeMu7MNo0978e4TqUoP
5VLEj9mHn+nIGlRFmrBel/jyqOVOnILJh2G3Trk5E1G9U+kqWwc6/p4fRp8tzMf/eeiX4pnQ6M0x
DtzcOsBac9bAXFJJCSyuT6llyHkzIOM9M+QMOuJOujnyxVYAZUOzC9Y+bz4IwkNvDxOlj/uISwRa
Uh9PzBOcro4Xzj4pQc5ASb7ISSqLemyfeu9Y8yVKO/6An+OaU9FLALkg7YKSqVijDwmrizM+U81D
kkXkvGVSbzAjn3jlxoboJYlyoTWuFlERspa0Qg04up8TBSKBKkI+ei5yomdUhQKUimpHSujIJBSs
byblixxvmrFqZvXHgDEZBTJGJ4e81Kpz4iBuQTq1aVe/5D2+sgDVIj0cHP0XJTgwa0JJK43ljtMZ
Vz34rwDMwGV/DuFE9iKz69//+28GZ9T9MbOn9B9FiIyl0Hnl9BxgkVL5ZxCJzcskIan6X0zMN0rg
UYSXr0eP1MfonvTQesK9uhq/Mcjm2KK4/guqWUyVChRCwRy/2zDfWkWc8rNt8Qty1gcUZcusiFxW
hl1SlRff8bMSxS8W/YBysAX8zdjO1wF+OR+OcupwJE4SZQ6w3Tiz4W2UqxQ4cSHt/mUy0rxj4e7u
mm1k/4+eg2MRfCjGti4Qpeh0jttva3apnDJOCWGscO8c26zG/oEdqQwZpW5iCc9ZVH5m4rj9qtuj
abRNoRwu5xIfEL58vWi0KXVbJ1cn0zgma3Fvs1GAXubki6To1EqTpkkrCLis5/H/iYY/JOBNCOpL
F/aPukDF0eH4eHqoIuvq13u2quI177N1h0qoruFOA2OVc/dZmFVQ3beDp4uCtRUfZksqsXLfxa+V
E8k2prpTcL5k7M5jdtLWxVI+C8TB5a2viScsKeweb5oxsDOwwjHgeEYWtnv8bPWWUS13oGgGsbYu
ja1oFzQeYVoHTZt1SLV5rFz4JvUzEZRvtp0kb2BmRGP4hiULk3rWDakUMkOqxg4Fy7gbtX9/WHR7
7H4C8HGzB0cQRa435JdFIOyst54j6lk++bQUYb8ttRTOMWuIR+eH9PLYwwOflvXWuBYtoI7ZjrjB
W2SrV/3B0xjGaAFQwXEZ2f+5Rq5f0lxGeuu/O4mKEzE0iNT9g+Q+xsPPFZU0WBQySKdKZW5Y/yrv
cQWpLdWlHZCCyl9GGVVz2vc7hgo5eZG0M3ml0nId3koJ874tTsirpHIGgvTSDqGmftnxnEbdLlym
9iTrMiEfldh0+I5yGtWuYdhtGr+jBZKQ6sW4xjOGzMiRA/rW6OW56+TPEByDJNDlw+qY2WSJutoT
ffj5NDEzciUmT92cqBsdIu6/twwcWqrHvEXWx4Xk8K1HDmT0c6g0RWxUabTOX6uUU7HH3BJKdy0a
d/7D4KgWhtlxClpIoUi8K/RRWLefurkIfc9+XDVUhV9Y9MoPZiFqlVUlxkIhv1yfP7Dy5NU6wy0r
HM5h338ZpbvvT9ouG5brmYbdRb64UpMbZN/qrwAS39ljWCFTa6F604ivvBhB6mkx+GQNrsEqiwqq
JlCU4bHuUCLANrpUW+VsyI1fs4tCnPfLivUwBiOCz5yuPTNd/4U5VLdFiqLw+9y+T/zRFi04vbtM
wdQPt9BkrpY5/uU3Nvd/yGZNBhAKqY8BQm1qymqttzG1gHp/6kPiWkvReeWjCpizxcR1FGutQOQz
ypmnYDHFkGQ/5SCcxv9AVDmDNhIsRkPd53eVY6tKr/qU7AybQTxDheCUfXK1EC/3nI8U8c84VcBP
ZD3LoJicXdxiwiJf58xFnhXKbEmL6U4Qmq37WuUAVrP5FhatCMStPbbIlzPnFqV1mMuGZgwSWOkP
WF/4aT1BnN4ZVX40Z7QeIHC84aI6zNYhfRS7qiIl++e5EOS+lyRz8mryvCK0LsTlo5PsfsJPXF3i
ok7BwsLuYmQpB19L/n6w8uYDvqc6peZuPXenfA5rjdCeN/YN3JCUqeaBRmlsdSTSyRkOMqKQKXFh
wWkKt25K5kjtemJl4dkrsfBH44swzbxQX0GPnpMa4TjKUy7EPTPUTcjrZsaNCqM3rp3bCxPP5xOo
a1KD3BRjsKZRUC3NiRidKFvIVUgh+XjeL7MTjaKASgQdTCbtB9WvBOTT5BEZrJDh/DWh8Lq60kcc
FHN5/ra6CTvcu7Um2NDFQJjxEszBn2MkKFYJk+8NCVyk9Dpio6YfJDpWxAipffcLW1ebDvgvXmzg
FMttqZTViaHSZUk3VIuarS1FKS+1duR+5KMk4GLsrGTJTQDRORcTNVK8pKvZxo4rCYC3eU8jU6fB
NWCM1o4M/C7AFDpodttl+fYb9+EaSq6Tso1RAIO8AE8qCqSM7ie/X5ePWYBSgho6x1W7vJTkJX/X
oWfui27syOJET3KYaWar8Xwr75Sia0wGzxSKq7UHYKRHlgeAY3ExKfCDHK+XcLWZOhYyUjmaQBRJ
BXWf5ybpQkkdSwbHAu3iJxHICt02zCBJCq+PLnGdqZAeFZPYgFqVtXbrqKuhgwv738ip6SOwMUkq
Oc/H7bbof5DhLHJSFOqXLhkLp6yn3K4BD47aPnZWFxwL5JltsZ3B1iRSsZVN7LMKqrheIr0gHNDj
IOfyKBN2fMJ+R8D/D5tInzYlo1HVfPyHqZMiU6IB40waKGjmzobuqf/Z5oO+S9OeQ4zJR3Dy/fR4
yVe17Y6DhT80g68ax1use/Llmu5JCabBejHPvv7Sgvcsp8biXk1gmivbvcFtM5578CR6EHCcDzdy
D3xmU4ax62LeKqPRzw1fFGcYhuHpaf8bmkJMimklUaWkEs2x+ntsm7BxOFC3zh/AYKc+ZDoMU2Al
khPwlMXnhxa7X5RIGltYWGjx9w5b9vzXi4whpDIYxMQNKnlEu2jCN3ahQ1u1kcUamj+BD9QgWk6B
dyghaTNHfI1b09Ye6n1sQe17lGlz2m/g9vgGWRGd0Ulrv9dHR2dPqfyJYocOT9B8nqq60iA1Cwfk
1jHKp4p5guk8XkwzQH54TLMswPtHUPVhZ2xYy0rVZWEQr4focftjg8UjKwvJ0pD6g1Bj7IZGo02r
8MZWCAnfsd3O0iLSnjgEFxJy2u4M5LH1r9cqrLvTA9Q+uJz8AqVW/2PmAAzRMyiN5P59jgSGt6WK
5wKgrWQtOPlozdX+gyVkocWenlIwJDgNiMWSV46mVOtrnychJNeA1mTycgalyXvOjNMRUgOoYDhP
KuWEq5wLuLfAplHdS0BYnqQu6Wf5yo+/8Mh1j+ORFQSHDidN14X59Jj2IuWXToqrT6W+YNjipWtI
+6dqsni+Yo6eBdptkq730Z7S8ICPXvfz5eGnq2SUNGXcJnWeUduG0hl+7x1F4z4SWKYVBDLRyZ4d
oEk9aD6/G9AEr3DAkZ4//FJwevMh7ET6oNf4uLrrRQcH7CepZJywV3ortAaR8SeWH+8BI72jnowg
ENSztQCMop2UA3X4PbNdLAnnCwvDtbOqJBFMdiH1+QpmxFW5awm+zB5gXcw5ymz5VC9Ow1DNUU/8
WyNIF3+Tja7d3eqycn2QMoKKHFVjn0ViVHD2+NrB75s5ZV5sE4Iu1LYgrUvh3YQhWCwt82/npdsE
Et8V1LTYYVzPuR+NSUj30QnWGXV1DEJ0xfLJ5JDtKrlQ9/pGRKpBzZTXLdxdFXoo4OFXKGVUknLA
jwINEAeLwpsLuBrIqfTIUxNP0dd+WKulSbzjUu+BNyQvJfGk5/tpGfwvhpye+CKTuEE5yoMJ0XCA
UFTA5hpJ/9hCEoIJBC+a+SrABkY/GJOtI05I/AMLjoC/EAxd6ZJT7cPRirmDgZjosZYiQDP2Db4w
yUtU2qg2ymid0aTW4xR+xZHpNp2k0D60rM7Ao9d8VBo/bDaSdyuCprzV7OmQlAhzZEDqBg2dTYgs
K0oFcV8Z/TCOWvYDAj8gg6FKTU5jZ5iHIMkZQLU8fqiBeo9m4X/JhRnyOgNMUSKXZErYE5Ls+MFc
9mXo+GikiTumD1LsMGXVA5lX1S4/nvmuR57gUZdatLzgTzNu/HrauQKE1HywjxHTd8C4uFdpZj5d
trIflhBR9XceC+9Tz9LoZ7OB2FjruhvwoITlYf9KxC130fFX2dTucj52Wh7pGhrN2Wb5hi1uPHyt
oMLL4/P8BktvzD9PV4ot0iHU1yCLO2eexjCPsRB/MbFuocEYVaDZOhEPrAcch8uhNHViPO3RbYAk
ypM/Y//7KN7aQr+XzzCzwdDAXQ4ks40A2EV1A0cmvB2tOCVYRH5+dUIx13tQmTXMToAEM+n1dEBF
4m81aiN4dui81v3O2FdF6MMHKgkvXV0+gOzQ1QlZw5UjjNiJ+xhHQGSYFQ2UOmq4FXTlDzClR3UH
Cui+21Du4Wy7Pv6ejuYOIqVV2vNoQdUmEJIABq0EO5AnHXnXzuX7NcHcLP42MEZwS3V6YHGN2qY6
kL2TxQYjUP2sXk+tK3SfabyLZB98Au29BbzFCwBfW6EJRLE+IBSVshASP1l/tx3EEV/N7VUx+T8e
AEqSDVK4fPF9YDJuZDgRTrDqlBUVI0gY7pT1sszRUfYfnGXFbN0WbDVF0YC0NzRTEdpBaezi0RNj
TC0o7iTyDPeww784edgvxI2ZAlb+YYj/7qBCbfyc7f0Rga5tYIp81Nkrx+AQaM9edAqN1D0YYnAk
4eyaohqmJ+6B00LNsHUcfmdLlk0usAKSkJdQNBsjONpRTuHQB4f3O9oqN+DTT4ba/Wj6JYT4jmID
D5tF3BoX4M6yeNaFXAM68gYyhQGNOrgZ76my3uQjqk8H0zJq10V7p78Cm/W55lBxAHSxetFWCds/
evpXF+ALhpeiofjOi27xdTSyXCTj6F9EajvSGG97CkuPTG3dd6odQX/pJzhUFQXLKEF5pUIafO2r
cBJqM0786ohjU81pPE4jwJMc/aXlEqlVI8pFd/6OMdtAaDjGCMhet2AOflo3Y64zBAaxlhq39xYu
2lCKlRgqZ9wiBOlj7F5XDy9sOXU5ykHsBLW22OSMrhmEAIoeE+TyLOcRH/YAWnJ4Hyep+xlyb9zr
OHMCeZyAbio6YJo09FR6SNGmmwSGyfGr8/onD+gFoGhe774E23MaC70uWKIPu46HZh6bxzo4diLc
CdPGqzsUFGjYsaXZS/fwPEJzFkPg9TUGfvfHBnDKgagr5btlWzBU/h25voLJYK2qokp5pX1uZS0q
inL0craMuVn0ynL7pWTpL/9TQ0SIR/AhfY1AaP4WK7hypcjch/ZFPZuFm7bv8m0WDfglASpHJbmw
cxXPoa5NpzvtVoTEC15Yhe6clweJrWdnCnQ/KrBn9IFSK0g0u8V0apGhJc4tpZ/R7Szh09MgmhTw
fHkJY7/z3k9B/MbETZgo7H13BEpbkA8fqlzGjmYtSpiyK6O/Dz4zGM4ikNK1ipoIDBKsl2BPe79U
DpB0osWigYCRM3gUYi2aQmPxphfg7ezvsDz6ZrDVzf1OAtf9h3LF2netPphLQ2NDO4JJNs6mkOIf
M1WJpdBlD6Wvr3nUUeUe9YrsSL6u6I2P0kdTr/jYPLOeYKg+1FWi6WZ1F+3dlj3DZpIGI6t9Q9zY
Tos4ML8ZBtSR2apOomFfRiFPHfpzfpleZGhGks+1mPbt5CbyEdU2FgQxQaJuheVuaWZy8I3HAfHw
LmHPLLxvkNIfrLZTTxSwY4n4SKriQYor+sP/3bm9olArDXbMCSpGYqh4xTKqlvLdMGc7oisnsOdB
x/JBrrNc+y40wcx+91el+Ksl5nuI4fwugPmoCzlWtbZzRQ635JlzuSmo6NV6x0YNHOZEkMFHYD9I
0MCcG4Fz8gH9+c0BezvzrFEfMbXmwuFkQmE5soTsRjtF01MlnVpRv3hCG8msf6S7OCS+mUqbjMkx
/16x8DJ8zxDb5jG5Wk9tj0DrhCNUP2qf+/IFKr43/zdXcRE/5ccMtMzw2j4LpqYSoF2u3OHFCdUb
Nw/doQc2tfFKy2INI5p5A+k/gDIxC+Upq+jxKbfvr9eKLBh684mggVjzI6WH0HddKGijPs4s38GA
xqge36wZIMytvwobwzK/4ZP3NJW3uiI9FrqbvglKv40nJBuLwjWumKpPFtqp1jmhI+/S9qRut3lZ
ywT/WiVCOb4J9itcUg5Kxf4kbGEOIZVgjD5IfOmBTatPRxJOhH5isqelq+C0B7+lqvgLnnHCtYVM
KRZ/JlE7wvJIq6p7feEhrGoDuNx/4Z1ih+K+Nyto+XAKTEzQTHutFQnJzU84sXm/esnDL/hcfk7y
yPvBSxarU5km+ScY7gVK8f6m0qfAkg9kK2rJX1yTADstxAC27x43x9oT4xOHpzVK5GZzBtfJS9C/
kccnJMZeTVsPbFAduftEanx+iJ+2ShSuGmOCHq7wVHiFu9jD4Tvdg2KIqASMHaVWvLf1poeOY84l
Th52v2iTQ4dNF+pu8630SBBIhwkEYlnlOcRm/I0CuYxXoxMCRgKLGR6KUXVZM5cQfbvshBZjtRrm
muDrQ0Ijg2ACco1/SzXFBtDZDNnGjJmW3vAENPPt9UtedO2O884kN3IyPTuUjDXqj5uLGQpCubN4
rkJMiTQXSvMFktNh8k8v13/XyIa+3KycErElZLvdG0fImEeS4kKhQ1MMe+RN3G7V/OCnNJ8pnNij
FlOA6l2U8EvCRbFosCl6Cg+hw/evZvquEUozRZU2h8x5QQZ6nGSQD3HB0AbZb7m6hy+9HJKOvdpA
HmIK+24RDSRk7klnS6bFYhN36quVtjFxGpv06m+puSudY9vSObsQGgmvKcrfex/UnO2zLA7cQMug
PmhL4h0ePo7bOAEM/YFh01tP9C4rrlpqq3/Dg7tYf24IeiWzHzdvZLZmbH25kMLCUUnalo4ACroe
5tXjAX3DoWEMUMEmtgHnHYOJYCDwTxc5QJntqz3oiF+Cufhb7K8YoOmdr4p7gcY5ktZeRcKIRb+f
jbtzfSG2loWyx/nSd1OXY1j0HID0pqxtV1qcovd/nERJbD8UAT7+gr/YYUjty7htuxH1FFiYqaxK
VUmVMpyBr83M6P+ico1NyVDPFsjz93bc/kVXuwT3Ul4dZKkTFGVhWpBk1B9+aLUVtBKyJcPHWArR
dWSynyH31pIq6RB8T7Se19o2jA6kd+6hLmT3Eiq3ELsenp8amRRWySglMUHhbTtNoHIsGui0Cmcd
Q78VkuhxuepNY/wDISAwyvDMJyTKTxo5Y68PaN4Z6ScSg3um+cOdMxvFGc7I9HxsGMY6zLbGQWBD
ng/GWgybPiIqybY5kjMuNtyYzOKbR7t8SkAxS0+HgZFk/FcJXzlJy7ohgS2KoBF/VZz86NWXWf15
m8TsUhYul7CYAfdL1+W0otOtufl3M39J0Tp+JBg+rY2wpfMT0xFuukoKLqz8YjirzVQ1W9BER4Jt
GdeQo2r/AFTkfXYQCpSPz8ZD2WtV/ZNx/CqOcv7M7uhDOrjBm3mlcoNgkyzfmL1QuSslTwLWd8o9
H18WA3IA4L5tQtW1pvY/A9KLeqkAPfyuuiI61XdBcb7r/T6UXiPgtRJSfjNBd7g7IaTQhrsipjVx
UxqdleKinaVAuC0XNe5AZm3yhsbrC7owEw5KklFR0rUYwus8HRqVAucEc0Lh2lr92XdVon1cK044
9eOoJC2VMM0SMBQcUS3fSfJzGdpM4EduB13pkZRp+O/jyfZpfQYu1OYaeCGFUwXXX+D3koReCeXw
PyCipnVqnX3jLDlg48eobR+KUwr71rtt7FvMky71QZeTtswzW6Of9WX18Tk2nQOamE58ybRv8xDr
V3AnJXkN/uooyG9cjJkepiQKfZ05Ebe5wL/1pTqe2h3NcwxnTCp692u4ct09LuVL1kCTU5sphWc6
oej2zulC7728tUdXPMvJ3czKKr6suxE30B9GUZpvujLapylF7s+a2eRUi16uv8isVgNMYBuC3IIN
uhDAU6GrHwT+RmUbyA3a+EZWmxR0aNFAFhnsZEt5Zp9Wr3NeiQi0NG61QqjyKqZy6jpuMcBvhvg/
iNTMmUtQXyEwl6KYXKh60+OTjuUCEy6BJJtfL+CWlzUdZJ4rgqaYyOdHiLertoJB8DesfK7mhqUL
VQiWOG4r1ZskMCQTPcejl0i2Dk4uaCvI46ckjd0MKCLUwM5fuFdIweQ0sSbNAbYO1tZ8ARB+E1Lf
YeCXiN+wBLoLO3GRrw3iSjJ3sUxILM3i7bdWVYkbuDWL8k/96Qp0Wn4h6WwHcM+y0kTOA5xRZsBC
AUokkFLgSJQz/JpXv6BwV0ZZnogp1yf1kmaKMw9Jo0QKtkFHolccV1FkxRTuJQIKtZkW/PeXnfw3
mNvejQ+lgqbUeE2BjVuDQPLmsLZWa7fLZNQR8wPg0Ar6LTnOCzt806lMbJ8Lt9nQ93Zb12UwQiml
HqV4KaFF48VN963zB2+EhdsUcKiou+KVDY8GtbpC8QzlAi0QYq4zwrrLQd4L2QGNvQboTPwmEMRg
MLG9Y1N/Y3inU3WTvRaArgqvuDktMEyPrkSR4zF5WwBmWAfU9HoDGB1WUBU9qIu61SI4SLzjFA1O
fsiWZluzxJ7wmY777PcAE0HvWxVfkOsUCjVpbOrJgkKT+mtvyOa3SdydpJZt4TaCdhoAH/QTp9xX
Dx3wMEGTGrv/JAJl637Rsqx2Bu0smd7ufW2VHh179i7SeY+BIfMmtUkvnCaO8XywCllCgqYFj2G4
27JvsYX1HWQ6gOTnnK91b29jRW9fUQatr5rDp76J7u9xNaOp0G6cgzGnr+9iLCe5l18yJbogqvzI
oTduekD6b/cS/JVDxvlBZ+fL/rNn/UQGzFpzmpgCkFecoLOqSizS4J5ot7BB4h+VUuGBQKsvIHJg
f/db3/gqc+FkLoL0klFDV7K/ELYPDHy3+K99OokD/ePcNyM3vwx7SWphxJi6mOo+Ry1y9jl2mr0B
dy3VfYWmxKb0EcG+4sbUJhl6ck4gixiQpu2Sgq71NdoZFYagm+TFIsWUI2WpQbhYd06lfLW5Sb4r
Iqy1k7l/aSlxJD4n8oqxnkoDMTQdzp/CxvSElHN7VDFvgKi+dYo45XlYVB49ZYKcFj4VD+J6D7a0
CVQRGobgKp1m9q/ctfR0Cb+RanIIxrFg8kSakJuQ+iiBh0zsGZItSdSO9Tk1OLCnCoqjjpm0CEI+
I99wR7rCenwsKkmEi76AhspXXAFP4bzYEEul3L18o6MAadVEVjKo/KyyCKWgkbXG0u+DHvgY+Nei
iSnST3waKIY9f0SHL8nwGr4vhEZGGFjtKWF0OORUhod1aZMnz+wXSJx/7/bLPsqHkzXW9VhcwtSl
aB+9ZvFUxA6K1NUkNSC481Pf05TN03OLUX92nobFj/8M/OoWxP2a2gj2qucc+jjs0Y1GIHn30b+2
rmG5kLSVQHbcsmKnnOqfCTF6QENSnXTwZ0nHadZj0Rvg42Ih9EvUnP2usc9QcURkeoyGm93Uy9wy
I4zGJZPARK8K5NW11Md/A+nJIuoAsLe0QHLesR8LKvr7UCpzwF3ccFaFeIUUE5Z+Eu68ob+bIwou
r1mNbSPlLWlv8XRLeDI8jiwEr8dGXGPiXLj9wduYb47Wb7F7sH7FOMHqxBj2fmA0G9yM2z794Z9Y
7BGX0yqPud5QOPe7BG0OdyGTsziPcgUjaKeDhkn1v6qYHwGL9rpJITm95hGLXPlxRts8KtRsUPaj
1AvQ1q1vN9kRmjZFlAlX96r2FDkpaj1IeO8x3rbHfGozwARcsxKBgQDQ56X0f+KPQFww/YK379XH
SjAMc/3nOHlEC9RdkH2EFbSyiq3EaNEBVaWLO4XZg/xWclrz/Bl3qf9WZfZcu4tgOvG5yb5r8u9g
9/7gh2pTrWKPazIMHdl7f09jRR564fNz0hJXZCAjE83sU0Fa+Qrb/R/mcBOJ+qbN3tZy1/o/DiPq
T6UntdLdxF7Xklm7hKaoFItCF3bTFR92jej+pokQPDulxPtIbZxFLpOCoRvUkz3NszHLOIcPS+Zd
jLjyx6uDu0+tcj8hhtZbbWEQWJS5Vdp6L388Y4+nTn3U2s/VnFYr8S5HFONp5RUQCZ+/gknsd5LF
4gfQGXXEtE1O5ledDDG0kGnyc3fv8xqEEI39EVwhW+BAOzoIC8p6kSRhtmGQWv2WPDl3/fDOkijK
SEq0NuKalq+r+I42xjH5pI6HALdIqmUhItdZN+3s2tBPpoyUnKfgzmxWDD1PrscuyogwkEGRlyAV
DUOOTr7zIH8xNqKd0Xdoph+Z7PsbfiGs4LQJCJHUA//nlO6zz5uVuIOE6iVk4M0nayzjHcqFet7q
ylrZksyWrw16/D5wV5Z0D5ijH4DVu9ju8QpV0yJFFwVw5xkbPFKnkLZ2h1VOneXH2FEKXFD+xcdP
uqZblvfYRKYmDNgLPXIZ+6/O1JfT0h5wh3xUqRi2U4v0JdRSSve6gL446XoYi2Lai+zmSxWWhI7t
Gq8OwS2toQ+UcVDKBRevq0CcJbJ68CSXuNvRUQWAC6pg+mEz9RHPJjo0wjE1yzyhoN5GNtYja5M4
Pe8+xdGFn1DJFBYQbO0FnChNtcauCllyy8POHJu9MtG93JMjLRC7LCsbXmOeTt19TbTL4LXaPEGX
sMAeSu/ntgGcREFE2xstF96O5nfAl0Ka0L2PAvN7byvcCGDiJX5H9BBDlaRryOg3VI5NZrePu5iF
+vJwyn+lQN9xE+oKEyernbVAsLASCKC3YJ1KJvvpU5a72iv+yZbI+CbnWFeSsxbyqZSOXpBFApBD
mif7YIp3KnTCBXriQYHZjuyPAkPF2UlOkNVs3rY2NtKlQAt/u0hRFRc5JCcRfhVRBVzQKHpvqkKF
L4Xzu9F0yCzonx4YTt0gTQB3EYxPzyA1PDfc7GWqVDSG18W/gtP7tSb/lnqRywDx+s7CylcWDO7c
3pN6K7dZAMn+JyYjCYYGZYcgS2gWY5KWSRLAnAGq52paLLWgbhn0+LaPwsKWtPZbluOKNl62hKY4
opP2SVM90zG/ZzngqhtcEksA37UO4vihq+AebTa3/Ke00C1ve0Xh98+tzOI/ovsET+gs1BsHdxyY
vTTqxe1aEd5M3oAfzuktXJmfLJSEfpWtTjfXBG2B5DeeRlxs7ZE/Bi2SyzcM6VSWwlPjKmxDI1Oj
0ttVnYEb+9KvDxhOJt9yonQsGFm7a9xWhq4eq5L0Ge7653rPciHh2F30auohN5bkeQtxRHUG8B2L
/4T1MyxWkObU/Fbka3gaghafMvSIXm+Hcgl0PjSkgLeeL6fdpjFFQX6g1rQ41pDxRbNrJp97W82N
fA9KnUvpdzzD2is6VPCoTYHWdSqJx13SxAYW7M92AUQgNG7/Q7PsKiYNzg2T0eoaJp6klyLbjOd9
zoKQ4fDlrssZJatLHeGhhWNkQLWHrcUupA8ga11p2OHbA1yhe9UD0vAZ0i9dIhxBhUcagEbTyBZv
NoBuEUq+TQT9szIF4zmrVEgmeJPMDcpgKGMsh1GPQMDua/dFh2Fc63L1Fh01i3DVD79hk+oAEaAx
WKTGWUsn1f63H9zRZROE5lzDVPHOqJVcbxUaUaR6OtiwW+NU6YaQG4sG6PN4wYdZItTmxEPvjrH7
O6fCw8tCx1L7vYXTAwTtF+PgifoyqjId+tdG888cq90LwInwM902j9rdlbm+eIm5oxlwSi+s/RpS
bGHh6yZuuwxVdkImJQjp1BnRj+x5u0t2QJSKKYe0WVzqhdPDRSDvdG4UaKUprqEZz6qbnSeDWrP8
eiqUBlph7Ie9tTftprIOGwyl4qhxWbZxZCyPVPZdKrLRpfQQTUcapDbfcN5WxtDeuysLRNExLMJa
HBB4GVzQWV8Tqs2Z2GwlUUVdGPKzKWiRLlu/o7F1OtmVoXKxhT0jteLdtt5LwNd2BagDVvPFkOrd
apCvQTNDenQSeGRnYvH86IbRc8clDRX1yhBObL2Q16Bsqn0e7ui8KJVCftoB1lV0o00lAGh16yMg
a67PkxuQcMuW7tU18d1ZQfNIZm16OO5p1Mk2govCZt1tKlVhAK8yLLsKnwSYLwHeH0ndAcVWvp1+
EZ1UBjPdGbMgTAF0nblW5CD2zByk0HI16DH5x7dCc3Fuw2jSkkdw3X/zhUhGoqjwxC4BAbKGuTx4
UgcSHs20x13OAjw9n+kyq+W6cXVgbTtFQzgMveR+uRniWmMo+TLsU1/gvvcbuyyAFhMplUCT0f1e
A1y8oiJoL7xjh3Z903mUnnZ4v0hAtEShzyaZPrq8y/uFm7+qykMr9Z0DYXb1TWPWw2wY22xMnt5K
C1Kk1lDnhfqAUjAlOE7n5g71Uff9ErYaXjozBQHUmGvtrLQCn9OO6B+47MXsrdQLBjVWPrY/c9BI
50juAosYF6XzbERPF3ylRtqbHGhkGvArh8L+5r+AikN5Kxf5ziilr/G1WxEK9ECf4V0fP3mbeJMy
/zOdLwZLmgyHtG/0nnFIGg/fuhVGhEN5gH8H7pAetaNA48jGvZ+LW5+RNbebXqGpM7WQxCL8yYTG
7dx3+iRKhQOEoihmEjw1Lh9fOdXPo0wLFI5U8UVzzGtABA6+Q6hnKGlf3twwUbxQvRYP7JlZppM2
zyLZLSKrN1BvYH/FsA9yy6NhNCCTkK9nwN84tEjJFhYKmvB+TxdHvQoSaghkKPv9+daKZL3YTmdE
rLPy1L8301/bA+kXYCE4wsmaoICtJVvrtswgZ6FAVF0pXD36dZ/B7XWnxWLVVvInf8PV86eRoVMn
ZzUXscVcd31ql8868uNgImVV75xdtsiSHPM30GBJWfXuRyuBhNnNJpM8D1R3ZS20OkvrE47SHKIy
otqBKVrci+K75TmHTdBO0g87/Uajp/MxlGXkc8K1mzyzDOHT4VEyt168ojgzVAXFv5D+U8VpFAPX
MZzwYv02sle2xPumJTPeE5FnLsrsJOKAv0urjyyFUWyiakiKJpQ6f8LMi9hhMmnoHPrEdjiFuBV6
CRIW0gX1+V7IQORGL1hIY7mJn/BeZrXsoULX32anR/gOVWgmHTu8PdpHWF/EeTUx6o9DiYRyNlpu
YxjJG5KSK0aAKbYAzV5IISQMIua5Pr4tXt+S5Ouu1cu/wkOcowukfFsxyEybTYfZy5Lgwy/Z4lPP
IZEqFIhqa9eNWSbbJtO3hjsDthrpeDbD2W4LunkzsaNqgM2+4+KoR0Wk0vj4rrmly2Us7r1v3XBW
t4XJbiN2T0bVrG1rMbkFXX7IVeGL2lKUBeAoUKlj/2JfZ4VAuPdJQ/xNqZ7ORKSScEa4pbccsp8m
kMnbSRTgeIDL553Oc2u1RptVPPD5eb7mnhecMhVvCItL9tJa0UbczJQllVNFJWmweR04f5+VIbTp
G6YeEK+9mrEOtwi9/hGYT9qNqYLl07mI+hmw6W/ui/QN4dBMR71Cf3x+V/9hN3G126Nv/2R4ITs2
Q5uPuOIPzjmuFLSXIms67Sx1JYoQrYVZ3qZzPBo6asQv/8yCU5pQ2uGM2Kpvtjs56dr/FSXpk+Tr
usQuat6x3sp20tIN9hZovLCWCztVRb0enNnbbx64clZ9lWiEWcChxOK7ncSmjdVYYCRLkSk2Oc04
Cg5vCmYGbDxrp4e7ZTx6m59kgq7C9kPqcxOYuUdLQxum/4DIIf693mt6EBdS05XVoIRl6dt97k5m
koh0utSmAvslCsfnQw8OPs195zQzxGjcNrUoYwQLuRQJCP+5uOwf0lLUYyGzXr0w5w2ESU7aEvWG
Xdby0S34rB8HXEBy+OT5jDYyZbbqMlwCUo6T2RvKcuKor0nm8coLda4M2UR0OiYgOGYMqtjHIJI4
1iHpS1sxoXPBPe93cEEZtBiqfpiuE2G6kygwrrhcIuJxwIX45VWRZFt5ePAiDgcnM82Lhd2FDVw8
Z2znTXK6BA3iturt4GYfTPVSaX+mybe1QJRbbqsiY6dRW7mxEMBlEPGm3DHqtZzCPLSJs5n04y1S
00Hf1kxVqzcEnAkbmyWTWK6DUxRgfoMnz1Q6HRPcCcPtBiqr/9S2tM3Ct8afXE04fcMW/zXKN2LH
qdvi5NumAH+0mEqC2FQE6TqhlrYTF2jL2ycW4iRJorZ9/My+uaBiKuwOMs1vOJZr2VQoen/PzpUE
a7sXDLBh7difsAebSirbHxWpOANgCiuqd2KFR32PLgAUGflPFPyWUoIHJdnsFFxBB/CI95dq7l5U
yxoF3hLYAZLCrrr29UvQ3pi7pVQSrDWXzhwkPmOrQLJZM8JU67oOXvhdhjLT8U3jkJCANdODMM27
9wH6jqTyd/KVAH8L1rj7NLYeW2dBKVh7z0yK1NreZAvIBjALW5ec8RZ2rdq/9/PVS+RmZLnRSOcf
d5eB/rKmW5Ha+wcwFqANTiZKTQSecIQBABIK/xj9jkG09JuW6hkTfXtsz0oCQXz4YaiyO1z/zUJu
OpTSJw7qAutVs+3Lb7prfPZH6Dgv4pt2cGVBnvTM7cNHPRsXOYyMiuw7Lomm8+NYCFk/cE1wMlaw
DL1gf3wmk/0gAo0AjZePQuk+dNXl3LcZ+wfEU7Wcx5oaIf1sg1suwdkLk4YEdAenl3x7iJ9iHVNp
JWeNvso3G+A1UwoOGZSiH69ak8QSrqHHDo0yRJFDSXAMmz9XYro4ZuN+h+sN3Y0uV820q7jgHbap
jyTotH21LP/y69rkkB9DaWZ0i4MDvnKo9RcnZt1f3/BBY7yo6IRoYAnEulL16T52jRusZDKXtsTZ
B1Lkc4CgB9x1qaalArWS/3TbTxaqav5rwd6SpzVZ8HdilgKUyWHS3YY56QGPQKfez7L8yvafasoJ
BBZRyLWQvSFRO3MopFzLHhPv/PC9PxSlVu4R6S0ijdBJOTKI+9obPqK+ChGMNcrnNitjyhhC3jRT
c13zdXui75l2VoZQgxoTRgOn4JhJvMED3DinQnPDaGIlvtY/fv0ALMpvsySzIj1pNbAW5CVcRln0
Z6o/jvdPDsP3izcgle03R11IS3zeUUdjcCveEHRvQ31gmDtyCHmWI4xRUuHxHszNLSUVnn0wvThz
dD9i+m7TcGQpasAMrVFHnJeIAeSotbk6z//wS8iz8lSPAqfyrG818Arz1zOGl8huqEI7TfhZ17bJ
7mpYE+2UtxFXEGBxuLtMp17NoB4xY2u5btNI6Rm72QdUYWu+yoKImxO4+NAHIkLfmAuISEs08PzD
7jWYOXA8w2xljmtNRO4fNd1LlQuqwdGwznOp35DxQVRfMcMjI2cCq8/mEURDian287u7g0Ejs+UY
As3NhpmoxJIXW/Hfl4H/I+P9sJe9UcsAZz6B4EEEp067AKEBjKhNa1nc6VLWoEE4tG4vPN3NFrk/
s/ozBRsDNvBrX1HdkhXDMGWmyNfEPg8DJaIRKBWN4+iUVKDf1Awo2/uUUH9+1DwYZlzFAQGJptPn
tluKNb9kdbWRU3r6/hUgLyY7dBWuBZP7kVx3sOP2VFkNj7sfK4qokq6DyRSPKio8+EupGYZdRXsw
9jTYr/MYbxfOUZVoXY0if+twHuF3DAmGLuO+HhwiFrek6+iipw9MeLQPSSIUf+9KndDlxETUxTXg
HbXeUjYdsNz0hAAKF1vFthO3dvdyUJbB1XttKcOvdt3THWUenDomnZfeJgPRl6qR5odMPwrnEqQr
etoTN4GrrP7JapF07ClXZLAKOF+UEVq/b9T9cp5sY6fklJyz9ji37yowgcKv1eCb2mqVwo9ECAJR
2bOdnYtrZJ3LScACkHWJZNSBh7eWM2ZFYDVvgM01V9P3swcyjUnxEZC51vnmF5TlZrpM3fNI258A
sMt045e+1v7hqEyyYj9bkzzIgIax547xWt3i2zsoQeosH4e0e/lFyx/XL31XKy7zgOksWkUc/WuC
OXLvzTS2dZwh0gQy3pkMxmsHLejF5VN58kIVwpUBR3fhdbyh2zz2a0V9AXKZXUqKtQ48v/Z2rt7Q
7lvTmKU97UxsVu9iOnChdcN3+zZdixHZbwgRRMeqRXo2aWtYz3Oa+BV14pK9HArKoTsHt5S9+BF/
hzYeodUAp0awzgBcpsZa7wfeHN6yBsRUD6ufFq5jPJJNrTjAg84Mx7L1V7paWQR/xiIzfQjv+EzH
u8nqbeyZQwCeGx1CFvNaFLAfElBp7xn1O12gwfg3eA15AgfzQwftJC+e9CKG1qmoaqqBAl6kiyFm
j5Z1KWloLsH2OcGEwgIZIpprxV1PLKo5DCIKC2UshHwunaBonr+skPbi67arxv9y+8/ISDPX4S9w
IxEYc/LT76pGVH6rSSIEbaXQYZUHuMcAOAhkGa/H7snrKwMbG0WtaWUj85w21JyJaM0iNwybiNgt
0gwP6CnDIKR5vnGDU39yT1dJO9r3B97H94EZ2nNAUG14qZY2WbgXWq8vo6SbWFOW/L8ALi2lXoT6
bNOcWObh4AQ6OIvY4TKO4jg6bOLZZchJFtRUce8BZU+/aDHjV7YarS0AKsta1TRbQQ6Z11oY+sIj
9YMGiIF/oOtirxVYWCPG8RFOkU7x6KOmanEljXzWuZwQYvG1E1cxBxZdg+Ppjn03FWzafxYr6w6p
zS3gxLA30TiXkdtGDXLN3IWLJe1YzuCYUlSx2t18stSrvsfwG1moMtBtk5tndtoRbt3ZvHIRtsHu
M7I4mwITH/UB8Jynwajag8euQNryIjgO1nMvaTm0a4UML+vMCogHce6/0YuCqvSqPhF0Yym4T/64
1z+DW5J2mkZp3I2CKlS0pZfIT9a9jBhHiSrIj710xtcxI2kbL32dvO5eMozgxvgoCA7AF5GK/oMo
fW9CZ2aMUP129DRI9ZSVbb8982egKE9Xp9rDFO+L5x8WfUY5YyAkuDi16JsA955J/9MDpny+Qurk
FzfmtcGel1uR4WZ1Lh5AgqPfhHVhtMLej20XmLUke7N0kySMguqf6SuXBY+oFShbKnCFjpbHTofb
XE2Qd9mNXkveK+STN6DteCdYlkj0X4kUfjNzDj7u1bC3w3YhV5i7ZmuKeLkj0Wk1sIy1BxVrFnzj
XbvNLgr3zKqfe8WWYZscU1N34/4vfDgqilodLDDMeC2c1ykiwkbBKW94oil6tCZgOUKGt4PYLJYO
ZuXDccrQWHlAoajPVS4C17MQIpwFstm9OxXwNpBJQyqisgiAGkOHIiMRAvTQa4L68trPqhUMF2TF
k4Ssc7wn28ntTGwxnHhOLdk3QRShE3wUx3KKw3lLbi0/9WYGSyDJykEg+AcvOSUtSEPb7JWHoGlD
OdwWAZNGJnDF6LtxuHs/fmxXon2d7XZFLlQ28wqpvdP1kNmLbQYen1T6oUfumv62hOCaKV+7Gdw2
GHGTjHuiVohylP8qAFaHV3H7SNNZ2kukbUgDUROZrVt85bKeofdsNZZcHy/dMYexBLrUVfiBokwZ
tWyTnpQJWxePkCp8dnvISskTFpINxT3aU8mJJu3f4rE9LETc8VSDxPMG6cXZgyzC8yATZ+48ogKL
eF6wDc2mUWIf6uK7/+Eb7OjuxvS6j5AjajiYCKS+7ywArCBbYNkdo/6FdCpttrCqbhud8PfFpc/8
gmHFR2AAyvGFRao2zI7zZnOPLyW2yceCPtk6vW7e59NC83V4mN6iraWjWa5+PISW2DYNznWiO5y3
G40hzq3NbG/1jFQJYWpDEgTRKpKqAgRF8r5g9+Z24rMJC9h8JmwOk+1IkkM4Hp58/5s+LoEjF+WY
wkME95ruiSLvedSH0q/QIiKzBNNsXW7VfuZw28iki4gUaYuDm+sXZS3wskiQCtHOhUO8qPMKOOzj
MIevxAI0GOKO2mMVNFLhOFbSSV2hJfQ51PF9iazBI5WyN3kyRlAMVKw7I2zyG2kqZ3Czk/FMfCsX
SvcIhwXqRusWngfm8JklEgdBfsUMpGSrDIHAsM6QsT9LzF94/9AlocbAh5iqD/lmuuQCZes9kn1h
XRBICxqwbFLaFcGT73v/XRL4WIcgDgYyBiEdoue4ZPhjriswhCxznfFVzdVBOe/x/072ZhH5zkVV
xyyKpe1JsN0GWTBySCMsAwvlQp/CLRSGYq1Kj5gT+1NCdhfsdnWR3AAFoevONegfeKREGmfF9gn5
Fzb2hSif/wVePsnmLWGLcUUBENMnK25m4lEsAo25gHMZJehtDMYpwrWbtZtbZKAxDoWsbuWsVE8m
7lF1owkNutdCKR8lJGwG27fm7axb6wmhXbd5/G7pAn/C2GdtFQaWT3pt46tb8i1atmi/iq1zHSzK
VyHScjosbfTRwyoS9h6aDbfReagzr7jVVLRekVfPRf7qyjTQkQdlMdic5uotfaCrRNaMmz/LK/JC
QwLHyuHrH+sXAk1iU/Yzjwq/oO+Z7M2+KjwHOpcnCpSiB21YUGB1WJqzZVQOqBeqKyVRmLytJdt5
S8wtEEKo9XaiyUblagdqjqV2J0xJUXoUEyWMs2PKgXC2BGCOdHMoUXanGTfHvGTe8qc6Tv9IaQRP
dZs+gz+bjgj2ww6xc0qE+0sIsu0Z6k+JEFwv1C9WPhI3VEKt4Z6NpVRkq1c5oKExKgL0YDd432Fm
3vYY8kH3VyP+W3pkiT/NMkVK1Z67ZR0Jgnj+aYxnG1CjqG7rs8IAhhz6XEq7CowFTMTRZSCZbJPa
xmQZFJn4G7RQYzV/mSk4/n8ZDcHznc61mK7tn0d0OWt44QadepI0usioLe10f4e+68dCR9+29Gg3
QpM/x/SMQHpM9fPaMYqBYzzhGTJNUsUfKn2fzyWZkHS8PUqsZvkNb3Nh/QpSa/OjeV1V2F49z1CR
Z06on8uuuSKntIYsoUykYX1VRsSEAIS6pQh76hiJL5Ay7dYWIQlfLny6TlmxiIira+XNFcQDQxZJ
gX/AAxXsQCFCtTEV9U5IaF12x3A3CeK+yojbCBEt1/QR2T3Pbp1adA2Sbb4oIJnJBpLzfM4vhbQj
6wrG4TwBvmqDJS7P/2Ygv/vGzrICj7RD8ADJDS3WqN6zDVf5mvk1wZFXvjg+fDRSe4/5cejJt3kO
kU0VYThNC/BUzyIGjdAgF9W32LTYipf255wvxpuBf4cVloDGGPG9dmjJVxVeBrCj3rn0+F223M0S
WsBGsYFGRDvC6BmLR/qIY2x0UP4F5m1HDa8OMm2KLQC+gJA8yenyVMxtQ63prXDIiYMo5lCWAKRr
xrEjnAR9N6CB6YxuS9yF14xZ74xzzxsSSBGQ9hAhDCKYbRSzRgmzOoCEhFzbcy8Jwk8HqFc0olo1
LKEKInrGZZSSXuSJ7251mm2fH2lmziIIZF5GLCUsHnkbO7VdmL5kuQphqqlRbv3LKukBlTCoXGKC
EfrV6uj3A3QtHB4JtvCdHh8UJ89WFXQGADsquHJorm9iMV7n3fJ3qT6Y1Mt5tlV0utK57m5o1XTf
bFz1AVILc0Fla8/zZhUdrCS4UbUZiBiuCXFQXjd+8skfM7DwqHnSmXJk3te6KU0V9BP15f6jOw99
Q/RFJqrHq7xLy9AB0qB43AgVeP+CRN3DEQt8swiJxV7DDX8sXb7I4Q9B7chjWa0mh6jT1EYN9FKD
W7eQCBlRLj0k80QZbKblm98Vs8v+3mXqWGlcGn8aBf6FIQK+CrYXXJJI98RnSa/lOufCIbohncz6
AMivX76evayZmvOMlbhjqkb8DaKzWDHoGBYkVpiO2kGA1GbY4kLQ7jfK33HSGzUqf4uSYn3nnfuX
MidwOnInAvG13zB+hqytOmX00rkXEacbbnZ8dGKFAlf/S8e7b1uB0OBvrc8M0ZuIowIBD0FbOjat
XJl8Y7SdxHgnWizg1T8gXwc99Ia+bJvwRSGC8QI94kdQpH83HSlw0go5lcN725H7gxAJejbQmT4P
jOoz/UN91NQEigBnflhmD7NQ/AubZs6pgT4AQ4Whq+gYgYjtcApkrHz4avWxCaw1dbJ5oHXv5QAd
4Fq6Z6AZjBjNMhfNRMC71mKqEFfFuZ7l8HZzWWzpaX81VmloA070zSX4RqpdW8u8Msw3ClSecUax
hpNTFyjtVBCeiKxpVS0S6lwX7K8KGpuVGSFb0Ns/H5ZwYIop/JGthCHlNeGGhBdf48vj6zp/hvQ6
w4Npemvb4y9w/klzj6QA9Rx/duRC6fnlD+WUpejfc2xF31DQeKRPNxIebu+AVOPNIHLSA4Xhri2L
SActCqrDjWh5JlKpCOlrK10QOE5BhdgNiTnbD448/gFGTAhHS6fRJkJlZDrEu6qWqgx+I5UKF1XP
ThMotGDbmcjla6fYd51i3jqfINv/WZSEYpOjhJ5ir6Uz3OBBnbunsM8+JCHH3ieiMPa7tnHcW99m
zE4zeWzzdV4GvaQ0hcd6XCVKKD50qbg0mcSniTMQ2I+8nH1nPqLXmCwnOR0QJlBqN+RQaBSJp6n8
4UlaYuryUQ/tT7siZ+leSA7GtoF/UVTGqSrx5DlBXJDwQvs1OjCtO+QMelaAHYPmdzngM3tpTrkZ
3Gv/Hdc+CheoiczeEI3alTNZUQzncUjdcU1HYPlibgWqUp/2BEuEfhoNQDV+BOhp7Syd+bFcRk8n
gOjuJ0ljjqdAMd67kjaUFZ+IacQr/VeQbplL+hHaKG34ZT6VugFwsgB7SQAq8XM5joTqKFlVkhSm
ra8y4LIjYyBhpRM4Ab3gd1JX+6k48ShgqH5VMi9CEjw5nFmWU3T+T12/evS19VwjLVTMwLS6Up9Z
020eeW1mi2vBfk3zjRKgrQwO3tnYZWqESrh5p+HQwT5tNEqEqiGErryxyf24kQn7pUfJTojzgBRo
/8lqOLrkckO9vUmSx59qYD1SbRZsaIRGoie16y6YQRbQ3ShwYcklY8Q0lO6Pz+kOcurORQWa9Z1e
ffz+QkBOzNh8iB6tD4fMgMwBri7eLBkBmUNCLrk4YcE1G4oblv1vxXD/OZrUixEnu42N5K0D2Eek
SI7/T9D2B6ejK8lO2ps63C2M/1dEQGAE1ONVXG7zjp+pJmSI40/wBAFWFC2A26fV36SeDem2mTSE
qjp1hAUUPdp6vnkqfa2UGZ9lq79/TnqHna4en6D471HuT7FXB01KvUuqy7V1ze5szH3uVxDTBoMO
qfRjY5ddDDFb4CjIsRxVgf0yUny1tQAh0jBqJowcR0MkHQ7TnXy0OneD2vznEtGGArl1VGjn7+YG
Z5Vir4GO7rpO1w5vjFfC4437PCATuzznjwEQj02HXCFmENP1AnQPCxTtZJIkTA7wt2zGzYMbD1LV
bnsSuh5uWgt/92qD6qxl0KS8vMVYfdSf7mLQvS4HjB0o124HbrXBrpmxPQymvJAIookUgERx12ow
PVuFySR9HJP4Fxd3gotC1WWfWGmflP7RF+VmCLlg3sX3BMEEcCLcdGaXB/QZ/8OQy8wIVj5OlfXW
sEUoCM16smkxPnYScTpv3isv9FEXyObShVxTr23SDLqm1jWHcz3oF7Supaf2heZOhCrRjW6IQLKl
j5O2D4RzQNleray1ISAdBQlxRwR/Dov/3LoyrbmToW5eWdRN6/fJTIjtcgQwkY6n7P1/nxgfivIS
tx6zFp25uMDWZHE5hXm7FIZTrLSRhRL7tYZawQn+8HGw3qTX4wRICCRmiSM6tvNsSBkyGXrxKDIt
RSXASj2KKiJVnsl/CChakdlJ+U09oy/AeDbgP/j+2bIpvG9Moi3OXluC0wjrEs4RlFQGIk8cN/RV
qSdFN1zUBXStHFIbmySgkOb/QJnQR8djTJKcHcnE/WSy6lP37M291pUHnLDC2Ks+t4Aos2dPAONf
C9FyySsaP8WUdt3/lIHXBdHWGWSnjmrP/tHJdlJYIYB+BLRjW5Kg5vwkpDTbOGnMtLGO6PW1GDAt
q/LldEUT67YIA/pBZo8788mo5s3/HE2W0Lxpxa6En0qwQSpyAgKULrtv8czYydCkpzb89x6jypJ5
AghpT5YUVimLEj/D0dZFrQAZNR7Rqy8Tkl8PEd51+SycO17NdZGDv5hnlID9ZKe4OKxaMdIpYLZs
z5A/7Y7es+Yq11MYsHjY2FF+COWaFyB84EZ3Qci8w9zhgPE/n34+PpmTaTgT6Co99MgxRZeENKZI
MCtJ5s9mCmcgt/2AHlLxFJsZrcCGqchGTomco22zC6BUyhVWYPzpl6AVrW02kZReyIgjx/lwxqij
zt7fUHo4Eadgmdq2+UBon+1JfIwG25iF+EQRJqx/DX/tI1GunFKBCt0WdTJ5F5/C+mDT4Se5G2AS
7YdgPzStZOE+2PBS9Q77M6alG0ByvmK1RsgoCMr78FNbsJJ1KMfAo9XP/OPPUwx4KY6uNCG13R0e
wAvGd1P5KmJXDjU4LaST7bqWUFL0J4aPUCPh3SSGuDkktz6sP19WAqhSNNCAdNTXY50m03YwaZ1/
OAJEx8HB9UTBErbz7KlrjEIY5WGhxyZiWcoGzbZJZTXd5HamAmu2rsWfoAIey31W7dpIFVFH6rrQ
S4Jk1y2blFkUnjBSn74D0nmYMuxakL9iRRi6QJKCnuGH5okO/DGiIHvFHAv1KyVm6a5lK/x+Xa71
+wGfnl/tSZk3jHOcG0WXGXf7iANDdoKjmQtz6A5o+dJxSJSfqadL0XV9+nnFEYUMGecin7Hie7VA
gaODFbxnJuRjcQVVKZFAc1U2rMcyh93S1lmvtkgzHNXjjlkX+GUFDYqG9zVkT7dr37h9t5u3UKhY
2aQ9mJAejZXwkfM+I3Kh5mvUygKYmpiiLlZJdXQq2HcxF3BjTPdt1QsVH6vVeDDQ90PaE4l5FVSF
B64YlQjJvxHa6qg388Ev4E/huXcwvv2PlFAbTc1ZLeQpiIGlWZ7j3Wf0/bMrKk7xaBmWg7sbP82j
GU/Prm462VUCEfm7MCUoB4phU+T0EJjBOqpkK21neDvP6rWUKG0p9h7W+ZK/HvDrzBmkTJbUU27L
tFeghSRhuMJINyPNyON0WXG2bFoG3qY+CyxKY74mrxaXAHZ/lSQmTIu5iZy7ctNwW15pigwqJypw
ylTA+clzvLjdrgnJNQ7xFCCpumKPDiO8foOfT2PsDI1RV8MMDhshqeifZAXzA2+tb4EyMAoJAntk
W8CpwD/XeleCiKci5zf/NWQT1ZEYpCw/CYbZcoyzmESneuWJs5iNn4rWoD2v+4ddrDO0mKG+zukS
xILHixB+QASFBgOyE31C+r1XmARY4diWqszg3OvBBeiFtDEJX3yziQHLcmt63bNU2M1XEW4/78dL
EHEnPp4brXwFQH8cj/RhQCLSSEuSDqo4DQallhXf1D/CHNAJf4q0+yFUwCcumGh5t7hK9OKrCgai
Cz4Z+KSFIVN8pTEmCXQNs/CsLrd7fr0xSdDeopu+X3kye1IlPqx/Vjb9k/vRi1U4Jmd0LoDS1S9x
9/4gL0hLWBaOqyo2KX4advLCDkuDFzwNc/tEuwIzVS5AxFGnxQLjSBXq+1DvAEn/BF5HmskS2C5m
gehnJDdI0P7hch5UqZVX6vEilZqARqZQRGW+bysNPc6Ka157PYkUHLmCWUy6ewfvAp2URxBfBrEo
tfDILYwWM6QBt8BLlmW7wsRbLMSsb6uuskAli+QpHeIn+89raD65HjrfOcdPhF4cVKxlzsfvvwYs
B6kcv6IYj23tIZlq5gjTNISF3zZ3FykQeCtT5j6cp0IzpweyjfLwursmTQFQZFotsX4ST8o8PF24
/u3Y5MGUBFTjCu7800c9UNnoQeV9ZCuJ2B7ffNsA1Ua1VvzibFroiCExB6EQT0TWxWQsS+FMQjHc
IIwU/g3tKNaLE836erX+yGCpejFX+XoxJTk/kTOvFJ7kIWv+Q75x08t0b1RqeuP3K0A13GsvdejR
VC0YWMccfO9ms0hborIlwQwXre768kdlZkNbZPsS9Vo949kXtxX9VQIWk68hbvvvUtaHvGbjwZVo
23RK/9QRpKabakH9iU1xsHH7aVvHQDb5sz1qcvx7iEWFYUl7UYH6/MBaWKBWrKPjEF/c48zEdX2j
nY0JUS8MnotTCCpJKpEO0O48Uq13EFQ68bY2WS0zKzx2y0Vge1WX1+c7M6g4/LY8flVrSvCNUXoo
wcU0+ZsrssKUnVRwAWIYcwx1H2eNEgWAf3p93792aD3foRYFmh0Mi/upBV2t+wxJ0ViPAtSAwh3J
FO4yMGiPnBizKnu+Ju+Y9kr+mXd9Fk/DF2+bfPasEGjA3Dlp+B7bQoOW9O+71cIYa6Ji1OxAW2fR
11wpSxe/H8kIdi3bqho7K3f9H0KItSzMGizoYIM5qZ3Jlrjp1wLw6d+69EVPYcyi8hRVw6SzejQD
oN5tI4lgunVbC3jcFFtxD40kGXwzWp0xtEXWRQQ4W55h1KZKriAcUsVJ1nV/sxaQfoP/bJLefdYi
k3S67Fh/29AwUm9zQe1FCi1nDhy2PokTV0eXi2uN6AGJLjXByps1h93rmL1LJHs7EjgZhxRLJ1Jj
lp7NKjI7/K7S6c8rU8Vmz2nUfD9eKki/n829KAO1CVFOPpjIqZ2leghfrHTXKAipABAwmiTvSmF5
SSUR/r8lVQni0GKBvfhQaa3tjEH2yrSAYRuUUfV76IcqEAmf5SdqqfTK4Z5dIlM6H6VonpnFxy/f
/1FNA5ZxaZZ/utCG4xRcWWYi9OZ/wOikGi7tXw6J8IpTafGd42wrB4K5XAGuKbp1mhqs9+bUHxQ1
XHqVHVNwlhYa2c/y27LQjnniuOJ6/ItFqbNpiNafr5tMjT442NZjah2FhpM8Zy5IKyPfnwWPtoY9
yyTN2k1OFDRZxg8shtagw/ewD4MqbmbMIbT47elxNEfYRa3KOYE2tOuRZNhWOMbxk4j1Cg/StaGE
xmRKCuG/sbeevH4auBRbh1svYCpAyowaH5klfDhT4LUZvr+CPQje/228qaM5W3BGzdQz/KxVmF5E
2hgbHdxwBqf2LLdZd/ehHyje3YPA1BPNbGmBnRcNJ9FnTXxWDcDK/+lVUo5mO8kS5KWvUGVmVA/m
RovCXk43j/kneN4zJzu/3A2tfYZ3UwXYlrSRrcNDQVJ5KwHfPowcl7wYqut6kAOvTHRK/mskWvhB
FO74PeHdKCAwH70nx/Z3pg+cREjWge30G+Jj8XCQdv2S70IKXfppz4szxfYMR3PbDIcDoKY2zE92
aNVy7bisx+IJiUtKW0WP6zo9kIIc3f5jahKp/6wWqXwZ1hPv+8t2A+ndy8AF9cSEtUooMZi6E9tC
QZTwZfYh+bgSNO/+TGn1dbJfy9cFh2R31NhTg1JbmN2JA8Zv45tNTejVrZA6XTCYUd3IBnuwaaS0
6iqTaUxirQBxKJKTeyqwtB8mliii+LbQxU0aq+4PJSu1DF2qQXc+Gnc4KDUZ2ZjqVtLDmZxSpFmB
u2tFQxR/3/W99GnJFkzA8/OQmYybVRbiRkNAkikiTPLm7OCQwRVfqel3KzZ+g9rT6di1/9fKOZUH
3PTyrcHYBv8E1ZOaOQ7p0fxlqt43NXfFrl9e5cShR6GPuhnt7DkBKmPlQbH1qhefI9qqRdbh0p1d
Axx5yXAPOGrTfCjfhh625C6VcSxlxtWQjBqPuHO671DpagRsRdtstCpkgbh+LoYTeR3BQddA7yBi
8ZdJbw0L1BYzzoth/HcEdNRuG6EXWdpCz84szemgZA69AqYGVi2Ws/Y19TJLpSJZDKUI4YLjKOei
31M4XgNOBEzDtExYkxU7jjR2B82rla6WcFNii3boSBDbvkrlmj5u331XEWPSE20qi77bx2uGeG60
kNrwA63+Vz/jEvIelOTMCepTy7v7iMhhWYNkKtqLVLm5gJ72doaaEqKbsFhupHiUXTmhL/fr+cP4
/8x/UqYkZPO70E1XrAuci1lgU1108QVe81VDIotfDJbHgVy0iW9Olahojg2aaa8R/pKKmewoB8sU
DcND0PbV9yHzERNOQJuMxR3W9hf1zymNrj3CwZQGig8bkUA75d/12EWLgkrnxLStrzozvXDmq9Dl
USARKz+Wd7hZjD1nxozKLAG3OiZOmBhUAa1nTp3OeLT4L+qOOVsL+T0D61NJFJlPWRh2AeLq0wEL
evWt9Styg4KYmOZDrJpUzS8ii0ShE6sqvVWYnsbuQ3W3otRZVPXbwnmnw3Yeu4RyrKBxdUq66HNW
mbrboNmd6QA9Awv4/19nMiQvmaw2R4Ttsx5BRl7YUKwyMcd6/trYMl8UASrVbYyIfZYhVncLtbAs
9izpdrHIStA63e9AFwVfxRJ19gRdN52xWP1Zgjx++sLJ8q1ZI+d77WxuZolr3ppqN+sXsQS+ZJZs
ESBXTdTmKMsXKl1WQmdhPqUIy1mAI2/wyUPvf0QoCodX0udv5opTdBstRUuIbl5rMmcZBWk20hms
44Yj6bcXHnjVU9ikvRXJra3uyanKPPFhjQ7zdyf/VWplxO/aSxaDZ9BCKBhB/3AUqYrED2HWMm4e
8K+NaS3hd6Vq5XDse0qjyOcm0KXFQIs1yBJhl+Vd2o9KrFg9guZ/GqEezhgE/r9mQ4an3NAu0TEx
olDOZ4EGAU2ry/c6+XGCJrjcCTWSSk/yxXiIhO5rBYddCfBqhF5lpfGsX1N0Lm86EWvio5TYPtYa
1EPmZjb+l+CpiLSv2KBSf1K+j66Z/AqCBh1+SzRRFCRCWsC7Mciy5JVlOsg5C7Nt1syUELEA74DF
z4T2/dSFu33FOd5Ypvkmb1CTuGuPsLus04SxdmUgJv9imqgdhSitaSuRZti8/X7+Kl3R0J7KsbiP
EauxBG9GP0gZBqLPDXSNwC78AZouoLB63tj4lF1yIXfqdCfrOVfVi/Gm++esYf6qOuE5vhGJ+ym8
vF1yWh1r5vq+2vnuQ+qSnRB2zEHsyZZh5ePe6+la27QZZKvq18R+IuYpDNXI0+sMIU0zCo83lMrq
hK3bvZYxGZCRJoT4cDoTmKBS3U5YHZ9G7x6YBERt+MyxEoMZwVT3wOBH3b2bqYei7SIoC4GdDkcf
5Ze9AcKgZYobvZlcicZMA7nLrnJ+krGpbaG23rkoHN4vjWF3Gc9tH6cOSbeu41n8m9WDbl5IoNjL
0ZE7XfAfdhZeo4tXyhToSxlhevLro1gYzT9bukLcLRibpcyfkGQfAbgU1XDW1GKYGTWJ3d0LjUHZ
vlkpG2QvfEhCF6OSbE7ToXRP8QPFmWzNw+Tyuk5lzX+vqwBOus3+fvL5iMUEi9POs+bCbTNOKbFf
70ghRrnBAUBSkyP7Uj5e9HIwJ2ZUxCRyUCYybnZ11uJTvp81kheJc1eR7T4OqYC55hXxkOpPcJkV
7oe34tFSoPSfdHFPuyJIgKgnZhzPVU6dRquMGqi8vpPsd/PSWfTcdeQbNzh3F0mh8DU76W2deQoe
73cx6WQjCQnpCv6sfPPfPy7FO1dRIHApgVQylo2NPtF+bqPvh0hiU7JJDPuDQ2fwXAi/ysDmSaFc
J5aWByrd0UBPEEKfHkYMv9sK/G7m7AyfYDEifCZTGna8nR07dAK/4FHw5eEwN2ctu+OMAGAw9kSR
2s5UGZy+ymWYqY93BgrPWIFKp5hpbVqPVmNcT8kwT3DaDS+2XX7C7k14r8gTlLLkv8bW+nALsWkH
VFKx5tSY6vY06H74O/ysv5cUuQaHOh4AerOfc/5VGrI4y/Gt3YkUlWxrgAt08/ggP7aNaV0GPPGZ
pv+0aGQHNF694XIi5glCKpugpHvISEfDMzwHC8IaJCeK1uwtWY1bMiEVd1K773rc6jX9xo1q4R4V
tFYF4FzKGYh99IlHT3JFLo46VgffWacbB1Q7Bh5S8pIyzHATg59NyumUr1fs2nTeLe0Z1kdUapYZ
tTumXJIC5S5Oaz83YTb/RCPG+BHbckjro9FI64YQryOBTeE2huphre3esJEPNdnaqBonUChguG2J
r056DjPcpDfkVaZ2KyJO9dAuxwnTPP3KkBzhgJy5QU1muEGagvkrs+TAdT0zyEkvBrRcSyLdTRqK
QsBK7VJDqjj/Y0RpnBYYP4P4vtzjFYfDpcnj819kW/hv+ZAclf4N957jGGxwK9oerXfPB/dZ2Iwj
3lw16czL2OiN3q8vcNbRFWuXbelt7YMthFQ+LOz3wA8NMySN/LFnGabMdmwS0+kq2iuKut0kqmBK
zrryxoV4oPqzchUxxm3JHP/1lej+1zerEIjtH+MsxzNjdivPAkoQE2jyuM2L5MjVAYuKFNKzyQjG
nF62WmPdHuw9Tme+kwlipWWoW2g43GiZuat0VGe6UxcV0upavC3XdHKO08Jv3UCSqlBaRxBI8n8i
n9y9+iWLrKYCxHS5If6rer0Nkcyy4O1I28lgNgUbr4eMtEcEUYOsdgedf1fc/rQcVHHnphjVWr7o
tJr49DRqlfxkQsHIKMsvsuESzRARoLvUfA6WOda95u5kvEInTaGm6Qo6JgNH4iImgq6UgWe0IkWr
srhJfoWmNfBs5kHckROM9fkRxfOlDiFSiwA9UXLgSfOUuCj3crfQBMqvgNt+qnynKpYptLfAWOam
IRGKATAdB0w/tg26+elcMNbp1vv0wznvixrqWK/f+0tDIhpIQ62kCYZIjqepqbZnzxWEIf0wl/FB
/vRt8Y8E4I7PvFc/RRTGGPCcfD9t/WyB9CVJ5LsM2HFEpQJPcTsEg/Tz8sKwqke1MNxLeVSMDcY0
Lce3W4UoDoKTjzGxikQU80CEmp7oMnCY1BBlLKN4sqSE2Nqk14+/aROH+2ttmRGaJl3wGoBKTRMg
uW0xnY8U1I7NH3NpB+zwt/0M8QYcdLjZaJz/aJcby30AgRzwGRdRFFcb9Z2nlkZsQpfq6f8b/8Q2
YqqMcdVY7Jaygc1H2DgU5EAjOAqhJrmNY06axT/ks1fGcJoy8nxhqUnLYnQbpTw9uawWDStqJ/IH
HSgRtgNXTePFOq2P2CbkOvkX8NUOl0noqXW/W45x3VVVjjLfdRUEzoVfXYC6nXMAaU/8e2D3sgGT
fgewxaqP4Nu4GgH/BSS5SnsdtaJ1nGutJHWeqO0Y8+gbF0z93KgDIRIHWdmQJ1RtGN+iusx1a1/p
yHX+176PphnFgNeYfLmZWkCPHsPxuD1LEpY8HDV6gyXJ7hANbhQS9qMbiR1pzymD7RbAY2zItuv3
ySyE8Cgs2QrQXHOk5HmAOQTKRj0MhHtFATnI8Jf+qb9u3DthMzJVKCabOxPwmkyqswDhJVlYUu+g
m7bZwr69ryn1ejJNQkidca9jnUPttpdmFHbXAVYLzyks95Ilm9xZ8zpYa7iZ7IdtsC0Nhbl2Qaal
vWvC2ta35RcN078kVSahGCgYfpyHFfRPjc+30BleSDpNW4GaZoSth2JrtpcdrTsfX57yI36+hpeF
Li93pDaBbWCI+3Fie0eNWnos8qsfNhtFY78+8zjxcN1f+Tvp6xOjJ192g2fqTE+X0lB0qFsfyUqz
9WXT8sWHv9ay2go55tUKzT3Jy63qRGFQAA5JFM8rRvi2+x91UYbfJJw52AHuFUOYxK/YgVWZwCu9
gsFauJG41UyCAKLTJp9LU7eN718coAV64E4gwPM2vYlFUz8Xfmo1DoYqA+g1fo403hySiSP3epbO
GmlvrRWLtvzpEnKnySXUF+8HRY9XP+5hiErb6nouzcIZk+RZnGlAnAMk8eADVWmwjcyPp4ymz8aI
KwxK55kkrgALmUwl13lwx0Og9Xc7Phbtykgh2Il8yxCcYp4V8z/GNBUQBRmCixCpB92LOrV9ZUEs
HAwbBJehhvRwTzcI2xATjKTwdPdyiHGwBfin+5MSyEp9Bsha5j+4hOaO0rFIb49Jc9dCDw5YQzL+
L+31AF7/+sKbRrsFV3W2sR7130/Tf6OIbpFJe7SzC6ylmr0l8joy0FaK8bDTlK7OnQHWtGql5FfS
/Lc7V96J1ICtSK1PyhU9vKhlB3fOvbzI6J8LPZk+rxzdIy6MKDR+s73kXQkzC7IxI+cxFVSjLHTP
2cMvLTSBsIrjPpWINhO/VbACbHofLK5QToi9eIJL6iVkvJE0bV3zQQMRqNGR8GZ0RfekPgTiRhrz
hYuO6Bs52+jntfTuwzsU3xg8D8DgEubag9CeRCH/PagJHQQgNGZ9xTn7u4Am5chiR2dWZaTG6C10
X+q/6SMJbAIhIYhIJMqiEdlaH4hgGp41E+ghYgY6PEJ19XO8UDoc/sJZ61DdCOsrZsfpXgjTYOGG
yRpVfEVguZhthUKB2SpgOtl2vjIBBXOezSB0NPgSpDdigoszpfJ4XwnxJy7W9RKVm5bWecKaiDRw
Rj/meqg9MGlmv2Wso68uPqHildeDwcAC9h0x78tELgjQZudpaTDCzW4Zlp/hC1djyZua7lDwRNh5
TXQt9wfQ5hvAHy+1IiH2YAOgKIReriPmzvbYWSbhUPFrkjP0dE0p5O80SHrD0q8163T8Wkr9vRIM
kZG/kmUlyDKVE51ueWAt2DwAcYJ0LUyj7NDQM9xBh6MIxNN8ne1AbXq9A/o8zDBTCiMKSVop85WO
DMJq4ETj8c7q1p3FXDbJ3yKsKejqIbAuGUPDV61wKPT2SFZ+hfir5bRspt0SKCsbvmG/paRQ+0dl
+KRX6oz7iVF9kEbUTVPty/8BDXzrWThATVZ/D1iXGDChRwii5Vj9cGthu4QuGfNnK6b6mU2n8mzI
Wpofw6u0Cd05BiebCvs2hUj3V8hVn9y7RVi06/S3POxZsrHxWBt5aJhx45u+GBRZQhGt2l/fA4UQ
5u+Ttk0+1c9yIDRpccjrHJ0eHn91xY45ySE4hsgtq3+dqioOpwpNUOUvkq8bb8/ajy75FMXTgDMV
HsWEnDXuQlA4D65tfrgka+Um+Vgjmwms9xIUw4FUUjXmkAUGJEW/E9FYKnbUHC703DNbHvltbHkm
Pbn91B/kx54VZ57M27szrK04duGUTwMMSyXvjZUs4+SuW0+2WndC2BEgHvOEt8QFTCpHR/GCLYW9
ZbFpRoPs5RwuZyo+ASERG8UvKOlPE3RTXD2rVGirA6gVHaI22PWZ4hrCEMwg3gd4XSjSOPVRQGCh
lPFOzN4jTZxLVUUUa53ZWGQoXnhAgTJarcE398lR8cCep1CLn/eu3a8sNjqb9dF3zibLf8NGCGtk
rZR199dSjJYDLnemb0hpnLWBUm8ZHRaWL8eXkQZ38Wi0OxM2XtP4Jf6TcaiLNAvbYlBbGHQxRrWQ
p9tDudMYT1xuZoU3t0iph/Wa8nlJ138LoYlP9tXoxTdbSEEHzkLUsLcz5aM9hPZWUzguV0YCCSbD
n+JRyzcCxvPct6UmtfaYvCRd90qsnatVP2rz/IYQUn+pKfc5xlYvZA99sBe2GwSDNpK28DQlrcMM
ASTbMZ4Hq/JQjCGrAolEtQYvsKMJ8BXULGuBUZQtJizNSMzbNMaTXi2k34Mt3fJAHByWfOZB8S2C
3Jysbl/KYe6diKlWtIFZ6XK4EeX1Ljt08nZiiB0lz4dbx7lsXOc16fooexGvbAAOUr8qrM2v+/I8
ErLUqKkeK4BRj4hdNTajQ6ekIBK9M9W1kCLNc1shzPo3nw5rvcd5A8EqP3uuVdzTQca9+LNYJjgY
5sAWBd3K6A8JdpLmbJBe3YER3m9yP2RG3wAP5tcOhNwehysaiyINOq7lhsMB1oXFW2wBAWSsgEFf
S8+KvUwo9kKYcResyOz25a7JDg40DeQnVOHo7v6IGi1LjcI/snxKgpv0R6u4q8PBs36hNISWGRRe
uCGbpXfHQi0cOzMxMSJA4BcN4OWWsWeGVCz8BsBOXekQk6vFmrbFsW8yvAZSllEPQuErAOorSvIj
M7Q8qTuxhh03kMZJ3mlZJhe/TFbQershVBejicMNLcIdyxsw0VdyfZS5Gfic4ckgnfSJekV/hm2U
ZxzmCVoE0kCecZICNmnQ1421OF5o7G6PXcZs4vVpiesLLk0dJIeAP4Ra/K+rE4K9ASwae8e1ki2Y
d3m0cfeNr55Ho24HHX8VsTYG9kNBbuBCLE4ye56esnNt8GojFv2I5XoJdprnWMaVtC9IoajsP2dh
/0WtxX9VUSmGkbz0eLbKY/uSIo9kZq7Zjgvr3g7fDMV9wF44JrrPLF7+Ak4qtB040Z1H3LCvwg+T
8V92hOw2byLLh9anLHDlbTbEvferM5w04V5fdLC5izYjXI4vaMqAInskOAEWoUhG33nLfBiiSpXZ
e5KNZ1iZ99gP92scH8TlFUC+KW4S83ffi17KYbzgmDv3BajVvbO5L3JXqrjJWQU8cLA9mbXYGY7V
pAw85AYIbHxQQnSfILNeGhvnhJZw6E+6PGTQs54J+Yuq5yNf+B+6v9Psj7n62kb6Sc0e3XYFyCL5
EOVb85LAcgxxH4/khpf9Obyl2PainraZa4KGzYXiDQNzDNEq9M8rOMQtVquxPpNkrpsB/GSa1FmM
uGamHiUEQGFgSkAvFjVZzbLFNP+rwLsdIVn1rNeAqdlXnrcdlv2xYONHcu2RBEGJ852M4DCD/SZO
frxN+fsrQp2IHJOvB4sWRybn1g03h2WBzc4RUYpRLiiA09W354PM7k8FHd6zxJTU3OVb6M5n/kk4
psu+kl9mu1dyQjfYCfXj0WRKAcH+2LcMiFrSef0Gr8tyqBshasmGqrmKQfHPTdWkYdZD9BNSTsES
5HunGQzbLZr4k++veZw7bIPkoYaLRtN4VziiJVekN+QeeFAGXTp6f6T2tZMbi485rcOlaow/CWNk
SPGv7/iMtWJV7SaIUV1uNYIUBnXyEVzsrgq6dAqraW7zL3RNbK9K9TpM4FeyAp2MRb5lG2NFRVOA
6d6g4nuLAz57J9aqhKitY12mSREJ8awmOREYMQFtRuPwWUzaMJgD22fhQgphSFFLV31fl/H/JAGh
6tanwYKzDJFGMSPaqjFnh18DC1E/Y2l0UHY0IbzH2Vi6siy2ndwtdI7X9AV3VRpMagnLkDUfKeqO
afdYlqEPKAUdUaW/6HK1VIwqnlvx5hNXpGBeAzv5q83aGkxcYn4gSLmwz8CxIk+ywibWUs7mMwI9
Zqc1ZbdgOnQhpWhtpKc7zDVn5cDoLc9bSMS8oNux2kwn/IwI1GqRv/dOEFDuhNTfcW0LJq9YBzYC
0SqkZ/ylRQCDMtvVO4l1loq9VRxcl1sc9BZe0kJFevmuiiB5zC94IKFcmO4/Oo2reyEiMFALriuU
xyfSBhuu9JBK3IE5NjKnkTIiORglmJfRM5eY1ztJiBGaEmtk9HM5zVW3yZWsyku5j1TicsxwzdKe
3uwW6EhMwh4hi01AvMFIoxaHDcrn03q8zdIceJCN93LDX4hvnJjKFKiDK3I87xxvU7IUfIDAddTk
5yoFaBl/F0zf82zstl6+E0iGWRhgipFpVyAfYK3YF1l1hEDWa+xONtgSFd5qJewAkEQC1YeuO6gS
DSQGAETisZWjHDTKfV7PP3RTuW0HoB6xeTmna0VsTtKzUJqFUIomwsxsUS63xgBuLKQ39+8WkoXK
lA9ClKrjPqbBkZ9NyBT+cyf6+/JiLT4Xfvb5HQQuel+5pHj0PkvxEFdhyldQtUigfR7Ve8cUBN5b
wISlO+4v1/zNEsFrbKH8wOZH2ObRyRRs4f0qKGK+AhOag4FY46ecv86ZZ+iIBYViuwCaDRLZ1fZt
1gkz6FfaVJe6Na0gZ0LYSZPsux+twLHGGJy3FREI3cPByOuoGwE9tsGCq2+lyhDNvG5j5lp9/U/D
86TofP7ZI5ood6tLQwM41w0SRiIsslLnQbWq4TckcdiZPBaTAE/JnsGXsbuz/bDlm1YzqVXKvv5w
C+6UmfFzE94EnMRDN1VprbdaZTKXUZuevibU3q8qw/RDrcKkXGwXkFiT65al2ln9frWQG4KrnJK3
iIV6QHwzwlwYUsEwvwO42by5aJTdx0NaXP8G5Ob8xrGQNb30JdHdTAgGrQWVYwb0/CX9k4jiEDZb
MYb0bhVFdurUY9PfBAX7ufqJXPfd9XP2zY5S1Q+/8xXHaM9sp2cJBCQ5IXPUqsgEogIIgyuPb+0S
THE70iz9N9lZQDvE2CikU7EONyzZCQqiZt2BiUXJeNzf/9z8I0Z2c9R7p+DZUsvtPLBQ/pgq7K6X
7DekJhm/hG7B2ERR1E+jHJ184MPSYy/4e7Ba5fBb+b3Al3Hc6qkSh8pbGH0Leeo4ZstRGe1s56h/
ZC85uIbf09kaPZlai/ZIxx1lNA/RuTJh9+v6SDCnJnzxnU7DuRy+oN3RUa2aw1yy/+DKIsE/Zn1l
vF4nLFtt/1ObLfdzlhy025Bq5A+Nltj5ACJEDVC1/YNVgrIuu/dhZAO0v7wDegJQFP04Ltrz7TsG
6ErF3uNkM0cQ6OjN2Jj8mgGKc7LkpIMf5XJwXHfdLijwQeUvszHgUcw9Zue6P+UOdrTk36+YHQ6X
p+BeR1OEYf1kNW4ItDcRTtugubYk/JHqI8ZUZgY3Mz9GNZg/5YD4nlsxlvFXCBR/F92LyHArQW7g
vtf9lLK2l6CEcSlfIDyoeUQmWuCzQeDzl1SyRgnJFcUl3LHRIizKd1oEMMOOfdO0ggkEhtf7klET
nmPQEqAqwi0RfLZaiN0UwcVh8N32+GKzPTdX4MPJ8OGa5EZVxAJEyyK+3oLexbTCTZbD32mOmB2B
agRt5dbcGynxCyJe2s5MPhzzVTDpEYsxRcVy7eIwD9ZGpXz+dUUyIT7k+BBGqIyaUN6nQMgYn9Tu
2cxiVdx2slf9dEHGouDTMyQ6YngwFFMr2RqrKM/MnHcYg+BX9m/Z5FqqjahcwNcVYTJpoZzjz5gz
etYL6WqCLtIXPw+x4YRgaAKkwE19jTf+TsbWM9dleqRU2WVBCJx6hTtyNHTy67cXPAgptubF2CBI
8NvercLnPbPBbTTE0Ek4VMqeAJtsH+LeOemlxyNY3Q8bkNsRktOrJkcb/1Oo9swDuU9M3IvPd0tS
vpa4ek24PU2yYRRU1dGSYmYm3Dy9SkuZsLnSSTP6ElA/Hq6J+DHmtQeVVBaqA7ozl8H587xZzBkh
s/BrfGhSLGjlZZf525YfzqHP1eQ/TAG+Ys86eP4xv4JIipY+crlqzQZPoNn4CiCmcMKz4jAs9vN/
Q5vFI0k8LzDbTjQlTTIYq6VoEineL2yz+mJ+Fz+RkbnYbdW6IJ7XHiEiQPk73w1PlDwp0aTVxmMl
3YSVtlCLqw0Ri1Getgt+a/94NItgAwl35HbHDSWt8ZAVZkLnxp+f4CKREGBZzGUAN4TQ53iB+joJ
p22PAtcYihXowDeC+q7QTw5xPnaz4bGl0U3/gaLSC75cQtyaf6ulBScdzoUKCamCokegj+L5T67z
l3hfGYFF7o94//gdPQRkXNj36tyoX51RK4FltGt1A1encOSxplVZE4uefJVJc/KnrkAnmcq1565f
Nu9nGp3LVlDxgIkff6BCEfo0gcCJWyxGOUijCEndyXIhiF/a26DNHzlZob5EjoKOhGBC/FOSyAjn
W0fYQMQjYymhKfqKvAp3oQDusXnQodnymsXsRRKQTjVv2+CE3Z2Rv6aRZGdQoRHu2EvpdOSY5+ls
p8PdRArCkImiY1WG4NgYjNmyM8hxijx0aKtJZ/Af0+ygsCHcuaI8HpyTLwect2vQEWeZJ0ef5giJ
7bSXS9LSoCzJ4fNFCqrvMQUIRzKPrXQMPcMCfe9k0JFm9lmQoJvwIOJa7IN5UwCvlby+D3anDq7T
ycrk1UOa4gkCcdzdXd7zC1Vy63ymgBygyVPiOAZTU74xDu0PJaFBvmicy+pXRw8o4tedo9HYwdhj
G8MtLOHj28rSLW0GsaX2hGHax35jjmQijnpyTweSeaLePLfL6rcF2nuNzPA1o4Loq3lsx9xXUn1b
90D1mwZ1kXGrdXTvxfAP328mDLKxN4A9n9qbvGyFHpILbhBeBDabHPjyDLnmBpmo8DWbolLPzYrM
vQOZt44S6D4JtRRLx6JwtDHocOtZ6QGIVSFHeZBwg8RO55cENw9C62NLh9HUHKAhAMu+dQBvo7Li
2HUaosLzwx27bLdXFr7YwJwyVI45FtYJuKM9kHqdtNtvHMH87dKrjNTHB12GlIqlWxYIbS2BoNWs
kq6GqmBKVLAWm5MFl4QL3iR2yMMLovUlYKM39iWRm9hCKN4SDGIh06VM2MqpAq/Uaf9JE0gyOS/m
uvtFFfuGnlWzciw8Vb58R452CY+cr5/yQGEaflMY1irs43S81fQD6nvqarW/fXrsEwCfaN60IUe+
vdRDGlMdiambWjLD8US3ZlINwrD3g0v64arqSXu90AWfVZlLFbz2HC6Q6GOY8jMmc5PzM4UOXIzz
HJiZoLv+KcREIhZyRbTkWzCiKh+8YdmmXNEljzB6yjkgW3F3dLPljIwK9D4WNqg/O4dKSGhmCTy5
sTsAEPJ4KWPLBHDa2yq+pCK4U82rI+NrHkJCcwOJyPg0PoryelBAF/JbY73+0jv6vAOjUbkpugFB
awjP63qx7/84mqGdFIC9Tb41LnwQjMI0CGMcARgpWBIk6WdwE4JHhLL8in/EkTIoaOmhnzCYmVVk
YSTk91ERjseffqcl/vDUP7LmONHc9vwioFWDiUZfDPAktu+Tso6Ytv7qQObrkyga3LXqW/K1O3R8
wlXsJ4qbvlMP52I+MaVNpZPr1Z3s/BrRvKhHhbKAtAvLoWOKpSNHD3K553tkUOYlS+w/1BFN55s4
qOLqbpoAgcRVfkytfnyMtLALsn7BVZLMC3RrLrnvB3PUcY+7qIyO427NjfCvUOLpgN6pxkYSbmSt
wza8wNfmy2srNJERlwxHa0F+k+vQPCwcd3oH/3y9rSqFdrrcyGHjwKolPyH/eVOR9rA3ASXtMXn1
DhE+5r8UkvUbV+SbiAv+VA2c6yo8dZqHlWbQCC7fhlur+7pcLGyQrtt3NeBI+fvqrPCKjp8nY7fm
ntEGOpoGfHwJNeTONiBZT7ayxIfwseCjTKTDdm9fkODMkcYYW8AgnsOEi6IDEeRk9tjdVIqMOgO7
K7tIhlIQzmpNmTvTAmGuzkrD0e0XdMflqxorH4wCk5B70N9soEwqc8pgu3cWysvKP6L73MUNR6M5
GP4YNAqa7EgoNGcR/Tk3RA3DRvGHoLSJ2Uq86a9LOudT+3go9k3ejYpZDc5ogeDHu8Iy6VSfIr+i
g+M1InVMJjrL+tYoJYcH6sietdoWdXKoveYF7DcbOo5LWeOmbrbdnUVYEA6UWnaiIulnTBuHwdWz
rmQYD9uhz9nGHpE+uG5m9FmCl6AZ4ZIKzVbI6qINhNwFmyI5xb62+6/jv4IpKPf6JCZWHKM03Vqb
+tfUhMHI1BaYl/fwkC3TlxMCnoAcgY9vwpLooTgyAPsuOwlm/lDrJ/i5Nt5ZvQbWeu9q34cQfFY/
+VBE/XTW+7OaqdmVH1jLmxu3NAHopdPkGwdvkloaTTM7a1E3PqK3c8RJG3hRpzflfPTeNZiV4oMA
DpgBpMZV+RnM8GsZPpST33M4S/vD+yS6IGcwYgx17X2GJo0qq+oqmpwfh38ZYdXWXk+Qqmpd6WK1
2Y/jtG8WwCDs5fZ0NHOmc+okz6GITGSGWyXl24gB+ptnuTdvJe1PwxTK0ZA3gYkeediOhkqc7ZtP
sWDwi7cVIkhcv5mr4CviL8LQLUoh17DXYw5telBQDJgtlBq9u7yZrf2TwZDZRdA8S1/JPnGBSL6r
TLaSC4weL3gjaTze+evLgvToUUvgGZBYoqHFSZaZiw4HiyWOxToLFmqQy4V+Nsc5y0zeW2/zWzfO
PHm0Ky4pjVGlJEVBfwxCwNp22HgkfdueFftxSR7wgQU46NN9omaDnkYs/OyYBQlyfLqyL9eMAYBm
jE5E7lpvoGWy7Dmz/8/3YMD6zeppi6tydPkzsnWFJk0+1A5YR7SJjlkoDOFdweD0hzOEW8tOgsFf
rW7G6hq5HomM0ocdYSHYClq2rCoWm94W+inIRylYbQhEUGmlZr5tFy0juYTPfD3FLlkGBqrydsoj
1jWUtPW5iZ2NeneorX/4o31D+GjorNB8cQFGBxmDVPbsxLS8n0FnDHGgxI1kgk0f/chEkpAdxrsM
miz/bw78TkqdeZu/eZ6UOUFXfkDIadvoRA5fXzuPivs+/aRH1dDD5faB/ItFU0k3AzHUTMZ9RbWH
8jhlus4qcpgrf3bOwD8JuK2dqWP4SU3SH5GaolBqkyn4FNap/9JPcVWwY68gNxUhUYYeVqPK30u+
GiLsqps0KgTFJNUih7V6+lMLIE10p9dHpgkVzW4roQywhDlNx9tQd8DANikC5mhQnpc0a6OM/BuI
TUlJB154F5GGKYBB965H10HZKhUxEbzu221Z3cvcsVixgmRsoxLKxhl4aF44hhb+bezpbvXIcnwB
jqkxboY4feXUGZuPvkNruotzYk85crjlflVk3F5OekzunH5woucpdqAyX0nGu1TK0xecjRJwCvnU
roxfhxfkF+euvB9mfg6fVWc46oM40fuPbdkKSjiRsfKgcnsx6RHQVcFs6xDZiK3OMXSf0zpEvzr/
iztGg54CwZ9oP/0ZQZDXaPCC3PsnTof1VUjUzl7q6k1fBPP2/gi8u/TrIq+XWxnUfme0cMrNOpDn
oKBX6IddLCE5ONkcJ9XKL4Uq2cg3xteVZeeNhQXu42OA1mGTtx4ddJ94EpfITvvGba/rqutpSqqd
UxkH6Q9qXQBQOs4Rg0RRJ2Xm1/qE+3H9dYpQu3mUZTAxBgY/Oa+wwRzQR00emBVFYCeGj+Lw2I3q
Uw+eYHcPmtIzHaCJoETgcV517wR+QzYG1v5l/FuKbYU55A2ZpHelTd65iYDNsW10IrZ7U3dWzM42
F57D8evVkpn1SuHFl1en63K41OUhVP/OvgPVio761dzedPlSoN2x8gp6299etxQ063JgVFXCKkiq
QBzZWehFD9aSxgmmrhjQonP0LXTEdYdhsl0KfvmYBElhIL0Fp21Llm0ehf1zxgrGvB+UsnCnlKcd
m52CoHVRu2LTGddM7Mk4it/KVzslI3lGOKz1XcTrDp+7X4PPtCEvbhAvPvd4nI33emXASlj2AJnx
KDB4IVfj80WLCbcVOpcgQ9+88L/EjVTfltpNHaW+JJVn4vukpmBtgoTSyQBZ7vrvVCB1StotCCTM
2Vmj3Z2uuS6wPySiO9LxzX8e1trhr/oc2Vk/k8KYcEYzIFN8xsZSf34nt6xTof725EUeYoQaX0Q/
O1Am5JMCtg3eKnHL1a6CWaRUDEp0SCiHFSjIReqlKGpsyhhbwNgqcKs4cu5eeQqGZr5SR4ADJUn7
hyczQUjPZ33rHI+dXYNLaDQ2zB1ygucOWAm/WpjlToP/kmMptKnd2BUeK9mBp40pPF/dDcHW9RDG
AvddAPnpARqgnnNuqXctIt6ZDKGw6koeMUn5cYBBqAFWXYfVrmnCEmRrw060c8XPgI8jmIDEo/Hs
Z6BnHcsjAlz/ghU6XEz7YgDxlD1OS81h3y0H9zJAqPNN2XNCzbEMcsb1H0wIlKI9XM9iumdlZqEf
tAvVIdXDBkDMPDh74SQ9p6qc3IJ/O4eML9ddTguDzwMG0T33QeH5bF+Ikf9H6wMiguzSgmEPFuZW
Ua8hRQ5qoYtm7kotcgBdpLx4by8V6anep3SUWLzHNihz6LkGeHUzY8BIrSlpn58RsVUt3ahRghr9
d8e4JjahDa4IEO3LiCGCHH0nE+q0jymKOHfW9/NDm0/7BXaNmT9caN6U46fKOjgMhJMwh16uSVoH
ltUjhLJ6jcfCOkTwhbkFN4YFDk263T/m8v0NzFd7KBHeTtynXsgUhwB1ebkKzB+nk//ARdDtfNYn
a/ZAz6ZisM/BKsKCQkEAQO3QRda4GBp2014+G4+uDcmPjxtauOYwFwngufd5LBPlkf+Qp2ma9g8K
GPEcz5FFWX/Kg0n3AWB46MCiKp0gL9Wgmqk3SxZNVnawQRE0LiFNEH/xoh6tq28s3HdpxPtzFoCE
yKJGI6PsC2s06RLTmC2G+u3Psk2m+RLUfNbxNtbGD/pBzpykDpBzJtZtOFDUmtRucO44NPZG16wR
YCgHv+I7ekZVz6Z5tkUS9zVkHfGRvxLxjYPM5nhY6yyK1NEIUttxew8yVGslbKvHTLFU9t/Yix6K
g/BFI4mJzoNs59ZmWql7z09iZJJ9OYfltCh6M3vHGDVgwQ5qCS73l0fWIKrCbU5QuJs1NWXlZRfL
p3Kn+pFXf4jXLke9xOCFaLhxC/I4770zR7Ho/9S2zXVEaqmhaCvJO12VSQIgq7Rnt+LnTsc3Lc1t
qxWatXi3LAqKgmknPnyhJbaNu/x08ZEM90VZGEYJ9w6QDz0mGDhxlb9K7BFfwHC7MP/JZlvubU5F
NldIm/leF/ZZAdXAQN9/KP67fX0lG21PXooqYlyJlzs1WJfkR1LhOdmT7RAq1e8xgkjzzvaSWpZH
w1VTBMlPiC2IIuCB2y6DlcG5q456JqPy0z4+PCzdD9cTWKj4Jx18rmJybJIQKRHs9JOUJgkpH5nb
7WxOyomkYnLxXADBDtID6gOW8bl+vt5HJI8vPbxHVJdZnVjh98MjubVNKRwC/z2Yp/4tG/q9SpfR
/Z4BUMTfgT0XZ/KOQ9x2y0HWAJS0AhfigeSPrqhjPsWWh+l81EXIN8w4k6HWGjoHbttDfQQkMb4p
1N88Ys0y5uskc/+duO/oRXDjgTuLjCwsSv7WqH6eOuJgEGHu/akQm932hmRjZj2BxkmW3qieuJ6C
UQUxma18F/hCA36ndX8o4KDiR9bdIqua334V8r4ikTqoD3LHjEm0XQ3up9b1vUBAue3DZfCQ5Jtn
D25duuiNw++TCsPfeeTYyLgQhXYrKwakLqcNU8GoF/SFNxFhTPJQLqB2BBUBaUJ4Ns+6t19iNtP0
rc8zorCUX2ziDNTlSs2JsXit21hi3vdI+0h5hty+YDZ7uSvlwJ3nM9iP7kkzT0GPm2D8DDrLuEWL
AgrBT6B3Tns4lajipIplZA61rBibt1t/TaOrCoo4JP1HbqAYe6kRqxK7ExowBDeWiI+Mwq48Z3B8
FpTgXkU9bqLPGRiRN1+i5nBmZGANymunR7OJDO8srK4aUxEw+vEG1WTZiOvdYyvIZ7Qn1eOBXLlQ
7O/+vA3bEf/zdSxXRbyR46HabDKgnjoRwGbruPjE9laE+ASE8IXIQxId2bsie6GiiX2gfnYDMW6S
aytJ5J8vndfbjRh7pEJ9w45PW0yOJVvQRbqyE7gz51nRoFiSQB0qIqxsKpMVs/s82MAMLaVJxcSR
ZrRpzRbTpxnuX+G+zk/AwrPpsKzTUopo0uCMpOnp77WKhsRmb7ldwCQP2jKAR62CafxOvATYdhbm
avjbs905JlJXnC3SELub
`pragma protect end_protected
