`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2024.1"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2023_11", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
CBun6fnRJNsVEowQ6itVc84tr3l3505iFxg7fFUwZ1APlKwqrTKOO5KKNSzxI4YGnoSBaZTt7Qju
ReW2sw0IYzgVLyeUNg22M1NcRFuxwTqSCUJZaYz8+yj/aLCr2SGmip8l2/2X7hV+r8L4twVlEYTM
6+HPevqfNvQ4neFhUnMlA4f+O7Kgsb0W2u+wt2Slxyst6PIFwuH+6ylyNgR2JvCBnMzEEZDC5Rfp
R9rMntE/OpLS4+UVrpVXvpW/Zf2sPs3pIZlVMywg9J/s5jN1TSbsiO76AAeN9So299iLSgyzNPBi
xunvGakq/yHTQQ1/YvaXKZzICmOoikT0GjAthA==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
Ei0EmtAWiUXM4JY4yNpqYxUSE5uGzfhHEl36nk60HNFyujrYk2YBFHsXEbiuXl5Omq1n31FIlp+z
UUA+rLU5+3M9rlDl/qKee7oafKiqNZEYfWMpH+viClLQ3ZNJu1+i7dy7IfKPmkWKHChIJzVW9QSm
8TZ7BjQBs4WPoLQ6qbY=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
KZb/VXjkXyXy3RBoyl/m2R9p4x+fXywjiOc/deZ+vqBB1msKIU55xk5iP1vrzbm7mgl3/xiD+5Kf
33u4rHUOSfg7GOwKddPtaKadSW0YQFh52LB2iz6KWHdlP30VXWMBSKeMP58veyGGA2PgMs+nlbVg
VvIOTgR5AkoFt5+R8VQ=

`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
nV7GCKMYXT8xz5moc4rfmq19oyNEfidhR4sR9SehP2X2DdDwOPhQWqme4mT6pc6waKO+Sv7RpxWx
4Is2092CDw==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3136)
`pragma protect data_block
JV+7KRULSFDVw4qi0oV3onCkUu9dAe+pi/AYNL/+O52LtLtKksuPmWPQhYJ3gVF/njq7+sfUnx1x
5VST2TRT11+qmt54aDam/aaSuw3unhXZVokA8mQcrWBiCkFLh45ae+7BDnaihDTlBBIJO8lC+VsS
fRRwjeLVgrjCAeR6SlueaEE6mOCMK9RYnrPeSAMRj6M3a1ou6d3t1vuNm7gz8BNXqmNC9MqhJqTk
BDdc2jSX5OnqxXjl9mB5mGRVFRi4+awGQyaeGtkeKCA7QmRGg7P1rYuxcWaymD3uMs1eaaQeQq+u
TTwxbaNwd3l6aDtPf0pqzhQxAR+rL/FpfZgAOP5+Vh8lM1X2p+4NbxVBIgn0v5nKdjj3+8LYjVuR
4GSdY+IJVcjfslVdSD5PpHlD9hGeMXOGx9ZykC4NDYPFcDheVJJvNzzCnXgTmWNhy5L0TJ8QYn0J
roq/xJbHGSO/o0D0gbeRSuymyZ97bI7sALsmszEcc9RDEZt3OgalQUSuL1RleFNnD8PcpVgFU/Vs
ALD403Lxy/FCQ7/EOjLIFamj0tyWheGDzJvG+BxlSd0rqh+ozuOO8wiHEQuGyELxXNm+R6Ova45p
9ZR8Ee+1pl4AOJhDfkrkG2Q9wBUC9DIpY0LJPKAL3ydeb38ZtQgXGLV+h8qql15esX3T3hJ4g2ZX
PrzO1jHjM/kBXV+uXck+em/1M5y4MF3vqsE965+E1leVJx26qkNPUw8MQ1TyK9/MlxcC2NtZsI5j
hvj4KbSGeoMGAidJH+ArhYHBqaurWf8Ku6QqxPHqnGlx8UpThSuhnlkb1v1KUp8iYBOtX7AGMuQn
RxiyGyPZbHcfgblDEzZow2OLg59kkR9zd8hZOTmtPkS0tXM+d0Ef9/WhDzVmEEinoOLY6WtF1ALt
m2GcHfDUafWsCay8/r2LaPYWnBFhZ6XwXhLi5rnXtdgqaTPGakjgdMiI+IXgTAleQI2Wqwpu316X
wPyImJ72bwg59DMVOd754i8D7lVoqkPg/QZau9JoOvyZ4Q3weuNgz+VTQTDj6PEWgrCJ8sI8sHvl
vEDpPVAX4zrdVX+gYoCk9V7tnjuaU9HNyCXdHCdeKo9pJNY3mgXXycC9+wfRRXvQ5PRvT9jqZt5g
fAby2ssi1fTvhUysA2xO8uhLyHMjyGY7fzCJGjvPEPDyscnzW3uqdLdaeRxlIfwTXP/inNDdwdDK
dImLPVthBSTqIO7C/yKJJpB5OWPbuM1BiFH5uaPb+tG2h9dRY8LxS1ujebFLrh6zuCK0I/phF/Ey
auje1cwtzWzdns/gqUzpYZFEy7Trlwcu+ubqYa/HV/kFrS5yFN8zhLENyD762OARAGNifX9vgW37
UCs8r2bmjA4Kg7/vsaTBnvsuqqR/RWigWknG1t5CuGMG0J4KhXnD33MtvZcOeAypm1vPzIBiieJb
dPNxobkgrTkRx2eFVfh1ENUdVBcBJwTLucZItl34p5Sx2hpgwwevroVf0vwFST8u5ty5g6ZLJ3Do
UFsOkWxv1N+v9eQ6/uXnjWbQwj7eljTInb1kxuRVhtjSIvtAmpkjBq/pMsDhwaJV3o2xOyEhArJv
mnX/Z+NXuangoTU3lPatwkG+ydRdx9qwl5gv+i9K8nk4qy4/vRhQRhe6j8Ifr9a+BRfmOOWE2gOv
4zqfW/kIq1VaY/qQtf3PfyhZbR3A5mBTQMrpkIzQ0ZZbbNd0dm7irkv5wOdZYUAuYMKM66jV9EGW
VT+ZFbIFyo73JUKmE/RBXOCHCS/oW6GGd1pxnTgIkSGSPHCd/56ZApmys8ClmVsYG8rp5QDeBWu3
vONr+CC2Ay6i8S9eHo/llyDi266qDtXJv3P171quT/KmTFR6eAu65n0mcoPJK9XEmn8olhB0sIH2
BJaswEIQhAfKFrXCvQ+NUSKTviPWGAqHgrCyOZ04mGFpPD4Z3SqpPTU8kPhqkqVJRXowSMhUMkMZ
ASywSTKoEKsRrZnKvmQTrFkvC/Q8UYm7q/Dw9sjSuij7rRxYmVhuqWDtsKqIIULkzd6ssCxbVLir
bcxFIYHuGqAD8nzYRLxRcYjP2NZTJOMjl1UmVN2B7eOr+ZZKzeIZfTHPyeM5j8l7p6FZVH04YCjx
c3Poka1V3dmsdU+qu42V9Cs9Bvmyh4NIopUB7gUxsf9QpyZc5NhN0JOzDwejz76/o0dTQ0Cx8unf
wBdvrAWT0otFLSL2l6snECfnoeIY2972zPREDTa/LzyEgu4O97y0ukV7T9+Z5WPu4TB9nziIWueb
OOmpCft5Vwi8yEJqQo/6CIG8agbuzLzXXlhRoEKnrgY6jjzwIm1bpBYQTI2tiU6PhUXxF+cmM9Ee
pOG+QEe+wI4PIB74qAToLZ/C4bAAW+HCXceucTUrwGg5R7dHVrMSS4P/hdXbtqQF6OTxfOYzspE0
ZN2rlNZornSEKhoDAXCl54wMzeWFvckRM0bpEhepOPkzjmjAA2ytLPimqecUoKw/JWH2/cOlKspI
EyUr8HPWpFqChv4LLSHEfEIY8cK9SnoIUHMtUb8cxt3wYWaa/8llsQRp66b+W0vuRLtkFtzh7Xld
v51+r1RmK1tBSmGDzmTIJT9A5IdNzlKtDoZJTDqX1ez+l9Lui0HCydJkhF0LwXRS/4O4Lf6mNc6R
cPjYiN2bTD5JI0snRQvSV1aAbY8ptP5Dj5bggo9TiivN5/JLQ8/d8Fx30uIQGhtf0j7XsSuFYSG2
3JV2nncRJB2co5Ti7jeHRt7k5KUMvcBgMAUyJ23dIHQYvEWFrc38aRLnHtSSKyUHgcbsHQDekQPa
y9e9YzqwYTIoTREmJfFz/uy91caJuly87AOnJHrL7oDAS/m5799edYOT1njcCn4VSEYeIUQnvMev
C+v1pfNKt1rtJp0U7aJHE7avpP3MmJymTbOtaE1sKU83lLzfJLxNSRA+CK9ALOMEOGcIGzuWn67w
+aZB1jwKQYGQwlICA2I6nKdDBzf3zis1/ZhNPs3s32gKhRh+G+7sWz1kbEdV7Gmeu3EcnetgrsSh
fTCXA63wywhmx+kUlNmqRmyC14iXhr1nGsXdHybZx9+L+ADr5QFOTJEv2ohNPR4sBzxDYZVhpraC
Sf24wbSPKxtZB5FmBPokVUcyOhZViv7YX/EDvUIrNi3DH/XHnkWHfKu4bxTWtnAPbNzMzZGX1rjb
whYkSbQKpfZxMzPOViX4jQ3iNNuvPBIgMG0kP5YtnX5zsGzCwjCCjDtyLrAo07C6ANSdlyBL2w8k
JXzE7V3w8fO/owMzz7vjjMM/gCqSDVsAD2oBDZUbUcbsko84kH8qoaT7ZoNohii/aiZajxvDEX0g
SsXEJ7+fi8hWNdGhuxCpITROwcWaUZ6uefkzWTGp0VMNHjaR0GPQyeqdkfN8t0AJ+lLfod+ZejeJ
OC45LBS8Z6Lggo5v10gfMJvPefd2UOpytj7zm7ujyeO4t5vXC/DcREAxFvBpiaySnfY00ZuIY3PH
PWqkwpfV1RSpV+3VEY1MxxteDmtZ1/zq10yVGcjW1t3aa3k6t9CH7qOBi5P9VlK+dTRatM7gE8I8
xnKfgo2A3KEkWflvm2+Lo5ZHeNfrByr0d+MM80p7YOZ8TU5EY5P6lf1aUChDnkdps3hE7ufZ8UEY
VzVGecHrBOolODenr91Xxo3L1xeYuFn/WJEG5DIYHPqz9eQ15/jbkkRbmfPU/cBpGz8GdmnqlsyR
MMT/v8Z8RqNt2mkKmhT9QSsOTuVEwWQlXG9rR2+ffjUMU7sCBpuBDoTA8YdnLjULXiJ0Qxy6Ur6g
geDdH2hPbp39Ms+LZVfxhVUPJUqRUQh3ytVRYI1CbwhdsY6S+LDHJe8OdLH4DtGrwveYxqRZtlet
jadxJOJ2EByvOmA5mYENx0FYlsAfZjyZEZz9pL5gJWkQuxBU0EXUJG8z+7KHUE/uC+6GmbqQbD/g
m6zysuQPYsUfbyZ4Zxm3O2+NinD8SuquAd3rqTYhpwyxrY2nQgAHdEMiwXvHbiR/2hqQHGUUray/
qa0g4RtoUh+Jiip1XC9ylI2xop7lQHbcAbS8UygHlrg1TsQVTrFNHYkruWtk5x9m8iNbHCYq2oTn
0+aQNz5S6p+4vxusEMN0OqCHoF8jPfnVyOpWMPH6IPKGijroAPoYqmBssn4K1qamPb3Gf+oeZTam
dw==
`pragma protect end_protected
