./../../../cl_dram_hbm_dma/verif/tests/test_dram_dma_mem_model_bdr_wr.sv