// Amazon FPGA Hardware Development Kit
//
// Copyright 2016 Amazon.com, Inc. or its affiliates. All Rights Reserved.
//
// Licensed under the Amazon Software License (the "License"). You may not use
// this file except in compliance with the License. A copy of the License is
// located at
//
// http://aws.amazon.com/asl/
//
// or in the "license" file accompanying this file. This file is distributed on
// an "AS IS" BASIS, WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, express or
// implied. See the License for the specific language governing permissions and
// limitations under the License.

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
qQ2dt/8Ka09Ompoek5riyUjmDWrffdrJNe38hM45yBGNF7vRmZwPuC7WKBHb1PioRiMekzSh+qhJ
Pigt/ewjo3ceKnMkMzpv2Xm5ZNDnAqVCRcpcSX4bE7OjxBXsD3SnyReDrogtdBToLn2ztocsCPse
55JsNzHHfAHNWezgZn08I2Y/bRqx5OuSQz8EJAd6pvD/7jCwYKpWKXdaeP1tuMIWn7xeRdN0+Qf7
GR5xzcnarVaqFs2gCTEC/o4FKrSpdd1+fbUZ1V5UdwLjnIiA5rjccrLa5Ma4ImKEyvVzCkmNGhj4
9anPYNCMYI5TUfaWd9AoNyEimOw8EWbOOG1Jkw==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
YjmgKv6WcEFWHhhWG0iEu8RgX2kEwBL5mZKx/bGuHocoku0vP7GuaMasD+uhAFnOgfO/38iNJHez
baH/+jfNJYRNcDIyCUseTHmFDpDEqOWzjOXItnPtoH3WOT45VawdJeNvzIq4KRJXPQ8yFuJMYH+5
PzSz8mq6j0a4oT0YRK4=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
a6rbR6JBnkC4wxTqHQMDElK8UK82D98C984iQMk3OgI9UtPnNUm1npjJPj9Dh5NjJx2AFugFTXd0
969LzR0LZD4MUUj/HMFFfnyLcG3DsUwQjSQNprl56j5CKgMCfvGmaTWEGeKrN/2hjP3gLNcxO7aC
EWqavW2uYmo+LUEAyrg=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12208)
`pragma protect data_block
rtlGyVcFbidvecBeKxyiPiC35qr+4UeKAzuYRvg8Ez3WK7ZHQ97mGqwT8o+rFQNOlbaTq8Ag9oed
xRSm8BJ7BiFD9/ctbH2ZeqPSkxQ9D7zd/dkHGj735UOh5zEqHuvra1Z9CVnfYqYKdtu5+pH/nEHF
CV8NIesCnF1O87A7ZLf3sb6Qv9quj82C6fYLROVBPqKAdWCpSusDafob5mS25VCrbTU3Gj6rqFI9
dHMkbRD7pgMl3qCiFzy9VywEyFMN27dPQXZIDHjVszuS1cAET79PiB9oUWBRc80QvDM+D1sq/1hL
4HbwftgZ4Cw15sV1sS7pTdw18ItcMN5rSaZDZqBuqmsoB2xsHTxfwSLvgaoB/9Fpy3P/j7ETIlxB
x7qPRJ5K1TeiHTU0MkIx7wm35L5ol+zwi180AXQaaeNJosw4aPEBa8UQ51gU8O8Eyeo0Vq1BhCZ8
TxU6QEj8aZ5ncMFVpYNympDqmrX6Z0wQTDMbNNTdyqALUIJAX42tDMBYfk3NRsZnXsV2fmbbG0s0
3zZgAvKM6wu+FXlbRHD5bL9K+xDC9oFcw1zOa/J807xddCBId+olw4QdIovSFMZbtEWpU1nv6EtP
3eDZ7DT9uy2mCnvaWhbUr0vIFZBxIaacE6jYe1NVYXrLL+UDm1IAPl8rBKcQm9mGxeANfr8ig431
hogJJ6L5gN/R2lMAPD3n2uzh8RgqNP5sEV+VuHU5HofndQ5KMH70B+ag8sZ2QX+1ZvNVpCJVScKX
WDV1QOOaQn1PByAfWnJFANRfjJqn81k96FOZgpoqroEvaMOU1lH5oLyqhLiw7A+Uu/257TYJ9S9L
KXTdlndu5WNq2S66SOG1suvALSC2xEzms4aJDyH7Ml5rfTaDQHZiYqQqaDUwKxsLRViWWzmMx7E+
ziANlUy0pvTY0nQR4DnJ1fnIsE8wz97k5ecd3HmX7p5qg4+DPlBkpmyfhs+OUGGXtADUt1cvCWuN
KPVbkei9pV70hOsd61leHf5vPbyyPMS4F717Dg+p2LGit1Ug9EAQuJrXy48nbYpgrYfFNimcwQMF
xQsAI0dxsnpTw+aiiXIthbNzKnspPhmKXy4/bLj8HOZ+8UEOgf+g6pzGs7H92HyS+0i0DlJU1n2J
DVF6j/2Fi3KeCzOMxo9si3GBj+2XcXDYgucvaugEtEPbDHmEvoO8T/N1JSWZouOIl2aqyq0vnaKW
tBSyrJ9grhiOqE6SXjXV0Ds0IifCFADOfv96RxmTnIC6V0LS4ngbJsXQiYDodnBoVVw69OjR6vEM
WABlLuF5/AFf3LNi3+QiGzyOCbzNNtItDTUGshrACKJlN4ApMU4JEpcWtzFxkpuYWeWZW4GQQPBv
xZAesBDy2P2a8pJKYc8Dbz7MDtDf8ms7sgg15aFtBvcCLk0QWqrYQFPAMjFB8bSTUhYWHYmWAIqj
z+W86FqUS3TB+m0p8ZC1sowbKqEQ2ClWnPRNEwWhy3AmODWb30IeG60mqP2t1qMM6wAMn2CYjOTf
bMYxjCc1KEWLF/m/WINLeJoXyOiAquc5Zg2OYmjtw8Z2QQ86X6hOhLUbzvr0/TGWKkLKzKcSauuK
+RP8Pm9MpBi/14rryiRHIW10Yixa2PKVD3Dbdq2WXf7thl7mmIDGzD/EqOUo+6RRnL74bjuhlTF6
JNW99AE0F29YeVnAsyLoKKzFLgFUrSPZMvXsZ5735ThD1mXWaWLpnp5Gd8rfOFsz+xY88CnvfHGH
Dfs1t2ffL/nh1BjEaDxjJSp4IC3ObuFVZmPy8HFIB5KetPJYiMduO0lJToLwa5AdW7YueRbwNQvT
pCY/1FZDqbxWSTISPe2sZVLyVhJSLIbNXh9bJ9PYxnssT7rQpKVhsMyxa6WiDUhIOCF1O2ObDiw0
278vtNSzFJ4xH37jx7dIGSMDXddz1ogtVFMKy/ic669MI+983kSYUUJsfSx/ycoVlz6gWqD+G9DW
lYnGT/Ep5dktvRBq0tmg6u6Zxnc8bio0bSRNwcXjGFv4XpUy0zRj/8+jBPWKkJZyhR0XLaVeLSHl
rAvvJr9Iai/eOi0JOnp4tgOG23gXNo4yGlfLnh8pBSdaRD3sGfm1vSmwHKwI4WwTsaBzgSrlZ7zk
gI8zdo9aovLKem6wvRj1AKlaOVNbJ3Bu2eXzQPvn+rxrB2IFvox3PHlgGmJnh7FVoACESwA382O6
TySIeehvbFfHo8JQgWZaE0CYKcZPaaQmnGbEhB/z91f4Ppa60HJfE8PS0EemwtlaaLuQfgr5U/Cq
T403J0C5w+Mxfz5RibwFuwD+9g8SwTNK2FqL8pu73fO/DAYmMzolGEhPAhioZU/+j2C8MDFXR0fd
WR+rlidl9NzhEUvaKeb7LaZMFtkZ2m++Gn0aEM7LR01ZP/WIrIbrv4NSTzQ5S9YWq2G1CDdw5Njv
hWsdh//Hvc2A12ro+mW5fAx6Btab3VqHPesE2lKAYfWGRWHKuTtrAZd6D4rbuTrAMXkbdilnmog7
h4MdnUagf35zN08XK7BMMDclkL9kObukFBMYU9BXuyy+EuCBpgXc2eohTWsHiWqxS7h9ZwPItyVW
vx2G+AYt3fU93w7KmUcG1WDKSht7Ud6unHTCX+RLA2c5KlV2h0GZ4jSGZvyOEggN7/4VWW+kdAOE
HN47B3IajXJjUy72RUobmpgWtL4WfG31aeN3YY2ZIXIUI3GBQMQtvPHg1E/pH5LggNoYkyGgBMBS
Dxmr8tCgsaFkd/m89GFiNk3i3qWqfesp/a5vAMH2VM1U/ngXGyvq+rcf6U6fCKb5xXYnZV6nE6vp
c/nEtgA6bOpYPvNtZ/YFOFxQ3ogBGfSn+RmPqGOymet5exZ/iB/T2UTYanCtFeB1iAMXRTbJOuft
p25c9tyE6G8UZNOkwtJnYjKi5seus3VuL/O2et1WHNBfsUu2XLWz+gLYoQiCF77HmMDN3xRGOo9B
KiWlHdrP6EL8e6h8rEkTOTDeLhF6gjkc/2hkHpMKkAtH4PX5HGeHbxv6VVR2qehh1eg/wt+0kCjk
jiiO8UFtChR5eHhS1a2DF4ZVNhIuIm0jB4eI8KlTfUG+98ZP7BvkxgROVbPDEeipV9rhHVhogqEK
quRaI6oril/8BBSyCbIHgBlK7aZ8Z7Tk8RlGU3O6kExaC0rmr3issOdbPW0/uWHJUX9rVfqXnKBN
aOL/JXeTFgcPXNmZgCuAQdqCQbX6uwf/hUIGXiHdL7cnFaF1KRi+7iN5+4DZEkju/ZAzn5Tf6tvt
azEkt6uL6u5k9Q+p6YerVUVsJdT5hSsxeM2GZW53bBQ2bGsMb843Yol+9J2rRAjHWr0N+dU9g4wt
6qPOC5tELoV1+QKVYLeDYBNQj5JxnBtzimlZn9Zf7o7AGk3Z4R210SyOIK4Ca/2sfSpwquIwUoIt
otsm6AQTWtNwPcceZeUHq5EO/Q79EH6DpXd1BgrI+qwZp1TDKZiPAHQ0KHZYU2lvYnPe4JaMFdF5
3Vk+ZQ+N3oVYF+5ll1aEP7KLBtaxX3FdccR8IyauCZy9JQebk0R2Xjyuhxm8NZCf4B+TokxnVPoQ
HDgBRgQIc3UZ38wmV7kUBletr4R2YaPt254nlq3pXbjmDpcgazbfqjwR4uc+gzWr2eGOp4yw0HCL
PERb8hYujbqWcumPqtua6UYskf9Ydjc0vAZpy8igVFe9nb/RaCwueoF9qgRZ7eTDe88KXUYZkwEv
fur6vO3Ft6Npq6vWA4LsKGoZcRlwfnKK17xu8GiSa5f0eK33nv+Phb5q8YIPNIg2JJtq016gzL4U
rD2VBhnv5b5YCSXXirjvdTSMXxGIZGUeuof/dItXUA+bYfiETHFA7lb0ZaBDxY3f29H94n44WGpl
czOx1FmCBButxmfZ713A4reVWaTzHSiAwsMjD2gVIMTm7ylXBkDmXedNlqOJCb2lZ6JuOJ3BmpNf
3oFYLYdy7fTB5DxuwWJUXFhTsbyAhYslzuI/WhNUt4v1ybxdJ+FRUAsj+bErkrx3hPtiwyez0E1d
m3BJsVZ1H8TB6B/5vP5AHNBqRA5zSFEP8A73Kpbt/IPbQaUbDAuOYd7ogOAe5GsDaPv4FqNQaJBj
9730Nw+T9U6FRHr51VOtNGIXDUEO6FXni9y6mnf9Nc3yV3uryRX86dkycUQsn+ECxvM/F+vntjFX
7lSQDt2kwdvbSiI+2ZSstgxW9To1twM6c3LC82Yg3zPX609Rk+GgVAHJLMEgs3JxR3fgkeQk6csm
Vq1+V4xbQsZe+0wRF8OMZ4416VOr8NtS96dV5lPyg9ifYaYNj9eo440qkrWvmIkV3HkhAeTls8Kb
X5jtoVVZlP8EBhjMiJKf1oO6hJOAxv4SXz2BAfeM1O8bYNZiWS16IXfVZcr+MCoYFua6F0XzacaU
eDKRyGg5WoYYBRJ8IPXpL/9pglwHWbMtSmn+MXdAAPl0QlmGzBOW3EXl2QNOC2kJ4A9HltrLx3FZ
otisvPC2aBjvrfqvMsZ3gfeq8Dz0/ByKDMEgPPe4BkxjgGDkSkApIeeOQNcxGg0wXOhZyEaoA+T1
44sspNE/DYBkBtQpyB51Zp5rtR6RD6fn0hTd5f0P5uXW3iU8Jk7IzeIUOieTW5LlYJqTiJFNrlzC
n23SORMziOHce5KHA6qsGLe4648fpIyOMxTqcEvZfHs2y9w7tAS+d9dsG68XhM00E3P5KFQ0yRQc
Bf+CK6YS+ihEztQAbiDKZX0+3s89JwYKhaO20VosFI/R2acR6KxNITakfktfHuudo/v8nUjAvnLv
yUz+8UQRmDm8yvNPQobaZi71ZYYUW/ERoLSZZdC9y645VekXKkNsfCAhuNaO0IcFD03oz2v9ii2S
jFMB7P3oXBK8qKNdeWvn1AkRV1Ncq1B4B3gQEhXr2EpIW6axhbXU2ZnPEx2BHi540OK7Ix47Is3w
4IfSIekrDhk6jkeZd2/HPGMlpUUNMnjAqUlmCOItZISwxPrXQrbQvs76Xzqhmyxwqq6D2gakl/ww
nlthHTXP/xX103u/XOkJ2P6meCgYa1iFl4umADXkW2uOBcFDBTbNV3Yff0nPYrSyiIOfKbOrPQfM
rKcbzc2MaBhQhHwCxT3ZK/GmIJRx3oVx6cEOCcq8M6HjNAh1E0BIDEr/yjTFX8KltD4X82NGf4j2
Mzb4fPPRS0UhiZxJ2QvxMZlX04x+6sVbtgRBlzv1cEHG6yglnvdJHgRsGlTuMQrcHkJUsDZkd+oU
9AVmlXVQsHXxEuLapZ85jaFlyb8vIsPK8m4H9iDvQtNZL6/ycRaXS//iJ/EUHhjkHURWfMtNxKy8
ksJXUP+r8XRA30mgyZoo5W5ckE4cJgJMQeUvhjg3+AEtGrsacOVKu1jpRQX3LrYLsuqY7CAKBakE
vh3QZtgKTTNJrFrg8F1PU/srvBLRU+KMGzlBUO+0SMyConNNsVFdUFWI2sVsuV8No1DJSt8QvWOS
Nmy8VibOiAKpjgEcGr/fXPbvMZ+6YkOUVePs/2jDKMIwvld6XqHLCvSZoSifqlNcaUY25PimihrX
rTUPaYv2Lf738pmn9uR8Ut08zygFD7pXsl8FQ4tsXOsBsPaRmLmHmFXueYzE25e7JYUyiSXqFXtr
IIXiPOMQ1aTDnm0P3q65zaDsEGNvqLrt4HP3uHDkNDI+vJYMn+vKIUdL0NYRxECxr0mQLxGxzRrm
Igj9PJEJiMOR/EzGnWoXY8xqwTmiEyxAk1gqtyHn8mNji20DoAq8uo+48cD/mL34xs/NutWgP8UA
Qw60snx7X+oOW3/yQywL988jCOSz1uQ+bLwwKNcrwNj78DLEaInorUHyxjJAjS1Op8CNhHG7CKMt
9pMPIJ1GrpyIHrdJN9hcwBhtB3sJQWswh9sMeQ4SE8EAeSxrijAr4f/zJWHiBlihMxAGtH8E0WWm
mxbAFnmJMnm9LP9iygD3LqLtCAoMToYkbFu4gYGLgA011K19yeTwelkdXO3MN0SUSSOxruI8TnA3
TjyxsHT47dj2QnRuskBLb3Rb+nui0eIGRAZJk3BPj6CDnvn/iDl8Bo12/kG0FUnf0QqiKxy/3VaV
GPKfC2dv/5/ta7dL796CEVtifJY43Qgl4FhKSkpCI7D/4EJRme5Bs/159jJgWFN8rggOP74NdjBO
fA++6YKgj+dTg4Rat0Arj+SqG6A1TjJv7uVU+I3RTlIzXMM2qgjvl1L15sPrv69D8u0TsURaAR+W
8F4Sg+F1Oylk1/PR/SF+GEnToTanCSFfFCQQ9qkK+PjP5CptErDoWe+lE71YHbltOigMnjuyeZGf
DajsDLI8U5YLcxJwdh2vzRwWuFpT/5v2HFvnBSp+5WIA9/AA+/8uIu1OMoASbXsuH8XrP/HHTHIH
BuwXS7q5aVOlqx9EVReEvv+LmR9TNyWgVLcQKiC4dQpkdmlCXeA3kqRboLV4aqjlJK3jM4MeDRNX
S/QM+Ju+YY8B7r/3E6gtA2BwN1hnmIV5uvyHJPgFQVHAR0XaBH1woMlf0k3AvTp5VzCajvv8+VR9
VXp30bLDZyIAZte97Ygdd6Jw9WNOWexAuvCaL9W+LPywuSGz2/h6CvaOt48wkXM2fGtRLq1bRXgR
ZEpLW5MpmYfwHInEz2WKepBbemKJ7f/z0IHIuNJFiEQ7pFiLpFxT1G8EoAeV5mpJzYPVIei5ByIs
krloH5j7FgNaWhABBNEqwqw26lwwVC3iCq8nLjarEvVjjQPVanb2ZoAPDfQlCLYwe2FYALZ2yyyP
RIkXimwECCwZUdgiXqROqNYTd+8lwYo0eVx68a3ynLOWkOS7Gdh8n03bhy4D03UXYz/bSRnPuqHp
gu6FAM9p4zkbjjOaCkYaB2c5PKl03OnzqPf9WDLOgBDPMPGVrU4ykTh6adbi7P++rhDmzHf02gpD
D4TEsivBZ4y63NLbMvoQK/a4zXFAn+Uxa3OsZTekcrO1MgkxsVw1vJtPe4pXcHhHVCSAhLFHlGeq
fhjrq6wcBr6HUVQJJWHS7Goeu46qLDUwN4qcESeRJknQ3szdpSUsN2YF+kqJ6PnAH5Thx4S06f0w
+3OWiHF6L4eS7YolHCp+nehqywmEIT6iLbmPoAms5tEyiFgiUmrM5bzDyyb0yG/L3q96ZSh7iy/z
0xzyuFBJCNEXIivEg0NyhtLyQXe/o++abUbXB9+y4j1akg0JEoovBuW5um3qLR8FKMAcO+D8+8Gw
+l7DP8lSjtid9Xy/KQx5P2hlqp3kU1rli9PhvzMu6xMWTmXz9kPCUYaMW0P0qmL+KkzNEhbWKr17
iG3yVdFyo89nTkqEJ/jCHncO95G99+9jAIzyOrZB2o9x1ZzHq3nMcQQ7M//Vq64tXdVA3/4o9Yoq
QWk9gYiB2o6JI93k03So838YJE1cWHwz8MJVE8l8UBjdGjU+0wyfoym1RTq4JQUNw7tUuGgohK+Q
nnzdxYUVHc2JZZCEyC6TIFe39cLJDqWZ8ihef9zb3S/etfS7fnXSuGNbrx3UxwNg7WNnhGRrfF+o
3VZuqWgRGAy22C/iZFi2EvNmS66iAW1+wVejsfPf2kG23jetz6y89mkz1UuQCxa9nbnNEMmbiuWI
ctd9Rt6cne2UWiISarg900tCrrvxlL5DoC3WH7sF80WdA+Ere9Q9Qm8fMRHwR4jVOTWnBX2l2/3X
vXUBZtYZpFn+rByhAQmp3cA24xI7xL8kQW3TyMrTcwD1fF4z8vIJGQiDbeiNp975MN5Kj9pyxzw+
lN13lB+k8/mLELHtRRFe/WeWWJuE/hyLeo5W7zsxKFWxCeuzMkUHQBjyTi6oOzDdH334Ekvz0tPn
c1+IkEqehkfiBBc+TxFvM4/B0SY3Q8KJMKfz+xEaKlpl/hqsfEl+NmE/qzVi7Yg0xx1ytNMNfBEk
OIuCDIPM9zCuWhV30kBFbrsECyH/kQZU5IlkQprnU5AGpypJtD/72Juum6ceUgc5AxD0M08PZpm/
LwU79v2ZKzFlvs8hEJuSAtWXfUakoIfwF04zHoECEJE5DR+PvXZr++prt93J3qTcI6X3D4kNVeVv
dJL0UjWd3jaBL+Xj2G+cqxYDQvt0y/XHskEj0DBdcnacgdhAEuMdr3iOQOdQKu0CQbadzzofglu5
GXUyo9M4zUTzO/wXUKYhpuB2fTKYx1QNqnKi1DfEzJGVQUomOGzxDdm1wqHDajCD6PHmBGL9YwtR
Jw8ILwjX4SrDefZL4lnpfJ8fWmIT/KJ4GPOa2BjVsGE73cUVxV3GHVKnTigK760BL+Nowf18n14s
O8CqSuLczpT2gkO4BxxKD7yhRM0Lz354W+uvxVLoUh2ubVHLdBaAifqH1OJG5HOnnvGmpZH9dZtv
BlmHZpKExFfW+VNFBB+a1ZG/3s5Csq8zwn++mp/DKSmWynmO6cDiSzTaB1vGy+AFSn9C1e9AzaXR
OEm3AlcLnkamf4A3STv5vxCcs/ccL2GMFnYIA+3I6rHpC0+qIFi1uF/ZigkImTx4fZLokP+mAUyw
cBnFqyvWSjx2wbviLwq9NJYFLJbAXVN+4jdNJy9r/W1xUjjsdC02KCKL36RypqvG/w919V/juAdc
tyw/s3t+TUdDdugp1nwlRISufXtrUVcWHDCwxuUZPI8FDmYQ6yHNKQ2rgxeJ1LYoweuhXAZij1rL
CiZDYZUvtyYoiRcGh0yR1FA7vFzAACVHAhjgfiN+K4fCzs7niUaFDdFpqJdJkyQssmD/VekJIjCd
21iZG7SUsHVk1Ff9eVZx3AIkU0ys3X6FZQi0xpLa7Bv0SocYbuV43djIpBgXIWpuO7EofUXQhAtD
B6Lsa3nIz8FJMr8uKsOc0UT+NQAE78y3Zfcoq/mo7uFCG+giHmF215vgtaP6fP9uOigYGj9XR5Yr
LPOvK5j46UAmDm8qtOLIx4zvIfxqKhPqAqh9GAwfHdDb+7y+CTSBWVMd0hc6hWzO0PRqs4W9A+S8
ckuDuZ1FabmX8xEwk/gNWV+wOMPqZitIl/LfCqg9IEL7KODHBzs5UPlr7lc6gBZh9tvMnwM7uPjC
DCfuAjJRYzjujMafE1ZauNDPABZRkI1F1rhz6MjbngDCjmUtOZzsbtZyq2vvpCrc2OLSro7tESnz
thCHgjKZJ4k35svdwC/e3XEhw7NJ/WbGbg+13FH3hDkJVzcXNu080r0+RHlj7F4N5S42WieP1bnx
g2vNPY2w6/lShKv9L11ye60QYSsMUU0c+ZO0Y9uwOO7KuFFH6bjCqI5AEWa68XD/u86zZ+sOwtvq
WUFI+JE1PdSB1qcI0KzXAORqJPeoMi/ZpYtqGhIeKev+WpT48BqMqBLPg7QdkBRfHzq39nlsmETY
UDYYiNRkgyYFyqZG7at9EpI4H/gW1cKRrl4YoSYH8b/QgT4uaJq4H+DgB92uGTAyUD43RHlvrPCU
9b1oi9KpW2ZK3hKLvRjfSYttwHlG4RZJcenhUT5gT96fhfzSjC6fK0Lw4JXoWTZTNnXoFuLGGK0V
4GyidNt+23oJv0XYIs4dv0/uloY+2aANPE1g1iuqSGQgwex8ELWhFZFgR6Dip49M+VQjxh81nxef
V8UslbmaAOckF1lYcGa6XoNFGi0qjSUIEqmHtURpoKx5i66I3Er+qf2FvzyX93gbKuddXB47HW95
xO6c9lJZxvY3iFrbEhqrU4XpHwD0ywQmdEtnzv7AYhsqSbDtAu/2NZU+2X2sYRxMiBrVe+hJSejG
zXpjLgos+UOlJuJQGsu6ukZWsoEpHAXKAPVS3XKNv8kOZzIFsutKhn3nxMgj58GyxnrUDRIJiLYa
2Wa5Y5Z7z3rpNyEUJDRq/xLvhPr/HMDx9GVsJw5ehhhYR+I312bwJwnFGheX5u1nMw16yflUxRuz
Grp/P3a4PzOpnMNexRb6nRGuklKil1kZLBQZEclJ0yZp/po9eskO0O5bXodQFgBK5vYv03jRPnj/
a6+mPFCoUlxFzST6NuGTCFrvWyiMQmvuyzaMqXo3Ps56RdjFhsKAgtuLv18ZkBoc4SRonGMBCdU9
3R6ICmTaxNhjTgQ7qtH+aOsMeZm792vUGL/qqSUSZlsjud2AIscPKLxnV09qDkZ45gpWi9F8bXGK
/zt+fLW/B4MML0lnBEdoJatSvhn0UieNybUj2sWh1vcLM+L6ksGpLQFCSjq2Rl0ueHLoeh4LaOd1
XzLn+VPFq5VLw8VRMa6mQp93HL0JUZGl2Iye3Rm7lUF7nESENHRDsape5+6UiwvA+q3TdPJIpaCZ
7CLdOhQU9EU/v7VrOPSvumaxKuqgW81PjnejSPflChLhPoxVpHdL7j/10N6DcUSPbQeHHFH0H8RC
a0UKqL8qN97j8TKb9gHQvV6DPjYe56hG8z5/BD4sNVNvrV+Gvjzqd53GK3vcdoKJmmccH1wUhA0x
UH7tOyFlDxc/vkngBhN2XdB59/tiD4zpzPX4hAP9U7dsVWge/0CPLpTfYG0711Phku10KV3jtfm/
Qk2UaqFrEaXUL0LNvOLBi8tMGLw8N150wX2mdvqX0ENyjUrb5PgUfVhmQmSAzssV+1qnE4ZHhM7V
W9k7VfkSo6298zrsqB0PHSE/m18G1Bx/N5u1dPm2u1+m5rpgNBt/NgBYoD4wz3qc1+78gOo92NSM
SPNdx8+jaTK74KOn017V8a1HpqWvchR/9yi7WXQ5D+TMRSwV+q2dLZgbmmPfkIh/pcA5zMTsUi/d
0d7sR/Y6DGlg+7n+pi/YVzcrE0RjU87vBGXF8GA5NDDNbDEkwsO8gIDM6NdwwddoSSoCsDQqDa+a
2nmYk3buSeow1cbyYRqG7bhieCWIuAgNXDIzpSMyMkMQxCPZvNyAv7ZSmTwloX7IL4T9Ej8zQpPm
FzDYRTJTbMQaNBXhagqpOWlrzETS3SW3ia1L6n69DmOlAeX1GObdEfESkMTJ4bIznJTWAzP5ogjA
ziasUgMUQb41E9eK671VejQEx8LMrbLLabpbt1crST6wvtxgjoOhMAyMguJCf86xhCtzMOvNXfDv
TnpW3A0Vj3r9cfJ6l2ElTUS27yf2BW+HPKCFSKXeQyDF09x9ZburzoWlrqXviYXMPFBS+iDkljjh
GtSmBkhjnsnthzjJHipDts8n/JcGZtl7UhjOFZ4UGgQfK8RI0EZ3J/1DD++QKr4p5d3Zn5hJ1FjH
Pd9TFGp5/CY6Mu5AkmBfybU2ei0VmUg4hIWFCDkEkvgHpoLMk5UvF+0iFhgN+UMIuteLKgkQBBX1
d6EV0dbp4wbDlVPLWp0nS/5aOqFeO6IeB6WjVdy2tLlEFDEFEWevz6i+JSpHBHCLSIC/VVMx8eEH
qJJP0MXQMx2awQ/ki+a7yysho2GjsFvJ92+YmBJQ2mr2TtkFZe1rWtSlYD1evz5p1Y0MShBI69lf
YYpqN5+5eitVLWVDpmaN0JNtvGfJu1nr6GSDIMonyUp+LfTQXpI5xr/UpQP3poL0LsCJn5SX5Et4
pkL2rBt2Ov55jEY8Qi8+CP9lXwA5ZFGIpBZWnHuCLnudL/hirNSJdOFfBmvdraJ+NJ+EAQCHhyaa
TkZ+mdyxEBUeE4LrepktIJ59UcqvvaJv3Gi/tqQRUWTsAzYtvuEPj+VpUML/p9a9iZBCSgckEAxQ
IEb8LDxeHa/xccVFCUgeIsACVilTUsztTR3c8e4p9qFXhRhKyDVYkD7rK+H9ZTCtoGDeT9Nd3UtU
iPftk6B2HI7tNpMMe3QSnLlTDbs3deTiXaedgE39+9WRYuLMqo5D+j+fx8KHpgiXdKGEgBi+aYpc
s7aX6CSqCTW8qgKH8pexg4qb8s8or9MtTAYv9+4Vqjq/427fONYpTJP8hQpRhWLh+toeZyIFzxtK
mTS8584nM+89e1bEy+9+O9PXiqzsDyvtN94vLHplvKxmuCF2PmoZd2/XGaefjegcj+IjAgPbcMGw
IU0UWxwoIJhsX2ZyadrrAeVj8Pxuv3QxKKJWPhj3aqFwE/nOKT3VzMBs4xaEJXSsdvj04BJuRQQa
565Gte2rUR6fY6ulczwy7C1sHL+y+h5xoVe7tUn/7jEHOdQyoIcqLkadq/COJJbpbIfU3cQ8Fmvi
88lBZ+UMw3TTK6BClZ5SplTkkyYZUWQSobsn9oW7Zt2NLz4U8icaP3F3qb9k5XWv5QcKU03uXUh8
eodNXQZW8fJntSYpdXJJKf3P8oZtflwn+/E3HD+7QW2fRwY/O0fK9GB6pJIUS+YoIR74BzKFdBNw
y2NLShyjil3T7hmYUpN8bGGFb8FExNVnT3ChmalbBEPTFmiDtAfM+IGjmcUqNBz8U57/YoT4MFXD
/dQ3Rcceh4sI1oHQktvUFrOdB/LoEXQxciNpNHIFjAdiIcsY/m/e7ALhGyYUxPyOXAobQSEWHqfb
SgD11a0CqoZD4pupZ6gl79TF/xBuL3n0ChwdpLGoQJOkT4/y0lKwax1aHlt8bYoFWbQu6TjsMtYf
ROM41hfCun3cm8yUGLWm3wBTA3w0PhRy8mvyNrcwZdzzRWdTzqRdWOqWXbLmmiWj0W7O3oKfle2l
SI/XlcKCFgZO3yW3Ah10uZWSHl3IY2EYuMLPTLn061RBpqJ+9CnSfw7EyrUs5Bd5rj5UMo4hhwBQ
A2r960xz0cg6sYWIa00Ui9Bw3tLI1jeWoU8PArVGl+T2wa+ct9TzKWc5EL1YGQacs/UK+hFpTiwA
/3JwaK53CvfoKvwgOagC01lh7eScS4xnjLIIPRlBAgY4i7HZ7Uo5tqC32kqsmOKMIeoDprdzLNC6
LtunG6mrkLx9pMUy9U1u3YgrzFklQHRt5mD45PS4MhSzSJFgQ5Zc2vqiFe75+t14WC85PIu4/S9H
sGTMNQV4Emnr2iMf8hVXYU1ft7cFcSj1pXUnGZ9sJkx8SxA79nkTx/63x9wbqC9SynaFoKQzWCE0
JF4JA8jmz0MCiQi9EC1fhQpHxVVlUEqWwuaSqYmuuV0lTHz1h8Ljcc1f6FClHv017CRUhEi+8grW
+AMSlTawGWTMH6dwObpq2GT8T+Lo/Pft+flspiUJZs1Wp8oXMQpEJ7+JVCsyHfizQy08wJOCvsWm
+HKRZQ2I0Fgc5IbUFHhNfnFR53bC7AOML9deEfUyXbWfaaMHGKvy/DOuapYrlSjnwdIplsOX7SKN
aW2EUQ/6Bia3jdURtxVnL5+AjTYI5cAl/tELoY2RCWC5s07NrRjYG+y+GBmOPwsb8ONXSpfvoXRP
K016y98OKiDBMgspxYJ7sbwrQhfmhzBjcTPD2U6VnDglsqNeeA2kwmOuLeolg5q/XpZNjOIS3iuB
RoK/rY7mSx4l5iSMj8cB8n0+amvB+m776qShNvMifXKtRSgFsYG03J2nB5bVvD7EiotOoCMlLeXW
o35hqDcI6oQ1oRMSsh6u5EeneTEET11HGvfH0dm/ietAe2nqL8B8KLSiDV5x8GSJcAh7REAvSnHh
jDRo+L/uxJN5sIEmWLSNKBGT3U4NC4kT2jON+i2ym3xFxgnQYRFnSj8zMJocQC7+AVat41bRlmuI
JARWdOt22d2BW7x19LX3mEXymW5NPN/51Z1xG9kl87dqdIJEazGDT3FPVeoOmrActXWznda5mVHj
8hIQj2MXNl6oBIBDwUJPF6GLa7btdwg0SkNjko5d/00zMTkBoeBGvW85+ClgoXxW7vaZHc70kLXK
qNPTWXE/aR6bmtkIPqkwj3LkvrlYUU7cyR6ckWXGdbxbtotseZG8Q3pdNgqGhuMPH2PWahJ6dIX2
RxWmoD1w69gzCWOlWZi5RBja/0ZRf24z0PPfKeuEVgJK6tdFxmO08JZpmttYVzpNrNyuK7p50FgT
gyk8X0n2KAMuXjjU+trLXioso04dpbF3JXAtLW8gGGqDffhYaoqpqoMkXSc1+eluQ0bvdzGIB3/z
qoMg5XpVvWoB8+dRbLTNgtsK6ycqw0U6RF4a1CHBxC7lylq1r1uL5KuDNVJnL6ED06f2+Oc9qWLo
8aBsQijD8DC4O6cxr6dnGLA8vleaKpF5t+3xtJvblTMn7PeF4dQSmyOoJ8M92LvvDa8DCyV4kOGE
ljzTl/eWzV27RlDz8qN5uVNHli+uNYPl4hHsnfHZx9NC+yq9twKZXR1tvsqr+qEX4+ioSdbK1s95
Kso2YXmcWnBVVjO+lGw7JTR2Bt/4U+I5ynFxMHKX1LADvz3bfjqUoCNvJPNRV/XrpQB9p8qSElCU
KD4leOBq9Cx/ynOgbs/3OKyHWZ1qDq0XOaWxwRQhOHju+vZLBpK12nmpuhm4pBHZhfpNIeyyXtWs
k2XLnWvyZnjksFq6q/v/uBE/oln3dPAcShiYQ4ev1602JGDfyp4Wvtp4ABQfepRLID8Yru2Uuh5L
j/KJnJpSULzd9hNAjL6dCNb3drQvfV3AhsHmjX8WHPmEGfS+v9Ea4DIYLJCCtglR8MRQ23eSSL97
hV+CIvyYyvr+qIfNJQMfPKj4sMhBZ1OQkwJfWZ87NcE3+CRTis+p4MDW9QFjXBwfavsbI9pwmoJu
w1VRobb4J8o3KOE3ANRMu6/EQNm4lc1zkEJdjF5JISBRjKc1ovUQuDIhbVwtBvxtQE+W3jtTzyCR
dSwUZlKFgiMVUynb8WAAy/Ze0lHa2vzZI2XLFJ7Pjo95Z61hh7zncsuO+SqLHu59X/Om7bQ6cG7L
8ID6mJ+IbIpD135x1fNYtpWLX1y17hrNPM+as0P/VVXkUI/DTwHZmlwT9A/u5+hwl5CZzNZrM2Ov
WKhe0ZYTXkI5AbivaKQgVNHGmt6Q1PuD8O1WzavBdGZuy5KkHMRw8qSX3zAFJ/2Mv++volg8teWR
wt7qboHi6aGxqSB4BxNQwDKMwLjQKF1E7BfsiolS9++Ul+KkmHQB301MgcHdpyiYK5ncZqQ4zRe2
ZyZZKxo9FfFEUNtZuCeZUlXFKFBfPbpDR2Frz+N5MLe6twqcgF8i6KnYwknREhUBJT0qGQSPQl8U
DzXsfIYjlIbkqaEKW+wN1LOuGOcD6o6MXpvDicOjS/ro18gEmM4FtCExhR1j7b84PuNnNMDas7d8
UPgS79o0QKnBFyYbJvxPdFic7mTKUNw0/k+Z2be7lvQ49ubwp2JyaUZx7S7oFhFny5xFL4HDTe8v
hMnVgkBuZYa2qof+gURJd8wDuhdwWgfHWQ5JPPIrJ/MnPBLlmhPzJH8f91aDISPukqv8BfF8EpV0
MDXE395Ztg6/A8seVm2GZTiLnyTMTamA0I27qBN4/p8lmjbjIRz6aZyfZmrvDikbzO2+5ibom6UJ
DKKDsYc1gkAbh1ZhFlBhP1tTI0k9xX/lgOSPiHGzTK/n7Ky8HM/uGm0aLJqtdgVT4w+Y3SDyPlPl
e2Ymf5O+KFoXe1hhAKS+Wra+ypJyXvwCqZ9iNtQnQxm8NNbNiNkjmleUICUt3JoIROXo77mv+4qb
880N62x0DT/YtSA85H3Z3y6+PJJRQzrA2AZH9VQiAHnMzUSycCIL55rMaInlfEY2PNSWmrZc8dZ3
Z4wl1VXcEVeHTQygXfUiZJVxuvaytw352HDQEriGpGNKbdpmjEsNBQ2pkR28K3MT782pm43768XG
zgyOEYNrDtmpgUHsZDloRbDeburToIRJrazzeCtyUyCGVVkU5W4zAo/ECKE37OSXOMfy00wwBmo0
j2y/DK7DE1g/cvB1hHIGZSAelLPleUYjGft/M9a50wGddSxeOFkvwRC84dzHO7LJBr2SIEQzdLG4
AnwJcvpAXu+gG7ZVaQwBWBZNfH4ICTmzfsZusSO+v1TV77panLt4/3m2zfLxsjKNlggN1vtH8N+r
BKAu2f1EE5OtxPzlxLk+lTM4cjm1xMiQfnBdH7MZWm1V1ExI/p6auGwGP/TzrTo5mcQ7XU4t/R83
nkf0cAyfKHfa/w7uZQPNBTnDOYSB6+YzHtaYvE+XGvxTeNVwujeF/wzg0uBYByox+Rt1Etf/CUm0
MAg4NLOhfapk1Sh5y9/OxzAIx/uauKvhj8edirO9aF0gbVxEokurFGwbht6s2d6t6ZkHVYRxYrdy
8Hyg5hRoGPqJdfQstmFTAlGwEz3riT7WB5UZbQ1zGyA+mgIdjgt4BmnmjnNHvlZD2GLyvDDaQOrY
zEs4fBim27mYL0RCS8weCQC4RSE9dPeRjL4RXk/cvtIfyE9x5v2A+hnrvmX0rY0iB40QEdHysD20
azSBaBmNa9AWK4LotjBJ3WiaQspo5yehkyenEVz0qyrgAI2A0GkcwDh1lMS7f8GH546oIo4Hv0Xi
f+/MfUBcsdVYVA==
`pragma protect end_protected
