`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
BKHAtT76jfARMqWIXDiB6jv119ZlGFVGlzNp2EC36MkKeV3zJzEYk1ks2Q/T/Sc68CgtWxagw2ZQ
PVN6CYWaxU0iWFGuu4/kbTOk15FsGmAzFZTKQrSEkLzaOipSpaiV15DSYnqgAILqhnLtv/jrxucy
KU9vCt9JWG3XDcT3eUzkpS1EeYRgGE2vDh9sLblnGuHY1fQ9nmNT0XWePpkZjJUJGk5eRZSpDeaM
6S/UjpZwqKQXv4g1KK9thfoKWW5LKK99i1Tyv6hQFZqCPNUIDwg+KnhBeEuR+NFA+nk5zi+iuDpF
8gM28xXMvL/axQQJCqwDnePG7OJgjkvnijxR+w==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
wUmlH/iYOsH2r8+9bWg865x7975rxZU7UKOEEmSsIgx6PbGNNBT9gtORTpiokPFh+K70xGEgrzml
eJeO969SlqM4kKxJ6biaSGvgLde3PFZrVbouYRa04T41pZD0R2EIDjl5E58RFSj+bzgMmZFT/Ssn
wcIPJqnlPkS7IaMEdr8=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
fkCWHa636QrFW6CyL3EtIlLXirvtCim0FdmHZilWL/TaScHrdGm3rxpWWtOl8eevz1pjx8xS+zyf
xwpz2qW8w4mfXgA9FnLtZycXuMMNydSITOqi6BRuKHVWUcz9WfyO9JUP7D/YVfEvcf6r8UPSWFVX
kPW2nWdqfNmYkBBIjec=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 37184)
`pragma protect data_block
rFoHClFBvoT+KYlVSrc/xciJc/P75G0P7p0Pb8bpT+Chk4cRYbbKrJW6pDbDaz0RN0VpyXnxY3W2
Z5X/kFkJZqgqxakO3OZ7rqVms0dvABqa0nqMHKMP7RWMw+V5zhZUFfD0/58aM9a+muXZqlA9gYQg
RqiTPshPbDZT2Ow6TbdIxlttauzKdr0eXPDmOTi50bFUXl4TGOKU1ll5hTrEnKBT3dtZxh5C/ggc
cFL2KDfqMib0aFwwHPN4oonxRnosDwukJtjmmFPyM5KEtyolzMvb07uFN1ncDzcqPqG1wfyQ5kgu
SjsjCpoK21S/emyuAivWolGR1j8yX58RKTwwgpqVUJBrsFH4fOfVFV7xySFKJ9QIWH4YZ0L722XJ
NLFUXAJ3IAQ8AE3CzMvWjvjpEqWxoDfaTEab9Y2Mn8U2XvdAu81AmQTgHPflBpdYy1nhLd9U/7xk
ULdb4jdnegDTbr9jECWKdwogwWLy+9J3Dw5EKqDIHAehrPbG4x0WsUA+ot2JAQDZwOWtFjwsu0wu
7yk+nAx8x//mMFQaEPF6tbonjzeHDKoWz+6dT+1R2BxrhHythJr656P5s7g07pDrFEZlCGGbnLzS
8xmWGSWiFC4X90Jb5hEip+U6rA7FWz/VZuhP63m7Q9SiHr+/OnNqBiZPLBKzyDd+SDf8kv4y99Kb
DkJG3Wann67PdHwbs/sKnUbsfKuK/Chf1tITqudWddfFocp4RE1fBXq9WvCo0rg5Gzhp4b0RujmE
eoPurTGnlBfwtV9dCBuXBTLPXbkDn1bds/gu04SzMjJSzCQhRvbom0nfPdQKNDNmTlPIcUa8OOmD
pLXwQrY0WQVo7MHaabvNbEglwJu+FvZ7PwotHCObgThI/szf5TU1peZNVrdutFYaMOY8vN/C6ksp
nb1H2eQRbP2h8llt34W1jBWMXVtSdLLTcmJZ9SZa9uX/dCuULwRvLaD4lHbH8aPCo/KKgFKtEBX4
wu1NCjSpat2UYi5xwnAzUPtc2ckB8qnm1lWg7FXybENoJfPoDxz/nxkVos6/IH2qgmZs+voJ4Qg7
z6je+Y5YBYqEg72D4e4N1brshXqe8bjPwGYQxe9yYtT/41omuhqGWAddMnlvg85uV8WSUfAcHhkI
WpEEHbgRw+xIyt0PQxFHrVBISunPSMJVqC8lUAQRqz2+1f5m4BdLpZEhELuHnqY1I08NeTOiPwGy
WAzUtUVE5fqzJiIwNoc2bhI34hKZSKdfqGFSVZ6YS3ePsK6pvYjG7CKMJOlSXoz5uB9xUmQzqjvc
jqGg0r3Rz9oI8Tiiv/n9hMH3Sx+I/HH9yHDw0/EONt1UxBpEfVNulcpl5xH0Wuqm7g0YBuHAARXO
3/bpPiPohA7vqI87/8G5hy+6uBiqOtbUcbnTyM3Itj1OmaTX+BjvQRHJD1e+InsEMscol6w0OW6R
1suJLG8ecPfFt/RyU8rTpjD75X1JEVAU1SdZ0NH0/9v0fABJhRvwA9VAIMnRzIjwus87etC4v/3M
NgP8LbG37ftE/AuaYh6PxhstzLl9BsxeIWxM16Rs/UFzRl7KjBDX6l5XCwPD1JwtKkAfFIjMGI/S
8QawGY9JyvX42T8VceHyxHZkGwno+bo1+Tp4r/14nci8Mhtd5h7hh3r9IjVwIIdlBSUFsdOfYQgz
wBSA/N7oxoQwUHZue2JIIRHh8nlkBwJB/n3dGWxcc5BCQrr3Mr5SEIAirhC1rIc2NNgBpVANRnw+
qDpNN9cT1Pd00BkRzmObicPk3voaSgIu/X1+LnUJ8XmMBKvD9X3aIvSRU3t6D5ldfrLXFDXX9QbC
j4WLQ/HjkRm1XxwW8p3lq95ztiIPX14khZav/tM/wZEwbGSudEDA0yvLuiVzYS/J6ZUDQBdNeUbL
kAyfxt4+yFNR7blscKKivVhnjzoYdWjtl9G8n8oDOLXr8i+5lRQGy58Qr+pmn9dv3hmcj2AwPXnp
BIHpSz+oNmWOy6kriliFMOW7JMf9LK0TsBJy2fntTDfLAZ5CPFtjFPrtE2nsOqZZVzNEpbbipmaH
9XbY0G0seFip7oJ4KSxhTsvzQ+6/xF3EIlTbMlpaexyRoH06BJ8+2SlSQNCEv0ZhUkdfW2zEKyfp
H/CWlngjxKUVx4VpzdcRvXITbS98H2jwz6FY6x32wUwwJ6Zva9a+L80jqbKB/gGkzXusM287OQm1
y+vPDgO9yxa50geXPdIL/DaDHXHGFIqsTlL9cs8B0NE/a6FpKGtYJ2jAJs+ClcoQoxJ/OcVXBhDo
jQfnQQuvx8KMIkxngm1ZA4LCNUrnPraVtnQLZVdchsdOGlT+hbV531nMZAdUkjOldJYTEkIHJnIV
882PWBq4Yo1xLkkWQi3dpRMLTMtV0Ok1T2NpgR+4oaA/gl404FP+6Ozty1Bk5XHC5ZBLDYK8fhcJ
mUuDy4uNCfX3KwS2EdhmGZNP3ZTbOquHIfvcUJ+swfugvlnBXcVaukjAgeCFDaw6CHG/Bj9ZsXlW
WvsBcXIjZwGoWkyl4Nj0wD+1q8P7E6wCRHxOH8HcNoGqsMUzPisJ1+6lVFBPLaIPPwGitC2yQlJB
egTRW2KEsVW1ZvND+NwdNArv0+7ieJ44rMC9W6x8JrjuJN6DqqMEOXN6kaN6kPETiHDjxo/78uAr
o2KjjuTAV0E0iE+ie9Va/pf0ykvvwhnrxmu/VtQ+xT/1540tuVXCaveMRHpzlvG65YBGYpDoHkbd
9glOoVwO+bW/6kn+UbUaY89FyEpi75h/cGCHEwCzP24jccOQ4jsYu3lQF6Go/2wGpDFzkrYqSpjJ
/wSar6j9pNJ7GIlhC+Y7GvnUCdCVEfqC4/cIg6d7z+JR4byqRmvkNb4JfFW7BkdF3HMKronDtYJZ
wxskB4JxMmH7/WtzI27Q+rMF2G7gpP/NKewkkGz586jMR8wSDT0/+viH1dTq1Jni6ChwU279FH04
gMdbRV63Q4GPSjlQnMGz9NrhVPLOFLS5DdCu/ErhupToD9E4np65rr1/gIhDuSLggW0maMdhyEY8
3ZtqccxLwBa+40mSCpb1SnRpTs2Hipm4tItjK3W4MAPBZ1Sv+1km0jETwJ/LlsPqrj2DwPM232+g
NPDDJP771d2YqinbF6t+EWDNL4kwGxy8er4UqtW0N6/mem4OaoArYWphSn0xPBI1kpzI+whodIHh
qy+mPhfhpGnVuhykSj8Jv5LhR0cJLTPm9v97DZRSmIHpXwCco5/neG1dWfxZE9J2JPxCW8b3wvSx
jM8+R4ae19SE2Ew1iqRyxSv9llVvvmxtl16eimn414yKvOKo1HH5EiZE7RWRU97XGaZzy727RvCP
0hv6DzeWOGxDybzxVMyqygtu4RwLZdJnSn9DM8hm+2jnJrjj6XXdPkIqI27cXdrZ6PJaqsaf2ZpE
Fjglt9xWqHqNq0YEDWVV86vFu4YsmoL8+DE3kqzCjmHAp8sdzYGYsv6bssShk2raqU78I1d/dzqL
AIWXx/tVOZ6bUQy46yeNkY0mMc0f0yRH52QOUF0MgMlD48uHQHuE8KFUL9Fwx+fe6zmpIhvFjUh9
BDAxrn0t3tpCGQ3754rauAqDl+zTT2k+9HF3eTCWQh8+IWzhYVBzrLWYJpnaAxXB/u+riXBclKtu
Et3+ZaT4qC/LL27rjGeKxwY4n7YV/cbjMqcwuAPdPEwLSshhWJ60FQAqYA001JfDdKdTsDEWf396
qB03uW/X20kCB9cSTjlRrHaZaoL6HY1NM8ckxRcExE+1IDf+kI9k++Df8H6cYlWsSR7Am7tvD4gV
MmDJ7I0+HSu79C9e6/feisvuUipeTnvCd5WNlUVlWPmNYISNtiwbafliNOOvzTdp45qEUwfMrq0t
xVvhyrGjeO+w27ihfTuWEUwtkfDTGonU62AJTy/DqwQe6C4sAukrKZVwqIFiBmU/5FdYoiWt62xv
42+rlXM27UxkAga4YDxSf72g++56r3gJ2KgBoPvFu9px0zApbBtgRmjV5UnwEqYVD1UUjZY5ph3/
acb1WUr5hrSHm2KTZc2pNe08d76STdunjsXmvFnbhrCbCvys0nDU8S9mbWACIX2J46nkf8/K3qJM
On4xCOtEgMmGdMlnuSa6gjblOO1Lgbbz5SqmAs3733HKtAvz1TtVAUu9Hxrvy6sT9iaHdvHf7Aoy
aNeGyGK3ag8PBeIhqD7X4NMuQOeuKUwprb2VfA43YauuhTT6rsRUNZG9Gp2QRe+Huqpte/o9B/bI
/cuRReDpxtnV4lZwjuu+zIsnbmLaAcGhnU0aQxNprigZfNpnCXOXHp2I8opk0keVNagibdAzs1BP
0zCIPPwwQS1th36IXx4nEuKkFUpLVPuPhnacZEWj9zFsp6k9w4NgsSuokCfYTFnsxnwZmPe3HM3h
vvDLE6+ur5yz/zO2saJ7AzdICOWbZc1P0lvdDNLkze7EPF57Sw5NJXFW/42rEnzBxdM3rVxjeDLu
/A5vq7W/TBTCXsloO30nHGI2mHEdaekHr6fLY+1dnSkPV267QiBm4FJT6djzPW5t4HpkBvYj2mVq
54sEHMzYqceRH4sTJqB8rag9Mqn8Gmd1BcUwLq5TsRfMbsq9bzNsRXx5fgkLx6eF+zbf+oB8t1Ws
6qJ3RD/3ejcXV2106fcRfwQ7+om+6efSWu90U1Ryy6Fdky//mWFm8V476e1xL+bcBAiB+stMF1l6
84ex7AYxmUq5mqiTUvo+XWxfNy2hRxOaBQuqEl/hzFfFkGFMgV/HJlsnEBOrPbENrExrhxxwf/aw
cgVXoZGY123HzCPqxUnKMwvnt9GcJoFgj0QmcMh1JyHxzHmVgiMci96iLa5hRq8LryOCIJUs3zIZ
7tAQNJcFPDXc31bW2zdhsD+hsmndxkrsu591YCFYOB3e/4n03lwAoDJY+i9bL4sBH6/R8jd5VAUF
8z+iQD87wRNCX/0pFF4vN49JOxPMvFv7l0TH+uV4cVPG077ynaA1fisl4etr0D0zIv1R4FCeUa8n
9Se9p9LbinR7koUBrswQ5U6RSr+oEnQFWbmaNeqeOb7MwHaf3OajQ37gv1ozBFOfLjqMzcXDgvfT
RaYr97hpL9yGRnyDe/GxaEXc094CwZr3CTyfZQQm5V/FnvH25/CzaulE3OdFplEKKDRkUzNYIoUz
i2oRMTds5+VMoXARuzBUFECQGxeKrDwX7AUouSPeUQOdFBUEt9ppz5JLlrU0c2K1Yjmov+Au/Ca4
byRfYYlGZkd5ezXUTmo9eAywqLW0ZRqD8p+bhDLmbufm+L19vc38KY3rCLjKZvBZIG3BrEwlT62W
W07jrBJC9oluE5cZetDgeoyIj+AxdJgbwps2S20EDNzvZJm7uXoZxwGuP2wHP+WlWqLRIy4eM7Ec
uVbc8hhC4WYudpIh++pqqeUWTM/siGHOU8kIcV3ay+FkG29q/5DkcX1hWILAXY5ZpUT/oSYo1AQk
Vdgzkys56gO72In3W5gVIWL9wX8n0CbbK5fU1n8w2oXHu/uP3pK/+hCiZdNGYKWD3+0W/URZ4nbe
+6vQd9NtA341zYNm0lOzrqmqqTOrB9D4Xq4KXmMkUn9xgm0uR17GGWC10MIKh7QmCSwbAE3y6iYQ
YpJeIUOS5lmVADgQPHwM0wqS353wL3cnM4NHMhk37QbvqXQtfF22Rl8IqvpxZmnnc94M28jA3V1Z
wYoQ0+QS8F91bgxcmzOC2Nw/KzexP5AnbLkARnomaO/9JQKaCOyGkY0ZNY2oiZsBL9jE0Ts6BI1d
fI05fSJi7IjpiY0Xt0PwXboTWPlnxwzOSkaacL4bFxpvd17G3eH0XUXguAg1jBcyHqsI3SYRmc54
zbiCJ63HGDSaWGoAJjkNKu6QvXglP20D9OVfekZskNS6wlIkLi28c613pmqoX9NLOWW+5OBTdfQB
Sf7jRMbNACEz3EVi4M1PFzfmvPGgasPGCFHGqn1DGsNYnQ+6kyi/oiGKhhECyEmtYAQDJocDDwPc
mEoWYld8+uTJ7aASGfDJfDgWM31j5aQnej7CKMx8r2qSTqSzzxWGzviq0+wqmbE6VjA/uOroIjzn
+4hPKD/W3LMrmJOA1ilXbcQ7C2DZGEg2j2YJbTXSgewTTPdlnOXGnbIAkFE9vPEWg7xizG16wScj
n2C7DKSBjmXvWi/IbtoGaikbEiD7s/8sShuZHxtevwmOWkVSaE70OYEPs5On/8tEl4Iv4DPvsnIQ
+/DPpuSwEXTwKizr1LTlwn036clE9grEq0gmgJ1hVFEHGHQgcOozG4Rop8BiUbcB1KN5J7tGwfz4
yyrk3kP4K3G1x/2P1YyeiH0qMdAowJRMj4CkKaoL6WsrO+ry/eC3GAxY8xS6ZTXuSR4tY3H5Zk8F
sQvIWPBxrvOOG0FiH+GOLgJN8E8OjUkghuv/0PxB4tIKzhvQeEb4PMPi9x21WoZZvYRmiI8UZu+8
iTKivfmkc0Y5HL/KcvF+xVMFu5KeUWSksq060pdmxgq/pxY4T1UakHxZ6RnFjPeuS0QErSjkgl5b
lmlnGW4rYvaZZeoNd4DbTrfS7aqTYO3eVIBtZYndlg9IUxhTMyhUadLuBYHqlV8Hz/wEiI6fYhKu
9sG8bsQiZdAd2bC3mEXoA3DANGdUk2r0XpcwolVoOIps2gWD0KjR6M2mY7deCnLfzMeDxFdIU+uW
/L4xATPkglV9UCfQE+LrlhKKq+tkCzN0PX/SnNPmKvhFLzqA4lBvtAnlTCri+FyLXkSmL8sDsIo8
ZGJ1ffct+BvIKony8g9WJEC+QVuLXkoP2uLUddE+TvPFaPckmPI+n8Em/c+A+zb0ECriSyuDpcVW
+gRVZQolBi1twhcAVChq+frwj6bOh72VH75NHEEA2Xdb1+LmqwZzp+A11OrJwqJMVofhCa7/8i2S
Bc6luJ6fLP2tisvUQGyUyC8qK202vLwbd+frV6Iu9YZBXKuK5Zuv2iLker1aqNq+hCrWb7UM1oQ+
8F1hv8TTBG9rEDyPkYNs/Vn15rwTrtZOUG8lyG5s0gOD41NN4c9FYUs82iMeeli+BN6KzAPgUZ5f
hpTJlXF7dmvCPAhYbVjLGUPRCoy45MgP6ehJRUZh0sFE+qM+DpdNxPWq95W4iJqAT1Re8O3Cbg/h
H6qfCAgYeQusq6LHaTY47NioPsdIUeQnGJGg+8IS/z51DDRZZ9/N187ti8BRTglH/y0ohm9w/I1g
4AUemhPf1jaNn9lSD05HI6h2p3Tfe+pAba3tJFXNg5avmUnV7tfdKnqwEjhHMBAyGn1APygKvxJW
FVHu957EVjZfibh7UauR9SqQPsA/qB41PZdx7HV+17DTXavv6QgoVCNlp6K7/m7usAY3ibH56enR
JbkahLoV/mLNENcJSYl00E888gzYaTDvkoCPGUuDkG6OKETLd1oK32qp3BxV0o/jrXQv6IANKxTp
HNKmNqFJZjUonlO+nMt9e02S4guA9RPHkwDPJrAkf4uR6ig2OIKND7KYjJ1thiUoENhO2Nu8jegu
e11GtkUKP3vJZwS0lv81dre+9qRo4GMOvaTBo/z6gGQB8PR8+3Tu/YTPT/2K0LSQbWN6JsK5sFBD
BeSMSR0v58DYJ5dKQlO5ECj4/AKjAkQlYVxYB6cUtMAOdBCsJ+jfMsYKJNHCfoDqag6R9Oj9PZko
1ARy09RpSZxaQGKoF6PgTVd7X78lLzQfrqJrXmM0XInnm+OkEkugUbdtJnUsQsYx4sn/elO870Xq
wcsud04x5nnMlvcMm0cDSogpP/T+Ng3iKYQDStcRrhIxRMzioGgy1gAeooe1rW9ubx/dtPguPuqU
21GTvIqZJI0AgGaMqUXVSTeuHUBo0JuNw3rJF/t49ktOGUzdhU6pWf5c/iQXqwBUL97CHBfFy2lQ
Ym82i32/LDNfeCiscbKTpNyqsKB6iWIxmh6XbIKTJplMJ8IccHv6zKJ7+fH2L+xH1jhbIJgFXsP3
a7Z698p1BC34ZEvwFYITch9bNIDX7Y9lq0Lpbq0TUw6obRlLBr5ffe1A7CPIAIF++a8egN/mcLFn
erHnbIMcFx7YXuFhn32nP4fzlKuTuimFB5oAPJndVIE4uTfhcxLXirqCZ0kpHebVkcdEy9fb7iSt
fzzK2+dbjzJxW88L6xUMQdEPWRFsQVrPi7dZLGQprmJ0d6c+LeKn0mzOhV7fy9xKXzA+HvlHVlu5
Z9mlS3CYET1W2lR1mWEi4RV/gy+Ui1QiqG8Lmfh3VL0XOGrJkBQKqYeYFItNkV/LclabAPgQYYTQ
F8J7q3WwlljeTWGRsKSNk5z7CGxu4gcni/Wt2D4eMur4zfjWaexIBrr1G6d1W4MvnB2kNfoNO5Pd
HrHsN4gIzdsTcY6MnUCLodArIO/UKoFI6XfX1VB9yblXjitBuOBRFlTJ5k6FcMNhBlkBYoKrTDg0
nLxlj+QBw3q1uA3aTVc8JKXWU/cDWvRG4BkuPsucy3Ye7c5KBLbc1DuILvY/IyBCp2wwahOEbYJ6
+gFZ9pF7+S41TnkMxmtw29EgP3WE83uD2dUS+xsQ/V3KDtJpD4RjyseZ2hLsOvGFA9rCOmYpW3wS
bt0nNTqQDF6Q35VVXyOI4Qw0qBlbNYrF9QfZ0XQDB9AIqKnAp4hRkKJhpBMm83eVI8dgvQ3WOsIs
XbVtoyT17BBETEit9L3Rh3prUL2jpdG4gaksjXtB+tRY10hrK8dALWkwO3RsKnsycr+JjZlTMJHK
oKhUbQfE6k7wDgalUFr5rchJQ0qqeWbUV8+QOmFmN3exC/tLYsro0T7XDyLmEDYRpH8rN35145fH
qt/TcJTE6sfAXyu/qY7TfVdSWS+9plREBX4Puedv2H8S+krL/8Vgal5h25o7EkVnUF9M2znW7NSG
70X/s2J4rhWCU1LeXhkhhQQxRbyO/K85B27xWg616EedV4DO/qg66ZN/MWBl3PS4ZA+vKifruUMG
kmSyApC+UGGlqmrPh367svNSp7mOqdocaNpuAhrwXbDIsvhzwfvYl2oBRDnrxIhy6BMFQ578I/SK
RfBzb9zi4RE6YQWTlGgRYoBLceeGNzLJ56OuTlU5F+fkgztAj3FZ1895AwHXoYITVGOFbr+V19+k
b5Sg2HVVwxO23lQ7K0GdCuAwWKyzek3XPbE0gQ1O96/3gX3Kr7dkieKyaw6+mC6Wezn3JfhIqSSV
iXip/0wLAzG0fBVPm1JLUkzZHlxgRBN1fkV/fb3EFsudm5E7USSv4k3qqBqIzeLpd/CLtXpzNnnb
tQlnv+bBT5Ge2P8FDaZQBJqd++gceNkFYRyHgnmCFs3bzAlk3R9UWUyLbf1ksWtB63Wi9sflweYm
NFI5SnCCP7uqaReRvsQ9Jwf48+NuXq6WiI6ZeK0bhmmzWJokaga8dGSuQaYB9ZsYC8PA4ZlpItEF
8birT5+siypDNUcogHlo0AdpTP16GJUT2ZzteAdZDlAAhQnmtMElmUF7A7wq4FqRLEbu2vM8dwsk
mHe3vNPMqgD+SNhU0DpUexwZhThjRzVXGAOz9OuizYJjveFV1AM/x3LMnhdVRjKWWirLdgoR/7vD
y//qY1OT2iIrAKUKE4a7/sG7ujwk/e0ll4bi7XOgrX/f0GCrEI3s/XVOLKXNC25ad4VMiq+Ddzk1
dsBO/h6hBJymYiqXvKjWaJbDXu4L2Jc88t2ZK3m7YBrLll0Yw5BZBmhpS72aoUrD24zhE5kYtIOO
h00/mYnipvzS6FoQ5lMqIUCQRZj7igzooTAA49BRRVwa//0bKX7QYJW1S1pKkwEv1FXKwH3yssj/
jwwk83eLs1vCZulcO9hMeT+pvBCE1ge4EXaKpJzUko6kfas6kpJTRHr7kDEDZXdkI67CY8QYVNVc
YKQJb6+9bp8XA6N5oRi7beyOmm4KUQknvvtVmKflKIoCZX5m9HA8OtaLIQgr7e2iSKMc78LJuR3/
mF4RlHSKiWtioA1EH1jT1CuobikAIx07sxpJNGuOoJZsIpzPB0/yMbyinckEbGf1PPBHhW3z3NqC
mlhOMxzGzLQ32lO22m6Wn5MZ5Thpmy67Ss0YTSValSlzcFWKWDNa8CPxsQ8zijDq4HNNf20bP03T
kl5QMv3r5l4rdKUMOgUHezT5I+KrdN2vDL6H7VF0+kD8zwwHOfA8HlGdguHS0YKaH+Zx7yz0zbYU
VaQK0XVBDJnj89BVec+/a7DLU5k2cvTQyujMFAxnvoOIpciyG6dm0Lu25p0veh/qxXZViHUHV0RR
3gOihDEVxEft//AnHEGmgwtZwHcskd+2EGBVqui0/8D7Z03Vj09G+b6ZpYUGsJcw1waVJqWVl8qT
no71Fj+N8v0SP6o30Ok7EnIjGTBGvZ9Zv9lczC8wiJsEx0Y1R0LOmk7+CUMzBBPXrLqTUwzuU6Aj
Re1JoHpVxLF8CfzZukPz4cbQc+aKTj4hEDcrU3M2OCtY0EvaoVgZjE7Fd7HSysDCKkVG3MVtiKvb
0Y7fkL1NsAGNVrAGsJBbIh79okx9AMhKL+q4wZXVB7UwJ9Toqd5tOLhI51Iy7u9dV48KegAkUPte
fPZUZTXvJajMd9qb5HdXiLnZMGF5Hy28+lJO+WRUXKH5zBCcj75ddrmRhRL/fXu4TpYZkjMVteFA
B64jHZl8mVpxEFXdV9TBTeMOxG5X9jozrzTcNOtrThlgPFTxRVpkm8YDqOBasdU72ug+T2A5nGBe
+7mtYn098ffmD2YG1LrwisswBPBThtmyqyFBMeHKYtjONfJJYz6k7jXjuPPdJ8+VV8mrh2pYSFbu
BWIlXaHnv3ie35EZ6uaEGoIIGwnL8S9gh1GuIwZePxbN63Eq9G3MOews43MCxKhTTBFkMKCngDyt
c4jFabBZ0SFH57l6w+iyy08S0C/aGkZLffh3VEnSu9OAgQYHyb6TFI11fTusC4jQjO6gDcMwUSV7
QeZSNuanGV26dTfilnigDA8nwvhFzrg9s4QW23JsS093nhnjR333F1ExZVJ8b5Zl4/GvWaCl5OHR
sV3KTRwRCXmAJE8ywFrBAvTmQcrtw3uh2IvNW/4Hd9AXvCNbfxBp1YmDusykg8hss42j/NHN2fTl
tgEHLU+0D6gOouBpZ9riy6HkqqouqO+e33JXkOE0CfpcDFtRm35oIb/d0Krk+RsGWzcHSVF8Qm9+
kk3M90lyc5T9WGVEp4AvkAMVfziNrmdaSbXlPrRSa4eAmQ3ZMShzUtMSHlYagOHoYyg6mO3D76Kg
KFrKo7lpVpPxQtbbHH31Xy5RsKyY5+rz+RnlzSzBtabgmLaMqSiwzP9y0kPYxz0nVT4zzVN/jarw
iZr4Rhp14etEddnCham7rpxYPO9fRT/GSIbnsB2WkRlunaqh3eDChb5xVkbnSCDE/0Df4KTlQVbo
Ypt/pl66H1jN/KI01D9H9plTHgzumVRWdOQbl0q0tCU/CJMmvpZ5CY3XpJj9AE5X1FlwK4aajIaQ
GP9/G7DPKp0GgQS7n3mpWE4X/1EdOwY2n6BTl6ViSVA2LB5jwHMiCWo+V6ck+94FyqN1fgI8b+NP
/qG+v7HxVX9n2YmMXQ411L3Z6S2w9KPw6Sr2ac9kpw0+qbJW68G53Lma/eeZWwnB3uGssFV6dQPV
B3l/s2ijku0yOsOM5VJITJfYv4yNkWarIhAIMsI+wQPOB4JGJCQhLkWgFS9wgD0GvrXBShHkAaml
luiZRHDDueGE0tBkfAmzuNfzncxo8bsCWdQzAeyFxVPTSh34L77gauqOET1ctGB0XHeAyQfsVbu0
OHQaF3ZMdVxwvC/dMUtGCGjJXhgP2Y0GNa+48fdk+CSjKlKGi/hHBmrR2XLQttHrUTOKV37IhMbk
9SNS1JksZaz9++0OhOyLCMTvz1N/tTFyvmbcO7QhYLkYi63f2n/OMFqfHwUvmA7eXD9ijTeY7bwQ
G7YEkAaVFdbhGO6LUQrTpH2gQF62Rn+gbcgogoO+M4d83qSO5XyGC/QNGby/OcJfZl0tlKHcRcC5
eVruAUyQ2IzdHVQtOmMivp+EuN4Y0/9utYbAMelhRd1MWnbRVOU9Bu4qyIOTm7OCBsJyS7gwqywJ
tfqP34RrNuP15oh5q8UTPuwqexf4ej+PophMzYUSQ9I9hn/xbfO78f6njoIUamr34YwW3fq+ZrZk
sAIEn3oQaDs/EF2sqYRQy+G+1jbfHp4dM7bPpUPwEBOhRUvTlK775ZxmGZJ/1hX1R14mUU7tFfOX
PdsqF5qpFvpyDWW6GwoPzdAXwmt2YFVhS4M57LoNn7xDYOOoSWTiPV4ce+WJicyCh9XfdWbxv6Fz
+V1e0HutjpImxgemgyz2vqmSgWEP+nR3zuEMgb2gXNEjj36S56Ij/+o2qPLkTKNCcic8nvqoNTUe
lga5fAMZqCfBZ5Evk5YaWmrk1F8ULp5WoOfz7ZcmlSf3ZgA4vu/rf8iSMkMJvCpD0ProTWO0dnHB
OEaUDE3Rn2hPnvxEsDSoud35oJ02+3CnpIlSV8K8wsA7lK1RKKBdNfnoUA+pMpRQWL7Hjft8IG1I
yEkBblL9l/J0X8J+JTgjCMafmfbkvH81Iqj9A4iCyadhDWZTBTr3ATwn0hHig0TCmTvEdGd1UyVm
bA6wrFwmIhumWUPp8GKXKkI0n4VbhQ1LjB2MOn2q8lYj4IY0agAFlL6hvL/2igXVMTx08L/8UntX
T9IOzh09qAyve4NC0p3gbR/Q503KJVyOkQG/bfgowstZpwYEeU/48HjD1hSTlWYmF77Pa8/y/5st
wf0d9CsCrUfGtxp5cJDKnuJ5aDuBLGVBPrdGzgQsBjFC4ehERuegdGVeLviaJeq16um2GiExq+8Y
NIrddl05JdTXgNlGSvXdyFt+3m84q1AqeicUUGaxUEa7MBGrOSa9qq3UfO7GQlU16weB3CqWtZYX
EzPdpbBjRGvgyk8km3ULhHzVrrRoVOURjfVHej6K/JFNAIHfsbg8bKcB5wIIEdE9j80VWnqPdeK1
2DNH15/zy+TyjQ3hkaOrGaSxznJJrjNmTr4n8vscUVxvD1XQz+c2XDtIPxw/94hLhiLdXsyLTkex
b6C6bTjW1BY5Y9gHupgp4Dn5KWpE1ZPSUOLM964lxWp9gZscEdLSas5XW04jGzoQsy4a7Q8SC7O+
Ik/urgCBUZJ+P0V3p3eZbyr+n0LgZK+mm0l5NQXcMdjLoWZqmqYvgvlUU96+VSL/e83ao5GKaGVM
ZQwVAkPBKAnfHSVfrA6mSLJKnqtrd9x2+/1pj33HO/MjON0v6248ZY3t9RPk8P4woRn8iqMqf8X9
55o15oizI2mbwXRhKCFgi/yopkJaCc6jf3md0kxh+q0r4KDVnWxDgQjVWk90WQRBLECW6IphbKFZ
UlsXh8X+9s05MKvxD0UVxmZ4G9sKq1pZ6PA0prB/SZnYXEwR82eCCMFabG0MCBUynHh8RBu1t9Hm
gnPqds7OlN5zpJBMV6xpvGcQA6IcqRxmuZpg6ANNvD0W3HYMVnYzc8O9eLZTrqqJEjBt2siFZkVu
T8KkF8f40U2ZK5z2ZKLW4j7+bjbnoaMM9DR488wp2F9dFIHhTIfA1+4rnLBohZWsp/ItQflx1ET1
eBE+42loRCmR+1chluFo8FTfFZv+vLAGE4UMmMaBhXzgAymAi5UcvlPJbHVPdOmrno5FCKNlnHaO
pLkvnXyymocFPgM68iLs3M91sId14JF0B7zrMN/gYck2D+IurqZFONo/eDfwZF3BYo8uwYgCsCXx
YeD3x/8rgWQdg+RQRrL++2iHWscYjVRIQiK5Dc222wWFsts3RjhjGipFckrB5rMLvsAZbZQp+dt7
T4u8iSYCUwWNpeExCMq5J25luFVkgZFWlIk7idGwNqa4Nuirhojp6rLsi3sVuAwXHGZFQw0b4scY
xTqniUc5dLRMAWGaK5628viW5aYNmP3Q9E53gc9Gslk6iB40rmdutmPRGfOTI+4IikbWnMvWx4Kk
BzgVpFs1STHaF2zZQX/HXPwj/AfS78W2nhAzqlJVAt8fOmnKvZL93sJMhhk5vp1cWfbg5huuWxrc
5+KxOxjAu8zOU2pEN0DgNkmNsRxtltWzTpu1DLFQfvyBHoAXbqHiN10q0w44DJRVnav1ZR/kiN/W
GDBYmeVfffrl/ncfkNZNQ9AH72lCfGM/BE7l/GNuonFDISJ/ZhZ9nL/HLviJy0d+qihdBHEJy5oQ
mJB2FqA4ZmnA+V1BkUu56306e6lLIqWxrn+xuOWgHoL3aubBdOAnpCLpV7DgbmQbW6s1Jc39zY/5
90cpvAWoDYI0KJ6HkQzdUf7QpgMhOGoCjaen0Oki1ZFpPVzLr/hF7aXAyrYe4eAFJps7Cu6QKGir
gQHccERjR49TJzbyJMzfQSCmUD96MmmXGyicjfvnmSyz2MPk3CwsfH81iWrNgWTOd7rKiRjN/NvX
FNZ52UpfDs1TdQ/BsPZHP9mfvXf3rOCGjAIL9AGGk1+WrWpUeeA8YRF9+VvndqmE9ziaubE+MEDk
k1USy2uaE4xcL3eV008FU860Dex+Rm10wp12fxTR4pF4WMBu0eYnO/9/bJ1BPhlOM6YBpYrWrfZm
7fj2eFGnLA6uZI7ZKr8Kb8gZHgegVudPL2LaEAxwF5YFjkRekhwOg/URuEj/b0Dw6ojVbeil1vEC
VTG2k7G1Iuywq752EQRie7ebcfEL12UUBC9jDkP6HDSufxSxeCDXW8VcvB/lyt7taIigDYa6Df3B
Xnb3furXAaXBif0FHIC3QsW0dBs8N5rbfJUwXvX5XbxFSdnmhWM23fZX2CetaAGV+2BKhv+/1Ofy
avWtWyNOS0olQpKu/1NHoA6+4M1JC7WUfpTmObS9sgaaK0Y+l13TJT3QIAA0fGZ7ytyF4OPWhqUe
w3b4pggQC1D/YAV+1kL6R15JgxtVV9JE6TfIrzm1Bb1Ju/vCl9eIA/BGtxdmwmY4hXlbKlQMrXwA
Qa2KPo0IXxx9tWFe44nA1L5UzM+hWDZd/n8jgmy+L+Q55hkKHECP8koOghMK59baPxxKFnv108Q7
1Tr4Qu39AzewCn0WMMGk4CdpR50ySWzamBqgw/cYc7S1Z/HihjHRzbgQNLAWVyD7ot9pt8mSMrJ8
q8h3zLxtfuPA84/2LiENJrw7EBWI3hD3go8dvSiUYStgnvOHArJYQl+HYsfwAX6AxL2HiSANx2NY
y0lB3q3NSNdWQ7NP+mKcSyjYigU/WlgIFjVxEc10iNy33xwPY/7hqIHXqkDZXtvBhr2dFVkp+vMK
E27kKCYylud3FM2HTNG/0MMG6eu8dOAzO4GCk+aOBCDQyVPcnwOcVodLGjZzdmkUzfhqGpH8I0Sg
un0GoenPFztj0E4IEZny4azCALfEfDaUshQt7ZnJZ1mfCjaPaq9jwaqcZpjQqEysz3Rk9G7wNFB+
R0iveYl9P/1NaQQPZshKKgcij/sCzWstkuTCTrmYjbXuosRHct2Sz8JjH4sMpAyfsKhc6ko2QjBV
2A1aSHT7BNBWroq/XcLr/XLUvyS9yvzrCiYVFNkveC2b/eDPOxXRfkhx+ypgpaFAjYBy+5Ip5kbc
1MwUmfAnHDFtD/YUdxk897SFLuO/MWWktu8VjFrOFnAKBDEBGpzzqdv5mFR6OrhqX8A4nvz0rYg5
wBD2P96fHr7OcMd7C9tf0vgUW9cr8DgCnKFv2eFXwfcMbKxOy3acQadOGt73MRtC4e0DkWW2OA9W
9V6wUMCvDQ/VpAb4QSfZf0Oc8UK+dA5nctXjroJWdvae8bCRQh+QLb4exjyyUwC/flOCaGSZ1Rpz
/Hs7IryJzwC7nxqjxpT2+amQGA7sZjwgCq/6kKaQ7ArOcHweuPMTqd/6mYcoi5aYK3CyDMaz6MZy
IKTxcimfdMNru3iJHda8oerXIDwE6edtdYrivm3QsuiL8kOk3a052J2HeSiMkqzE6Z3RmKKcaKC5
cialv/7b0IRkEvQuCltxCqtiQlsV4GZ7KKleK633nGJaRFKIti6BUJV0vUdJ4nJXRQKcjZVMpjxv
DmyM2bzQyjyvPg4HlKFt+U2HZGuig3pXgPAcn9mpTfwuWDHQ7cM/LXfDkcfdPIokb88hf2+20rkt
q7TL28deXZYNU7Y62vpow42nq62eHcrGP57DIoUT8O0D3BIBKhwAdkHMZMnBUVbXGCIAvEFeK2Bp
yCqk4sBYiy6ITIuIT42aENUpn3yIT6P2wKS16Ai6Gbpcvd9HXhoe8kTE8It8aj/5ke5bZqKNeXDp
RzPmujSArygae6wHW/lck90rDoaTykN2M5UKvfHaYkFQf5dSQJvz0/9ay8/yoxEgXIbwF/y56zDc
LuRxMNuVkWVQFEaFbYjSws3D1vdVYihIW6UEgEcF0u8kynEjq/fl3b1jnSsAH3su4qFDpozYiyji
ePSi+GoyHdcLgRR6RyPfyXy28pkvMCRdzMyVVZymu6JMW3RRdtpJ1j1B7vVaYexL8muAnvVVperw
t9zPsFQqePlXK0J4kqVfIanJ9XUA9jC5J5Voo6ASH2Kw+0nNKozQWR53ijl3NxVpirnkhaiL2BwQ
GvSmMM3eBaGiQHf6VClh1yBG4ScgDpo1mWRDhxvJNDjQWuD8jdc1PRPLfM8fiBI3Yo1HQwnwHvOi
scYIkmU7OIyCQoCSmgpALaNpJrNr4yRgWaU3cnmKcspROu86dTKIYyn+sfyDOSgzqXhetbK0D9JS
aKGH1SuT6rRjkubifgJ/r4SNjtKQeGhnZf1boJ4F5mwopcVWXst5hxnAyPIj2XmAnQhVe3ybJnpd
cc11nwrDOLUX08BpmMJuFv+SSX2To04eQI+zOmgnxTWulPQadSDbch2657uLgTt0GkbJ5YJnSTRm
Bb5jp0ly3n473Po3HlBUuLkuinhclysdMMqC//GglMLJy17vd8sAIa4316b/UlQSk7csrhSkhFK2
nijfHnGnxMWjv4XskFtl21LksKB95FbFyTQ/zhigXvtTE0DmQJ/+/+v9HAUnlVHafwREVtv5Flgf
MhP9yITtrlsFjNRs5h+HP/gTDctyae3SoqP/N/8bKe6gXHo4OzOOi7OYAX8zQLpZxqwU14RRHtja
kROnH+GrC8JEMrkcnKHs6U2HzdwsB9y+hd3MORRJCurDoZBGFUD8XFX3ZWBnPFIVtypewIOLIdrn
0yrCoHfq9pg+7jTVRI7yRntvNFbZxNdCXIXw8Yib36Rh9zds6LghNWJDMCOQNORIbT42Yb4TKn8U
PVAIY5bvCjw0Gmlm1nFBlZOQD5EvmSLhEQnfta0k5552EvPne6EMDD0cgt0nsKiNXE4snLkUBnEr
aq3Y5b3OJpQbFCkZsHyCal3paJjbkJZxlIK8+iwUgZqDzSmzq6PYUIsczz8H57aab3qUaE1PVlHp
7j6Ef5Dkvbutryw+38D87cGLj3XrXLOfKQQtT9mOgWa18fwRyKPZEe99ibgM0uhCFEGYWxeqojME
T4NFm2rBf77hazU0x5v8Z+4fvjLaS4873U/Bj6qF2p4bRamcYA8a2Z6ylfT2n0DoNRGyyCZCCPkY
ntDfMwB0tUsMuMqBDPykz37wSOm5qOfYjz5HqyUkJBx16WAKZASKImY+qhOlsLG7Rnour3Qsmnon
LkM63FjXbk3CmJqftTKgsJGa4bHs4rCKov3C3cUoJUt3moXsRyA0fXdbVT95IEyOdkKFMLTxAi/P
26nNtbLjtgc5rg8/DDOWkLCadn3L2c3quCDefMJBCd+H2vuXV30gc8Jdw7cLPrSyg7GkCHyRfyH9
PRGpNAsqWMlAw+1x5XIruRUezvY6XBN2HmvObemuZmOHBe31+ZGqteBI33tFbIMKRUP/5cxIxUlG
bWXAnHk6tl5h15dXr415Ilu+NYm+Hia/RGyAG/Ig9386pQA7ZFsaaB7U396EQe/BIvizRBYwdBY1
ahbbkZR+rXF1vJvimZ26TK+L0dwV7k3mgDTdsEf1iAZs3x4W/3Hm8D7S7y6PpKcoF9zQBGke5Eaq
edKSMSxzsobpjLvccgofTEm+VgXaBNT8mURh4dMaI80C99erOm8KnGLD5oeQeH8r3Y4J18nGCzZs
ZO07PEk58wiwmzRscbpbOr4jzF7y8OuhNjgVwBoK1DBTKwNrjSh/6LULjwoGoP/GskEz5plufm2E
k+N4X+OlZMceV7ja9bxP3R1TN8l3UNpLiMAwXZUvGwD2pu+zcxbCzkIVl5pJaeWRDvMCaQ4tpWHI
lzvBLNOSGsu8ZAnkjoGjQbKuXuV4QutoQnSfp/TwpNCkrsLemjX8kx9gl5G22YBjQ4cDAEAvfQl5
uME4N0x3U0vvmNyGSoLNiOAT1tfb7DAGuIN9x1V3YEORrk4gRbNBZeM8OvYncGXBzM7iEVML7iRq
MJX/SW009TsQXh0nqzQcPvQd2yy4dScLiz+i7mgxggPwJcTQBTx2Wq4SeNzhvqQiK3IuNYF4TeUB
oIH1C7VRQ1bt4xE8Lts8WI6tLM5XU+IwrGR75vKQDHG9d+TBpCo+mj5zBQj3Ttm4ZTRDpB+X7SQl
Wlas+8GuSKzYUUWAvhEUmoV/oW00NiEu5HFxAWEnHAt/PArJzh/VQL6Py3f0OIIMpIGMoXmZvEJP
V6weXCjP10lzIrbh47vL/b8SDjUzDge+aGV/7HH19MF3KvADNdbKJb3OssMqpdoyV61rZ8LSiJTn
LkzaY+gG4zsw6Y+EHVgaAkjINsi+UkSfzMhOj2kpYw58VXR0YAOPbaz0ch6buqqZ1mQlMYGiHaih
4B4bFZGeVKdn0r+6e81U4nxquZ+FI25g0w8xSnDlTzgaO8dmBnP7GqAdEGeR6L7nLVAv5O2kBOLi
TpgvNs1zgeCkmZaa7geyM+X27vXFf4Wf8dfStIpcRrAIQ4731kij+6/2zXahtUJ1eUh59Y6Q08ps
vbjaTeOXDcwlG8JxyEaX5//TdhEXCK9tnFGN0SPZnO4X7044I2VXh0THiUQach8MIAEmlQzWZsMQ
mZIVVj69ostlY8e5tdHv3wJVxf3lV+czQyIE/VO8JP8EjCHvqGJUF+4/6zkrrF0yNnwdxpfv6NGP
/OoTItCqknn27mnHgLbi4jWHE2bMwhqXmT47xttMbY1B+CgaMJyq6aXvh6tkBdy/URJAmlEyN6r5
8Lzt6TrnhMCoI70vUcDUN66VTY8NuPe3y3DbHfJlSIuhgNDGGNkqqeYSYNZBLZaO7wxlMIIDxv7N
CJ/RJy9kwLxWQpUx3eZGqioCzyzN67EE6LQINnThVt/S6hocyxAXvJxKEHNz4LkaIyUN+gOEQrgb
CZ3d8wYU0si08WdpH8G6NUcmRCho/mQf+G/3V8Fl9QmLqtg39Pzwl0HnyLshTxPdnEdIaqoUvs9a
lH+mOQSImDc43p6sFaw5tDjdIEU4JWFXOrDrI38ycC6RQ/jxGUCYDBxFPtCJCo4Y6UCo160/AHQ2
fDnfQC++fgx2vlF2+VQIhKEyPsaMzgFDKEHkMU8B2A2Y9Env5tePpjTcqokQ4Z5kclYHEfIpJXM0
PEAbzXx33g9knBVeNOAXpK7JYXBzq21e9EB7Gf3FsYRMnLKIogtJUOnxxpRcGyRtOsJuiWtpyakO
ilUYOWRjV+o02cdNFFdP4GnLtY+k/clw5QIP2pkYktNqqSZinDBS5Uy2bh8I6VlanGoB4zihOVND
bq5mp8jylQTZW5agjcbzQUWhepS9DdVdCQG8QrwKzctjeEFZB9FUfUniJBn5gGhu5XeVV7SdhinU
uWeMoBcoABzsShOw+D7a9xU3WsGNDPNcvCvP2Y9HlJHxigmP9pJOhmIT8mWPyK6lanYTe0gDxGZ1
lQOexudGQI/pQlwolK8VlNIo+W7B/dZbecwVOjbKASTna9nvVpeA82q4Bij30Ush+IIhAcXm54qA
8a0/flNw8GGOsmqlQKRo9aBaaXe+M/64N+DPTZaMKaRBhh66dk1MXe3X8aMYbZjOlDqNo/1BPPKb
zFwaNrm2v87dAUitWNY2gPgjOZJlp/RUnQJY1gNigpjLEH3/Bzqin9v0t3qB7GB/EMGXGz1T762g
uBFCsiNzPs3x+6X/0ActPqtsPhw/MttzkFcpXH/oRNUiZ5lRvgtSFyptFPts+ISUZKPXx2BdntpY
SrWKlGSvVF3PCXu4PSQqfHhsO07ir21rOkqFJmOw9ZOwlZBYODzGQS9Grq7f+lCnsGZm/HjZYvCb
sOkM4XW9eoWcJhDCtLt82SkgnhGLyV7bG9zfdZFK2xGFHeanLiKoE7gX/WiFoh9xfLhJAJwgrWND
UGmc5w/SJ7xM5RSgxZe+DJzM0zo2yv66Ydpkoniivyr0ARFFcLtZ8ZOXSpu9+I1Qldt6EddXg6Xu
7ZEPly8nurXZB7Gh6zBUhoI8s1odiKmbKBFyBPqtueOFFz0EmqEn6IqmmfoUJ9b+1w0J710pik40
quoG94E8hJCQb/ApRk/VXEyTBZiHuEQzd8v0LnhIx/rCaLf/Ob5Jx5E4nxJKLmdQ8mc/gb8aMsw3
QPRoCOjZz54bqza6psrPgmsz1jOxQuNEwvIDfxrbiQOoP9sechd4r12vLFSzAmynkRhb+EeDqnrj
ATfMVexhFvm0hbN4jjHNGUeWuk5Mo8Pci4VGsVgbtQ7zjmcIpqmCEepcFwD0JnqQky07EU5i3lVx
7Sp7XVR8SUAErAfsN1krotyH7vB3EwI66Az/9+KJNKCEAYHJOtc3bAnJDCNamSSIg1G3D2bCbhhf
q+tjs1b2Kb51BZuGiKlLfsPbArdfnlaL6eib7bYul29k4XNlLRjhGCZxkmirpkTZSvjWyyAX45PC
R2Sp0A77qsObEeRVWuZI0BL8YlYihEalNL6aMSOAM13vfYTdiZpNRg492D1Oaqlk7o4cRW+c6cRI
232Ob+DuzeWmgnBEm9hliRAeJrhtlsLqW6CNluT9VM9+hjt1Ykfyua3xjC/jn3wf7/CmxhVxEFXH
MGCqqSxkhzck0Jous6g6n7DUOYGKDa+CyLZf65rQEv1jdsuY7xhBthtq5yeD7djg/Th3zbdx0pUu
0CGXqJNY2GdVeg6k99iIgrTQ3DylW4YopCpaBssjKgiNWmCEqCxJMFbjn+PP7UmD5rzQjVL5OFTN
rVBYP7X/M5O97k+YoZ6MaTGQvTUAaKtKbNz9wqSbYNDCd38OrHe/er/LtViGlxQ2no27fRjc6G1J
HP+rIyzzG50fDPVR9YUlXyFB+m8bbpXoe2igwL/gtNTzgj+TZH2tVmBUWkRy+MVQdsx8YJ6T7ZoA
nGVQKC5KZHZCGwdsuMui/ugXjdrufB1qGsw0uQUdL694OFjf2k3+wWV6GuXGnEuSH37BcMdzVeyj
myHrAhF4uUtNl9Vyuiq8LtqfhOYtp5QQOqAE50NH9a8k/o8mSWiZX0xxogorCJG56iPO0nMrpDrk
OpdMtPG2/DWl9VWgZdKDUhb2yQ85kbNPa0ClhOB2nZhbWDNqTnxSksZDLKY5VP1KF1n2kQfvI7BM
J6y0berlk89HS2BTm69TMCoZIHBd/RtmV9ggyJ8laCo9Gp+KA6faHEI36rnHXoHmU+pw6nyJrWgT
hvjpIqn/CQ49KfGFIAo4XDAqvzIMIm+V6H2GR0pNGONRHbvacdJKNLhSdoHhfftEGHcE1qh10k0a
0PkxiqdgiD42mX3J9LgYm3BthwZw7tFbr8S4YMs9HUZ0q/L96LPxbdJO+anK0Ooq86E36rtWG1c8
hsd5QdKIj9FdrxxBgDR8rqDk35Sa1e0swn9A1ypsMJETNnQuQSmu6ekoR4+3ZGJM8NingU/NHgZb
AFn1V8CAgzy+LkL1VgR/WzwGf9YIrDsm0EtObFvGPyGEtR263IGH2wOVVS1DunGRSxs0foDaRcsN
QrriIsrp3/MFTlsM7dd0qhBiNfpxQ7PoliQZEc6KzMVUrxLVrLjO0x0wrb+oRUvSEXr7qBShVCPw
6tzlssALNLfWIOOoVylCFVx+MpvKCi86AbY0Egxr37bch+3Gf1pTDKnzD7z2v7Y4NJT78SY2EQEL
KT36r7JOq4wbVafp7x3m4Us1hJHMltpLtlmNZTvEl5KTOjr2lmXAd51TAQIV1sUfD/BL1MEga2fL
h4wBit2vDAB/5cD/hAbHXOE3qHrK13WUvLjBqtWq7GXdr8FF95AKhoi47qrlAa2yrvkhiCCOogof
yOkuJ/mcQRsUwlZznu9Zx+MqkxVgrXdkiBA0y4nkQZPlkYCycLkMyNZly0KqkLXmsJqC0Cy6Uu13
tBuQAOsraVqBWclTfVxEnlJ1/MX5hk8S/NPN86HGjoIdIidtucqqRdbWUGlYKS48Y99zpWlfpZGU
YWIMugqSac1Jsq/Li0b83Qo5QuW34dCKJoLdefo/gvebCHKuRiRurKUVe8+HKIMuTMnXNbBFlvSA
Bk6GdhLmr4rVvpzPX0mcQwbkVqafAxyWFvgneUOS+YJu5u+wycnbC8QApfuMWT0RETXPmOLzF1At
QASsmthpFisO/U8geQxv8nEW+kYOAiZNzrTwdA9FY0Snvg3dCrDipyzEVeyCU074zz7NXsiEZ+WQ
vwxe5Xe6SYwtc/p7KFVXmaXTTMQc89anYMfafYRjON7hbAOVwng8v+Uf5pTWbQmtgkyIXkahPHkZ
7GADHucGZfkdeswl6dtGyGRECqG3gz583Y0fn6Th0U8tTFk2JPcOU241xFoYDLqWrhVjDO0J8e0W
n820p/oVxAdYPuqjlyvJ556FL/g2U4MiIo2qQw3NtSoHbPtx85pX4oJmyUzdQr3fFlRXwtqbHhgI
X3cw915ZnbBJHSQiLcNRH+h9P8GD3ZGjlvq5phcYMTYE4+3eZ7pw30ckCuDDQA0X8rwxapRpXPk6
Y5iFcGJRM6D2dREbR7axYFg3M2TYgPbDVAX31hDqvZJQmrD3PeU8OIhYE1BdrqYgW2Ee2J/DOCl5
cUZGVav+k6vM5BswqoOeAAd82aDz49p9dJUp2eZHxs+byl00p8Ts+OkX8DfkB+v/3dMm9+kIkkYh
I+FiBMlgCCP1JRcE154AtiqRS7Bbjwmg7sZEMfFTVQ8wDQdIx/qElU1yV9HWHvzG+1JxG9K7WAvL
tSiBg3pV7C1ppQTlrCMZAVBaHmPwVLK0Pz+saNlAHvvHo+KODLwhrRE2mTvUFaOT4E0oflkB1wv+
cHuO2ZW4EOt+MFhNzxrt2oKzjr7S1y19k24ZbQ7pDnGEsIHD7GRYVviGJhftMEY9h4KmnLGLiggv
kSDNmXISzQP5+gGiGbAdDBgGnRxrbBMh57a5WQE8tBs2F2oDiL/c1EVlFgsIa/Q7oB6lwl4mQ1Z1
ESO8Op+cpeS+t0SnFTPQixCPtkgo0tfcZpPHCMJxw5cFLGJmU07fztMmgrWFNVrFXrpnsmnrk9aQ
0nGTVEEB1XHofD855554AIHruSDYtU7Vksucb5wbduY+GgqrUVa4/qSDo/7IezR/JR+H5OKlVxBI
lu0TmS8Xfb+E33J6skKiElD0a42Rgd84gQOJHj7mE6QhcHdHoKXFOpp9DiOv734us4gwvsGBS4OG
Cam7ZW+izkZWvpCDV1eq+hnVMeqG7M8dsBQyWYZXPw7zCTV0+WY9o/fL8Lt+2D9pD6DB4H84SaYN
qrXmG1GArW0fNz86G0PcFWTIfiwroiuaKBuWd2qBGYy/8q6S52ja6QLpO+oE8+L7a9iBQRQWgIo0
l5Bxp9zn56a8R7fF+5W9Ck8iI3zcZJl0lcIC6osQq0nsC7Ms/UPP+R5O0swmKNpjofIWwFit6p48
D43JS3Yn0LyBs1q+F89Wwyk9RIx4bc5QNFKQPWJ60WrfY1+hiGF5BOKjEbWenyp9wGLnOOCmDUMl
Hg4N2YWIxbVVk8ayZZDjJ+RxBWT2aRq1LVQ1/F/kBBa2ebURusUhvPwXc46iqAUFP+jzxehdX957
L54gSHzcSo2wCM8lOHeKG8mwvHGH2ydxXes2Xqbe7Oq/l0D/gjr5F+6poxelNSEBIofYGKsyS3bl
H0I/dhyLPpsYxzvxgbSI8q3V3cg4/kOavMSMifbm8qN+VDGoSQrwjAuz1sXM4z9l+i1z8cSNlbLU
4QQvsroMAALUvHPGu6hlQdYoDkJ+3BHE88o8Dvn2jjXWt+bUEgQUIjEAu6OZ9FXYSDXqyRYi/LnT
Oof1KW+epAFPtPN3f5go/f+95iK3PmZmVxj0IvZbuUP0JQZvAL6KMZsck08CJuRcTABXHknUwdWd
N7AYv8KlN4VR9lzZJVO2ViDa8ljuxShpZZ+7EmEupMhHrlhSiuKnjA9XJt3Stq8xgHDEsCUEhRm6
HcDdAnJbWcHGY3AN29U69jhHuI3ieuxK00om/lR3MZnTpXDW//k9MDe9OpMA7AkLBU2wPPwG2b+T
6unsHFS/hjQOYc9PHASLBFyfZzl0nQTogy7K8sMsEg5QdPk5VBpqIEO2Kg41ej6BVf2YX+j17RhM
RsCNgq18XCG08ri7d42IrtU6CNxvve5BXRRB7X6D03JBYdgYSzKBlO+nHInzXXMruWb7DeDlCF34
eNcHFfDe0AOqNjnamWY9rliAVrtEupvlGr51ZxjK9zODFn+iTzMNr9Lhj4VVODBHF1HvpiqJisXq
W7HZw7DmS6zFAJoGjKgt59DXqiEikFYGJFIf/L3eForo9eCCJEZjQqTJ4z8stjkcTaPj8c/8SV3o
Qj/qMU83deVXKpfrM90+mGl6QnjZS7YxKpO5t63a4wMpaIvtGGcPKY3IpGofImOxI73KT92xwRFm
TG5yJ+eyYVqa2Nh6XALGH08gC/xtbak2VUZnd3+Mg9Gcay/oqhdI3Xpy6NkVdqhF0yT8kIYp+O3s
Y898yx+6Vsu8EUGCj9lYGE4f0Dil2p3jZu0kcmODVj6HJ3kS2eA5O9MIe0LoWqNMTTbRzxq0/3DZ
WoJMrr4lHKQrHMiZX6ExQInxbDUjlpoIFQ4J/HkcKK0s/hrLpxjKkPDx/pwUH+xwhb6bQdHisePW
UatuUEyySht6JHhnA8d5ijFcAR47RUN1JNWlOGzb27Zb9ygmDaSkaxxz0BpmpbDerxVwrvwDiCI8
6m53K42rVyqCm0dfMeP/RfyDJzpI/Tjzy8gKN42h9ZWufLp2uhLvgNYb2oljfshXHrSZxKN0S1NG
cnrGpGT6gF4Fi2kPi919ZJxQe/5Q3SIDMhCav9pnll4bWns7LZDFO8snyzlgHCG/tXy5yrMD0QqY
w2gNRTzW06WwBHLoqR7n0TV5qjzUxmIClzTUccKeJ9cI/QiDhFlQny3kfN2yexZQ+cf8NvgwNIMi
hp6v4XJ3IRFehT23x7EIZiFAOHXG0eBWd2fwk8fd5rYSlL21X7zNoAWv/QUh9EFrDMmUEEr+WrF7
kbIj7YoieYPdDikHa/tfBjjvZE7pXNnojjhYGOo6LFIMBSO7MBVVb7g9AmCaZ8wE1mFp1IJ8cl4M
PprTYG7lMrst5R4Ei9lK5g1LFoTch5mxLI9ZYhDGE2lFs8VgQmia663ZD4KLUm+d0H0PN18VhoOn
lCjVtJuEcQdtiMEPFnwV31DJl2eltFrGwm8YgM4SJirjUTnZ6ZW2iWHX+LC0Pr6NVq8zj1Byc3HL
VomKepsqIlblc6PA8dKg+iLn5wTSeP/qtA7lz2BAKEEejohF7CVjIC054zyKEg+0TO4fg5nJaJOR
nLYRV0Liih6x+A3JEmRdANXIK7/3eXWRWsMvQffVyJJKEWFF8P2D23N8pILTIWeRhs+D1m3xlM6k
f5IEY2WN6a+zjmpBj9g/otVLCZjVSjPRR0dzZvWmnUsGjqky6pvPOjq/5zlPhg0G4xO2rQEe4kaj
BI1R3JN4Jt/b8PZ35X1Np+1vlHBsMtaefjr2qKAWhmqCZehJT4xEXhcHCjSprhylNMYBi27vG4DJ
uNQ4cRfylQTlxwlf0GI+R2yIL1lk7cSO08xmpBUCrXPBmPX/FY4lqR4lAJH5i+Los5AWAQ4Umvq+
53M34nebQjNMVxD2Trz6EsCvDWDJsDIhXxrUYLZ26qeuwQq3EginiK47yQJlLHMZPf+Avsyyv0mS
UqThL6ClLUyVpYZZDDUHEuiC2A+ayHFcoI8lXrjTRQm/VVjUuvrHpxcLjN6CpAKHASaUwIQj8uCj
YfaWNKxsVox+jf+9A0Srpt6XAeyBuEx2N3ttrGIJW8LIjs/8JrCEEqzfdS40VqRLdZ1NUx90RE1n
Lm6oGLNfYd8kTsyoPnZPffP1A153PwJrgiR1EAqcqk55ZlB5W2Sd3zpCAhbWK4UEsSBkN0gSo+o9
YzjPTNQHAV6Fk9JMpcMuVpkXR9+1kB4gNJNg6J8aj4gqNQuR8Rc/v5G75EWSYzMk4MM7wrDObaHl
c5yha6IPATc2uG3nyah7VgHISTGfz7RxdpoAupg1GLSDDuyjC+AVUjy/N8EyKryZ3Q3vuZxQwQjT
dz3LhU1oDUd+vfmHMN4m7iC/HZeye0S2T9YsnSO7cmoIGpOmhdqgoIqkliCivn4f0QklM9xg01/R
iPG5eaemeSxl8nJe3vJLk14sgw6FRw5hKH8rLkNAFH2JXv55UzjWA09rZIQXn8enkKYXy4cdV6em
giaXLvoKgBr/Sanw0Ajl1LzKoNqBPTMx2qm1W96WdMzNT+ALwoAzTzcQOxV0Ja1mRP/OF35Sw5d8
Sz1TtXOWld4uGjhJbgXFymayl0lCyOs2A3PsISNVcvrWpfD5+vh5cWNm4H+n9gCSSj2AcvGSrPS0
vwJFq6JNfEr4s/kFXGWUNqLnubiiszWOBcoMMd2OTU2wy+AcY7j8F2bQjb701Y4CmyYIFaus6y5X
RK0gpzphp4mnyT4pzvWYf8jIXNbnFTXsFq2KjtqPY6k/RFnTOFh6CYhDc2gNo/4J7I6DUZ1eYEK7
wdzjzSIkqTWFfGTftERnDvyb0tHfiT1drOChu+UqPh7wqqIklHaDOhXLmnBinHHsXGQd0kRZ/7oF
Z2LY9DGfuFmiwaErH3odMbs00Q4p/KgYRuVlc6iJYBdXnViD61fNMv14TC1/dAMlO5VDl35vUr1u
yXb4qM2UG+VBA9wcogOep4XXmwF9E1zrXa6Sc1qjF2GHkhWN25dxTpFze9SJ04oDg/HmzqYH/LB7
w+XshIMCZ4WXwjb4+usdopxyd4dXx1oKsqRH3wEXnqaGlFDMTk+xt17ppncMAwit02RgY4vnr1ei
NTHbK2m8kHLAr/YKPO+5O6qO8mOTyZnKx37onHlxwXG8OMruss6JUDDf8NY4xjxYOr9YHckRynCv
Ns8j/rxB+aZlwEIbJNFjcInfSLL2v8eg00Y3ZOlB5YoDkI9jzJ87j1ZZiuWMVDlTHWvvNBwu4Gaj
iCi6EiMQBajHl/6CZM54VFTiyzlSB/0lJF+2f2rzxUVVgtMK2ZNQgebnrx+aKsGITv1x/b5iS5kl
NCnaU+Wr87mNvzJ4BJhInmBmedBrrBe2dbb1Tw00uwl9U/vcnWsTELDKKafGtzqQ2/Gr9orUVPN3
q5AskCevDoGeZl5e1W2+HwXuUUfmWQHaGead69G7bUZUUrXoMopyp/rbM2acmBght7svh1r0UfnW
J8GFbOIel3vJfqcemRgKuC4DdD4Mebxmo00ofdoBQllgFO8QXlwu2hc7hDBDLojfSo2a8PnCf1zk
ePcH9O8uBDBadVaxo+pjVukQUbTvJtBkwE7LGCVVEQRo7JwZtsUxLBCwqU9PrjI4RV+rpLpruVtF
V/TIUNb8DWQ0KKWSQ/ThAQQpf3ahcqam4vJtpNrRrFlQGeblh3GU0gIn3cBiCiEZP+N/qKkZ4EfI
R0lP9gvA7t1J2e+ZHmRCtg3FV2KzpEHe3TnGuNr7adWyJc6EtHET8U9BKNQQE0QNI+3BTzCFBnyi
TZS0RKG77hmD2nSvSB+N+BOPrjIgoAdqYd3vlDfLR0MY2jGT/RPHNwqfoeEIQlbTOtqt8E2NplMr
+e2fSxgCVl2/nXgDFPeGNOgGpL12a/hmIcSbokRh2YKj+i63c4u9s4C7gOPG0FZFx2NwImQyTGva
j5DJ/g6avUp79Uw298ciK1xtpZGHCkxHykYEd80sBhFr/T1BVJdzQ9/YTSuRBXDXB8Pk1mcpeVM8
Hr+ZNY2eFmj34hPFDb5mogDKHKuREd3SvonXMUxlWZOyqVGxv/9pxD0iX6bBeZXRuOHk4V+mR1vZ
vifqdBv8stAVbqziUyMCoj34awo/9CAVRSkH966LHqSheRVC0IlIu/bILFNNjsk3dSffFZwlY0Ef
wP6IcQhLBlqPfb6/AYrgsZQ6tpPoNSothXzHwqlie9hJxV6Rb8J36ku4mqI3NzjlREPAJ56/NIm8
DsPP7h26qHKuws226DDEA5AvcnlbgU8wzOMwGzXspc+z1rJ+nQi7xNEmNzBG5LLrqgPaR43QIQOS
808QpDXFvJ5zznSqPZPCh+/282s+e5C+umhw0/MLOmrtQ/AVn4Clgj65HIQPSZd/gm1m37S90cnk
mNN/2k1HBNj5lYBzbd2oKjt17Y8N6vAiC6FSKw9R69aqez73OQ/seOHvn7k4W7at4T0mSw51gqRb
AeFOHkK1KU5qW89fWfvK5/gWVZED6f2ISg1s4DRNzQ/6NnkDKCW6BnOxUfIWkxUcCq0SnmKmU1zA
oaHWItfpJhIGB8jR4BS1QuLyEUqWNtr2hauZC7upDViwUD+pnGb8RfVZhOb8VRY29uOWKRXdyZKi
V+xOC9SKMAe3VznHKWSSpYiB2erXAGO296mF1mI1QrfwrUgqqDnlLEuuPicqq92dtWagUDahv/Ca
KcOjoB4LxCY1EI+EQ0GcGmKGhRCQ2fElTw5fkZTHcBQ0uIkGQujHZ5mUBkQSJ0UsF3BtrNwH6hM0
Blw94tkztLK/zOLrQvA3t5mbGEHGLe6QdGhEo4u1qPnIX4ltBsXgf0SNSq01F0iuO81LKnz86eHL
S283P/FtrOcfbhqCb4jZWIGUfr9hv1DwHiVygyVx4cpmsM/56XEoQnEhUoTul2Z8iW7/O9D3NMXQ
KU3G/xBgSfTuEiuNMBg7DmEIpdE/qnyQiwbSr9+TGadfkgXg1jTZpzneZMt1hz8TeQMi1xXwe6pv
6rekgI9CrDrs4dJithS332dkfB4LM6IvA9F0rBQ8EJWztHnRbbTv7iF7d/JEl2EszvN1eSGc4Fcv
/c+7BXOYuFSisF+d7pFTgwImTMIanc1m/UQhJwFsQxZ1drCtBCyOze8zyPRz4iIZiLksOEqGhDjr
2M9s2JEal6oYhBcR2WI125HhaNOw5JcnGn5HM2zsH7qVD2oDIhmsZnTNogHda6wDn+IASfYFyFNU
Bl2vKjbIO/X8IR5mfNyiGD5cIT4gHXjTGOfzJxSY7csxcN0vOtYRqed6GBleDuWsQiZwlB99Na3P
6SSZp593ESw6ERd3R7srsPPGr+QqguPYRefFK5vfiNIAoTIFrk1AIxPUa7k2JTIXGnJjDfeoZP+Z
JYqKvpp+6q3X4/tyKKxc6YGU/wy8sluxNcWfdWSj5e049bR2dzJ31LqsR8xKiY9Mn7Jf3BkEEjaC
2Rz4zN8iw7NecftSBUIZud/7uPvLb/KOffGlz7F/3ATuikrgqc1TXV+vry6GOEIkmon+ddMErgh4
fjJTLj+v441GGw2mUXlkjvuGjLtuEQUiRM3z/W9jr7WKu3xqR1otm/YZrd55d9yLaNl1BXhnkJqw
Mi6xsp87wwP8Yw4nctN6cVdbCYtL40qOewnXnQ+OB+21U28Kj1//3jImOEociWBCjKwiDSF+eEVw
ooWegWn6moQVEDygmd/Y3ye/34wulVk6N1Wii/1U4QK5wrRXvo65MHiVExAb5c6ajnH1aP81IDgU
p1vSskENB+yCClDw47BBnwZbWlYiumxi3wMcMLcNHvjl0kKyo3/OFSb5hoxvhQ94gMhbmtKrInjJ
wYRIVVMMkjVE4NQRMlqR0cQ38jcOgxnCmZ/WMaRPEF1nAqQ2996yVfjiA2uwuPNbtJa1DK7MrB1v
XAvNEt0stSQyj+ShogmpP21QNdMMShkX7FIbINnSIjxTk2Vz0KId3nC1F7KkC1XYi3rorLeQckiZ
39dth25weyEUV7VDoZMynPUXjUXPl1/VTqk212OB+kH+Zni2xqjRwC//mUgt0FDwHzSrXwWij/qo
wS2i+4ThwfguKbBdqxSd0f+Q3DHgLkojjpvM2qWNrjtiUpDdWYfKbVuga8rxYnVVr+6X4QL2XLpw
fsvS3UtbMipXDwnUh+6uSvmStV03I+Lqv8UmC3ORd5A48ZQkeu4TNSOnav69gxmSN8U4f/TFU7Pe
QmaUDDUIZoTdgTT/nqSZKR55Le+fIGsEnL82N3grqfC6MD2XWTiyPRZw6n50/2dBMYjCQsA+RSF3
tr4ZfSUh330m/Xa1J4sFMfl7/+UEnmK7meYdjqh71wBY74s26svTbaPRMD8/JaiMgn2ueVSmcYkN
qnBMLpeRd3Os2W+M2MAKCtlosQEsdIpG8g80IR8oUGWkaktBY37tBYbRWX1jtf6BGQb2h1+mSRle
824iLO+dSs/TtcoyQK2DqVWPRDrIpEB7fbn42msViDY8H9EeAN1LItH5MYpD9N5z/n7oFZefap7Y
4ArOeQbpZcxhQTFpoUwL+xJMjOwRubTfXegqKxY2yOnVuUyktHTU9l9aNEZVilpvddv6BW3UQNUN
0n5LTkJVHzbNLmbwyzlDVKP/SJBkC7T4ja5r296C3fPrArI6bDcGlgKk/cypi4Vi7SJa3dmcdEcF
Bo0N6s1Kjhpox1Ru0zljxbz5GKqn39DtpkDlQyEChL6Iy/B2TuHqO7ujjOnutIT4zmgM/TxfeR1k
nU96DoxuKUF23V+rheD+EgHhzxuy4O0MrhhkF5jUaphkls5hgBFpjWprfymVoxsp/Ra0oJGx1VmG
9FnvuI82szfu8jnvGWhy3q4OGueGiTENNtxjxsNEhZ+2CZobOycJHppcXZKXQBZfQQ8+WkzmYDMn
zKBx5Jhcy1bRLtMh9kcJgktpuXLGXIHQjlnZtI54DIviLByr2kH2B2g29SY8NkPwYpyTzflmcygG
r3aBvkAQMBvkJoQ3HwqI7gQUU/aK9IGLLfokGy3kFmiHKfRf3fWZwupTHzvVsVJvHwA82erwa+nZ
6RtxfaiFTTITU0V/tgpsoIuU7QdOnJ7bzyR4cKaX+j3qqYoXIhguaiIseS3A7Z9oKl+JUg5YTc24
oQDVfoE17zLEzC4EwsJhd9Fe7sRNF7s0qDD++y5oq7OkhJb1ZXrUj7JgNvq5lY1RE09hjUOXw4HO
pTJoX6+KKrNh1y40ebrkF3GEnbsPVd7f4voxkdHVmWZsrul8IpIv7JM0s9OHPLFOQ+gGpwIn8tYA
ZQulcfOvhmPlpmohxgKV3LoWbnWSBRkye2WRWVbcpVnAvwGLByhr/eKeD9j+mgf45RtzYhyCoKWE
8dROiikB62cshCQGE4ThxEIxpnWHaFjuyIVKInU5m3YIAcSwKSjxSGrPkSgJDI2dLLCSFlIy5O3R
qK5zu3OungLJgSs6rK2o5c6XtctVCs1wfhEOCl8YJL9S+W+iUnYeIhwo1jna8ddwfnci7mrOstfd
K/x7UfJ0sBKhOQCzZcQ6pSDIA7egtYb4VdJ2ynlbWsD3WsY+GvPlLDviqgCk6S3B1IF6ndHrBLKt
/BVfc6IGIR3gb5vAhU12+D4+9cvxkz1i45BhvJNBcVbl8HxPXDz/vNL9dXyKIpuu21n/t6eUI8sM
cC92pQ/KTQVt5hUeQVFWYWe3wz6Pk9Cf2IV6+YWCQMYA3YTsN98BREofoL685Aa1ORazKQb69pW3
OrWwsve7XDve2AA/x4ZztkddUBTfMp0SdqoZYMRcZX9WdUyBZbfc2LSaCKjzVd6RDsmyHIbgkFFa
OdWThKi40ODUvVvtJn2czs0Ls8stZXHbGv7kzJb3b00YPCWTaY5mOsHq3ZtcjcUnbW2rOGhG9kvp
j4Kmun9c6MsdMIIrQfbv5RrxZ7wZZ7Ljrq9COieAJ1kj64/zTTNREvF2Wq5FjTb8Sa0Wki5f2G7a
7H4rwBCe5czwdIpHY4CiG9iiD8HTi/kAXPo+w/ybILLDdq6Ch/j3R0oVouRbG60Grcl3v+dg8cKM
jCWsgRA0Btl7sU6NdXlhyADT0UIMfMh60p3tSIeBeQMsvpWlIUTH2hrGmU8OYqAncNXVQ8YBjEbk
VmkGGpFMCnf0FlnyBw1JWCW25RDg+qUMYzv35XQj95Fb0wZRbmPLXxps3/Zij4tkzNMPfKx74YQo
9lPGBSJ2Dl8OUYquoaClBiGeo1yG+OecG+Kw2zyKEMjGIKjd5xg92yyvaPJw94hcSuGBcTfuLJZk
aq8uHskJszf2lPIRNfMapvL6CeINvZNn3H89rgF74LnPWoWdMuiZX/rXXRv8VK8ECElj+FhOqVUJ
RpyNb4W0iM7iDZw54wUnSLJ5xLtO4UmzbBDgP7jqStOtUSq/eYrzHNW6WceL3g21aGR6jvUdMW97
xh2Wu8UNdmbpOKYhuWFI+oW7JAFpPG+bPya+y37dycTD/naki6w9v18BCot4PvoGBSy/S8F8/KYA
ydOAaH3rjF2fYqAWFksvvVaw6PcAnaMFrl08CKVKIEoYCp9h7B1oXOCinAlBt3fZFrPL33IVC6yc
hVnJgLeG+4Cu6t1Bq9H9wDN+lN02yHUzGnIY84DZf6UfjNSTvlvL42PS6N+GDW0SIN3Ge1mcgxbo
zNkIji/7/IT2tn7nL9rVyZFUmkO+YRON5vhEqzJO9C72WrKCQW837VBFiRvFBA5xippKn2ikpmnP
sdLGOAWEsus909R86BiU0GrrexfY4Nb4ZVfw8rbxidqi2kYsnQMEWFpP9o1ATxNnubvBctGqMnmB
AauoXa9GOIJRrcfevxKfmnUcYaWpi4nJIPeAPiCg+RD5XgkheQ8CSkAwOWsl8exa1hTBaXegcJcg
eRIevdIbCUzSTPqL5VVsGV898suyvf0KF2xpq/rL51wH4QhqU+gzy6dvI7Bv4I+ox93sMRa3kKll
kbS6wa1DnwiKubCq4H+gHu4/Ip61Dt4Gf8iRXGUvyFVQ3USzfTTlUxQ4vLGYnuAS6QC9IaXnD8Eb
bPC/uVyE8Or8uHeWI3Te371KdxI5ZSEawlA7je0lSWAO9rzekE/49WAp/5ICSDTdyacSqWy2igtm
eHCURObXpL7+9vOOPfxns9kNTNDc8noa27zdE6YqH2rFmCrNQtuUfSXP/BWn0qBAbzI//unGQa7M
WRcd+1vin0S4dq28HdmfSnZiOuN9Jhbiep5Fxy9htcjgikNDC5ee+esPh5LCmddeZ48fKK6z2lNM
1Q4mSL4NYuUuJA4emw4zw1zTaSp5Yy1j57SEw9unyRZdO6omVjtT5hFziyNWg9PFTjJnV4hFqdkc
Qf6bwTB7HDcaHU9gmOn/bT7HR90g0BHQFgVwlBQairy891xELeoYPuQuTjpFpQ7bjWGaSKs7HmSs
mK8dCliLWSqCrRh7PIDuTGFYOOPW9KSR1irgwJVcX4+N8PgG93YolvCj6A9ZpVbTg0emH6zYYyLv
INa3FNZIvpo/sJVo7vaXcPXQln4End5Ke0n6247dz2ZSjsly961OuiA/Z8EzSGJD8/YabLvFurdA
f/b6pIEkOpccLvxidQC8xHQlqQRmUzXGcILtbobgzgvgcRQc79h/Gq26vLtNgE0VyjyWUo2UmeI8
muRaHj//ja6Pqz88dah6XJocDE2DFFsOQkpTAAwYCQjh0LCS7STStEKj1k0Peo6ENdwWIhi9AGa4
UT/Uy14eIYpCMO58siHB7UcxoI/PwSMeKmsC7Btvd0Cq71Rw6XXFjlJNB/MNQpOwYpKCJ5qgydUD
7sKUuuksBnNNTI63v0YIfUbukRxL6W4GPBbuxf1q4DUgBbUJ12tlbXL/EeSO/VNsUxaXU2vCMXRH
E5pGo13KKNdvDLeqUeyFCmvv3mzHqq219JiE3i3n9tJyVyJSnQlNcr4IC1Vgm9JyPSsX5b0EDjQw
ybne8W678vYeuT1Lmzwv+tzpKxmH5LkaOKolDuLC6xB+pfhLfDYmsz1Y/TKJX1r9C/lxMCLybFeF
zoisZ1+NFjLFXPNKdNQGTMjM7mtwhvWhQ27yTzlVsZfjyEIjHCLsSMMOtZ8UOmVUnLX6Zk+VF5Rd
zUtyHuoM+7cdw2WmHc9/W17oX8396xxXx/B7fcIXbFHl+u80htbyArmYEu+W6IWNtle3waQ0mtwy
8MGtRbXaOEOVH6ZKYcihVYgd65mxivGT/6QTBHC1UnSXApiuLjwcy7X4/tFqsRhhv9BArUfyJd1+
gpdCUmW/bqbySGmVfVlj7NSlmk0PQ2ZRvLJX6x9IifDljD5tiY8anNDDdtE2mXSGPQBjA8gKb3fR
yFWf5HnJ7FSdyYe7NM93ZgrCqqhEBGC4ZSsxCmHqv4Gm/Z5f0Pe8aMW07Mflq9JLLkPLgtPARdyi
TGB2li2Wy6XTm0pR7ztlY2eZ1fqSIHpSZzATQcSMlVYWXGklX84tlFzEjJCEWlAu6pEJ3uIPER4j
TKYacTM5+gA5JrvdtOjnO+L/klnUPx5Db0jqyJEqZ3JPt6IHuYJ/d9I7YhMleM4bRSd/Gx9oAfSr
bZ6KVzYMNJyf9KGbk4+JfbY4T/S4P13EF7tTvn+KJNfT5DtZ8Czy8X8Szx+V8BF0TF+XoccBnZsY
0/0rdMfiD+uwGqQYu/B0C3XpA4frnDjhHYhgfKq7D3ILTZE+7DInCUWtI1tuP8LXVvHrDGGdPvv1
e8DxdE6AE/QkGUGbjGHqdJU/R60RcI9IMewrnmj7SsML6ofM6u93Qu2+Nvzsu43Zrp/YIkBmfMyV
n+SaQsSFRMGxMabNLjRagoIqENH6PmEAHBbGwhNEDlnGzY8yMfSZ4yT9Sm12CaEbwo0O7SyAjHec
jPuzqocjYBCU5XP0x833bbx4vCXtQhRbgnGUTL0f0XxUTXZsmjakWiZjqgUfxhk46rsFMYZVzjRA
vqgntz/0xz6txWTCtxU9oN0Xg6vnaNCqqdH3Y5lSFXEbWHg3yNKKfFbSU0hFRLwfmvvv88TLY0Z0
ysBlgHyPms8Ac0IfW70osItlKajG0MbMt3EWN40H/XTRDG8sOikEpxG0vhUgduoOpW1XPyCKoqJP
9LREo/gi1MgvksEFT79jseDYwt2fcb7APCgrXivLeUGlQCSIGk0A7ZeBepbS9JyeW3+fgz6zqE3C
fajTqQ/ByeBGIT/GpxNyRJirhEXKekoDyw1DrwipWJJKak5SnKcweilBL+QYkdmlD4njcmia+oRl
1mt8bEOKvm9hOokneutPiVJMFwEPxvfAofskdnV+GLWnwhIfb0MrMuSMoLEvILjERpQjpv0j+uto
gl75gWa6MjUZzKGEkWOjzfqg9BjXl6rmqQtlxf12snQgJ66kSl1M31z1MEMr+aFR+nmslGKx2UEm
tH+aFPQgtzEkMuWVs72bWJI+fzc00oS88h5Z6dBqgVNYEQJl6/rhgxyo4lrPwZEUVIyl7AUNmiLd
+xvoDaC3bzOKb2FTcJvwpx4efgYEzJoQLAQdIB9B1DM3Id0joBS7L+KFcbdhIKizQWV/T6uGPHHS
YxY15m71Jz7PxvlZUITWGiEyHyU1biQARL5kff4i9GbpxHuhZorL0lSnrRBk7Z8N5vfV52o2WrxQ
R/tTOTb0nisuCAQW+uj7+gWo5WRcT1/2nZAOaWK3ULPDubc8NDtn/3AOvskIj2eyBE28T9xMvucC
n5aovODtu6XbIcLqMWeH0naVJblmINvL2ZaQyVcMPiTVQRPKH84jf2vxXvqNNrz2sTxd6i/+J2WX
OaC8M8UztYnTcET74ouMe4Uer5D7ssf/82oG9yhMi/QS8c283bLiYeczjIqz8/U2U1apImEGjWEm
wbbzVL3ycV/1/hdzG+8OmaR0ovTZ8nubFyyZnrp3fWnteB7fKf7A/zdhRvoBovxPtb61zOPZDu2B
iB4wxweQHc9wam1iTo3fW5H/IWNV9gLAhUS4C678to7DX4ASsp4S5VWRvPVl+8cHRH8JSLjpTzlo
GneOdPN4xgH6Y9YAl/NutODVhoIkoUM6lVxfUzXhWdRRIWkDcJ50X0Hx53zhQiTpktFyzxZ/S3F7
lr8+H6Gw0ZqC5LYgukN8hmpfVspiHMCUBqhzFcmwbrfSEKsXLgqLaDxFxxP74nIcDrK2O5boTx2v
LavnmoB7J+KkcksnQKt7VAM3M4mRY3DxMxahGhQs0YjRMf5IKSh30JrMDbKWNTjn8BMaf8lUOVvf
PQhTFVtBYskkdptgbo4t85s/jYNWq0QjN/648OLymzjnmAJLs4ZClz71Og7PTm4fg3i6v3aJ2M2z
IE7Ym41qmr5wfGYO/SfD4jazIo0bPkQnFg3ADDplPtxsmnb/ItbGNn5ZyPNZLy7/R17AhrBkyk7q
ehYao9kaw6pKtFsGseXsKYW6sUY5/CllC//dJrH/pzhg3Qs7tfv1lq/FWNRtoah3WQTGeE2eC9eF
xFyz/ME+AGD8Rol3Cjek8EEWDTdTwcqRoIQHN4AYdzPBRu6sJ40376bg8wqO2327NJzIlc+Zn85G
KQeSUoD1aqeToK2qoLZ6Pbqf1BcZB81IgLRQOWOnIts8xOTTKdEWofBhs7z1rVa1y56O0R+UDubt
RGeOAFhM8QW3ALolJ79cAc0E4DUbDpD7jZZiGtaymko4g2pxpBFC7qnRm3irxzDdO6R7sH1K3w6p
Hpfo4tkqiJvmC8ccUlaxJDBzKOCzBqhGYvpscCDKsyB9Tc49IS0vtmmNJzvSw6tFB4ij+h3Z90o4
URYZ8l/IbMEythTfjs0LNzMWk0RFNYfsCEHs31jnTMBUnEBQQQL3gMfhUxBhGe6dLfVPNyAVRmdf
UBuB1YhS3rYDjncaYYPzeJvlWCfcFBrPCsU+il0iENdVExSlE/m3lHBBUSe3xbbxjgUuCClZB4Pe
llhrERmX7FVz/8KLtfJp4JE3RYxXVLKAjeiyXob695WO5AaAOYFq4pbp+cgy1bM5ApjsbIuWJxhD
t+1+r1h8jBJ2Oh2CYcsRkDnzr30A/Ji/l47M9GI3z75WJ/vCFTTmi0hTJ3X8stuNUfH6kaGSBtcW
KmDXTBpoIsfCKkepiyQ2RYWhfxkZbj9JkrUr1EyyraP4aIREQqO/LsghhPnKgmmiWcFSM26RdQGD
Eu1ZEfJEy/1aAmibXtc45kay8zcvkKOMkxSW7n1NBQkzBdYlgnbXxIWNjH9RdC0tbGY1YspzSzFT
EhrRdNIjlUgFachhV92JR5gTvRuAM27Xl6toWZ2BuHSOoLdlfUunQgYihDCLRMKYTxJA1VcwLI7N
RM3CmPYOpyr0ar0we291O4P/30PMC15LlvN+ossc2NaVNdccCXcv+7MfSIYnCXbLhGP/uYj5Pz0m
1M22HMWXLFmEfJRU5lTtmFWrAOF29OtTrzq74KeIDIPPY+O2D1YQSAdopg2gGZtvYEl9UlknOrgE
9tILAqtb33OHL2jLS4zPcttp86A0oqBucVHD0xmFylf7/m0RE/2w00YcnPt2zczKdAJzaiaZXtC2
rnW0Jq7iN6OHK/2JHFEB2HKugv7NxaJKKuY/k3yoAInx7/cNnBRPhLiRkxZnE3lA/FyDUxszW9EH
QAe40qpYreKGUg3IvV3QpYXogidDOH6OeYD1yAAJIcl9LCT8ap4uO99yt66KRSwiuU6MQpNseU4k
5rH7jLvaCVkgQRBRnebo9TLhCed6IvjYhhWya9QA+5GQnJVe3nxz8xe8S7yIaHcy0FzsXbggsnRp
CU6Ek3w3UaF06Mvfw2+IkKyC59lL9CvGYUSRJhX6I+YMqf4Ktv+v+GAjau4CTKY6yBRtAY32JxCw
TbbZcF2iz3KvuonBeqpaZYFLJuiPB4tOq+jOggCaxGMsbiRWp8CGVndT1RV1ysOSnJrkT/+Qe2sq
Av19+2hd+bjDKtW5QS6/XookcwNaBT0EFjl5DqcR3KRekOzbZzzLp0zpb2ijcsnUQhEGw2odmIcA
mN92hrs2hg/XgXBaOeM3kHncWpQQEE+XREtIwNpVYyJi9+aay8WZ0o62DTxIJpX0O9pyO3eS/+J+
kCbu7Jh4GN0diuGX8UVG/OpFwDUipYjy+/3PHIuSe6uG4v+XwJG/3x8pWr2F6mEYdcHjLA6/sKig
y2rPsiU2Gp0V8etOjbhH4Cwzx1+rbO6gOR7d5Q/ZzBXAMFgl5zo0nC3BUI93IRWnMiCrAbDLLSUH
xNuz+1DFCeqAxMNzkXZNoZci+ZswiS4O2jLz5AzQ6idA8yAiP+4CjAULIqdK7S5tyPn+TTPKgsED
0NOHhILvYP/rk41XmKj0h/hWUktDQWZxD0Vkdmset3ybZauQr/sr8xFun3ur5L0nNYvHJ8LVEsPO
YnNGPxE9xLCCiXGFrZYezYAySCJniEiF0rkKpl7Ngtr3wKZ2Ufjc9x5RT2u2f/XX4YHCj215/G8R
3x6Mdq/ysF7mGjruzbOuVlRAYa0C6ZXAeE2sh02s35CBH1mOm9VqaUurZvRYJXj0W5o/sfeGAa8Q
f2kfYkzZp5aJ0neErI62yG2X3quNgdw37y7qGtoyZJ1DLylM/7iyxk6/5mABZMeY/504ckjZOw99
IumH/qa08vBCwxVtJsX2yjzmXXhytF5BET7iv4yQAqfYB+Hjul+6p7SjNOnzmfc7iO8x/JyMGO4h
5IA33qGQVUEHsoeHmRRKZptltwC3oCM8ekwHmEbSl9ObKIMIv0lRLRKnk0FhA4f/ds4CCfb1j7HH
FDCaXj2AThq0m/um5IPCFZLjPXSlTsQr7kx8Bpq6lutvoRgz7zZfJ4Ssc4qqdKO2DycDA8tjjPvv
KfYfQWvCftgLK6IkZWiLAfUi5LmKKUy4/buSKhs9XyD8iEMGF1tSfSqQZifJkQoJ8RDpKQUAlJh4
EzysHqntAfOsTjy1rywwbZA8+TKI9QmK+3AFxc21rphUo0lr1jd8ClWZUwO+pw9FzrTrjicoMdLS
0BXp6sNiesolirWWHH3gXaF3nq9mZLKKFoFq3WyNTXjJzYN9WdEiaFG+fCuUHAcEL99ARvdrJ5dC
J8L9s36gbIFjLIiZxqD9hEyFePtjKncyIpbIEx4ttf4Wgcu6TtPhlx+L9GWv+k5GIp4b5O8mN927
3h0OqdpcYDlztExiF1qTp1oYHJPHqdQNGS01kgOil9fqnb2U03DgN/9bCLPW3eZtchnP3zsczUgx
sFrCDaitQKihmDwfQTeJL6ArtYShs9ZDPFx67epjrgN4k0AaYGcZ0JChUOZ8fiusAHh6JTUMuqjJ
VxAt/cgaULBMXAxRLGulamCGrYC8nWW9FuLBQxKTiVRQu1Lujy+19tjGr1YZsp9s6fo59iPtEajY
CtuTQKyFXUHzXrD79RZTfM6TN6cXVZKiIhvgHH2oT4IOroVJjKmwBRb5O1LWOcBPaMtRWHGRk+p0
LLHHVMP7qifMK4efKC8iuzEvfdrVIcleNCHvAMKPJbjFv7mzDKhGDdVfHunjygyDEwycCxNNzGIu
aZy/doiT9GVF8XsfE9dhx1VIn/C0QcMoifUUHuU4YeuHXzc2Ckhn31hfj5o8CnDU7/LGokdNdD5H
Y8eTail4Ss/1CJHqcXIA8nAOGDrstsyXuG7Sto0PnPC9BP/btfHc++PzYNZjbr5hUcPApTUudIgz
4/S5UmSo/rO9xle9YId1pCHgcQv+3EmSspA93r/VRIIVcdp/Ur54RZ9pgWhmMGOdqNpJu+h07Hxd
W46XOYpOAPpQn/tay+nOv7pZnHiy3cPx3EKFx+bB9sMaBmXIPDBn/wfokreMPsQfn9sMxXsRRa9l
Y4jtc41UX3XxFG3feqrSQjknrh9pGtYef6VukxWHdRaxtV4EaS72r3zRkRIVrpPiEqr7sGBu0sz2
p4L2yPiBrkG7+qeMXxpCTd+a0MmCa7zqeTlZpHbK2vJzU8/E9erkpaiiryX1NlOY1COiyC+DVxhZ
sP34Wm5kXo81TerQ3CrY1LAJHS0SBs9zpSvRYsoEzB1kgWz3PjtIx4XLhG7xZdq5ZF8HA9G3g5A3
T/+DBIm5zoYMBuvgmqscEuGI9r0yqgWD0wsbzys1464ABevlM5T673obbdWKzaR3/wjqMm50lTcS
0f2+I24GWMDHINd1kYUW9Sz4Mp4N7lUE36yifv8NzML1lGdP0ye9YZhZBIEEAc73p52YYR44EUGz
UBoHFSdVrHSu2EnE7jibFgZ7LTEDzy6HBFGULjrwYv0r20SBI9wXr+Re+ofS8XxgUxM2xO7Ulp5z
HCBw1mI/hWWlfalhEaJkJ1vupY/L94edxAR8mbk12ykMwHewiOh8tWCGcw7dkwzpMgXqwTAQGWYs
7Zp3bwj/Yli48X0za6T1TdPU7sbJ41LrffsCdDOntgL6UGcwkf66D/p3M/rey7ejUfqlffxAki9o
SwdFpOnBGf18jWSnwcRH6HQCW5ZTI2CCd0O5rOC2t14XjJxsnWpwiNiDoo1MFSSHUi68OyhnT31m
lTvhQVCF+cPlBTW1QmsVyfqosSQ/4ip091oav/SSLBV+LQxmXdZRbxso64m5jbi3/UI4ZgMjkMBT
CBnlXui3o4OqOCn4xXyXGb4yt62HU3nFaCVW5WAIioEd9dgRm1K27czyiSmYarcyjJ/J0euaxYDc
WvjxFELKlkiUBj8nvcr2xgC/vYu/IRSw6jh5X9nTG2hHbBP2gUc38a97xgORSCduL5wMGGq4vews
oDmOz29hlOg48kRXgpdcCU22FLoZfSW0TYwiMN6siBll90QEh6JianVz1L5nGslgKfqyxzefc8de
AyM6YXUwfJumgDawlTEEZd/3kO7XFSLY1GxjLiDKkkQcp35zHZVLxSVQWsZCYoAWCiOajpFgEFhF
Jk68Wc+30LCEC2oN8rQtYeUcDagKdKBG1jGboodr0lmJiA5xM777gRlRoKjRjwI0p+WSq8OycrIc
ea/iZf39vEdZ3+pz+qpfJsovqWNGQYUc2jkLF+9Mag7GIHBnPSUlGfLqK1bnNuHBa5MEl4JLPDwe
MJREuCq5Qq5V5hg0epepxwIfrBcVivOdUdLVQO7UBIkH8AKjVrFg2m65L51uUwhbvjJGx2z7s2lV
swUyaCiQOB9ECCz/tL4Kmwc1Eic1AOrd3H0mTXDX3T2Z64HmJH0Fj623k0FYEVUscO73nbHz5yVF
Pl6xi/Qg0YGyQXx3Dxx82os1eAmjwwGrYRyGPXYBN2KztefUO59bXQ4QUMxRZYwdtmRamzyG/BCJ
xHylEypN7ZyEGTYUZ3Gv9TlMewoEXp5NIx/BWmyzF4lNfcFd0qBoi82VVBTGZJOJhkpm2OY8ByxO
TM7gPeYNYp8shZcHd7tdDhElUtDFEfWoOhxPy6KTGUNg4+M0g9JGtLIqLGyR8rxUD5qM2GsK6kwA
6/TsujuKu3HXax8BgPcB/h7k+WhVeTyqOdXThkFnoEMN0euL4HJ61A6m9cPKXxwZ9xwgWZenVqrV
5IycNWDMaQFKqaEccwLBoTcV3fHVGFsLgLWjrPkG7iK3TAeTZ74CPLYVexUP9Z7ryWTpKvT4qWH6
C7L9p677iII5AoXQO5BWM+36vpBXCiQ0l1+iLf/80SJKt8cKu4LNbCTrma0e6W6QaLBjCFLtxa7S
eMvMLN7shgVFXmO+zOvVCtopGZyo+F6ZdVUDUFfx4vjOVVYXNMeiRgwPm6QmzgQjac0IgUHh3/Uk
mMHB5mcd9yij8ZcccErTp1fPoxCOERb27GLjcnW1IkV+iGBEZKA6Z22H88Qb6JTGpaxwtuDkXcAN
a/WYAjv72e4Y7fN6quyXK/8uYCrgdlBsqacVi/c3b8R3fhJt4NWuc0Big3mVv+mVoLyXynno62Xx
THpAP/tCi2WeUmqM4oNkHc90Wu879+LDrrJL+689Ro8aKec9fcgCl9igxBjz667d6lSrVYFaVoDO
wlYoN4gokENb1V8fofJvNYrOmVcwZ6hRKdleRWxwOP4PejLNL43HDB1LjdLP3VOHVhxX7tyUgZ+I
yswrRB9sX3m8shAK2Wxy1QkD5WwHCA/EYxwnGJnZ6STkLvxYo+Mpg8QVV3BMBC6piK9IRjNu0RPe
iOtX4QahBmZfuIEj+wxjkAEi+XYEUQDWS9RNIsT0VoEwb+U5cQ//4AQyliYWLTUeQPxa04VnJrHu
xX4sOyyQLpoeES+MDqvNfFmYA4CjpPf3P7rlMozAtXQJY3DH7UK5xC/Vn/pEHEdYtGuYA3VIWl7W
JpRDxOkCNFkxmlBdkSVEU1T/3LbTE+ZtP8Ni8XzWwNRcePv7yZ+sITkuC2/JS7QGWbw9vRbqcN4w
f8IclnIK+okGIsgQAjT2ALuLqhrBUqLfoqjTiUy2irNQ5fUqz2EjdqArYyX9bIQKHbZmbTdJkV6V
JhspS2uk5AhOsiwMWEa/1Fq+Mg78JR4V37QY0pVlZHpOMo5Kk3G8XpsrXmZaSU9Q0P+nYMxryIHN
uEzCVHi4sPUCY9qDRX6VTaj+G8ikaI9XloDKRqbZgRJuCqfmpbjupSPKej/kR62nVmMjt3vgGOFJ
LcjCdh2f4s48QlP6151WRcXHzA5bBouOj0CBa7k/mbt66etiTwAQFtWGz03KOQ2Dv9c+6I76rH2o
mAEFtQSWh9sgfI9SkSsivrpCbjRALEYWefcjpTqTqlLDi5uPWMfkpEQi4Hcw7UVPJMZ1Fesnp6u5
fkOE48rXnIbE7ayEAggjSSUwc0vaqHkZKYaAJi8P5JLANTWx/29APVtsXPWuxv6Au+fuhqOufXI7
+DeynJG/Xyo23613rY4DbBc1bj5GDtU6UrM1nByoD2ypPru6GY8pk/Wir/Avu+KtkKVhwhuipDkA
f1BZrn2t8ADEoOYqAnwHc6ya8mKCrWXyseyImkFHi0b9qpS+k29Dd0hI7DCAJTF4hbZhIUsMNCu1
EdOfUCbT8L/0TmiupiEBE/NKcwCkPMxo85aZLCof9k753PhCskeTmyM57QOaZjtUrHrqTdJWlPC7
coD1F2yVgWpkK20K/70ft/WRsUGeABnbSmOrQv+bYX43mN4aQHMQia0e/0ZdG/iWz26C6aes4BM9
Hq6A7S3Rk7MPThRNSLLQep1MRjzSq7YEb3qfe3kl4zkR8scmme8Q+euoWLDtNO40HLsCCRX0ZbDJ
btbmhBkEv42eNNuIuSlHnUch+6PS3sLngdYU3sX68y6SbSD6uuioDz5nKcmVIUdva8K1sWsacQOc
mRpmuuXQSUqqicNxiai/DsNjbdrX/5DWWnJ5eghwCdIEl4/sV9goC2OMXaGYt7R45ZHf2MijKsdo
i5YgzQp2J1glYewCt8zu3LxFz+YnTLoVESPf9x7W8K32PsKh5qGZ/EJYNajZr1n1hxDlzY1JPc8x
WtMI4nW03ILYMelCVw4bzDZXoXVcdGBNURI0JeA9h3YJ9xN8MaLmy88YOCVSHZb/c5CZgeeoQpdO
NOruNB1lZAgaZtaTHoEt643ZFkdtOu6wsuRhnfqRLqL7PcPv2MUzapCmCoafhLkHOro96wF10CRF
nLWj7uLBnjvcCQFQOXkHm/LL1ouEveBiSNxR/ikM+O70WxmwCemr0A/ZTWVSFav/3+ZaYWUwNlpd
o9LxRLJ5JkNS1+TwtB/UK+nAiFvpVXioCfv5K86jn2RqgXpSOWpzHHFjV1cHKLEIyKUajhJZUQ29
AcI7kdPsOfihAlAHJQrRLTSq0egYCbvHcYDWMlDUND4Tsq4WeEkxDWQEHvM0pPoNj0RE6Ln8oq1B
vMEjNkyvvrX79S45N8SOXxofHbvLNUgaBTD/BdS3x7ENiqUYBG1kwJm7pVmkgL4BJk7HHhIFNYJy
DyqFO5kFffiz/DIRSanyjhu7i+uKqPxyweoScph6ZwYIHra+xVLE9JxHfN8ptjT+wh7iV1D05BG8
MiI8KlBcgnFCaGnqZ8SIhG5Tu4np9MCLQhTuNFNmBS3BS6RD2NM9xtbAmMrLwjeZsD1kDbMc1bjS
NkMUkbDcXmFvanByXtVzRcs4kDxNDhj50M9yB3inDyazCDeK3PduVEPum9mI91HyHVz1Wr6+G53T
W22tib+dY78SPz+8KYmf4853vYpihgeG89n0T6OHQnzUAxJ2GNgRixC4dEJo0Cr8iBopAEb7ykxm
BSZkaiIM3ERi/nhJUkde7A09Cli74bp9p2C6QllAFdxGAKoZupBAUi4eky9WwaD6u/7DuRgZ6eG5
WWdICR4axJvH1lpd3tdcxAY95ZDVXSBjCPSgkgrqpmgvImt35kAiDflGs+KWN0Z1rQq5GzibQZ2e
mEdIFL01mspNp8A2CctwblqaMtmiqU0DMvyUE+MpNt/AhpWaE0zeH2D6KfVuzdfKs/0AuOHvR3nF
Gq9qYQ3ZoLByKgiwsJnwu7T4xcK3yS2MXbw7xfb4Xl5RccvocuRkt3A1eoh1KdyQuRYhqt5d/yRt
mjsMY9pJlHpfADmXSwsvWGBjE0d6MdwXB7u6an0ne1J1pNvvWRPHuJIIygMEGDgWDBUb7B+tQd9c
fJu2CysE8eHzkOcqMVqxYy4uYeRqQcrx9rIxZyKEs5q2qUayXFcZXzgL0I4ACl/sE2oWuvqxHP1X
2uKEECSNbUr8oddYa9gs9OIvA8Qb26P0DXlf23ky5WXlTw7B+ise2ajy3dd4ODT+YeWQQj4+63Sb
oDcbSeVmJQ4BqaX2vYu4V02o1kq4thMxSLdTL7pfqEywWqR3gjkDJdey6Rl6MJD282vz0ftYURuA
cEvR6CLTvZXbzZVysKJ6UiW3ZENKoucKJl+2EWsRe+e27tDspe8QKeKXAmmHerqBscwFi04Mnabb
qxUktkn2MZTaHIr18YG/9y+t4Y/XxzwdQeWnZ/J56Um5XCwSe2aEQ9kEZTFs7mvcfoNKXGpErAYH
36lrGtAl8DBXT/gM5XuWNoeJL5prpzZGHxav+GMI1c/G4TuTmoGMoEXfeaUqvn6hjVzqTkMvoYLN
hHHMMA9xVTfA36HRaeMg8e5eU4n7iQ044mT6uwPYFKLdiLXX+9l6mgAduf1HK3sCB4C6Uj4iWt5X
WRTDSFx9ptf8yX92Wqkqk7i+aGUcF2EdSqtGiNYXArVAAaiB2llmGcuZ3I7Q5HzHnwa4GMUqYMiZ
+l/nOYRE2vfsPijJVXOuU5rRiv0aaY2eVOWMHrvANQ1lAywc8Bkyix2FrKv2j3zBatOXWPeLpGVB
mlf/D/jRb+xOfHdhX/nDTX1G705wp1puUNjLuzwEdN8d3vO9KFYlMmlYeEl3ZHmXltI8cgfTMt7W
h9OYPcoTLzmOhkVlem5i9BY2+Yfmu66fvvGva87XTVJeXbX7sv6DPXUcvmn0RaSoMhbT1msgSElc
1n9XBhzEfOOa57Pjdah5LOm1sfolKSRGr2QtYswCn6vqpLgBI0oawGEyfjlVde1dRdexJYFv4vSF
KVW+wA2zdS+Ovs/W328RHBTHRG66qj+aTHcNz26S2UKVFV2Zqc+3MGNtdDBg+9XWNvsRhN9GhtYi
KT9Ajg96Zbz1rqK09sIUKcC00BeowPmjaV6AaMLNLPMhf9WpzeMw8sajBcyM+qlUWHnN5nSC4VZC
nHvpZXFzkuNSNkqMFz1QpngQDqibA0hNOvLBg/SBy8v5ZKliDgxgnGNouNz53hUikYt/EmtHKozk
Ix0ljq/KapSlRduGfDZ1W14x926KHWkuAKIlfip8ya+woT/FaHM9e+IM8aTzjlDhYgbm4Bdxtef5
sPVmP+aX6R3BY4TY6qy3rdCvO9LCXPjx5MbXUkfhZrWH8VJ3Lq+62UkPxcKWsnt3rdki1rTUVdTX
joYU1+03WbA8AupGYM3REGVWb17ycbCMM7bCsDZ+QEvRLpjwhOpIGpjVuGpr3I1RRCOijUya5Azi
ZGL/cUexlo3wVdWBAW5dFTcJ4CWnKwAysyglnoOCQ0O02bABFm9fm+eVRt96nUQ9ZezTG/2Hkz6E
9tJs2TYDBxrSr/NU9DwsKHEiHWsqBJ8FU1/2Cq2ZpNs0r9L+LOscbNCu0jXZBX7CQp/6yDcllgJy
qituLHMSQyWw0LecScmFYHvaCE1fgdeQYzLyj2gQWsuHcD8tUvmsHU2SFA3Izt4uy52n6fcgNwpB
D4dScK9VAfHcVcwIxbYPk2Y4m3tlFc3I6nWDn38f8G53AV+zunCK0RMyWdpWZipsIm0DKspmAMgY
LKw8RQKPnYy4RRRqZa4nk/cG6Bqp+bzAARJV41xYZ2G4mDm4WvPJURYxgAU+XhPnjTjxTH8JWezY
/1pfYkVZABcy7wDb2T0v2xOwbAwoiatO2jyyw3AFDyweJfJZOAgpqEU3X03DzQg64xirdifPieLC
+e04CiPg5r0EEO9u7sUTIlXj23okC5ntX6Mfln9Nc9APu1PyE9nxcUJIDezcdSnv2N37NxjfdHfD
UwvIUZ1jD2WZiqg5QG2kak209Ave8dEH8u+qvaEMz8ppugh4KWB1THZz46B/Z+QweeIMOzoanS8K
0zZJL8BvbcwyxM7Y2sPge9Kvub6bcqAtBBsdfkgB1/0ONQ2CgzJ8dbQZSV/Zu1pSikjdcXHZMMWE
Oj2YM0Huk3k39VxStIuFUQquRLXT9+rJDZ9NnDfsZKFErV/uXqu6PgijL19J1De+IeOjI4E3CM6i
lCV4gH2XgZU8s90+irc9kf1/to+z0nF5iWFUpa4BpmRyjE1JfhWpJzDBtZCP4KyFFNfFPgwgd6RS
RgstVNMQEIOFCU75dNmfpC6sN3unCg2QxBv32qinWqW+YmSEPqcyjBxx1W+f08aIJeJh4dL8FndC
W1B8Qt7dMnRq3cZ+k1Q21HgKATl6o297yItx6/a9Lt+zAkDWY+ES9fifRA6GvxTRdQth9SlwRLeF
1i4r8ECw8HO4SWtvla8aWBnSSzRdOl0dqdl7je8v82RGtyL0b0JD1hVGCJNtE+3q60mgdV9CLdWW
xP34FINlWxStUaN2hBnITw/uKW5smYyz4paYZrrLszCNsOxnR1Aa9NqOdkr/K0TJfMqPyxTHtDJC
ccxEbiCE7zT1dZ27K2ejPva76pvWhwoLK/d05qwgNJFR2PExTrZVMGMuD3tZuwkIZe5sSJJSF3d5
i+r34o7BKrXFOsc5frIethU2iAem8tCLcHjl8XuMkJOGZOJ27/+DnEjjmxPd8tLOyVCpk+ozWt9K
oXJDx6sJArSkQPeU2mAEI4b1uHD7CVGdwhqdsdoxsrzwOIlgaBVTcJSmM4CJqW+MxvRa3Vfx7FIg
PFbGVjFhbttD4JiAZ+uKTaURLl+mkvbjSKlrFUboXx3fbA0Nnl/7a4l5h6hgBxtREKz2HOYwTrgv
Ij+h4A0VlyrEtnkYfxpY5V5tB4gfUB5u/KluChjvcAyDBkJ/v03cNpyOsrDKboU7RotiJRBgI/k8
Oc2EKWh5Zfz4Wb1OoPZ7wDP11WgP/d1YLWhRWXd0P1BcD0w6dmqn46iMPJ+P6hSRYRjWcFizb2mD
jMwKs8LBBU6qIWC4J9rRyIXogtVm3sJC3hZQBOxrJX6/zZkMi67fjpRzFCg4wbRTbowSAKyqkTsg
YY272xvKUFxDZQmHlCZ+r0zKT2y90CRLmBHldeqXmTgKHObep9fz7uwoVjNZIgcXOxiUWRmA6+sX
WG+eE2lE1dWFBJTDxOM+JHe6G0srrFTrI1BDmz6REaopkDOuD2rpU+5gnHSLUZxg/sNba1gR8ITm
rEbkTjGVUKFv9cyj+wnDv88t5YkAUS6am1oQYZmoXxKMLL2kuVimEWgVAZ9wWtCagZCKpgz+FZL6
uWbJJBHcXL2NrgWISF5azY2AqufdkNwpUFEETFIlJ9VVND5KOVf6m0wZMh9Sgmp6nA0xYOKUGyMv
4c7rKl02LLPlz6d53WDGJO/SckSXtEdY972LgIf3dDs+GBaxwMdc+o5seBguwV0Yi8NHAUbrxZep
R4h+EGgNbRJAxvRD9BolHndQS2C7ffI7SMEARQUiLa1QYeNPgs+Bc9/gtG6eOLcGxafSSNKp7KH8
++IvtooFfEDJxRmFDKfxKUKgsRmnO4TzXovD8GAGTAxFDp+es94/h8My4VtCvtLx5CMTmjIkMi3h
lnud3rHEz8YhvMjMhI1hyxSNdMfqbWaHKx+C3pXR5Ps+YLz9pSLqn5iyDUZO6QPP3/ICpFkGCPy2
sSbHXuv8YefzLEvbmT+AhaARAyRbsWCaPjX0mWvs1pFKJ11d5xhmoqrlPiRcm2wK5vxebhuHJuKC
lT0BTygVzPlOzVxcfpegGCkTwY6P9H5SESRtrlERkx1lTVHafRwN31LTjfAIz6tJ1kgf8B9iRQg7
Z9dzPf/tnVcg4NJGNp3GAqeJoDUXru8QwSpEqw7A6STf76pKdyfqh+2s59wpDzl2vDfCd0jbXPco
6f3VBD6qVrD1X/CAXXRHZm/I5JxDbS/Vt9n/VWz4MwjjNoDEBouBd29cbmAb3o9DoYQDKMJs+Qw9
0oi05O/8g81lc9BFmhKUl/iViNXeJj6QVtGVM8SAFR5ir1vTkmK0CjTr1dSLxxbytII3/IZ19Q/+
t/iew882yiwrGnngHnZgmpNV6+EHJG5aJq9lURDIsh8qqaMBRQziSAtNrAUdCPwlzhoUyc232cdy
OIva51XqQ2eHrPhKw7V2CoxbmmSImsABZw7fd3MJxXB/e62HjSRZJBPVgDrRa/WCcFB3kA0OfIAD
/QZCNHA4lqP/4EoFodZDJotvy8CHIDXq+EqjYM5FF3+KoMC45MHlERspK58vmFFtUyV9YSv7aVIU
IzWXSaBpTHvGRAOeiA60VK6eKn8pM0fNM5d+jisEolYJrkrzfmJ6+bafnh+HU09pQ5VFn92Z47y4
GNaAet4TqFTKeRWqz8pckL5OJMQhDU5z+DKYh5JQuWeA8oZMh5G+H0H4jtVPB1KT4wRYB3M4Sxf4
6Qbf+VSH4iSl5efU+WH9yeoArel0gpVgbTeuLXimFLt7pe5PHHZrJOCsC+PNj1C75xUVSK7D3Wm/
CzsEjAqvVRCdkfhpY7vqBavCc8G8hXOEGpINCcXbJDNk+RCPnvIfSQuktAOBOzCRgsE9y5963liS
+WF1W+t//p06wEduUgzQSWfvnd5qCWbQfifFeYavQfCaVXG72ji/kZ0iGT9Y0aMQsdvYkz+uq/A8
HfY7ocvlNx2aM59+W2ZLmMvOB6L4SjvSQBzb34VHVEKWPw71WTM8b2g5QJsQFdaT1LYnYlYRrrQd
3b8Z8HRQZEoAJL6P8lTYJGAnd3be5smjMbdqjYqmk3u2szFRwmEW1bwgvgnID6x2GvF+1Y+Bv1/V
9dVUex7XekPPYN/HulnTl5Nw3LzIjmT4sbCboccBbUKnyUJ2+NBzyIolkBRKZYDYr2Hj7qMbDSi7
Ma5/j6Q5LkyqbCntphm3xkXq3UMb0QDoSE2AaAz+G8d2wVKkhIK0aVVT9vvI3SYUPi1tRWW1e8/H
dnN0kWNyH/FlOoXpdoTvmHz03qA=
`pragma protect end_protected
