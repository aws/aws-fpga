// =============================================================================
// Copyright 2016 Amazon.com, Inc. or its affiliates.
// All Rights Reserved Worldwide.
// Amazon Confidential information
// Restricted NDA Material
// =============================================================================


//FIXME -- Need to do the clocking correctly:
//    - Async Stream between PCIe cores and User logic

module sh #(
                     parameter NUM_HMC = 4,
                     parameter NUM_QSFP = 4,
                     parameter NUM_PCIE = 1,
                     parameter NUM_GTY = 4,
                     parameter NUM_I2C = 2,
                     parameter NUM_POWER = 4,
                     parameter DDR_C_PRESENT = 0
                  )

   (
   //--------------------
   // Main input clock
   //--------------------
//   input clk_in_n,
//   input clk_in_p,
//
//   input rst_n,
//

   input                       clk_xtra_p,
   input                       clk_xtra_n,

   input [31:0]                cl_sh_status0,
   input [31:0]                cl_sh_status1,
   input [31:0]                cl_sh_id0,
   input [31:0]                cl_sh_id1,

   output logic[31:0]          sh_cl_ctl0,
   output logic[31:0]          sh_cl_ctl1,
   output logic                clk_xtra,
   output logic                rst_xtra_n,
   output logic[1:0]           sh_cl_pwr_state,

   //------------------------
   // PCI Express
   //------------------------
   output logic [15:0]         pci_txp,
   output logic [15:0]         pci_txn,
   input [15:0]                pci_rxp,
   input [15:0]                pci_rxn,

   input                       pci_clk_p,
   input                       pci_clk_n,
   input                       pci_rst_n,

    
   output logic                clk_out,
   output logic                rst_out_n,

   output logic                sh_cl_flr_assert,
   input                       cl_sh_flr_done

   //-------------------------------   
   // HMC
   //-------------------------------   
   ,
   output logic               hmc_iic_scl_i,
   input                      hmc_iic_scl_o,
   input                      hmc_iic_scl_t,
   output logic               hmc_iic_sda_i,
   input                      hmc_iic_sda_o,
   input                      hmc_iic_sda_t,

   output[7:0]                 sh_hmc_stat_addr,
   output                      sh_hmc_stat_wr,
   output                      sh_hmc_stat_rd,
   output[31:0]                sh_hmc_stat_wdata,

   input                       hmc_sh_stat_ack,
   input [31:0]                hmc_sh_stat_rdata,

   input[7:0]                  hmc_sh_stat_int

    
   ,
   //-------------------------------------
   // PCIe Interface from CL (AXI-4) (CL is PCI-master)
   //-------------------------------------
   input [4:0]                 cl_sh_pcim_awid[NUM_PCIE-1:0],
   input [63:0]                cl_sh_pcim_awaddr[NUM_PCIE-1:0],
   input [7:0]                 cl_sh_pcim_awlen[NUM_PCIE-1:0],
   input [18:0]                cl_sh_pcim_awuser[NUM_PCIE-1:0], //DW length of transfer
   input [NUM_PCIE-1:0]        cl_sh_pcim_awvalid,
   output logic [NUM_PCIE-1:0] sh_cl_pcim_awready,

//Not used   input [4:0]                 cl_sh_pcim_wid[NUM_PCIE-1:0],
   input [511:0]               cl_sh_pcim_wdata[NUM_PCIE-1:0],
   input [63:0]                cl_sh_pcim_wstrb[NUM_PCIE-1:0],
   input [NUM_PCIE-1:0]        cl_sh_pcim_wlast,
   input [NUM_PCIE-1:0]        cl_sh_pcim_wvalid,
   output logic [NUM_PCIE-1:0] sh_cl_pcim_wready,

   output logic [4:0]          sh_cl_pcim_bid[NUM_PCIE-1:0],
   output logic [1:0]          sh_cl_pcim_bresp[NUM_PCIE-1:0],
   output logic [NUM_PCIE-1:0] sh_cl_pcim_bvalid,
   input [NUM_PCIE-1:0]        cl_sh_pcim_bready,

   input [4:0]                 cl_sh_pcim_arid[NUM_PCIE-1:0],
   input [63:0]                cl_sh_pcim_araddr[NUM_PCIE-1:0],
   input [7:0]                 cl_sh_pcim_arlen[NUM_PCIE-1:0],
   input [18:0]                cl_sh_pcim_aruser[NUM_PCIE-1:0], //DW length of transfer
   input [NUM_PCIE-1:0]        cl_sh_pcim_arvalid,
   output logic [NUM_PCIE-1:0] sh_cl_pcim_arready,

   output logic [4:0]          sh_cl_pcim_rid[NUM_PCIE-1:0],
   output logic [511:0]        sh_cl_pcim_rdata[NUM_PCIE-1:0],
   output logic [1:0]          sh_cl_pcim_rresp[NUM_PCIE-1:0],
   output logic [NUM_PCIE-1:0] sh_cl_pcim_rlast,
   output logic [NUM_PCIE-1:0] sh_cl_pcim_rvalid,
   input [NUM_PCIE-1:0]        cl_sh_pcim_rready,

   output logic[1:0] cfg_max_payload[NUM_PCIE-1:0],               //Max payload size - 00:128B, 01:256B, 10:512B
   output logic[2:0] cfg_max_read_req[NUM_PCIE-1:0],              //Max read requst size - 000b:128B, 001b:256B, 010b:512B, 011b:1024B
                                                                  // 100b-2048B, 101b:4096B


   //-------------------------------------
   // PCIe Interface to CL (AXI-4) (CL is PCI-slave)
   //-------------------------------------
   output [63:0]               sh_cl_pcis_awaddr[NUM_PCIE-1:0],
   output [4:0]                sh_cl_pcis_awid[NUM_PCIE-1:0],
   output [7:0]                sh_cl_pcis_awlen[NUM_PCIE-1:0],
//   output [7:0]                sh_cl_pcis_awuser[NUM_PCIE-1:0],
   output [NUM_PCIE-1:0]       sh_cl_pcis_awvalid,
   input [NUM_PCIE-1:0]        cl_sh_pcis_awready,

   output [511:0]              sh_cl_pcis_wdata[NUM_PCIE-1:0],
   output [63:0]               sh_cl_pcis_wstrb[NUM_PCIE-1:0],
   output [NUM_PCIE-1:0]       sh_cl_pcis_wvalid,
   output [NUM_PCIE-1:0]       sh_cl_pcis_wlast,
   input [NUM_PCIE-1:0]        cl_sh_pcis_wready,

   input [1:0]                 cl_sh_pcis_bresp[NUM_PCIE-1:0],
   input [NUM_PCIE-1:0]        cl_sh_pcis_bvalid,
   input [4:0]                 cl_sh_pcis_bid[NUM_PCIE-1:0],
   output [NUM_PCIE-1:0]       sh_cl_pcis_bready,

   output [63:0]               sh_cl_pcis_araddr[NUM_PCIE-1:0],
   output [4:0]                sh_cl_pcis_arid[NUM_PCIE-1:0],
   output [7:0]                sh_cl_pcis_arlen[NUM_PCIE-1:0],
//   output [7:0]                sh_cl_pcis_aruser[NUM_PCIE-1:0],
   output [NUM_PCIE-1:0]       sh_cl_pcis_arvalid,
   input [NUM_PCIE-1:0]        cl_sh_pcis_arready,

   input [4:0]                 cl_sh_pcis_rid[NUM_PCIE-1:0],
   input [511:0]               cl_sh_pcis_rdata[NUM_PCIE-1:0],
   input [1:0]                 cl_sh_pcis_rresp[NUM_PCIE-1:0],
   input [NUM_PCIE-1:0]        cl_sh_pcis_rlast,
   input [NUM_PCIE-1:0]        cl_sh_pcis_rvalid,
   output [NUM_PCIE-1:0]       sh_cl_pcis_rready

`ifndef NO_XDMA
    ,
    input [15:0] cl_sh_irq_req,
    output [15:0] sh_cl_irq_ack
`else
    
`ifndef VU190    

`ifdef MSIX_PRESENT
   ,
   //-----------------------------------------
   // CL MSIX
   //-----------------------------------------
    input               cl_sh_msix_int,
    input [7:0]         cl_sh_msix_vec,
    output logic        sh_cl_msix_int_sent,
    output logic        sh_cl_msix_int_ack
`endif //  `ifdef MSIX_PRESENT

`endif //  `ifndef VU190
         
`endif // !`ifndef NO_XDMA
    
   ,
   input [NUM_GTY-1:0]        cl_sh_aurora_channel_up,
   output[7:0]                 sh_aurora_stat_addr,
   output                      sh_aurora_stat_wr,
   output                      sh_aurora_stat_rd,
   output[31:0]                sh_aurora_stat_wdata,

   input                       aurora_sh_stat_ack,
   input [31:0]                aurora_sh_stat_rdata,
   input[7:0]                 aurora_sh_stat_int

   //--------------------------------------------------------------
   // DDR[3] (M_C_) interface 
   //--------------------------------------------------------------
   ,
   // ------------------- DDR4 x72 RDIMM 2100 Interface C ----------------------------------
   input                       CLK_300M_DIMM2_DP,
   input                       CLK_300M_DIMM2_DN,
   output logic                M_C_ACT_N,
   output logic [16:0]         M_C_MA,
   output logic [1:0]          M_C_BA,
   output logic [1:0]          M_C_BG,
   output logic [0:0]          M_C_CKE,
   output logic [0:0]          M_C_ODT,
   output logic [0:0]          M_C_CS_N,
   output logic [0:0]          M_C_CLK_DN,
   output logic [0:0]          M_C_CLK_DP,
   output logic                RST_DIMM_C_N,
   output logic                M_C_PAR,
   inout [63:0]                M_C_DQ,
   inout [7:0]                 M_C_ECC,
   inout [17:0]                M_C_DQS_DP,
   inout [17:0]                M_C_DQS_DN,



   //----------------------------------------------
   // DDR stats
   //----------------------------------------------
   output logic[7:0]           sh_ddr_stat_addr[2:0],
   output logic[2:0]           sh_ddr_stat_wr,
   output logic[2:0]           sh_ddr_stat_rd,
   output logic[31:0]          sh_ddr_stat_wdata[2:0],

   input [2:0]                 ddr_sh_stat_ack,
   input [31:0]                ddr_sh_stat_rdata[2:0],
   input[7:0]                  ddr_sh_stat_int[2:0],

   input [5:0]                 cl_sh_ddr_awid,
   input [63:0]                cl_sh_ddr_awaddr,
   input [7:0]                 cl_sh_ddr_awlen,
   input                       cl_sh_ddr_awvalid,
   output logic                sh_cl_ddr_awready,

   input [5:0]                 cl_sh_ddr_wid,
   input [511:0]               cl_sh_ddr_wdata,
   input [63:0]                cl_sh_ddr_wstrb,
   input                       cl_sh_ddr_wlast,
   input                       cl_sh_ddr_wvalid,
   output logic                sh_cl_ddr_wready,

   output logic [5:0]          sh_cl_ddr_bid,
   output logic [1:0]          sh_cl_ddr_bresp,
   output logic                sh_cl_ddr_bvalid,
   input                       cl_sh_ddr_bready,

   input [5:0]                 cl_sh_ddr_arid,
   input [63:0]                cl_sh_ddr_araddr,
   input [7:0]                 cl_sh_ddr_arlen,
   input                       cl_sh_ddr_arvalid,
   output logic                sh_cl_ddr_arready,

   output logic [5:0]          sh_cl_ddr_rid,
   output logic [511:0]        sh_cl_ddr_rdata,
   output logic [1:0]          sh_cl_ddr_rresp,
   output logic                sh_cl_ddr_rlast,
   output logic                sh_cl_ddr_rvalid,
   input                       cl_sh_ddr_rready,

   output logic                sh_cl_ddr_is_ready,

   inout                       SYSMON_SCL,
   inout                       SYSMON_SDA,

   inout[3:0]                 fpga_uctrl_gpio

   //--------------------------------
   // Debug bridge
   //--------------------------------
`ifdef ENABLE_CS_DEBUG
   ,
   output drck,
   output shift,
   output tdi,
   output update,
   output sel,
   input logic tdo,
   output tms,
   output tck,
   output runtest,
   output reset,
   output capture,
   input logic[31:0] bscanid
`endif


`ifndef NO_CL_DDR
   ,
   output              sh_RST_DIMM_A_N,
   output              sh_RST_DIMM_B_N,
   output              sh_RST_DIMM_D_N
`endif  
                               
`ifdef I2C_SPI
   ,
   //--------------------------------------------------------  
   // I2C
   //--------------------------------------------------------  
   output logic [NUM_I2C-1:0]  i2c_scl_o,
   output logic [NUM_I2C-1:0]  i2c_scl_oe,
   input [NUM_I2C-1:0]         i2c_scl_i,

   output logic [NUM_I2C-1:0]  i2c_sda_o,
   output logic [NUM_I2C-1:0]  i2c_sda_oe,
   input [NUM_I2C-1:0]         i2c_sda_i,

   //--------------------------------------------------------  
   // SPI
   //--------------------------------------------------------  
   input                       spi_sck,
   output                      spi_miso,
   input                       spi_mosi,
   input                       spi_cs_n,
   output                      spi_int_n

`endif //  `ifdef I2C_SPI

`ifndef NO_XDMA_CL_IF
   ,

   //-----------------------------------------------
   // AXI-L interface to access XDMA configuration
   //-----------------------------------------------
   input [31:0] cl_sh_xdcfg_awaddr,

   input cl_sh_xdcfg_awvalid,
   output logic sh_cl_xdcfg_awready,
   input[31:0] cl_sh_xdcfg_wdata,
   input[3:0] cl_sh_xdcfg_wstrb,
   input cl_sh_xdcfg_wvalid,
   output logic sh_cl_xdcfg_wready,
   output logic sh_cl_xdcfg_bvalid,
   output logic[1:0] sh_cl_xdcfg_bresp,
   input cl_sh_xdcfg_bready,

   input[31:0] cl_sh_xdcfg_araddr,
   input cl_sh_xdcfg_arvalid,
   output logic sh_cl_xdcfg_arready,
   output logic[31:0] sh_cl_xdcfg_rdata,
   output logic[1:0] sh_cl_xdcfg_rresp,
   output logic sh_cl_xdcfg_rvalid,
   input cl_sh_xdcfg_rready,

   //----------------------------------------------------
   // XDMA AXI-4 interface to master cycles to CL
   //----------------------------------------------------
   output logic[4:0] sh_cl_xdma_awid,
   output logic[63:0] sh_cl_xdma_awaddr,
   output logic[7:0] sh_cl_xdma_awlen,
   output logic sh_cl_xdma_awvalid,
   input cl_sh_xdma_awready,

   output logic[511:0] sh_cl_xdma_wdata,
   output logic[63:0] sh_cl_xdma_wstrb,
   output logic sh_cl_xdma_wlast,
   output logic sh_cl_xdma_wvalid,
   input cl_sh_xdma_wready,

   input[4:0] cl_sh_xdma_bid,
   input[1:0] cl_sh_xdma_bresp,
   input cl_sh_xdma_bvalid,
   output logic sh_cl_xdma_bready,

   output logic[4:0] sh_cl_xdma_arid,
   output logic[63:0] sh_cl_xdma_araddr,
   output logic[7:0] sh_cl_xdma_arlen,
   output logic sh_cl_xdma_arvalid,
   input cl_sh_xdma_arready,

   input[4:0] cl_sh_xdma_rid,
   input[511:0] cl_sh_xdma_rdata,
   input[1:0] cl_sh_xdma_rresp,
   input cl_sh_xdma_rlast,
   input cl_sh_xdma_rvalid,
   output logic sh_cl_xdma_rready
`endif
    
  
   );


`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
oYBUgI3r2bm/BSj0c7tXVQyGSAILqEz5xnKrqeiiOWf23k2p0ql3mXu1a0z/XrXs5LO3rdjPKh31
lq9gHVE9EtE4ttV4AFGgTbHSKuzM+Af6yvJHzNuWuPOD9/19Cei51FUL5Zz9kdc3vT2vJmBNkSdM
GnguI4+aADZCV0goXYcUuE3Cfg4uMZdEgJv/YLBP1haQ6xHQh2cumgV3/hv8cQzkdKeSUpgvSgeX
BjBMkWEvH0wH0jxfQiod6ql6tLsppjAxRqhcslYxUwWZdV0+ma6Is6ZXw4OB8elYC6hFTNbbY2m/
rVwx9kD82FxpSO8THHHwQn7lP5qeXxjMaVOLUg==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
BwQGqgResJTCHQzan+PcNp9OAzvq6V9vms1lpu8Pt+R2mXsfaP2u1ezDNTcLXRfvBgt/4HcLrPwh
f+KXgNsRV9NuTboWyqYmR49nnGeNDII+84U7gt2abwt+3Gbab2iOshcnTjWHy8j3yMyIMkZ8pO1l
8/CS7nkfLzdZAQLOowU=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
mbey8MDNbRNimjRt+kcmcf3TG9OJ1qsmJnmNCCIYFb6xTy3R9LA6onjxkIcGPmVwh8oC+qCu5xwF
82t51BAvbuh0zLGrwqZro0IxTMeiivgzJs2MclLU3OYBB456psli9I6TIC2DYCqYBk9+c0DfHc8M
1+QhoD9MIeAlRuMIxe4=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 119104)
`pragma protect data_block
wFQgcsXgapQt2M5LKqZzPxYFYnAY8BOeW+a4SJRrPdEExQZIG/9NT1cpKGF6bYcs3KX19QQ+0pp6
/z2GkISe7sk4QQkZWZa4ObK+udhKvEIbIp0J9ZQpoUyN6ZtTVjdlX6PX/SthOU+AcFuv4+cdfM58
p88R4FWrujyzzV6tfjxTkeZwArR4JaFBrj66QPd62iuLEe9MzUKenzGkmvL3Fi9lQlQe9WwlnLxa
+8I25FFb6+5nbo37v5g3eiGNO5mZ/OTDZ3jwbBGPS86KGBhs1eczCUMLtbta1IzhJjRqv/39tmkZ
afXTatg6Qnjwu+SQQSPAcwiPOVv0CMCwwm4y9FaylzWJdTIY1i3VVpuNpNXtaMZ7cwCnLeDqXT4F
dTzsWmz3+YfEjCdSMwa4sWaBX4ds5cPmQ/2GUYNnr3kGiSaT8jIx0+epa+cCLlmmOyEmnXByF0Fe
inCnKwcN+mnEERh7vzxBMnuwPnwqBzJqpW41z6yfxfBvB4M0qxV0+KOl46EOaua1YyBCodmbhNvX
B+Ovu6XTNZXiVyNMoQ/ZC6DVKLITvloaFzc9mWU5+XKXeTfAyrOvm3XLbU3g6lMnJauS7ASG6/3C
GzoEly8PvThAosJhok48Jhs7y52Zsopr8o0et3DI6ZpmY75wEodbj9Oq4/F7XUN/l2qySmO8ijgI
OC4grLqBWfHC/fAi3TDMUXobUGV3EbT/01Kg+7Vnoszo8kuI3UJ2Tl+cSIzcc/hGKLeMa2z1hYIb
BmY6paU9jG/bfuCoqwcnNTxA5ByR2dWsQQMfSSfM2HMZDgIbHYa5sBlQN+K0ZWiU/uDbSEevgUV+
OAQjh+4Y4L+uNiQkVTU6io0XxyzVhnGcXb9niCGkqVo6cc7XPru51gn0TJd0LYqkZcQ7emjHP/UO
jdEe0FkFtjXnJ8Isa3h4iVt4Kn1kSU52jEFcRILSdP4vBU3FVqrxyORJ6xkqYp28slWvf2IzTUsE
/SHRUML9x7amIIqzJNUcn2rKVFlZDcix/bG7/hkhfyjyKiqqwRqDoj4SdzIYWUP1lLNWDXdPrh5v
tvLMM7+Hx2tB5c7txZQG6KGjxS88oHGtc4TpM79gCxJc0HrybhHml9VuRtnD/9w6cT/l2jKQ86re
xfwB/awIshb288hsLaoqoOwZeRKb/TSHip9VSiEOZg81sO9BYBwhvDQ84UYhrLqj+tFchNcDUdun
C8s66YKn7SH5L+c7e7r+nvi1Tr1sHb6CA6VZz6b7x2txDndlB4byYwlUwLStbj0TdEXl+Omfbq/7
C8Dg7mPZqBBDDWHZ8kxjgxw5bk/ux0fCr1BWmwXjgA6Z5Mj6a9lLqGdF8Rl9+pOrcIfB2i64bjaz
etMJFkWv/+yTDLVC/g2h5C6mTlRCZvha3QtrwyNWUfKKByhUASNl596uqGYLNfB1ISn7czTU8+vc
DPvbma3jYXAHEjryCO/g6tO0CNeDSLBEzuAFclzWpsDDDpPBKa6RJ738SWr0oz2UGKvsdCCoWCQV
pBfPws0H/IJV1fFWOjQPvjyd0j+6elAl2HC+773+DuvuWUjG+8fByQ44JvHvaycaaPwx9gkWEbO0
eU+3R+5hfCQLtTRM8vDLiP4R5rSGRBv80ZNo45yvAATt7ZWsHKvOnN7vQtTWLWU/6ekN6acBR69Y
gDGWupz7AjpbUHX76MYf0EEVUJ6HdInXn3QsNPALP7b5mRBfZNjdB7qhgrOBbC46nezUQDWP7d/P
BsSfrUAy7U77FfYXN8U/MPG28Li/pq/LWcGTzDP6lIz5tQdwHvslx7+G67DY7GarRnAP7aorU61h
AnBM68imC7VRphGDbQiHuh4mG5AVKywjsVVSRrdHhdPxSJPVHl8da5XQEjsF9YRPeBvit022WL3Y
juiiJuYrYFQLxyDHtwXaGQDya18pUi5HJtgW4F5YtmN9vFgx5RgZdKOBMrszJSH7mQRa9dqfnCpw
FxhRKDzcuUaGYnCAown1q7WMFSU0xhT+5MtHTn+TVfpk6I8tBU5JOOMY30atMkcFZKe3FYOXnAQ+
5bA7Tx5irVPPLRSWonn8QkI93XPfVhy+BOY33OteFz6tCa8On2je381+F5FOQqx3atjk0brvtfF5
L7q3qiNmfLxxlM+Hhie1at5MYbvQihEf0K3TeX4oNfbAWIhqLzHNA+kGrp0acV/SVxVlvgBqgFgT
BUEc87cYvl07rl9z/du25zOcxPkATDvMXrwmJtR3fCiHZXQ9SYhNzLCxe0OomIhcKo124Ch8CnV9
VToswXsqb6Gl6Cfm9M7T5lrjSZwJQ4I1vcwq3+XjGk6KIIPtKcCecJrhcU8qc/ijom0+jjM/2k87
buOkKOAy4MZS0raUXVWAP1pMNLGOwLCjooNYqLmhUhRVWH4o3s0N4ZfjP+te8zQ2cjnJlbJRzORd
hBYtRHjiLW9geaGHz8PYd8Rzij0Lt3rJxyumyJLy2co7tON5vNSH2xXrgTp1V5Mud8B4/43cPiYx
7iHjrZoDi+YQwkd6kqkXTOHRTaSUnG7wki9ad2dn1lpClubKonTZdFfzGbpKIX2b5feae3b2SoeF
DYzIbE7Oy2HYfpo/t+oAuhJ5iUwtO672hB48QXj5nABUQi84Gack0MbZI6U1SNww3dJy2Qp+GNJP
pO1XtTTtp+ggOH4PL5o94Y23LtbyvfRroBro+Uj1e8+6dHfwI1GyC2pmJshCrtxPzXI9GokA4aX4
smrKOs3QzhLHx5ekTdIBG0b/dQ28irlySPteowwdD3j4+a9DGH7qXC91w0F5TFMbgH3LRxjPTa3J
l9J1EC9HYWDMsOlmn7Pc/lf5fRFgSQxNOUHR91xvAmm0p6BP8Bf3787LNDSCkrKvzdfEVBTMAv6X
EP/mGbjnDMRtrErd0mggJrtAy2L9KIW9PYMasryr/mdE1+sxqiBHDSXRGdooRpq02C1tX/IGdoxb
d8HMftRQjelMIhEifjUa9vxA3NyeBmoPIN2qSykZa5SIjRHpl1SszHQ+LeQDkhdaVexsHdub/NkP
FN99NxygZ3ERPN0tTH52wz+xxu0wkUtfPuIw71EFPrC7TWgsomAE5Dw5UUwu/uQ9949pSiH8uYKz
XdYKoGinkqzHdRcqp/LjEjq8TL9CL/7YeeLV96owNcg64XWkGkn+GneOWOxfkDKg+NKjyTPhisPe
HPskfABBXokbvgOzXkbYoRy+HGnuOfjfslk6f4EOpxDHZYxYYlPkFYF2NDq88sNW7kGSM4pL/C86
PBhxwIKYfpfo3K6YTSCH8PV/BCwcMFNoEyD3PR/P+k6acnxBiELNTiHe4vlEUYrgZw3OLHpPxk5y
JpZLZ1GViXk8Rmv9xVuuRz1t9ECtNkilyADj8fc5BteIclwJkQG2Jo8KwJq6raSZCgy6EjLpS+wE
0UawXG0jipFWzMHYJSxLmdoWNsT08bDTq8SgKiA4PAhqINBaEViBdfpSAGC+hAsJvz73O/IcrrXP
j76JmuTLkWEryZzNiOxLhskt9BVAmrXcmvr7Rbo8+divsmIV517wogCBypTyHS8RiuDNdN25Q5oG
eNxA4i4QUD50FBOWcy43zQZkpg+K5EQ6J5+KUKXsSl/29ZMg2Jupd4mdn20jPKGy01uBL9PKfp3j
ddp4PyshaOilWDAICKSaHxnaRxJShWuQ90UmAxZdd8+vKOm4bi0aQBsSVkeUKotEBVfa81Ha3jpw
aO4hR/XQ6Dm2VOeFIeQ0Zi9hf36JxXYlgR30WwHnh54DMJv14odzj7LMcu8rVU8YdCv2hE55QMDU
VcBDJOtv109cIJn+Pj+Dexs2fRpIbIS+ugRYqi+SveZuHRQPDEoyxWJRaskqpCdE1taAMFzckrQN
u5GjU9r4mt9Bd7Q/QeM4GSA00pQZFXkvh4EEsrOdmfykPcrv0aITPIoWiDF1xS5Cbir+FklnobUC
r/WXbRfXQBOUAOzmG6aTfM8P+N6QRS4EfFymkmIjbFMi38b8hjeZEAxHI0VTRjJLU4gNc4CA/CQu
W/PhzqnBMiFkUEiRObkHYev5p6oQvw37a6rpm4rB+Ft2FbqMiLIGHkDDZXR3BZDGvj4RzIId+oYK
GK9UlPyoH/bfTy3QKqwlMmc7+CJyswoiSc1LnhBZRwLIcYSXK4NWjwWY4H6rJlEkiB5LvpZZx28+
pJlAxbXNAXXCFoemAu2zdnbqWxZGwhkRRkVQhQGkO60b4ohQSq+uJ3swac3cmKFg1dxGdFRJAqH0
lPtLa3a+QImj4Gli9bXTnSQgLWFFmYtNJ6gBWVFiUg+79zeOqUyFUiblOQq4OeIVJvtioyCiVhcU
jB6P5Xinof651CSg3kDqhePRV9shbo+gbn1tOU3NJh2hiy2Bct7aSKRBHVD5zH7CzHF6paVrDs7b
+vMRWH9MWefFXcBq9OOgMkOmiT2snTt2CUYaIizxO4YFEaukLTsvE5/lS6A5uvExgRf9xsa9W0sY
EpRu/lLQWGS5i4Mfl8a/RUM7PFDxjWEZ7z6fiPOXEeeqlUSd33ipc2mOs8WyaVX9SHBLfnCY/Zg0
qD5/GfwEjatOzl1yYU4TfDHNtVTGe8i6AJ8+CMUISG+UjgWFK16ZGIOQ/d3R1cugRfmPmF0+bD/R
9U4+doH6ML+crhpFR6DO2dBVeFNQ6h2DWq5J84pJ4qUWY1zfYtJyeihrFfLCPZjfYOdCpYjuz7Zy
0AtbA9OG9DGsnzz06MIg31sLhffsGn/TXz7ksTg0HEIFRXkN5pmNSRT8r1IjehBIdOw1ht+q9zaz
pdQVdjiGH17UsF2a6Toschoz4zf9xoqzPN2ihh13OKTO/QFPloRn3vn7fuQ+vugIXlgfJitwSxlW
uTbfD77TxW5hZ+uKu6a7cwPcjjIFAeYikXGzyfaz+gsRwvOW+wBNrkTbQ96IR2zx/EWvIhqgUR6x
66JuoNrgCfS3WQOCpYdizz8hHBb0Zs7shZEr0atq7t0eFJSPq6CdAIYFh7OOm9PzxOa3kDdDd3nh
Wq9qw4zsP89epmNCexJiSQiUbOF/qKkhz2tITZvz44miqVA6+OyMRmnlIbNtHR73gf5sxpWUenmh
M3Fnz4oHPfrMX+bdXBWJjiGIRBxjQ170iF29bkDiJQLfpQBW3jmn3zWnp4Z5FpQg8XIXPmeonrS/
A6FZ0v2JQNHt8GJUMBaKi8042rolROrhzZ9r64YZY53zLcK7kyaazkNJsHLSqAN0hO3T18AEDNYh
LIa5lMDnVeMkl4tQG5akWFVsg3lrha6brggnjc+u8dS2FqpgAhlF7w55A1fc2N8NcHEx2+srjX1g
q4wOkYPY5qAhvhf7w8FEC9yNdwL9ferzuJaypRKzxRUbvm1+oGIvahK/fdRlFUMBqzZ1nigq86Ym
Yq+v/9W1HKFuIVcUm2ruXWjsrzEQXioZAS7Mif86I7c23DqyLgD8M8fIu+VZ3ovKG4GLtajouZ1w
CRwamMP6NHfAkAbg+G4DNcZwv7TQvKo3NjvFeSA5i+KZTeZwqh+SO5ZGWaU3CFLmiwy8zfOuZWnw
oS4k4WXSZ39lkH/V0VxP61tENwiNYgAbMUJFfxNUm1VGtRHvYRmlMBUVFyE9Ck54Bw5vjrAM1qaO
kr2dVCdK5jhAG7PB0+DcrEQmSlzC+Z7ISCmCHwkWnCi99xQNL3nkFin507XNFCHo6MFuRJgyMVmk
m2ajYIEm0M+hDLkZj+o+9/HiZ7+RIaJphzoZKJmBaGDLb5uj3dkMQQfTBfXfkv9z3HDbgkEN2dZl
iurK1+x/fvltUuTs3KBjxywRGdE3PAUOVRZ2Hxo+1OK+tuqzJJOiUKxcBvZyfcKQe/jpdDaQ32r6
g3ATQoQcCt40msKYOfG/U4DMyX0PR2va/v5BBHCcTPcmDzfBYTZZpzkjGa/4LSzaIpMrLwpRTmpU
tieD78cy6yEBjPVGKGFlNFZpcXa0t2/ssCwlxuOqF+EvMD9ZaRXPL2CZSSS/2xHYQ6bnHeRUiOTe
lM7iRNDFjRAYqRPCkw+ngTUTbVQC5kCfQC+c5qM1suc4QJDX1ByghCKexkbiLfu5T4AEh3LUtsgZ
QszxO7KZs35QquCj911NTebE8zWvrTA3ZxSULPTRM63xg/sX6fboBWZb1NzG/2CIMOrTt6LsoJMS
faVCU1DBP0rDsKhkW2Q6BbVLG/vSDC7LnSGtz12hXuJqdeLfWYSNpnfUuE65tTJecPHd3UvHf9b1
ECLrRU83UyfeyUBv7/VA13ejYqBXu4bTQ8pWlXwji24hgvqs8+dSEgShcZm8y1yklM9DEut6kNPZ
FH4V31/CQi3Bd4rmjF/otGG/NkSXkxrRRiUhDkoLrEOkvFc+u9LHomAxRW3xMpee26Rk4mwofSF8
8F5LGuOpiIp3ggvnGM/iAADyNax+ourURfKzrhejhr5rAbtvgJ4QZlotcJiQ2dWdDJGvL6aMpdjz
yZlybnPzyW6uGGq0+m21OGwcFWwj3v3XbQpDbnbiNaJMRusHr3L0pEma+k+s0fgkJJtLULe+rea2
xzhA4quRJ6rXyAb4bsvFEmo4tIw8fmiiiS5/i4X5ZQq7lEIMzJdp02cFZTO2Zzn7i0dXW3gGIHcK
pQpF9e22pmm5aqnSJI/WUAznrSdh7m/xxZh5YqO2r5QRE3MuINuYfKYYNfnLu9hzd3DUl/XecWOa
AhCbpWYuzzpgY6bUqYH5be7x3iLPPkgbDHkXFprkZR+ZWZ5yIMuRPd2TvuxpRB/FQ4OQaP7gBiD3
7WpNdvqYrIpSbZTVENAwieb8YVIeQNKwtgicYnURhukdgfArWc4KhFyHpJ64wV07CY4V0n4h3Ojh
qOI0latYh1LYh3XbvIxHu1ciLjnx6o1U3oPMEOvBhuBuO0K69pjEtduegTcZcGlvM4PFS5UBJdW4
fPr/WUCxnJr3HNWfIE7+af1iiHVTHGZmKIm2kSg3mGZhFz30uuClhjfWj9H9b1+MV8Ybb4RTn0Hk
17WoY+krPqpIEqA2BIJoZ1hQY4fhrIEa1lzHKrDsQdp5f+VnC/ac4rg12JBuKuHRs6umdV8IYTBk
LAfEEkJILsexzGvb4C7Se4NaUEbhtODWulJnO77ddyaJc8GZRupTW//8RAU2lAhWtTbuDvSRsGSz
yhL7PZD2b5j/33od4CHVZOKFFlS3xNGIH2ARkehNK01JgfyCfK5SM9XHOoVIvfRoj8ro2O2UHoYt
H8Cs+ecEqxKxUcvJSQOZ523mKa5iWGuIw8VlJXMgy/ZFcKGsJo5cQseM+DiyS/ss4N0+C2r1GW/k
2uw1kftV9VbUZlKVW/fwnoRx728VzoVe/9O3BMk+OxlBqva8kcWw0dPBqEGxy4gBqqa/lJrgXnOl
QZe+h5tYn+U7KA8/QhL5xwY1FsBrpPAGQF+wyKAHrSJ5kPZhde/dLj2nIFbSzCJaNrRnECFoWust
41uOK1ODF4Yr01Ulv2a7XaAVee5xwyBskTbb+r4M2gcOhAKJrD6kAy7kP2h0f5mhfStNi+nW5cgF
3dUkzlq5/SPs2fqoSh9KywAeAt3NdU3fBzjcFr1txGopfR38d5zShuSmkl8CYhF/JUJOJSRo1qKt
aVomkIY10pX8ZKy5Qo0vd21berVivmfSxqXUmIuo1JzknjPHMYfdylKBgp9agOVN5732FpUn4KNn
U0+1n3rojsHG9T7JSSQPCOORMSmTLLh3GN4UHk3ZX6AztQgacl15zEHcyKNevdkUnj4wPzU2KGL1
y4L9UBp0mclaY0Gou/Vzn07Ee4E8m+t4EBK/CDy9qQZmvmCq3dHoURGi0lWg1ZaGxIlpveD+bTvv
y90Ka1dEuKP87Rnx9FvhGO0JQH97QrplGDHJXpn7Tr/MNmRjtI9qjY347nvWy1oUg6rvBv/y/UOZ
7CfQgLoO0FIcgJAPfHJ5DtY0f3QHkWRHNEvCLiy6AatsSNPuyvnBo3LglEDqEnW3/dpwZn3nOjFp
z66l6W9gMAJfkpmXhXZ4xgBlSV89ogYhep0g/JZQpGeXfVoBA7adUbN33mitloBYihy4TPiNhOGj
6KodQcG6cx/JOjrOLctLAci34f+CnTHtyQvRM7eoXJ8ozVoHf/a5DWe6leI+Ax5hapxRwHNrTbzx
+A8tb0KHUNZQgLje103rwLXTNZNK1ASwTnltdtTPxqc81UuyypDl3KzB9oSwR/GZy+hYWRd5/rvw
NCKAILYxnkeNFlKjTa1dxHarG7DA/n04KN+OCz7z3N0L3OVFGYQzed0gsMdK8AXU7LxO+GXW+TVn
NKPG7WxGOrzZyGn/ow+fynbXT70HV+WwZIgrkKXKTirS75GdzfgbGLYnmdy1ndLZMwAlKPotcVJi
WAliqyx4BJ81/tOd5atOzNBuEiQeKdr4yNwQC93IIQazZK+SAvgY2W46aGM9Xev3WiCmJ0TXzd25
YsK79qreSYwG4GJt8mPb09rLtDBTwU/8JTS2v++zyw4bmGtAkfXOvHhPevLStjrhHn9RXeymhCY+
Q6IFwSxc5BhalN7rPXzfXE5gwJmxMbuZwrJirahLAmoAun9V9rICADpF0KMsQxAEWHaBYPtba4PY
GwxCM3XRuPKesTxq24Hpx8pZd2psMxRs0YsbGcZ/hNte9AxVFk3K97Kl0GPdNMFQtAkXj0RN89Ew
uLWa5xdIMa1rrHHhgqGwXPTWsL5LoVEzl33bE4BDe/cIwvKdq/08BfExP7ZTA2Q1b1Ga+V6uOKA7
EGHoagokg/U1isn3wD9wDGLJ91OB5K6fOslTtSFZofQ/OUfCRwvacLDwVv6kVhVslA53VLbiDS+H
G7gHuAB8P4oBvD0gBrbWgKNPeFfMuuTRljQWSlmpAB4tK7AdTYJNuXLAJP8/JDSg/rd2bFoJQawi
wLTbVgwUbFhyJqnDHwwPAWZKVHGEP3GJkEk5WBZVjuTzh4KR51Vv7CdvC+Ec03DT+mI4Nl0SwwtY
P4GtwXTgQLUuS7AmpqgFwr+aSVYfasvQMo+LqYgLbQXH3oyw4kqryCssRUZ56UQFaFl4pmhkXe5w
v1IHwPd9r7E9+tMN3kk1e6YTnYy59lahNxozYf9Yd01e2jvmcny7NwZO+WbOfLimjljekVGUB/JL
ZhQo1eOiNWPbCXvqUSDN4PpXrQZwDF1OJJqpFoGg0DNZOkqtn+6ii4KihiHnp6EvSxI4WeQGWHze
kGo07akbnqIvd44Vg+e1zBZ/8Zv1rtn5mRBYKozbeNpltKtr7QSrR+d84MnlShZmdmsJF5NhvJRw
noR6yn0P+Pw3n8mp7nqseCVBxvuSNTnEipEoeYejbJHp17R6doVjB7HrdgIJXYQF8DavVoWV9t9X
YcTn2oyNhlJknA4cfbd82iTL9m78jWX3GH9nSwZUe+F0nUwbQD2pSyT2COGdWyOwXZ4yZPUkONrz
OYczoK+es2I8q/a9zXOOm9OzFnympjxY7zcqC/5+Yi4f4wW878ibxytW7am2dPWGL/Ilo7brqETw
eBwr8sCDlIF1VVfR84pglP4PKrcON8RBzqAnwk8Gz2p+URZ0qTwEmTvGSfjgEf/hMMckvsF183zD
iVvSXVRYb5QkHYvHowGw4YUs52QCvOG2BT/7EkxyKtiUc/8L7DERXS3NxkxWo/RRtEtbHClq472N
W0KOyp4K0tnha9i223p8EBH2+Gbr607j816/HJ1NmmwbFAGY04DSW2ok3Kmw/Fx4Su2WHchgvJXn
uWrsYPnnmr6nJm7Cf0lVxOpdM7Nh/BELXL10WmiX4bxaONpU+5Deskml1Dx/qR0ASq33iH6REJ7x
++cUnmr39FZpMwQr+O6fCI3KWRPzBImzRToky+FX833ca8DJKKidq8qSMBQnPSpOVA6I4uqvHUre
KjAb0UZ2J3n84kjPmRCn//Zvhw6qBZ7CI3Utn+Pv7HQZVwadt+omOVOMcDeeC0YYrQtWrBEGNaAr
1GuI9slT/7FCzgSeGjvU+bYPNkLUT+RsmcceIbhsr1L/AhbFA3eIAWS8NASX1zA9YTIm5RNZ3SsO
xaLeK6T8+A0zpzcz/Vbt0yIpstzhhiyFjQWK/FqrXjAPmeAX5FKjtPmR0Kqkxpou2PFTDWNqWSkA
4cU8skWKJt65hBAx8wx8/te0NL/mTseZhbz5x7+iPY28LvwfAlJiuBkHd66UJEYpSRWvYOUoQ0am
FK/Ijyx1hQB53HymrZKh32q0Djxyg3fP47plAkJdIjgq8chG3G7VJEv5MAvcdPpAHkpUDvk+1LMv
ikOabzvSDanpWmIjUcvReYkQlDChhuQXxoAxe56lXAUOhbIewwfHyPm5ARxNTl9QjGwGXJIsgv6n
4AvClzS9DnzkMmMTPwO+R01MLaSyGNys7/9oxV6h1huTt9nY6eXGhevqXGZdg159DsiPrQ+HLp1U
4/7G4nJSo2yKvhsy8FEQWKbYYSjHe83ZltDPLkl9E0DoyA1VZKAtXHgGlc0n4Q6TmfYapj7hGBgQ
gBkVFzcZ1mXg46suXxj9vFBso6TH1q/c6PXI2iqRzzGmzIlVdXwgtdgkSEFhokIxvpcq29ef841f
qqV/XL9csT30W0vl1UO47MGXZQKRkBm/fLa80xjacNWqFTwc20mPm/sdUcQb9Rj9Wcrb2miEDW50
24+QLSC7POo9khcHHXRrdF8sgFlbXE22kloO+6QLmHoFyX8wMV3M3KRv2vp0YJhN2/M5ye2m1lRw
yqTuIzlxNiJsLQgPEQxQzae/yXRWwUY3SE+jyqvlIzunfgefQg11dierhx5xoEwEnm0tKF94JHcy
AtRtkRYrs4PsRKwk2JsJLloQYOK1HWLr4aN/5KiornMa+OgDkdrOX/0PG4F0x12F1Jkbzzraof1t
t4CnrydtFcRX1X67OwjwFRb1MJZ6eJXtTp728t6kG3YenCCDXBOoQ/+DqSgM+Hgm1xBScFhRGYi8
ql0dAUHz40B6Z4oVNMewl+pKSDBPdHB6GMskEbV8KNFxP0WKkdBMm1ZGK4rX0nWY7RDsZl7z9ywP
lewRwVartzz0fhTLkeXniLwCP2ol4uBsBgBsUjwe47GutWnQEbUuiNmpfyzM+ic729qHyMKCR/Cp
FC9VOzBAYpPIgbWledYy6/VuXDIczBTndDVwF0p4Nv1NQUfWLuqT1CkgcOEUfpzERaARKgTEMXwT
gxNfe90DEcb3tzo0LT+SPoykfGJemwb2wtzyx3UtbWVaQtf7pqfoc2AGxjKNGr0iSdlCatCQnVQ8
czDY+GCYH/sUIakjOgoMMw3wQloo93d6t+XNdiyoFJUVOIkoG7Ydm+eAHFhLwijOMrMKGXOb0ZbV
BlOspFk6FQjLGvjbImDm8Ty1R/BQ33+OntjJRPslKJiZ8Nr/l0unksNLhNAPeLKzVO2qCUqWZ4jH
wlPqE2iFMQpCQc5ZnVv3Wo8B8PKeIu9emBPIUlpAqckB5PVWpPfdVzaUz+rblC4geTVN+D6SzfgL
4M70ghtL+pGo/t+zAEFMJ6E4agmJMlcDyIsN8a6siXYhgo9n+ODQmxpK32YblIQ42YL7gvbSeVsQ
c4aDp4o0h+/awbKbV4OgjC/McU4EZrXgjSP7pr+i//8A0rY6ETMfAVSVn4XbA5QbsmTeZ/dvK2mS
GrBMyMnBpIgYUCKHagRz/ctcBEAGQMQbRY9qft1EG293s5CKuA/9quz45boQTRDQedQyBFZ/2ro2
r5GUaiSWHOPid/xbnfbWVN5SNiVNWT/C5mhkVxqTodLeT3la4IWOHxpj7xsYmffYsKVegkh2a1ch
B96t8ZgvPfbku9UXMRNLYQJmIg4W/nigFjsx4TdTVKMNSoR+g5GVD7FoPEkUZtfOXaqWMfEijOn8
t6oQ7bLYqnG+y4HU1QYgnYLGpM3+v+A5PfH5taX4dc/t22pMSWP32mXry1YtjLKQ/rMah09ChtlW
5qSUwaZdajBxHoJDthraA7R3rW5sUIM6jQr8pP4Ta1Pek7o//E2rcuA5GQ6dpVX89Rxr0Ad2vWuu
12esuREscVapAa3drQKF+9hzrBHZFG8JN/sKht4Scf8wJMfHAnoiIyd9WsvJq18egKNe1bRSpSu+
rPs3sw/obIaqT1+978bKJLDMP1OVZzWpyoHgKs5uxC8uY6kx18e80nVqz3vvlXonvrc1Sj+BU5r4
+c9dDfyQM53Hrljzvs84xm11O36NDu8mVbd4mVyDw9wCnSpb1C4fuF8tYVvjuqmTM6fnmZyiTETJ
wyvcbnxXgIG4ro9KuCjw3rUwsFdI/dg9dd0LlsmQKB8XP/qn5oByzGGJtdG7tHjHHaml1G1FVaOW
krbBdR7PFlNek1J2oSbuaVxHTR76/sJTtOW5QW47jnqDUq1j5ByZBmfmzNkAH3T/lgp8HnAve1g5
457oXt11W//kjQAnbUvHj+0JPqkfTEoJ3JIViWOsyKyZVsciDz9vajYgueIVJXH1c1kHGT4jagx0
Pom9bzoEeH3jES4hgx/znEZcqvVwgA0ovW3BkOk+nknbVAij0eClRtBM4SNbZ3NKRzM3m9aN3a8r
obJvBnMmZnsGwlh+MFjSgGaECiDRw8hiaiMp/iCtEyvDodRI35CtNGe7Bgcvgk/Y/Cc8o0dcNeRU
YX0S7gM6ajZe5rROyeGRdRj2ZMvqE8YJ528uhcYJ2a+CWSYdX0zk4BA4JNODYfLlOqRuVOSErAhy
JogEEFKuxWvnWTzKqjsp3DnPtp35SULFDkg6WwYoflySdt1GRW6bOALrR7+7oqPc97nnjx4TH+K0
EKC3B3j8YWOfNQAWDjhXyKRPSCcIuUbYkrBlso17+3ykTZ7F+SyVjP3Q7v1VMKpp9esuFpuHG2vA
qVdBG4Jki1AtWS8x30G9/bBrdEHlTfWSu1D1Z6xiK/TJrv3tfGl3ydTWTUlDIFxg6I2tEj0nwlOK
QNRj/ruaAGuLvOZdT5DcbQDLbAaJ9ZJgehwi+MWJTxlopPjpuN7rJZh/pqCLpeEyAffev3GP4ylH
0WDqHXZ36TL3Bv8C/BBsJ/4t5lRiGq3Jyhv5HRZGXysJijLyKoBhO7nqshCsOjri9y3DnIhlqBkH
xfHOHm3Wq84q1H3L6ZB6kVlxMVjS/syYwmtAX059Tpi9mPzQ+6GtCPGE9CAFA9XKNPXH+GzUuZnJ
vSmUq6fScOUF6JT8OvrGvR0jiSQKYQTRqK80h+bla3LNqV5LLHf8KR8RlqZDWund7C257mTgVLgH
vL34iEkOtEeZBLnGVw1qXWKv4jOrTlauE21Oh1LJzCJw0IHuRmYfFt8vza6LqVQ1LpVORjBil0G4
8EaPhMbTmoJ43B37Se65k0N2x811wy1zUZ3yU57R8DIaObo5R0xVILekqA2USpCT1ZNrXiTA/9O6
eAqK1uhCWLCF0D0nW1t3777UtTJPdnGSmaNMGvXAULcr9LB8z+5fmPgyiGT24kTrmHN4ePyOb+qt
GRiR2hdpvkhZeMWjYbXy7KyiC/CkIwZolbz3obnRYow5QvHGtSDOijGv1oFJnHwyHZukAccOqA3B
3mAbLifnDc8DZGbW0Z6yeVdz3wb8H/K1JgxZI9qbui3lis02TKauPfsg+7s/3jdyHwce1s8SyRKH
Akmiag5fbuLAePVVoEKBR2ejBhbRL8rQqUByTRy/Ofa0Y652ucYDmAzLZZWcP7YTEJ5AlZF1o6b5
Ej0Z3srzy0XOieCgoR0asWEm6UFospUdqT/j0UxCKVNeXwBTZTad1H0GkTgdT7ySIA9EtMjrXQ4i
xZW4msuWo2ubYjdusHoqn+oZqRWLFZziiVkO1rg9jUxRz67r6xpn3VMtXBGu3awJMtIeRVGQ1+ge
MHfDNV2LJXyrfBYzgKNpx66L95Nl9flRHWPbGIbHY8KlepvFg3upzvQMflrBfTqvrJyD6tdhyhJC
WQVwRfboiiH55RhqTIuINZPmF7QQ1ael301Ay5b4ORvneZ7Kdn+/qYQKHMsky8OZsp2lMP856phb
Lc+RgOok3x/tdZKrRsTG4lGxfiTcnuWSsoy5G60rwfvBPQZ2X5ZHVuby//O2Jq4mTYfpvWMsoo93
m6J00mIs04KTGA3nzTRAR/gUViruJdFZhEZoF/fSSMLet0EuP7e4oH9lK012oaQ0Rb5gN74Ridjn
1BZ5upxPhpx5Ha3/H5Wfi7NJ/SexN6mzkFLdkIgtmTsLjAdTWafcbwnVTa1M8Ix7dSVlOBiX4yYp
eUYq2qKST1EMkmrs+qeEFI/wcRFVEyXXN1ET1VpKhwHH+0DemfzG1cieZ/dgJvf3NPevReaMYCxc
KWoJXAIYqpPyTAIjMa+CaTebLnZMSQjkMu0B66Bv904nRAXQSwHrZbFY3i71pWG/N6dT9O34JNyG
2LIcqIlTL+CfnzOKzkwxs2r+BxskgKX33YnK/BUg/87v7JCPhQVZNlFdVlT5K28WwOA4y5qOLLy2
mt5+KOeLK90uq+9OknEYj+VvRRVyogO7lp/OqJjBkkEGH04vK/wMzfhXkQ7Lt8P6S46RTzY3+0Yr
G8mg5Ng9KPTM+0xzYGhPhKp241ZqxW+kPGW2w3zhbv2IaOvnFiY6fX4pomHc3p6FSPoE1xHFPRiB
qGRkxIrQY5BOGVU1Efg5IBuRC3maVecJHFzW+Cptj88sYOFfLd+5MS4l63clgconu+99XUr1xVtA
HOYwJr1HfVJ7h78G1cxAcpbg7XNrEGd+31vNriUAP4HnbLLRkUppuDFO0QhlPmYPHnf7RtGbGOYN
OJcZCYk5kTsN6Dz4ItqwzHXc6JblkZGOAG0sMoC5HPpWVazo1poFPRVUk4apTsrLMm5VCZrPgJug
42EVcMVbWk8DIkKzDRegZX+CiEqgz3ItCMgHEYIlTECgFYPwneUAZl2ImJtyoZ6EX0f5Zha+5zNV
tOjS6tviNJhEgLgdwsVXXb1HTfxCetTv0pPS9uURnt0wl54ny8VkFQDcr6GHHpeTlo8wyzlC6AhC
/fnPpIwHynJCvUPL+XOgj4IWmD4/gC6jWUO5oSXQnYLuVvE+UN6uQo6iRaPMspCmZ7yT1EdcjHSf
cB9apCBNNJ+FQ90HT6vhYZzk/yCFNpo94Gt9u08QMsQJBlMmMTk42ODDvFfQX78x6MhPritJs3dQ
2BA9KWCk6h9he50qjPXlzehtzZ3Mmsvt0QW4xhhavXOrU6mptZh6NKJsDbmQ0+93QJuVPm1KxmYo
QfeMaGRIX4lbGZCdR+d/VJvgdPisk99XhiOEwndzubFKHoTXZkVmNt20P7SWN0cpY5Uro30QR6l+
IDjkhIXbIXqCWgNTzPqWH0W6JoPYXXUraYk04qg367JF15a6SjjFjQSZNuZMpjA0bgTBdQtge/WM
SReRIrSZkWTI83VMZliuOZYMCBjxW+pFkm6zoNJ3ENj3eO/xu9ylcLs89IDcnxjvtjN3ZiWXNnoA
UVaK5EOzqynwF/PlH0k/par9QCwrjS6LLTOJZ0bv8fBdvVqFOJqCU5Lg13hQJyjFQI9Qqol9rbmK
CpBsmUYAesGWYZKfTXE26wX5apXdMF1ywcpDw/CUlU7zviT9UxJDejdrYVITaMRZxsNyfwokpCDo
0S2b5fhYHqvYvuaJ2hPJ/4R0XiO03dYzWyfS3fGoS7nsWlzvp7aiI+zn8O2fQfV4CvgRvOgZedTA
3ug+LdMCCo5SwfovlGeEfBM5kPzJUhvNBQtrKFYOpgh/brzoun02cxRH6V7D0/QBN/+lqhrDbsu6
pUfCNg7oV3zA5gAeg7a6Xvw8qTf5S2+rCdH0n00udmXdVjbQGlDNsw0E37yigGYnH0JJlB/5j/3Q
BiEL90zF/+MWcMqkDWGDeHcUNKnpdLyAu+YR4PIsf4Vld+3Y+/eh3/nJdWsoREw1eLU4bVgMIQJM
w3pzeGGB/bT24ERpPV+P+9MGN4Ga9pHiDgPb/QpC7RObPQ5ObYxoSYYJl7d0jwTqLXXAs6ufS4P8
+kap15HPzZnXpg56HAsSknqVyqU4KMyuSB1VxjUa6ExHPjOY9+OXkq5hZstOb70LOdDIiNxJjyaX
Gxde0w347aIuA+T3DW7Fsn4g7Ob+si+0Dy+YgJacfETgEOedFMQpHwMLMaE4N0aXm/0puV8iy061
4xjij0kqRHVRp3+2eKzsXAXGKzUu3XX+/Rn+3HrvTQWeYbQ+dut3BF9qnH8g1rVa7VyEUMqXv2fT
BsgNgj9t/Oz/TE8L0nEqb0kwIJW5moeo4gQAqVmg4kr83GbhJK0AYA268/QOe1FEVSJFNapqBhHR
Nqtrmzm7153gQW+frhdYWyDkFsigI+DX/8cwXWAIWiJIxknnDi69LMk4OGv0xL3MWxrxryzp1uIX
FVNRKl/vvrhzbipxAcParO308n3+KUTJHt8ibRyC0v3ulp5tWrw22Hl9VsR33xlKDpG8WkK7UGP5
FufT8qabUHriVbrx2QU2J2glHYUkFX0fFeTZUayzHelrGHbX2mdjp1Rfzxh+aMwuN3VKJnRdgc1Q
V8LLEmxlJUC4ZcbRGLGm3h6G/uq1IAAvNpJdojtOH0KsdoQOUVxhPqJM/WU63VeD+b1Qt+EIlSBR
LWsGTB00CCYytCDtpd+zIQ2Oh18gASoaJM08ge2q19uV9xR/3x+Gu6M7kV3LDBtjokK6YEq+Nk4T
LimDdn0B3rwhIBDpZACkwPseaCrYhB1rgjxDiwDjTcFEJ1RNlZiQ13KEpHMtnSa19c1fo4RjAtg4
9dueX2wi/9suXDx2Q9vs2+jogDVdCxnLL4tUmOHya4b4JssrQLZ7v25+5acrLvkMEbXt5rNFSfeZ
cdUk0VC8QTrFjtNlhsYP0Pi0zkBjvwkq2LZ6BEsyQ2IgOZxOWFhiTSSJPjjHzrKMNwzEhR7Urs04
6TBlOZvpNt6StkoIsy6OVuO1XY7PZh7ZW6zNt+HXZYCE4TTM05JHDJSI0xAarof3E3wKHVDQwTCa
2z3c6y3kR60B7aUcim4labSEEJU4r2ykni4+M74BV0KGW2ZrBzHYODD2H9BBp+j2a22QICgOnv1c
9BZ5lFwpkPO1FbTkqAoFsuiEklaO6/DTWUO7FkJrv+K91xEQjSTWRMjnXElagdcHNEsiVckD5pgj
fE4ycoOsz+dcZHRQm8X43Bd4W7kYnJX63c0m7m9U9IGJLtpr9Jee5vpWTl61r/XYiiIjTNLilH96
+y+DMkCjDgJrISk52rHGcXIym3obe9yAxwGMphfo/Xz/sQ7Ul23xG9QNpAZ0g7sCDjE+2EdIuakN
Av40ZS6NCruQsbE1NFuBY1kxhqOHkhcEJ1PD08Chd77uWHitPyR+58+x5CUvsN0XEJXS9NWlpa48
35Mvk5czbQ+bS/BVsJHKG4C+CCmRsTMxXSIn8e4g5lcKKqS+RssOxh0XDcAZij8WINRbcUq0ARfM
IhwdzgL05zVz/OKoktIJD70wQMt5wSdLWstlqsBHCdKsL7pnW0tJngUfKo1S7u2UcaAmi5vRgeo9
CWRkbP3xFQf+5aSxWDwS3LJswB53o36ZKtmmIunVNzgycmT2aLS2/9ltsfmBt7ctTRGKR7CdB3Es
BZtYoQJVTp552+1ZWfyirLwrAe/J/i3Fe2yQzpCDeu95bZgng11PLbvvvY1K6DHc1DoyU/Mb1/bc
9mhUAkW09AeNgTmfS3sWpCcbpeSiL+gnlECIDh4kUAjjuLY0icF7e4NanrYFl2bTGqQPk8bgV/H2
Pf9om2ZI3FSjbuKsj3ypxZBCTNGwVWwtTSZvWjABkivbnQWgZE4BxFiwODEoptWdDBfeHkGs0qDU
9kVAIMP/v3Iw4mrMlLHxAS2cSqrNfD9Etkw5EAdvMz+UtSMJmf1EGhFeZ5zEsmRFvrIiaJM0ZLpd
MlIj8yluMJKKEWwqwQU9h0eDZ3xucn8QbelZ72gtjRcL1vwFgxeS7nAM2dey1DHNm9Nh7aguXQrX
MvdrLltE6hpYNU2uMTG0OF9QYeddUKxlWgnW0W13MnG1H15LMD6WWRNl8i7foSThCykPxojYR3vg
Qt9gtGinSQETll+oQ9uF/14I7e24bNI15MrT+fHRVnyYvU7DIC+lbvaPc3pxQdEVZoMjv4to+QMb
vmlFf7jHWSOdDzhAJWaiAUSm3o1RdCya/ku8kNLZASxtlsUn6MQ2EVP/Fy4ebvHQ/rSFHlbZ+eX9
u4dXmziNFrUkd27hE6AvYr7LG8nJFXUVV6mPeeh/hbKL7k3y1UEGqcuJ4LUJVnDqV/52beLviBa0
ZdtnSsmyHcJH9vNZ0vRa2oeDX+Cpb7KLPFFRpzbOSu9+PIsulSsBbh1yVsG5aw82lM25mOvLn0Jh
eUdLU1OoVpj3Lvvazhi64urblYscwxHDbx4DizuE0YB9salcwzudedxrKJEPIsT0NUdab0ZsqXwk
EthSFJXZiRXl7eZUmuE19fQGirF/O1RWGxVaOisSXBMrETlJsskIBD2a93ZtzajDl95jX4SogVeD
HGVnBuPHIIKHWVDC/+wM+JsB4Nb2JqvawhGEarfrqiiga0CQDp0CyxcRWvxxpYfQvRJOzqN/gaLj
y3tLrk0bEmjGFDq2EEn/1kJw+4bEYlOV71W63GHpdihryMwx5qMjM+QuOy8VTU8U/oTO0C73M/7P
IQ1d7MtBec2HtWoR/9ctCyUXcVgUcNt52ZdDVF2DCjAz+ZrBF78xF2JYsqXiltU5uKTBiecd0Tz4
qYKNHV/VJ5yHpbvxapIvohFnnY5zJmnpgPOieiUw7GOtlzOBgTz8G5EpsAHhrHsngjb9oKCo9HVT
wt/x66K0jw9NiqIXFTUWnGvKXLuWXO09LmOKr3fzvdsruk4lx/hckw9ICZfllhlIKphHzw4fHfJY
EKzWVkcL8kcrBpeLmXfACaHjoKQ2fU1VFF9mYymN5cJOQD1C4wMBUR8PPb8Juz23RLT7ol5Xjuzf
/VSwmCbIixKbRhfl7KW6vOpf8TQsonx9kam39/bMfi9QS+dp5JBLiex1cq9LkMTdc0vOouhCrzbG
FsxTbgO9BBbwohRNApEWNjuJETWQrf7DSPq1/eN/rorHCX3afg7IAv2D3i2ZqXA7qe5mRV27vw97
683ha20IgPjlN9n0qoaaTBua9W0HbHux394WauqvLHyMhx754ks/0sql/pYoONNU621HhsXL/NPE
iB/Yeh5wEIblgeXP2RFOAQzaJjFeTBrvDiVUjN1wEbe6juD1voThoEiFS/+OZW/4kqUS9INFuZLl
fgti9o+a19p+Okb2vBXbNoiMIVSKW9nMLqiFfJiUKwDLY4k2/7Npa3TCSehs2B4O7c6++U/DYznx
6+m45ml3MFMwJqSb01EdU+AiXK4Ysc4MCXLHlsNa1ok4LTOds8pE5CMnPPNo5vStlcdqaYHx1Xf7
hB0ALUh/D86to1roxK3T642Q5a5R0Sd5my3MdFr95eCUuAFAzOPensdY3OdpmEkoyD92l5Uf/jBu
nE1l+EAglFALba7wHI05a1K54NOTbbS6XgYgc1FBWv1WG+lPd4s/cEezpO9WLsDybu2oyIPlcL6v
NtCzs+/oszKxnvmLkXRBrtP7vqT25rmVaCMRfkz0KSXvjmH7MV1pCtIyS+TpKEI2ncQ0s6VEHaP8
XVd5oZR5yzYP1xfFM801sbun4B2dmrIZ87evkcbObdhYWh1vzzFqCcOHFqGxGezx5vjAtfB9YGPV
aeN4CFtDLtN4zngeb+2RIQcTcYZKfNB9ndC4ghv/fxbgnL1aU3ZtaY/UyY3KlhxLKGs9sUt5TrTc
IEkTT54PVxT1BypLDW2prktfu6bfwf67b/tvUNZNJVEyH3F4rM7unsMGWgA6YO4YbsvEX/bFvA48
n+1eZNPSMe5agYSa6RbOByTaKHwsi/63HdL4vlFyvHplwbY5DZPRKaUVUPevBbWWPbKW9G7N/uf2
oikwyyZu7+H3eV3riqRpQ6cbbqr54Ymi+6rnovR2W8qvkuu5PwZg8wWH1kyWIVxhG0mzbdx3j7+2
3rz/6gZeyTfHqaVqLVNqYA8923IgcjCWNPEXZmiL7fq7LZYcZWi+YMxq6UC44yyRoHk4DmXOKmIz
ApPNM+xwL3vLUlt/6craK+U5EuAgfbqw7rFMqg1m85nCyPFEXiluPGO+/ELeXBYMnqPYVyv/lvtU
dhMdj5pBi1ZDTdPYFJ/QZiLxVnH1pLjwEz0i26Wr0ehlD9dJl3wdE4UMWc9+aVbzlZxelQoJy03y
2zOh+Eb6Rtuqf/BC6W94QM4Qd1gnfXf7JtF+LhlZrlRJB2CX7wdKCQWOAGnUQrSGkCBEk8V/u6y8
xD7y7Rne2hEKpNJdMkPTZAtinczGg+IlC1U7u0xV4xVPYQRSiVBKbrOGcefawG2fFXPcWAkaW4Cp
/tHZ1ohFZdf9hP5qvfzGcAkU5xu8hnTS1se4biRURNRMALy034lHeIksuLmL5pSq/3FsxV0Fop44
zPyEKlI1O2MjLUDD5DVzrjZvz6qsCKvCJO5eU1C30C5uUBGDd3VpC02UhBbNTeB259wFrv9G5Byh
oPFci7ZmuZXc7tLMfSmZ3kq16u2+hIne3R0aVeSnkahmBRlA8wJsqT9tyF7HZw7PClDwfZjpYIax
x8UTGIec1Yf8yOAv0wMhQGy+W78Cv2SqBp/RYs3Ax3v52Nrq4XDosqd0wTQLnbZ0EBwih2B8IbzZ
HgZmqa2GPJ/unAHmAIB1MvUfBr/Lw49CHD7njv1TFIzYPPRzjxDv7uwNnpjT0tub16ijYqLnwH1l
E6Zxx4eALuyE5I+Lw24/M3wr996CdqBjcMHiVTJx5jdco5iCLPy7k8ojAByPFNLGUSymJkYXPw6q
ug/SGoyFt4HO8NsTeSv9CR6/ZQrthqeDkwBVjA+8QuawDQzpToDkspJ/goKX2zs7u6K6+miU2UvF
YP+JcPYlnAIjlR2KRE4pVmcMZzp85y6SrNGLW1TEOtDuBDNTx0P3hgSU22vT3A5ldt4xBLQORfcW
aHot96KsGgUDDw1NdAKyx8BbggxuTN0+a772ZezW5NC9FCiE9YepzaIA1CZsKuXKQ1v2wDW8/XPQ
ZEE8Aq7cNQxMNf41WAUMensMWcvlkBLKoA7bLkko/EKNzR5NBSLHIvDJJiL0rphwRFeTtOd2LFYk
3FL1F/uBq3oLkuc6PRfK9Wt0/2NTwSyXDN1YACoJi4A+5tTKWh25dKfX4f2PlymDSFe6agb4jfV0
jx/aX6Z+o+sUteFtAGe8ROh7DWgKx65JKdHiBquqHeE+y9ysdIA14To0rfWyHJysa/lKInmnjsbw
rTHJtOATEapx2NyzaksZcWMUW5OTXOUHFrb8AwHdAMnKMLTXiFf3+ehW7uv2m3sk7fGM/oUtWGsH
FyJd2kKUrHwldr3qZ7I9qXcec0jYnQQ7ObsoA1ehnZ33rqJkVKJ1MdJDKwMcmIeE0roZ9G5CWYgx
TmMutGRRY5PmrkvR4Za/We5+YWO/+B4NlYx+LalVJF/TbOkjTZGoR5KA91y2NZnf/8Wabb5v3lKE
yLtJzYExJ8MU0Y02KjE5R+FxI7PTnn6pGCrcq1nf6Ipory0z6QbpsHjsq1caDZ5g1nEDaxCnykeZ
PbF7O5keGm8a64vr6CBHR1ueo2p7SMFRMUl4v6m2wRpupbP/GKsYdBdpy7oGIpHXoxMZohSPNNUf
rv8QJLWZhrhCVD46wGC5g3WHXZcd1J7cbc/zu6qFNGJ1tOB3ks3ZosgIM+6M1j1wvNJeFwye2Ns/
djeIWJM3v/ELLAfvknVUUyxcVuSlUe+GEFEcvxPlbFhJ1SSD6kPuKPRB5T4tHT7BeK8R+dffye2T
ZGgtL6K+LmyjXg4UJmsvKKhEGvl1RGFUq6L7y9FoDoO9Inmdn/GJ1zcHtF3Sv6QtxxDdtZDmqbV4
GB6RNj7Sj3MMQFSEfBE0lb/cYZOQwhLr+mZpvAGyI8W/KdQ9/+O3TbWrMgnp4g5fPEwtnhR9ZlLh
nWx5e6XIuR07LiuG1ykBdX7kljF8QVj3TJ7Pyozf8QYMo85Ol8Q8w+TiXr1ddTIFchBV24E0hhlA
7wvgWxd+7Foyj8dlBZcemOoLIzTnV7B+yRS5LMHUcx55tjtnzt7p/sAUByTSoIIlBbJ/1ZJonwIV
wn7SoSRc5ojMPoRckoFl5bHM1sh7M7nJRpIL3rP0oNYXPOjqsgPFbm2Sp4/oO2qcXWkBNHFzRtjv
XEzheBkucf4vMl18RJEVNk0PKEaXULlBHv8uBhZdaSo0m9i1969ApTGo3QWADwctcLZKTb56VAl3
DleFEYWGThSXZkr91b7ouEobej4JD2+cbFB6mWJokJCoYHb/USfdRspprmBFGFWSaGhjHu9HRVp/
N6j5RakIYWzGgrd80I/5UpdVk7O50kgZXqMfE3cCXykDj7rAav59UWFKGBqgjCZG81+zMbB7SJWP
6FKI7WkNcKcdVDJHmS36oRjdSloRG4bG+8Fp0a+NuGAXaR6PzwB1FwcTOuR6IIGDq8i4BUeiUJQJ
cTl1Rzr7oDtXCFfgOdxA5VJwJug+5TUzQn+prU5CjmprstfxsbLHFM1xFLlfV3neKsm7/7hx+cJE
oFjybpVepNkR8OWYOodAoOCcsyfkcxCm12m0vWS53jQgQ8vrDx88QqhpgBttxksv7ZJyVy9EPNwV
/MqrFBKsUanWrsYnpngF1z5tyEgnwIGhCL5L7VGFRpLb4crBWTHTMpFRpOY1OCd35o039GbI4IIb
QjNYcEPNSau/6xZrcRZjZicjaqpHpVhGAC1I7fAjolOBzNv6L3/mf/8cyUnh1Z3J7JYb462jDDRN
ophux9qxuA4ZJ1lLc2g7up/+6j5lOi+wGeYpOB2kgalMPRKH1Tbbs5/s8isBBXatrY9xIMrD3kHg
vfMFm5dRB2i7jgm6zKRqPA0xd8b10wjLWE/7eER6agsbI/DUPfMqMD/iHqIwYinSNyKgkBD6p3da
OBMzavbvAOnOlUbiTlpRaypAwGL7lzv/uYng1NKJjjdDX93I/jvE6OrW0KPKIuwa1IgdN3+KxBaL
RAAUq3iMRuOTNOODW9scx7xzvUDftzh+ni0Vovn++bkT5zRHWPr8HsYMXTNv7EbSxQnfAJ8IzwRP
0eEgwEt/RtGJ8A9u2LNEIz1BKTWiS1OVWB4SWENzpUuLD72p8OG+vTqkweXtj+WaHdgJPdVRbV2C
cn3w8NC7CZR7V4RffIPrGDWILQsgQ+rNtSjAtCF6TiLsbq9q5DOuole1i8xeFKuldZNBsMtt443+
vNahRwFGgnCnxE8suvic5r9lRHHpx0rw3wl3pPaJTtSeMuY2nqku/tHUsxDR4mJv5HlKPlHQaDYm
6pAHuNoHdKrGuUrcKRKVMn0MORIgmjTpO+nJXpiatXRSDHDAsgouvlGR6LAbsZot+LHZ8w1UKSdP
zh+NI9BzVnrvyPyffymlDN0YnOCgKLIaoSh/ekZo2ve7ixsG5H3dAw7quIZRBPUC2vssCBaTkpx8
D+cEfDHEB4AED+Ff0ONyQavFfpf7LZK7G5KyyZlgobDaaHZ5O8A45W/UfjBBG3XU+2P65I3oMvup
Vk1fD1ee4TMk6NN7Gymb0W0AyEEZrPRK/SVtTT1qjBCEAR3MOUgVEIJMKamq8O0RmqQerL64NLk8
KZjlCpxeZfjTaroWtc0XXdJv0g/Nmp0vNDa939l752ui7Oow9M9w5o7Tyd8nJx91Lky4OccFvM4a
R/8EsEkMjf/zU1DnEm2HwyuZ9ZKcFAU1PYcX3tHS2PrLtF22yPEr5Iyf3jWzoGcIvLCQ5dDYy1p1
vqqXF/QbvJexk3D8dmJvEkYEGQ78fzMhYSzQxUZybvQfusyktTqC4OLwFBrVp8Qway3Fmxqsotn9
Hw3XDQTPtXMbJiWfUCjNzMu9qEU3g8UtW84ETWOeCKYpTU09LKPa6gLmKOi7HJy5QKnpPEeFLWp6
EVq3GmC7ajRv4b+GTL5A6VjuvvgwCcyC6AZrUJhY+xZSroJ1exebF/TisFoPCkTS1HLr3Tw8oqez
v9hqMEoZPep9sw6sJpV2BXfIcZKE6UHZ3lKv//6MefOVbVUG6wcnm0ha0pPOXWQncCRlFsuDuZZf
keTrXAA8wFm4PoYY7gNPhG9dOhHRzl+NPSpEI5PQR0+4deePi0rllGUjmNBygwDFJWGdCon7K3IL
d2dfIbNGksfGKLIRK0xS5w8tXKsoCft8UP25ujGixtHpvhl8VQ22SDBvUjWXeljzGjFnww6O3YPE
r4eXvejksFwXFML/DcDY9JoIVe78xsKKIWyoLh+xJPy5h38fKihCaew8d63BWOj4vd0NX+/kOZu7
XFulTsfK5XtdqEg8ZAwU0HdP/cNc9s9LsO4LMzT+NRGv+0JX2MvraVoGZHzDeb3OWuo7MOEnIRgH
9YSVYdMLeNaQEsuV3wYwZWHcxf3OQuu7ev2abt6C7NcqWpteGAIEqieNgP3neuJf4NPKVQz3d+qD
KC/gTPLdFuIeps1G2OxqCslUD7TLGBjP6ndiaZu/OQ1gJddXYHE75ifFVD+LDiEKV8ZuYCnGibsq
mzeHI1eA9ogEx0BwFkiJ5WeWeDPHtyY3j9nNnFb8xLFW5QNMZEpYaRuz4T6eSEnfwqO0fCR+BxVe
qhIjHxQg4FQVMDZZVX6edCZs2BBth2t4KunnPYpi90fkW10cQKnfx/YdbWaEO4WHk5mbkzLsUB6J
94sKkKW6i6+roZr8SLFUlXj+kmlWAChxlhm/mK0JCdnY/8msIo9cml/KQLFgtd9WDQp/8ea807eU
To9/G2lUJilUQ70+2hBzx2/tAHmqJWRsspTfvJVregc2klUhuHd8mpb+eUHMp7M0vTH1/7qo2J8d
CnqD+R7fVNe6t4i32IdHmfc92h5h3jSMsOAbeA/Q279Tm5XIA4IMYD0vtOgfEixUkCaXQkiGkOQo
5Sln1oNA+cxM2FhSys2nSxeFiJ8QAG/y1Z1tJpxGA6SgNCJJkq3bF06AOeDjEU0Cgp+jkoZSVtyE
PL6SsU/Vu2S6d3wUCNYDSlypEAkH/Z1K6ilZK7ci2GTLP/IXLn0wroee60TBrFJ5Fu9gLw0K5zUO
vIYUk7vidfgcZONt/aC6Tl0Hg7VpaiivA0CuE01KoTghxLRXH6sb6WDsQ25ykTEuomYtz2KSv+dE
hwdBynOPsSCFG/MisdIjwQ7eI+wT7Ac7Mk7sJJlK9vNdK2N/boiaxuqgbwESsQIbq0dDtv4J4J4p
fJncb8zJYAIZyXhh1jpgHxGyKrs8ze6M4rzbN0TpyFBle3l7AFI+nIHYoAzy4qXtokkud6MknlKN
Zs9p1Ng2u1wqf9SYFbG6CarsIp6EaI+3dBeR3Hu/GIvcFuCM+v/VH7yXCK4jUM1LL/o1khhBE5BQ
x4PRHoj//M45+FbViPw9/iEZyjkRFp1ut8e6gOGAXa3yEyOZSGN9t4HCophByeyb1L5pJmm52xUn
yv+n/qsjqFqdhMPc3WGhCzzlKu6jiKpm/nHDO7lFL5Tj6UpqmG7uq7ZncR7zyft9bo5UPVYlmF4K
WUCc72zsZsB2lvyfA1easvcT4VBWhIj8c0V5xsD+MCDnb7V5dPzTltNqR5t69eeahpUYlTwpTfDJ
ne/bIMT+TeSZQ46ApEuXMSdq2pKMtl46OD+po1bkhi1vwZ2ZWHKOB45WBYidsmJjDrRx4bcVBeNx
VN/ELAjjK6Tc9hbhxtlFrbfYqcnBFZvZSJacE6fnFF4JnE9zws8nFo1FesveDeHCbMTUkP7G/8ZO
YZOx06/2uYiXOvfnGsQdQltsu7oiqRx4ZImsGxnKMc+RUlbQK5jjyfBjZ22DriHFPkMtz36rGyX3
XJl62F6wMPlQkrHOzdQ7jVJsj3r7SzRma5pGkWBrZgNAvFFEA5Z/lWkh+NxX0gvMfZ2ZyvJN6Hu8
7t+LsnXF6lrzCvtMTmuwPddrvkXWSnkrXbeh+GX3Fr8HNlCiVjvS0N47SCx7RxTubp+EURJyUcMJ
69e9l1zUdjWATGj91TSeYMGKjE0n9RWJqY1J0kBRI/tHpWpbRPfBh7Zz76Tki4xkk7UaT2W0SFLg
lCrdfRX+novMu8ngrw03vGhTTLX8815ZRsLZL5Ik4GDkXgJtGHQPYAYc4JdDAWV1qdQskaVz7VYu
XCnmdBmJcJvX5XbzbRzrdJBoBGP7H5YD3u5T6EaPViWYGekuJv60VOvx5fDJ7xuQ5EQHZZzMH+Df
BA+6ibjdNT0mHe8LMs8JNDCP7NmQ/vNUABn0OGi1mmN1113WTA33F1IrUrcgWJ4xSIjWZYexo2lh
1ab66+3fnI5wpuSrImx7S/98BQTnmQp3x4fx2cKn3UfqzopTO6YKZxLWHPZ5xKYed+lSqI15GY5n
43w21UedgPy+DNOVKnSwI3ogRi7TkNoXhj99FAawUPBWHWsuGd4DkaF/25mA2mYBP8LkAfld/x36
gYcJpD5oHil+67PdLprn4WPb22mEk9MkWkmZmCXPamyW/APzuyQ/y4CHiUg7d3k+JkS9qtg4COsI
RHuwt4BI08Z8pOERWImnwbVIX0MASZnaXVqjIelt/8vyuhCBG27R3DxRYhHuIYcHS9VRTWYWNNDG
IO+7j5RL7YhBKAlKSPUr4UUbq5LA3SAuoeRsU0oR4fVia9BuF7Oo194WMrQqO3lay5E3MuP/gXTT
L5i88KFYNr+c6+moa4Xsf1ChDLn7epLvwhbCjH60EwNUeC4vAV0Bzh8woqJGNFxONJZ8XS96MGNs
AV6YNS+vX2DXgIXLw3iT3AciOlLr+Zib+aBbJhi303uyB939cH+a2pH0tUnbS5wIWP8aY6hcn9Fz
Q6VFqJk13XpWBybeHPGqoBLPiQ7YfWj8rg7iVe/9VccuPPTjO5k2DvN2yA5jY/hqcXewYRj84lMZ
7anJj0P5Y3Ohp1fmAI+rkNVOZSgFN4U7ZZLBqF92EnkJpX8uZXso0HVzxlaKZ9JvQq44nb+uyV/i
JCdWB4HV1QqCwwChD9XYdccX0V9d2Pd5HQEIGsMqL1EtxesIhI40bfhK9qWDl1G8BhzINKm+al8Z
mrFoj76rxS4QwVqJVRIiNyEAfV/INemXfyV2c0v8CwYsAkRAFcHud0Th8W7EkL0BQ0ZgSMWyWFM0
V/CkWqJ9T+NYnlRjyed6YXbyGtyVWlApzydNFLsSoH396xu5++trd7YOxzTGLf7Na0Gxy5ynt/R0
3XeKraKj2Ca7tcZ8RBsgtxoSOf+3+eLNAHTj6UzbYIZVc0O5FV1wvgKuh1+OdY+BAeMSGHeoczRA
2o60835qZ7wuFvfRWpFYjdYCE9HNauniIgIFwCluuTgp0lQ+CyG2P6aPCgN1l37LfX8oopQ8P3v+
v700rDW9Dct7wagsJiBYF3Mc9vTWrOGeoHVqhFxCPJXQiOrzrxYTzNGI10trr1quxIq0Oybbsudn
mXf/c+ATeq4lNdC4Snnchpg8Rd23ZIvuwbOp8cnhD3T4ikkBoJ2AaGkp22TkNEO9ZRo0ai3e7V/W
DQozNrGZqYEk/qAyropBRLzRVLWQqQgpwoMBDXj25Ts+C952fjL67PPnTkpDF8FHaA/gkOM/s3RD
hIdDveAZf2MreK/mGqO4nbcD2ZYg1qNp0/72ttUOoyCD1tkIDiLS13J1Isv6A+X97V/Z5yAG7qTR
UIFORn5nEft6sXJaHuMBJj+B71qjuBqFucslK/TAIvb8fphTwaQgr+qsMsJ+DuQrYf7sYhDoL5bt
4IT8zRkvcwKKKzTwWmuKe+Mi5Pg1JLorw4Q58RbfUHgkjDulECDAatR2xWIwU540btJP3wbQlqDh
ISr5cE6qYvjbhncSN2Wm35ZW1JgtreFhTHiZyEa8JtWlI8Za660FHxzaDrcueYNtplU36nsXNf+h
uvgTGinWrHHmfFV5pmUcc8zOhX4kmTbG1e4mrCLneLpcrnLJnpQZY5umg3iaoiKqoeuKhQb/QcgL
Bdkma20DY6F7FPPkwF37PmF85RujIoB18hMQHFOprsb6IdVvAucjV0v6u8LVWYtrCDSnR/91Htis
f85p4vPhvbgN5tE9CVPaJLJPpOhHWG4nFQzHk9gW/un0pF2MideyFnRk5hpu4w71MbPdqSGCtI6+
56+Ypxy2ViK5TEp3U0LVaqUeG1wQNI/6l1yzyCRPCjQu7DstpcjZTsBch6cgWNON7z8+gX44uRuX
pYrVYS+qzJ/Er/VHykk7/DRSQsif0yOBgM1Zv7w20C88nOw6I/uayYgT/RVp36YIi6dlcSodTAeC
CnrxSIlfSvLKaE55lpJe2kaH4jiq8u2KdXJbvd8c2zgrk0VGbsRhLT454hF4g3/OpNclKE5Q1+n0
1nGdKkWly+10bb3QZClmO02QlmG2oB6wDnwa1IwcSi5FDVLcd3Kn+bEfttSzWKpx08/9OrjhSAEd
JMpn2v9e+4M4BH7WA8AsxzbSrySq/ocTjOOfLqV0Rx/oLTt6De4pBovonkHF20gQnu5OnaS7p6mG
d2OIhK/JP4QiWl1wBIJOD3Jq4CkFJWhzoUuY5wHusqQLTatsGAyKNzApgT3btQAMEZwTYhWvo1ru
XXn9YPsigIieBPx0QSkxRVMQIZwAbobgSqV8ZOjOSr+kvbRm1vYD6GMb3v6W3ioEaU8PIivSRWYK
hzfmCYviWMg8yg6aQYWGZ9nC2P6XiT0S+OyMiTnGfXlPXo6fG/nrRmiwouMjI7kWVvY847Co7FQK
pBm1yntzyHgJg+6DKYyXqp/Bt26DXl+GaShKDSw+7Qn0g3b4vEBYibqgyg4bfqdEwu3K79yYuq9J
f1ifhWajF/ifK/lQM6WUXLG+oc3FahMyca9gVS9MWxgVN6sFv1CtEOak03wFQXQmkR8S4L6wF+l4
RR3+93dAkshkx/EcVJlmA20wC4UtVrtnCORRwb4LSga/Ef4bNDoNCsb8tmnedidSs7g5RLseWIrR
Ij3ZzJCTkTW4HJQ2A9kHwXh354kmhcT7mvRvg8vK4m7z1RO3f9srVjUWHvJaLE3gvZWbMR7c/V12
p8DQUgOoIjvzJD0/egHgDeuJ/8R1/pduKMtKdfdpPUzZ6IbrTG41HKbpN8P/DknxSgMREQZGE62n
DHU4zuz9gheYlg0LbnrmFApj8Hd59nro79akGRjie6j/HXTKBAighvtSazdCgV14A+umlIJnkkHX
E/wtPWsF5MlTPBHY8IrpqsVgBayQ6qLvrrVBkSo8002Jqh3gkSprSrtQmVYrh49MImVpu3K8pN36
mZOWNEhKpc5veyZI1RndJgBF8AaivTbq64PA+pOGY2YpHH8wGtf3V8B2orRPVX0c171budOx0d64
0N+8ne9mdAwLvLl0337hQe5yCFsMjAVtcmLpSJRKY++nl4hw2lgVMuVtZjePJax4ORD1ZW2eUtRX
QM7UXvP4IjaAn7rNV78fjmi6000+8o3I3uqmXFH0kRmLBk4dPZYkDmC8mhz75mB/HBm/O5jYEQLL
AFt6FzeJu1G1H1MyOjehVn/RWFUd70t8i4vEMnBLBDrWJNNU37pxp2f2bjVqhd74jx9gBbQn8ta4
4cErz7pLMdrNbZHllCdg7BL8vZsMV4WeQA1xAxbJOpXvWM5LchOA7SLxnjSJWuTtEkLgryDzuGaO
JljvRZwnXdj1/E0m1/2XOwXJsaF6xate0OVYSuwvWwZWxUQksftbceQ4fANmYhlFx/j0iTc09afb
3RHivPpXy1CyTGiDDAPKxPOx6YDU3MlsfJIdUwk4Ne+emVcA4o0NfOcwvdaBkzHKlfZp/5kHwfR3
OV6u6stWJFOKorlRIAlN1PhMWTi/fC34i5eqAsPMjbs0AD1VR6Z06I4MljGHzZuHQcfrFEEoV5n9
v5+7BAowZoI2lt5EbuCfkbretadokyGCMxS8OsFz2IcjRz3Io730RP8pi0P6ix1F22RhbdgqpHid
5XlL8e/yw7D3vZnHuGotLDdOGD2DsGWwxf9+hMMluAZyHYBXLoq/l5OaF4BIN0BTf+gIWl7xAv1h
wxoovaZL4SpBr201UtmA7/6ZyP+Xb2D64iHhGZKulJguOZ6VFl2fdjQPFqOwQM5fivn2OuERxOJo
I/vijJ/rB8hoyF1LNcsUaarfD/izkRXKJk+DHBUTX1wFGULk5znDLbaO3/0cyKurQsNNPaPZxnr8
R4dt2x6c13HS53EVqrmyRNF4trA7PAfMcHjMgNJdEsDxJeRMWC+6nTmU2FdX7SbtDLQfGyGguVPn
Gi173jR8onS6TJb62bLngWcj6rPWeraCiq41XitcaVSwSXgupaKp6uf3HPB8YRpKAzxHdeLG8PRS
RdRBYKP59TR6hD3npca1RbPKg2DsN/VP3nchY0jDXzqtur0OyQkxPnlm3z5uwHLLvTJsKpiL0SR5
kxLKnNlL9tWZ2E/iuhFkIWJSOuHKXgMNBvHYfASrHoO0fRDWcKMzqQZ9QggkJa279zdQjWYv7GAi
2fzU16LI9KKuAzWvaNF9BphMYAfAJV3FGZUOlABoxwZ8BeeO4tYY2dF5LERTNSUPZlpTw/0twuHd
rbgQqnisoG+SLq5HbCwG1Vok8dvFOULOEF7KRE06c/sCLT70XYdi0GkTZXrF7MaPrWEwQz+Vk+3g
J86g/srqhvDaUgip8BVA2fMo7FbhOB5px96SbnNFxEOSrpiNnLfA0x8cojqOZjfXJp8MBy5dkkjM
ZIaZt7RkXRssZ+bUXZ9tnp8B4hAN2YFntpokGcJUQTnibD7nm5KsnT0KYUJseOgW4K+98gppbSEw
KYrT1WG3z5KmXOeW8Kc4EeXoFx0CF7u9wZIU25uSGa+44wfPl4w/IUyf7u9QRoxPrRZCmSeBg1sD
xuttDrle0zLoodrt8n13RutVRQRo1u7Ugc+889WhRHl9XilJLvRpt07r0Q+YM63+0jRvwYPtUAtd
BUNRatx/HX7jhNw5Hir1XqvhgEe9P5tAPHWlVwGm0WCFnmUimG9o1LeetQYE7kcXYPen/Q5pUjBP
wsabLpUh+VI1tfqlwsWHvF7MHAgGU3UWEJS0OmV4kZEwQxzRh5s5+Y8ICv0PxAhF2740XyOBXyMB
foPBP66LsyeC41GJ7zfchVIbbAUJhKTS6McUxVL3NMrRz+cJf4sHYk7FfMip9Z9g9IczaV1uTjme
VaTLsW3/Y8HN0fgGkxU5R2ZnhCKQ0wRfYHVqgULqVpIdh9rDpmjfGvlBF84yaBEvpANrYio9UiDI
p1e2npGImX07HnaTv+skPxorYrKCup+xq3rO9djOUAyulw02NHOcQqDKGIR6OHf97H2Lg8XE2LS7
/QprTBYvGpzvDlcACvmoC212DE+jzMI3XnmRsu2Jx2ySKoAt02kObl7nxUiWphpZQW8tF1FRirqF
YzVjArB2A8gFjC37JfLAEv/IDf7VI6qplQ+m6ED26XdfgreWX7MpSd3MnbpTBAlGhwK1XZvME9Kw
ueSjPRAxRYuvxa4AEXjqRuanazjrhkIq+Juk3oO6LF8iDrKfCFq8a7OwKbx2WAtmClYeEOgzfBYj
TjNApgijERxVvy9c+orB9zZQLRbpnMgiHi/ACWFoxZDc1OY1aDDj4WwvizLqgHDPwaPIrvtK01se
MOiRl55QsNGkQTomvqGmsXWRMKQyQOX5ZuQWb9FtL5DTfTIOP9z9pMLqaYlQqCORWaCp0R7fhXMJ
DxdbfAbBGqlwO2hbRX6zL8GUuFCF1T1ETc5+PLor6XILjM2h1Gfru4dTXmVgY4r+5WXZzDzQ/fus
nW74JLNBBpFSjBGDogEYVS/i/pZ1GAWe5qr+2nhZafY9YavGbZTfBo8J8qzzj4ZYMmgn2MvAA3kq
9FuAx15IaM2LFfJhAv3pnrnFuVRq140e4XR5rbPykoiikU+ZGM+03dcH3faxRVlWKif5imxTBQEH
qOUGeubP6455NV5AO2ff3BIY0mkgve9B9cCXmcJYdAvISke3zZB7XkNb61UEkDKbUUE8xU/7FQfc
T+z1C7YybCv3lAKG4IpwnR068Od0o8OhJ3Jw7XOnFbsoqibWltPrLqzLyfi8RMUwXJyp9XTG0ubY
z5hDfpYxIPByf5Gt1nSIzC5V8e7vaPnQAUdFB/UK2uR+nrLC/aOawwTBsRUQzMCz4twon8+HZ5YK
pOoGV57g7kqIxK0B0f5P1G/l00gonrBoIfFYbSynovzfX5/0DRbrZSJETLtyjS65xOt7BmZ57aB0
wIdHgVCeayQhwy/lLUgO7mrdaWnEVxp402EtqyLRXH0sh3IeXMKTCzcsTAXcle5ihhf8YzgihDgf
2jXQ6rUO5RZE7ZxYVUCHqXZvUNhJyOYnh71mkz4PuwKvQsiZc6lAHWHwpL7E0klrjMfEnmVqJ2bY
rQKuYeZeoIITH1RsDJEdgp8wflkPSjNBO4V7bGpqYauYhFhGLTfiA+9OYBcubsOzk9XjaVNmJEkA
LcrjTbItPKz8VVW0yo28TpASMtVH7+4EC/077RVExwIZGFEYLnCAfDdyPFOtCcXEIpgMh9zYfBAW
LTg44ltXRHVhie93KVyd8cyWp0kaId5dv1lpRXs77qa32iOVIws0fN0Ts6OIMXMEcT+5dFaTm03u
GRLNLnLhCsutCuBJmSQqY1hP3+qOn30TttGjiCtvWbh4GTU8SlUXRe5jqPG4msRTxq9Z2EbugyDR
n4Owr1Odd9sg/JRqEgygngSyzxbEAm2Ip7BQJT6T1OvTgVfyFggbx2xwsf1ggRjq0N0oV1keMTVs
a5QaSijiSY3nnxtN6F/Iqk0VJTeAJMTF4eLKIpWiCC8DvkxKM0yubDfhtttjZF/XMNCPeUKi4HcV
W1wdQLw6G7+ptaRvSt7wccpoNksruWV1G6c4K0+Mo968JDELf7Tgu9S57y5f92UOnlKC3FwXjhKm
LGeI5+DCPNygV/BkHSTEvLNGYVMijWVSOMOI3jilmBQMND7+F0Bl3dgBes8iBQVScWve9oxlPZ+P
YhHQJmB9s0kZIU3xnmEIJLQ5UDxg1nGM2omx17RxdV8uWUAkH4kK4QGnBhQsdCUlWVLv1STzjHVX
tVjgSt+eP+zXUub1s5I09pn90OGCgS5bx0QQqob/7dUSTacNGudEPMjI+SNs4EtS46QhrzBWC319
JsFVQ1mMkiu+Baz6aqUZQIQZbUF54hPcx6aqCiLxPJJE4O3u7K4ijB8p0HFt24H9qL/lrzzhzKEU
eJG+kJOSO30z63FYuLd4wNniHmtGeKKTupfz29TwFTWjDyQYdMwuP2b7/a7DSwr8rTkobWf7DfoE
km/6lOtYoRrqvsywnvW8tANmAQhO6+7PxI5VczxbKvnjHfOHHhlmyi+XOSW5Wouzmhv1HZKYcbiN
KQxNmAMRTNnmsTn2Wiuv5XYHECJrg2ZNTpPx7O3TtQxVlo3ORnNZU+y/azWrwV2PMknJUigsvV5T
fB6ySIk/0Nuvc6Hep8MY+pVLWqtCMWT3wmHJTcwU3N4oVOo8qqNdmM1TM85Pjq9NEQMLZm6KQWZv
sQDGwtdKDZVV1FOm4CBRw4Ruw/y7GC2XxWQm9kqHDiuG2DYfTOe8Atx4dB1yuY3Pn8ACrC9eTGWl
4GVgz8Rmqfe4tBjwZtzs3KHkfIC/ig9w+N4faW7l50FEBKNNjDMzHiMFNtJC+mFP8LKHrMy+PEoR
4Jd3JUJ8cHND/mCt3eAO5M2HhntJKWEmhGzlnGvIu0Fi+XTB14e6sv3S1rwuGmzn74VAYmDo4HIR
tr7FXCjBVHTJ9JUlBnDc7QDZ+sq3N82v5YTItvy7j4UP2DWpOUUxmDppY+4D+/413jQsgcXgA15l
2/7fhIjAOLVIRg2PafbmKOnUuZvtjpVJ7Wv07W0b+BwsQfX4QrS9kklVLzD3Ty9Z80DKsYS74dMy
Zl5jIWQIpvTQWlQdnVofpTnBM2Rwa/fU46tVvfNGa5OCSMiqTS+h6TIJny+ma8JwK4GRjua/ITU8
6/dF4vG6w91p+uDub4F+PJd2VfGxcUUhu8qZgI/lLEvyOWNdfnAon4vS34lzFfrrAUmfr1vTE5d8
vEdmBB6lAlCDYmY5Y2P6Qe9hEKr55K2Xo0MqyWtJ7+0WzdMPhVwBfRdaiDeLlsyEUiD7xjtBVdv3
JWz1ionbRHqiELULOJ5HqM2gZy1sjTNVlUasQARvy4bgd/uIOpo9Kz0Gm1UTujARP5p3XrAD44sv
MJaBz2rWvwr+ppdf+96cllu89HXwngAxdkhoJEljmwSNbyL0UJKpE7ZPU/1x/IyJIHHrIQKuAHBa
OXeWmu4CwbFdLxJVTN03QEEyx4V5P4VUbWOJW4hoU1rAQk9HFxdE5zXKeKnbjHBSZOEHr1dgtpIw
QepOYG5eglQwb81GfnxX8Iko8abnf7snIap7s5ue/SqpjvtoHJjmeGp2Jisy524P4s6ZCowLtKV7
XLJGdFw7yTUMWcpampt3L1KjXrUomkQ7BowgPbVlTdrGnYSODpcfwgTtmAKsZVXkEF8o8+Y/4sAT
n04dApH4l+KhhcVDe6XRGgrVG3eJGrZo47qMsWRtML+/EpMWmnB0kJC++g31ZpO4DImj0W/m9tJV
GSFi81ZrbkOZJhZy+3qh30lL+eS1mVOqvvGyC7wqGEPUPkstHlJIYd9amdDuUDWWP1lBsgvUvR9l
xGYQQkc4fayYY9OQAWv3zGPFUP7OGk5FVtXfH0/smUUrqsomTKXl8RCV2FuE7xOtNeQeECz8okPD
K/oFIXIMsS7d9bds/XEh9JEFyBk7zr6wjTkZaavIuV8QBDZ4eKeIQAcVtRk+OBOW4Y3c/lAcsUod
1LJTWCCPm88xFbTF3aCFdm3JIja+Z6laO6YkeT6fZ6tLX8tJRcgQXVcK2gUTArOIgiR4Gg4gqfMJ
6GPwonkeguGOniNpoG99yq1EZ8SI9TU4OnCOIFBJfAox1y1ieC2GVhL4GEinucH6VILwOKm04SnI
SC8x5GEgIPPyuG8VOjnCtoxOvB2kAnf/fMiSFPLOfUQ2gpZBaLkiD1ncgA5Ut45Pq3FRAXnOEvRr
F+UCfclvyWckJNyhVzkAPSihMD6FqC5FvcZ69nNFZQpeM+zBuYFk6gRQKr9IhkJmDF96ojGAyIuY
YnDh1pOSNhTnigi/rDxjpwVTU0/BEOVqOt/SjActYro8A9TwzWKYCKV7W53ErHHZh1w/AhjE9jhG
+Ek5jWVkMyXhul5z1h4XzisbGbysE5eNksJaTqbYDHGL+KzcRh2VhFaj6v/+Mys7wnAt/Tn16eAg
t7sAs2Nni1jN/R3CwXUmeGQwEe27dpvCOY2pp4yIWaJGMPK9T8rzH5eGFuKP4e58XqM7tNojWVgE
u9HNthAFRdY00/pueK5+w2j7Tt3hHYTphfcYRiO3wTS8l0cuqxtD3eZVJ0CyTFsyuX2i9B2OEoEe
nQmCk2qVeQ899Zywhj9PV9f6mQypd7mWWgvNrTKICR0cZO4MucoFLn18mP3GdjoV+GgO7ohZXzbT
MmuJJzJhP1iw4M9Zls0GtzxsFPNvyoJweesLONfV196nAbrjds8Lr+LtP7OwrjV733TJmDkkZZnq
dQNA19kkQoO7OmYL6LSezLnYCeX790mGaM5BgSX6CEKjH8wTRt7NzURBiS/TiKn/sfldxGgn+bHj
BGupH7PEqhfZq/T7xFj/sJMTm1rbXoJ4N96jDJ2ryCSEhEAcdf8YHhYQcd/5GtA6ZCo7VC0Drt7k
7XSBgqfkQWQiuZLgoCPLs5eU3t2p0yWICTqvrnJ+qb2Sl53l+jQdfZnP+MgsaiANSdXtJzOWHiDk
uA+EC9Kg85dwHQ57Bc5Z9BUMaxckWr3ygjY1e8J5DJUoMoVZLCdXEDgBUy8ForAHSVLkLCF4JHof
VOPkhX8RFoQkKKIz/7x4dJZPC7/3gfWHEUAloIOjpx1kVnzYr8ZyoMmGeJtDKvoeDY5v3w2AQD9L
5iu56QWc0+vxKSaduw55p7h9wlP17yhalz1xcjD+5u8DLZnRoc2WuFCAE58GXeTTzEOVrV1QZxBO
BQE+W0/DdEdKcn+ChZ0WRtUGwyOfoKCX7F/hcWZejW98haxbPmuNQicsvkGqHHrmCl3TxdYQB/ut
AeJbMEGjeht8Fn8mNBP5e1+tMPZAn0o2E5WVy6alafSmxqK7UpFEn+lz+8cv18mCweX6PUAbWOiS
hiZewtxwCCi/Dn2Y/Bvv6+FRU89yjZaLQ0+YkQr1dBUC43iVEI1kKb4Izc/Y3HF2Hw2C1GlW4zWz
lXrTl81Fpy3luFK0VPPLyXv5q9AOVl5T2/b+tMlmHzlSBnGIoBwU91I1/zVYH2Z+TG6vXzv4T3wE
BpL2LlP1XCKow8RpXmB1Vlcyi1E70wwAr9/OW2BgpZ9BRPy1R0+VVoOHgTpRk83112SD4PYoV9gp
d2seZCe0rNuIF1vssD3IwdVpgxd688rR55uv1qGjrImzwEqXduzBmSVRHMpKsfDCff6pig1x1mFL
NSgK9wiNaKzGJMWE1EnrTLxh/QVhl215mj/E4qyBMwZ/j3MhBwEUm6VqhgIfqURVECIvoWGe6NKh
8FUsJmlP1jk9BG5MfRa7M8H1d9c5kWkmW/nR+P4xWXYeDgNtrHEPmsOwPEi8VYBlzAjPIuiqcmU/
YyHF4LmaU4OebylJ7eSc3h2pgetJ4gpc92n7UVYBwxqItZHWU+IK7J5MNEvYEqJwJx4VsqUIBgrG
3DSJuVvWaBsZ7NN0TX59sfXP0zfUNS2mnRazS//tmzkq3EmVq657b4IVo7q2jaVUAt0/8bK6yheX
bJP7Uyv2ELHAngbh+zNmCtC6SqZTogE93LCZkUcHe/6ixfBF96NvzWckr0eYa/EuebtiDagvpe4/
TiVNITbE375GeIb1yLrhEJygIjekHp0dUTliurZULx1gAC337jQ97lmeyo9liGQt9enb7nX7eT4D
mG0FFvGCV5t9c6sr0wet1IJdwJ3cyWlivLqckVJxv8fYFgjAxfzKSfio/VTozZ0jz5YXGWfTuGjL
UdbQmmDuzIQZ81+8pCX1PVYlZr+i1u5B5tdziv2Cvgq0YobjG0vPG62srtYhQcHuaIPEw+gjBLFw
NFvgrcjQYoWmMdN51IQyJnS57NjYxmC+xQoW3NSQaZkHLFIqO2WvJPSIEYz4jHh6yVN8hJcjzNxs
DWfiwlvlttGm218UIREGA3YPHNnKpgcRhpnhbsRIexMgdTuW9KRvjubuziJiAefhslVTNROiR/ew
rAJqzZhRPGEBw+uNDMJ600DThjJVx8jj2QOboyCt+yc9EoM35jXa/P2CYArNHkxvQXVP3TeNCsX1
s6QT7VIgynCF6truqO/ReOnReLoJGkXZAjDd19weIRi8HM1xEgMIne/8riTKswzjaE0ZhjWs7Fqy
ckKmTJVh1jU6MX1/mSEeeHSSR7WZyrfK05k58ZOAX9boxBBNrb62qwbr6gBnxIFa733pZH7K63Wb
+WAS3q6iLPdWgHyxE1vrB9xCDOkoFxDSSqtPcBjH/D0MCcBH89mvd2sfxAg70c1fB4Uu4Rxr+IyC
gJe6+cqW01kPJXEkInRpON3x6X4ZquJFNJrUeIERgVIissnVMu/Vje3Gr9y5fjbE3WCaYbuTp1Wy
jb2iMADgCPWK2zL/Ryu/sv3QfQexNH2QlnsBjxFXLusX4QqvIy4d6xwabKU6Yrdzs7GS/Pjp2uAM
5gVuJlidNQBpRFACLnViLQjji7TGCmN0NIo+kRTEAGevGVhRIkXmuvuiE4hVza7w1xBsAZy0o8Qu
6U3JG+LsAoJD5OYg1TsaEv4mQCxCgsYcAXkVhOhVlI7cSJvcCh6zN6VWEEWvABuDwRkD5phOkH+i
6kmThPaX1Bn3qC033C73iyKQMJP+hSVdMi5ZRP+DlrFUjv/lEAJMZxfu9qTeBS58Az0jboLlgsP6
oRD/+m8x3GG4+LSjgMa4SghY9Ul91/kTKpUFCIzCwTRZJm05e4tC4vnor+WtrCRhk7Jhba4gjumb
j9Ta/tsf9BG+2smeKaW0X6Ru//UxwbmxLUAoE9l0fZfEspWjws6eFnNKE9jqub3ycqWFLnEvl53G
ldSjrOd+6Zg4c+/Azmq06kPvNDNqatw4yXjmZ2cyoqZGx0bHxHqDu8+UVPH/nOz9hEN0vBrwd7Qo
N5yFn/KAkfVQ/NtCPn6oPf3Ycj8jE81sXHfh34mINTspRyoj6GBJF3Yy4LBWXeGDpvKZvv7fa7Dq
XHpakXS+2ti3zclAxii9Ag8iVzroNGz0BKCj4rfp00x/npYnaduddSe8U/yO7mxonXWj7iOZEBB8
kkTNTuyf4B8wcfGJg4PPaqRoeoWK7BxHkdryv17ptUXaWHNXc5ShVX7AW7/8BX2h301m+shBKKH9
To3dHFNaAiaqlHPgRZ/ZW81rAEx9lT4g4YW0ENYW5xs5WLOes3xlD6FFKBuMmEE8/4h3KUy2ORZq
pfW+bf2Es6r/8JUX92aCv0cZjgRKAyy04pA7fjwilBHXw/UqUbV5ldnjmqGY15O9ZUtap4rM7Tlq
hb9ysEKlLVS4oXwJrh17qkDtJWX+WQeRvMwmXzZ5WpUWLUWRHk+KdO1Jn7gJAg6PjhfArP/wJZFI
OgDTR/i+6rDryNEP+9pNJtW1/SxncXHVo0UTs7ShzaJfSBQe44nDcHOpjPbAcsUuAVt2yuW52OkH
vZ/UUX6jI6KMh3HEKVXKYe6SnxVQL1pgtrL3teuOgTwwzMwA6UNj8fWZtpkop1TPH1MuXxK0PeEs
TFU4aY86Mtm8r5TAdLwewCy11Yvo1AetZ+iHPUIn3gD8TdEPxcf8W3aYk+ALPswVC7R9IEN1SYJp
LN4alK7L2tYkXJ3m9VWjrygeKlU3g85buAvh/uqNmSlImRaZZmfopsFchWwAGIoojzMHPGK7WHnd
Ihzgb24cqsUQ+cvaOImLss0bte7m0lKLqpZi1Ro8fXypYsC8cUNyVf9cVtuBJpQdFH/UuCeisNae
bYMdkiz+dCjbblEmD2oEkl4fBa5+T3+d0QW+ZfACGFS46neMu7gP+x70IeoNBR6E+xN0ISr0732+
AmkdgDfGgK/J9FdgzB/FtCE7H3lijz9QHgqVTNe18TylAQ3ujvk38zO/0eV7xjmThs4RN2ojtBOP
vwF0WSr1eCX/end+hzbkG5EkzD7eGln5XHSWeajurFXOoiCJ72IjNpDetPWLlNuXPw6Gw1QIuKBd
M8fqlqhVUaI4HTvLzF5IoRWyn5utKolLIF+jIy3anvDJoWWSM4RZFITyclskZeeQ7a5tepND/uk7
EzRn1JKq+87FO/tJKj7JwHGVwMidA0cjKEEG1OT8TqnfoMDJRnj51D2hEW3tx+gJCaWaL5KHkdys
qAeK4FBr02xLJU7R90QnvnmeietZy9R5BYfCcUponeNGKGTBAOfO1gRhBLn2GamC8QKBF2wwtxkc
m7ozSfYqdjXZqXFf+3sWkHntiCiFGyfQ/k+YZ2gsL2DjZs65zpzwUPyh2XyrJVCfRKXv9WNKYIlu
6gIKJvIk19N8TvOnyjjMIkPp1pXeFRXrleM/h7i4wDZ7Hyn2iONcpCphQREDBSyruAihQR3EEWDR
PB4NZqTZ9vNvye/6Ht5WMiSp/mhCdd/tQ6Gnc2z0PE0lyBfwLN5TP978aP+KAgfQg+DALqOg2dId
woSb1I3wXHiRxG8Ygnu3R/lXaShjSK8G0j/tldXQnBNA7TEE9iVltZsrsMhR8hKGErvIv8LztePQ
JvKkWxALFaLmXEn/V71CAAjfxxe3rHjToXD2I8Yk8gRgqMYY5dQZ2v3UwZ1W3AUAnJd/YlUcOVxd
2DiYLuSMq0QA1cRpOL3tbjfFayDdyLxlzLb287QSUsoYxhbxaXWkIyaQmjqua159cxJIYvswuXtj
tbeaNP+CJtTDKF0ze8FSaAk8AVZVEGtcUmREEt4qK8M2/+90zta79hjP8IxvJN+v3Fhz54qzXSH8
eEzisGPom8Q2fQxfnMKfhbYMCC+fvHSA+uR1rrfSWCbZkfyxqBlTUHYQ/jWQVEtOQEmD57dG9bI8
uZBZH9qFrXdoAa0aaGdUHqD3cQ3u+q5FdAL+AwBf4t0Wh8Yt9JFxzwetijnl5rzUmeFS23ZPvPem
GAouyxdvFDhAHYTZrR5EU67rTaFwvCO5dIKhqQWnFLxP5VU09T29BsCoNo1zk5U4ei2hHL9seOiu
LST3try1M7ZG+sEfIVJIMwbm+ICwXqlol5pIYgo8oTboUFdt+/+smdNQENOGy4/2B3QWJNYhomqQ
ecbjoMvOvTdKTetOP2S8ODJ0+IRMfOt3169a6zqU//Q7IMWoK8M/h8RuT0s4RTxMvIjpJcjIWmpy
oCX251Hx1AVRWWd94Q7YkrUvK82ceDhcmxsY9xLBCHDroo9WPYuz5/Kbw0xoEZY+jNLCBJ8Juorm
LaSc60ttfMYbEsadAoO5Rbjai2fof9SUoNmX1akWaaq3K2UmOjFPjd9CM3XmfaptfZajHj6bMUDd
h3fag8pcHF9hIuW7t8r3dm/Di/YKt7X/55fRHsnpqPLBjOtZe3SVfUjR7ojUZ9JqDjfCrhosbt5E
yzrZSjF9e9dAVpFKKK4Gob9VlPJ6W4rsTNdiacSNFs4DTUJoXh9IHfXMDJleTl6/Qkr4GHEs43jk
VzeWWVzf3MVLc+82c502obCvOBzisP5wUTFkPDTHikXPXezMxFbAxOxizkuhp9E19PGIaX8M5/kt
TD9W5hFDlyiaSjzyzOalBzepdNZie3jxbmSHDnhEsvbHeLiiDGwujB3BaJuno2jxd5/NHyYgGa6d
//ncES2u9Mp+ilQJRJhopCx8wWZD4OaWXmU0LVFWL0AJJcbb8QjYGpCi3Thx8+f4BmRoJhMbxpFk
sxfSbSMC1wMTs7hRmt7uwDa3FBb8JzMbMR0jFAp2m2tzdxIFqY2ensI2+pFo/F8iw7wsoPehnyBO
bv3Xa5iErRXo2mP8CvhbKOviB13NMCGY84Y27rjY0pZQ4og5n92o48yfnoyKuUSD14xvJhcmSggo
s8f36M6Ctr1Y63JRF9h9qtwcxNXljAayqD8IPrb7UIYTWs7l+zkux3iayW8SRwnZj75RXZ4mtvhm
pmN3xFv45rnEYC/cWagyzX5wfxTlo/txil7dSb6/FmvXkv3KCY/bzkRVixLhoQAAoxNur/JlZ4bj
k+V1Q3FHx4FFRAEMBqy2a/hKTFuQZEb08fts3u49w7wBBcq1btHtMuTHcl0NvmKS3nSBG9h4exZZ
wwsA9Y6NTrLnina5JNAsJ8G5P7jysocNAKeYeIIAoDxKHFWWvLkY5ODSljcIgcihDOlpiEQcjNOi
BKem8neQtXQO9mVGfk1X2u3Q06LjZUy/pk7n261QJezI0brMc6rDvbyDw+UB5ryBPk7FcbFqzn40
/CzK2gDwU3lTwlgcB4KIwJJlBpj4RfOFf7blhM8N8ZxPuigeRe5e1OA2PtRmJa4wIctvwoRPlf1m
LsobYcl7XI0oIoRRdayZGx1tdiYSkfLSUgKFYtaDBOzSK+0hYO/ELzuZg/P6LbzDJG7h7ppWjJ2R
M+yC3h4Md2Fi8rCUFMdKZl6E7purzAl00I50mpevsSp9ALDvE1b+IddQGihvrVJBiA+GeIz6chgG
M02xWgYxlCSWOE8EYTXF/38/l6mbxDkzDxfZyZlbreYGcTToPTT/ZAdMCwd9QEIAqahhlyLxgMh+
68MXs/9HmoLQYc5DENNXY6VrN4IQ1SNzLQXNyqXZvipwjERwSPbehohNIkm66WXpd6o3JSHzbdTC
QXYTe8CmL5msyEm9ceXIy/E+AGJrwFj4r/FDSVwBv/ph2vWyXGBFO41VR+Spt2XFB7Gtqy9rJVrU
VoDPxpb/4afPu3I1a1z1aDj8Rj4azqTp3FomdbVxyU9xTfcfbCFFrDrBG+wD6J1OP6x1wpvnVYzX
CRBrnEHYiRRfAAKEs/ExzoP4K+LCwvswAqZwhbX7qhHkuljqMTG4nrl1Wr6b24rK37KpU6wBsGZI
53+jGGq2a7/dg90L3CYA7mZprmo/jIlIpIWkgz76tY4WGJ/ahQm3q2s1zqcuIEigJH588mphG52S
cl93V/a7xeEl9n5SmOuOFduL3XxfRKSIfqWG/YChdAadjCy/B6Sul+uZdvbR1mhhuvs/bGYIgiH1
m/HjjEHW9OqIKMfO5uBa/FFcJqLVOU8PqhWQet6O8f0kVt9J4h+if4ddxb3yUA6htB9/KqjpEWjF
hcnp8rcWqzVPsgfD/hargl7KvKaVeP0eQipctyX99davnFrfpbkEcVhaUut0DCq5t30W0qgLTqnQ
+rf56bnAszqmIM5HsMowlFtZ4isTSiiLCuKv637Kr3nxt7+xM+jOS3YRE3AocG29eoYHb6Axdmm0
zBv3RrIkkhiU/L1NO6QgmI91JEEQqZkCmBNIiGd9L7CjYxu0novibG/8nnFyt/enRegkBvMsL2tW
fKvLhtNlYRo3woHhZurfj8b4fSjg35aqlYWBCnY/Db6aVWH6Dd0DG02xED7w8oDdO5f0j4ypVJF6
gzsC0kS3yzls/EN/5uctwA4mODu7GHrlS26nDPD0BBZeC11HjJbBwjjkrhMM9q50LPe8UYx4Hlxa
V29xSTqgRvctW7+ijsug19dMSFO2dgV2OjUZiLjFgysO3en/tO2jvCU8u2qLuiCHkm901O1F0LGw
d2o2vNang/wSKr64VZbuKTem9iUFLZ3nJ7OSDGX3shC8kqJu6lHKdvneySlvsBGn2p8tmrihOuSs
vo79ypcpmC6oUkkYZ3UW0OMtBSLiYqIYc3q2d1/ahSV8HCw+p8Sq6nEJjGgXxTYC4jhKn+Rfte9s
UqHrR1WITQ/RF2QX4lWqVLUKUQno/LZyRCsWstI7AYafcevqAdSsuBw4gH6O2TsAdu1+ZNkTdM/u
bPmfTBnmmOWac6DGQSB3Tyso6ydwip2P1Eg6tShi7aRweZxczo3HRSgCp48XxBeARtZgh4jsv6N5
ngsuE+a9Kwrxmz4Mf3+VirXhmg8WvQTLEpIbvGGdP707YWciYEapHL/P3xRyDbZa8tr9+0tEm9oo
R079Q8oWgqiEXBf31yPQTbEWZGl50lIE7yMq6ormbROj5W6ywjBgdRjFZGYXjSRQ4mV7et2HD6XG
evW1n0aKT+zeB794dxu68etKIsfwjEGi4L36MHQToifVUKJ4XhMtxP+yKU1ktnDlEOBhnxDa5r+x
v3ttDb+enqmqEGVXwATbcqOjbD1QuRpCaFGr1UHaaBTTslaUw6aYR907BYa8NN2/4oW82aJJMg/U
7GvHlvcm8yuYo8M01o1UKFYV+l591WvC/1SgNu9n3tjq4364iqME0hwAKTHixeYIPxVn2JOqPFq8
WXg7z/yWLAtDsXp3pm231VXCg17qWnZ0bZ3ycnpaTo/G+kjn5QuF7hC1GqrbSOVYh8xq6/KFNP2u
I9D3FPKwNX2Koywn3iumzk5zYPZ0pr0fpN9czydJN5RM8I140A3zg50c7GlqyqC7OFFyntMWl+51
jkk5FVzf9xGZE6S8AjyTBJA8AErIE7V/dYaqMCtIoYDYu7fa0i19zqWYyMpg2ZKKBY1/8+IwtOwz
v4BANGYPisBpkaC69DK+sUWFgCpvwyMSbQ03PisaeZhTvEN608xJxNkDuepqUEjRMHTEh2WC6F+y
3v7ch0ucuw5TGvEGOH0W6uM0mqbNdQ/i5up3ChvPFf2Mci0+LXjxjUVTqFh5Z3UksWzwfnUd08If
A8ixEG0nq+a3rCo81/AGe50PQRQO9lI2QrFkqF+VUSxrMEcJHcp54uYjXzNSgAlectths3TOXizR
tMjirzoQaWb48aDBwBRcIrlxyqGmaAOQoLv5XQ7zT2Z8vJuyv4jBoXzlhKPk7p/dOZ8+XGtDPND5
XunvmaIsSpe0EY7gxY+uyXNwMJiy5cav9ammSHssma0uZwOaxAcmNLlFcuSiZypBGSNPFU7xeM3T
2uabtF2S1Ja6d85rB5iJ3VJg1W9WZSzAh6KVuN9OUHNxn1EqR6kQaCjAYo/D6AkiRaYUf0eo+b5h
8L0p8nxpKaSU2IYIGtWiU37kLuiVnKDYzrCfDcQPcckWQT3QZqtr53qsJc7oGMRyvClBB1cSJwa+
20T3u0o0mWNToGL9IZsWXe1JwasmHa1k1v5m8uwCVPzN5dTohsNMtaRjoVwKsMC7t94U3J7tbkXc
++zX7RLbFoJ5/31MiMIPd623LWzfO2vXka9JRLwQkyIsWcKw0Dqtszy0ohsqnxkJWhehk4JyXPyh
bqNzXunpyNA1/ilkKDvSnHuloD+NBqj1IOCjTj8bKW2s4cNAUEOCWGSW02ksqP4rsR+0x1Uu1KDc
ku2fWgLnJiHnKNv5Jgb6in8T/7apNnumSDYfl3/MAzF3pKx6wqtZgLTO6kjpYIlLyhmDsCOGgJDv
q+bXEmoUhZ5bvg3YA7c7omGy6Au3pmoEDagldGfdIbWrOJiL8j4YT3HN6IKnC5Bnl34eXuBDSLNB
d3QdtE4hAXZgFvVGqHsayA8zb9FTv9CFa+UJOCb3DguvX/nnMQQKfbce6osaN8NtwhwjN5/So71a
DAL9RMG2BvQLSEA4p+Y33KGZmu9pW3FjEquOdjHC5pI+TPS0SLWG9G00fgg1hR8UWMUOR68Xyg6y
9H0qgE+2GyAn5CKG1LEqfRgeU1METqnT47drz1KIMF0uDK8H98NiNrF2p2QO2TNDf7EKqciZOeNs
IsXrD71dSyO2PrmcRVhCFu9Ui9WKi36FlsoWre9jZ5D/z9Fi7BJ5WzB1nZgKEZhZvHgHQc1t7CDP
Khtpo+XJqH6zTSnF5OxFWwa3h564eehsgGYklpx3GVRsvU+8JgSlwUn1bNh+Rw65XoerKAdO1mQr
09+zlp9/egMKnHKLuu5ul9S6g/DiFrNxfOo/xY9MnPpzLPsxJBcnNRD3TaobVlY+Un1LxYsdKak2
OaA3FxTmFDOIVljqXGWXvNn3lgvDdfpGTaAa93AtIjB3+d1vfVwvk79KeOTe4I6OF4mAfEfRST+G
PuaomnCzAzBUZY3bZ6uXmDTt1Yr7tyIFCoXdD6K/9n78Bblq2BQqZwu5V0ylzvNijmwwagAUv3EG
aw0Dc7k0wdhMkwvoTZ5vBOVGBH/V/qo/wbwubXv0SY5RkZtKnt+agesbCoUjEr1OqtZwt2cp4XkL
Hmk0N1KHGtdO6fdBQe/rOSMNbPUIPdnOAxwaRlsRYUDtQwPajfhvytxj3a3PdQRxkMByKw9/4YS9
nXKqgbwU9VIXgABNGL3wSWgpI1MJ+8sO2jL8Uz92T6RtNY5Wh3yo+t8sTZ6N6KkngqEsnQsCXwDV
m7HdAmk+6JTwurAEaYkAJ4njvYbt5dw1p04aOgHGeht/AwHa91GzgacN9JLfkNBJiFA5/ruik18k
h4rX6OTcl9Z1ywX7dsxyBC3DqocZ0coV+ViyGutF7es36Nlbyk+g39La780PU/r9iXuB34qMBrey
LFGrMHv/dJdi09PzmorAJrRd5NyL9Z8WHMBvqrx7PJ8KvqF7zGPiRjU06jfJHKfrwMYsBtgebap3
JiSUiSknVmPucqKxO3eEKD0KN0qB5gXQaKWtR47szdGpRUszGxcTNnvIwZEkoWgTpAuufB+RT4S1
0KN7WvLH8YDSONso1gaWemzEUNHfD4Weswg0Xc3On/C9ar6drFfEFLR2x6Tm8kNzt16xaAyIxENY
fxMZl2PMzjwls16J+ZNXsGdJsOWSqeL0fLyko5nJvqgPAvWjGFEuiROzn86gM1M1LydXwZdPVbH6
LsUqg6DZ7hKYk9BFsrp36jXpsWntpPOtP2nIMiYFtVoR79CnkSwEjjn9aSJtGxS3BE1iAS4Dwy3S
DJIcDezUuTIliDn8ixeEqDZv+nOoA70TazsHOxA0mpJnXFAsHB9t4L0nyKpGaGnR8+lW551VgShQ
HLZJ2MZOhk62bfev/j+Y5nsq2eFGDmtKmMr/KMAh8fVJ7qGHxUsLtAkv/vd/aP9/iRvGIwwZSRYd
wrxrQ22GyEGa1s+P309YlFDPqbAu0bUeEdWWbyfjq4m1BYbSpUchOQ8t43r9eAbNlHpRcgKNDeD9
opyL6nDLXF5wxdPXJ8+KOWJTBMXMlPVnRAyU8CE56K/40l+ipg/8QAb9atGtbbt8Sb1OU0Qi2yIy
w/ye0LPcLjlhwoSjmkPKUdeP4ZsLIWKuCXRY6gjlq2zMewTbDHFa7cdmUYn+0eXxivbW2MS/CnIx
0zGColrtYv9LCs7Xw1jnp9FUbNFXHHZb/IeKN+70VnqFZoOhgGG8hL7VfHAO9vk/PFtLX/ewMtnN
EvXLmeJrb+OSKcVLnRdllG7GeLOUlVJJG6Ya06jshqUHv/sNK0HqdgkKxXHsit/WZBAt17yqRYYM
MR/uPWWNgu/L7fQfleVjjylLrukb/y+dTxNJOdQy70RHLGDttLy+yoKNzw8BlIins24nt8Dxwnrj
bFin52Ya+dBMAZI80qVYq5DdkpFQYrGs1yXkzQrxsm/l4vbfICChuD4um50XgwamOwdw28L7dRhj
S6CRdt38r8sYZ9jLlOjeVWtobf65iWpzNemCTSyJS4xOlvuYrrNvlW1dh112Zxtfh5YIQqjsa1pD
NjkKxNfeGH5WiKcCnr5lnzrfg8qSbGgzPRMPagPwBBaHLGuHuEKs06Q65WIDY1XAs+JGb924Pyxk
ROGqg76YnKFTpKSGyHtGHGO/C94YyId/ik9iloi5FZYd5myPfWf2s1cMESbogwmhyZ1EfhTZW6zC
/wTQk4e43+elczDIMkmmb6ma4FiU8yNud2JTFIJb6ZlMRyN85OtyQyTpnBjoCDPuGhYrADrRR29L
9uP3L0FcqizK/AOna4iXW/PcaYAG9ln3ffQmzE7vgaQzvXVHk4zE1waVAj9tH9fYopWZofLoFMS/
WhChzyU1w/59AJ/XDPBSaNUFoKGqR/rw2Z57R+gz9pJJY/x5aeucpifHG10zYoHWUEsGD1SshI1B
rD9CSSFtsuas8SkkXThXyAEHhE8PCvX77pSkLmM1bW2Fr84vKEoKpm5jovO8f19BSKhtogvKuIPh
FtGcuYBpb2k1nOERK0cxBsmFmiSGsQj38+40qo7X7BnRkJX7XUmJ09iM+bDolesBafRvZ8IDUX+H
KO/CxnoxYNgR9XO5JU8NoVlQdyIi+IXD/Ye1QyReSr/cOwU7pBPj+xPvIDmVRcvezTfaA4IgAH/l
0Vy4FXutRV0LAKSq/tw3t5K1D+Uc0QvOzue/WInfnPP4Xh0I369Znfb8RXhDGZlBq/65a+lRDfFp
3EyUmWuckVAAzR5ggOt0CXI4YaQbbsv3VZxupqgK9gb94nKhOaVQoA+Ceh51EB02IK6HK0lxWvD9
+0+dscIu82An09rLWDsvCecdZKdjeHX282OwLHY4lcKunyvhDdJOBXbYnuOqUyneXPqIMZIJuHnZ
ZGnlatTCm+XLRJ8DDKLY+VT3Erxt+LgTBeRGbh/EyeJQeBzEO3AZ4gZCj+/hpPsdUE2uIqrkB8nh
bZFMnKiBRCTUJ+ydcHWwTpt3DiUE/tiHM0LH0I+KJycnNDkwy657XimxJv/nJwx3l8+vWSs6LDxB
s+6bFR2RVIjJnfOHxMtggxl/ptlL0iYNywn/239KOnSQY8dbB14lZ44lUzzINPa375QK7M3GUF5X
nt6U/TU7UrSDMBwetU13ChRm7yAG62M9LlWw4vE/EN5+g6BU4baZhqCwFPIIjWGkUr7LIaZ8r53c
mdpUVXrV4WJRx3JF+4IDi+GMwIKLC+hwTRSgz40uHy+pLw9a1pynLtr9Ktujm/fUijsMsG4i86qo
WG409gL6Mr0dHzTVfvyujiZ1cUGvWj+u3Bbq7yIuTbStSPbBALAuqmMLH1y570LlLbZOEFGHRw14
U7mwRtx8Ccgxp8jyjMTomi2RNpsGDQ61OpHE5vorYct26p2CK12e+F91hS8e9enn1KpVsqDIG+T+
pk3XKFQsdq+EJFGOOS+7Cji34lgTZwrQOXwLDIztD0Dt5vaMoNm1bHsRBQQ9t9lUBbvi1Fa5u/q0
/URI/6E9l/30WDmGbfNYTWZxjavnvpQsgiqXmbPWPLZphg/bJu8J6jVobb9i2SwyapmT5xkJQT+0
SNSQ1hvx66H1nb8otahXdSEuqmmO/PYhQvPhTQ7ZjUFLVxw9bySNusj08X/K32dYAWfNM/6cyFux
5ZJHj6PNpFLgfn3KB7jKbQQ+1vuHmqNn6LbuY3I62qvYOsEgY3z6/gL4fUvQWV99Cwqu62fZ3BXV
anz1+JPhNmnulTIaIddfrSxXmK1JEFwIs0A+gfEw2ljvWErV1JDa69wgHf4dAy0GY9QgY3xahqd5
IOX9a4OVGXfQHctqGrp6D1CdSPC/bdNBF4hAd+xDhgZu6wJL9nvc7B4IIrLZRSu+HGI0j1nda+oM
tL0mRDTb3Z+aOtGw6RTeGphqWsOFEFtJYskS1HvfvMItCWTpU3LWUfzNdgb8xyQgfpjQPmFNT4rE
pdY3k0Tz3PfYhEhgux+4sIuZ7Ht/jR8zx/tkbOzk5tUdsjt6ak6SVBRAx9J8kMtoMXfKQkuxLvNe
15HcYNscm5Sf70G5h3Cc7Sh4IHBKwC1sHPO1GS0SBGX1vg16enY9hPICmXOUTkAi/qU9Klx7eb6Q
xnHmYfupmY53VJSj5syuL2GbkUH3Le3qGrCCndR/mSXN0r0fp6lRBJQym4M4ZjgDj8cXmFZcu9fp
qVxDGD++4G79bJx/MiBijFudoDaGDVc13+kTACt+q2bT015EPlCSMurwGgIh4r5b2eYRJKg2Vxcb
lEpSzRh1yu0DUuqcsbnHRtqtxNxzeYX1bZCu5Cry0BqKu/Yks6spU5ihOtcwkzZOkDjgmDzRJ7/O
c0sFFLTAGt4nMGdhJzPGDZuXIstCbPI16ujMPWrIbhHrkSg886+sfQJR7Wk3v1IhXQ3XvsR07+5a
8Svc1M5ARZz+RN3vvDmtHjE33ZD/61SnU5yXmeZT+lupkPqz9q9WS36uqQK9PJ3X1XyDahZovD09
y94+hwGkr1IU3PTGKUhVgvvzmXMUYFKLNkLG0Iey1HsRVvGc0FO/4yIVjDvFQVG1dNWaBezYe+06
hlS5sCO3jwbE/RIwT5AOsX79MziyGmOumPPqMZa4UApKCGlZwW1NDqOCOisr9Z3BQGTCeWNKY9x5
CKAvWrJ0sqPQqD3Ymhl1dKgKpEIH7mL/dydzclNEb3XzBV/kDkJ+G/8Vsau8b+y9mbd9La5h7Lpv
140e3uZOYAFW7+OkJ8q4GIHTtKMll9Dux7YRwyoJ0EFImxi+BjUKcs7EhZJWq4DreX/GabsEgl/U
9dlH+oPmWzEDWf3AsMq2pvqcl3hycodKikfO90akSLH573Wuu/TvJGOljim5vlqpVNfYlubZC2h1
eXnx4LgXDc3w5YH+6QlHGoYUz4m2DMEHnoU/4yfblUT1tqVmeGbtRW6LKH/aEURBTV+atkNqitgJ
v5LrWMutF7vBwk72AyY/elBvZMHK1lmAuVnitORzP0JobFaRR0/VyE+X4QcilMR+fo2IEUq3mH9n
tyqk0FIq6fMvrdbpviEqnbdPHD5AdwSpydRRII218qm1p00t14X0p40K+DcfMDCIhpf6goNr5mmX
8PQcBnBP4uK/nTaNhsvjeuPufoPhQEWc5fPg/SKOSabJCmkV+TQKw0bkvJKwxy0D/I/4tC6nxmko
00pKWqIERlOibUglb0LXV3WqH9CF2o2tF4aJhR3TnyhEblQPRzSb5Y6VwTzj3GOe0KrCHYfMXpRk
dNKKTh5kojFNSL5w90qGNyxEBc40rXgjP+APYn53eFcbhONvWa+sm7cV4Iy9oo0zKbl+SbzoDjYX
Jw/7Yy4ibS26KKEkiEIYvb6g/Bfdg52n/qxVwwVueadAUc2nfyni/ND+Py+KnzjI9pl6dygLQuzS
wVt9TFlia8Wace2wG8B+84Si7/Cr45I/GRv6jyhzvDWy5DS/qdYL2bp0ukTSiVh+o+fLhTTsd9AT
V1xozXVo26MKd+jRLAA1WtTSJeV/2ks7Ghxab3KQwWpjT8+8y1y6NA4JBw9gfV6UNOgyih1M4FZR
7GRm9d9gnZti2lQtGgfyOoULHImdBkDkwgZRWT8RciYyKe8G1JJ7TTmd1hWpCMpWkb8WqRwCfXW4
HtmoGjXgXaDByXWtcOz6b/lkRuSRvnOVFpHe860aNkuZ2vwV8/mMmbAmpylTLQps2akgXOxhl+L/
gjoqgClH4HHfjfOzcxOJKI0M4pQUBpN9qm0s4YKDQeEvxePCnYtylF2oUjY1tjW2qsVhk4L4CJXw
+ZN/SowM0xMH7cZMEbmeJbBaixUuQeG98q9nzRUe1/nRVJ/Pi00mhDyA5DOjZyvSWv0ip3eP53IS
64nclfcKVdJs/qJvUwTWi8o1E+hbKoDUseu1gQQoYODdewlzyIrc4HkGLZv6hXpeK7JDFPdhwFKj
0Y71Ouh/sk4UDFF+qXWPnKdOcNeUbBx081qOrKCOvrzWvzdbb8vs7rWPfRIxcMa03vfRXO8NED/N
W61nBegfrVXKI4Fi09TE0lAL0ym0kAMLL4r3Jxok462uKr6qx7IIFyg+pLKnyLyDIiBRv82S3I+1
5qTw3zjzBZg9jfdJ07i7z+20rZTlDfldzWaXme6ozENPncoPHJBCHBgz0hvZqebJivXNbZI3dD8j
IjOMF/i2waeAbpnqFelNpzwvNGUqEanELNyanAyIuA4L0qfvtllyD8lSPZmNyJTphkvc26iwQ8jv
32tenw+OcEN3Kulv3xhrJeou0HR109BteOLhVVmGCosy6UELaw0BmvX2sAu0XimNXzEm/mJAlSnG
g1w81EAgY95+Rlj5T1Zj9uJsTNQQEYHsj6NZB1DULOInzfqs0ZFPlafzWUr0aR5qwRfEcRfkpro7
AE+lPlsHCWsQZ2qMz5R7r19EcM0K4fO9eOS5myuSloSS8scx1dsiHemNBtVvRTW+akcM3g+wAsfJ
4JAkIEodA8KMK90zgB5ITfkQuHoSF6aHi35QbMraCmbFGsG9teKMmHIH2x5BgZS17e2aeYnEx0kc
GjYGZQnjr6YCYrMBV/IJIPOcacgY2lDJ3pFu/EemiveYEClcz5e3pQ0l9ZNZdrffbGPDKSIm0fv8
iplMxQmSbMv1LCQl0qgQ7Q68a8F9EoConrALpDoM6rTDsOaLvozK4zxSB+WiNGlk85nCx5Mi9LUt
BIRrKawS+YyjV0G/+GnfCMrVcbhMXbWcnIq/YfWXKV8EVf39O5uBW+gP/0eoxXjJwkRf7nkSh+Fo
aCdI2qWmydFj0FkJOJUNqPgMJua7LGS047iOzoPm9JyrWfQyBDEUVNxETbWlBX8vU6o5//ExY4Tj
eE6Xx2s6zRnUGd1W3VXG3P8/Tnwrow1kqscdEo45OcvT+D9zv5+4h0Gcm+1w9qjbWM8KYk3b+iSM
FSkvJbM04/iliX42Av+oZZKi3+Z5hCDlLs+Y7OyDNsk00TJNvBVQZUmTBWjKEDv2Kq3UoWthJEvh
cghXO7V+OhyiTPA/F6qRcFcO3waQMv3Pd1jc2PYzJBBO1qP1VWndWyxwEBcUgeqkpcWrHkkZZISX
z5JIU2aqQsMLx9cplHiDwd+crx6pTzVLi3SvIqIKenshodZ1Zrf86uwpZa5GKbSjVpQMx9O6Fy5o
Mtk179uTrZjzqls9rI33Ix3tyb4z3ESG+OcUQGvgkHAAxWu8Ty3s3z3UK4T3xR1GHQJOEly+xz/3
nZm9MwAJu50JjC/aYrYehiSS4FCRfuXQUGiSSwhmEjXHySnKSICXs27TuAqtGGI3E+7mYqOnhtKM
zo+IC0wWsN3EIDdcTl1I9wDs0EVDkrCRDFCoENsxP3N6uWt2JqNHkqQjldOaxeucO3jTAavYWT2V
9jC8IepZrxEtxFoEgfN6f9dY6pN4zUKStbagDBYPMmYyfvQC2vJE4aGFjK/yNOwi5xR2V+F7BUCp
nXaJ2KlFmL4XuO43f5elTcL5hsZBYMZjqbIzg2iROYWPSQ8td62KAJpozNSJaUn2wlNKiuNACs+a
hcrSFNNoW0HePwwzp4anDfBjWFwpq0H7CWLIuEa2WFGNyU2/W/O6B5occ/KmzFnyW3EwKqbdWHbW
27Zy5B5+cjochPBo2IDFhPmHk0GcTOXdtOdWoesqn8RUZXheD2UHfr58AJO1gcxVOeGDA1TZWf/R
OPXwLjpQFjCIe6TSwBZRuS9viY9iF3DQ4FU7ABwRIiTk062RWv0my9IbV3Q7uDOMCGvERAhMVj9J
tEAHFFt1UJS8M1OECuP0S1T1kPPE4yx+hcMys+xN0hUo3u04MRTOJkytmARxTTpogBXyBpsVLws9
MV29KHbROn/OOoE8iNmOMjSxSGYf0UxXLc3r06lee0Dos1Xw9myX1CqHvWjxnabDSFI0VyQI6c/M
lE7SJd5uaaIJ6jFyOVBwhfzgVzRo1A8ALliszJ5jMufu5f5OmsRqRn9I/p/3EHhSo7rxu7W0l2/B
rJ8UNQWNWbb9tDFc9U90G95sR3RdfRiaYIU6kKT89p5wqfX4GBXi54agcZo8zlBOeYtEGXC+Wd2Q
Ujpf7YtOWYc/TFrNfEtQ3AM+GYma6uRi6nizhwRvD0eWTuo1PHQBt/mzw7b1ugfLaudM1YfvDXg5
GQ1gQsMovVMuIQ8BzDWk8Zez2U+hqbtZoF3CG7Uj/n0H7rrPyX4AX3LWecfZyqExLflF2jKM1XXw
t570X9NvkDZABFDCAM8JTqI5uxc7s82ErepLGmGhEZ7WSm3KY9wf64YX6RFqrXgT9Q6krwMmDxX/
tC/ENGeVOConkHR/IscpKZ14hvKOeUaEJWG8kqO7yo0c7U3IU0vDXK4aw5eZ2vY7FS8hFYtDwgpr
/2uZL4CH1i3WX2L/KU1ZH/Ijyq3kn7atcGavN2Dd92GAHtbvpH3HOZ+2pFCdHlTgGtf5Rz/p6HrT
uNCpccLD907JDjMnea9e8tT8ZR26eoRqoMF2Fuinrf+96A/L0X9gSfG6d1RdVaTPmc0p//Bqmqm9
Nj3mwZMzi9QYPp9yfkov1DDlVnV296m2JYHq3HaBdCmuf5rrBl2CyYvcbXNE0Z3fkBtD2VxbEHR5
MznzdREu9cycWJyFe/R7nlxPGeycx9Pu80W+Dl+BXmp4myeif09vlsNWnrfHU6SDDA/jLUJuDlSd
I3ViqvgVKkq9IdX6ICcRKkJV9vtMlCQwpK4R+4NVwLTcPlxh/zVfOikF8N7RA3/j3E+hi1MOBq5O
pYKgHEjPd25dzjN+D+XvzaLDeI/GkVTDJQ+vcMYDT3VQdfuSeBKDhXDESgGqb1YqdGRLPxajAI+O
IFDfN9YxydFFl5QW3fa15wVAldD1SJdIsdFAJili0wI8qu2w+FjCv6FnYdRzbsaoNpuMgMmfRhVJ
lWYn5oYT5ndW9cSCOX3McWbTVAiiYV8S23nYwZT/sgLaN750lUDMID+WpPvYUDbEnNYFB3+Hp6YI
oACYueGCE0wthuMghAlBi2z09NPdoNbldE12yg/G5DaNfwfgvkvY7FqYRlR3Kirsw0C1Ft4T/XXR
NOuQisIxZz9qgOyNL+FsMoVzM9mZgkW9UgYvu1s9W3lkzhj2YIOflkW2myIFWMVZgngpcZFAjH0P
jpIfOGnCGmayOqwQMplW0p81Mj5VPcXfKGBT88gg1UFLMjS2HgmqEZIDDWl7Ln0BFfB11zVt6N33
uA8iZdOzMyj044VT9e1DXuamOMNSPiref2MYf4VD3TcQxzHLjhYfRXTuw/a3GEhmmicvonlcr5XA
dflabFOqggIA5NV9KGeVNLbcbeonuJgA+bCPFXvZD7BLQQgefUR/HQcYM4nWhUbr2HXTtlyYnIoV
5MsR5rXnFwWvV0Xr2R31iErfe4ed+MT8r2GxqqN7C0audpLhu6nA+dL4rp48tkZf+BEPiOSsOjJG
gpurCzTE081MblIDRyJdyaUGggmn8k1RVgDYjkWeQBQz0qHKzMqztp7TSfpwmcqf5cVIA+TvNM04
syk5YjRAX2B5byuiu0EdG2v7NF49KOU9YGoN2DGKMqYQmVxHHtiYRNl1Oz45IaCb0PEb9F+sHwy/
kFBP4vM9fhGCMZ5/FvC86BIgAqoSSkqC8GadLEtK/g0HY5OmQeOLkH8X3/BwHpLExRZPUsnFecff
RipELbLBEUOTcfktSFms71nnOs9YAn6jQN374vyKtb1dE1QcPLfSw88vYRrSne/+QeBF/sEP+HiR
u4+FAHTNY3haWpcwIuJSLticc3h9jS2fPnvDZVRNK7vk+Sk6YyE4sU8WNNByFt0QckagrrubrJWz
+yzIvuHHK0UyakewhcG4jJi1oP9aLYDjNp06Kuz8ElWuWrQWKVbWeQMwbjPSvXI9Ny3/6Q+6+Nqe
8vRJE4MpRIXdsyeUunQ3d40h/KwEQhwjX8P3yhzgV6YlmIajvrXPyHSzz81PuJcd3UKJ+FrcWots
85FciB9DmbmNo3ZEOPS4EWS89Z8dYTjleNdii3JOxyUYUeYiUUQAVhnoa7IIThen9xzqWNGbsqnw
I2G8gpuCxNhq+I0ZQq0gC4RHXLszuADJiYRillxX6uN7VYvbx4v+2unlhGoL3DuHm+J4vD3Wbgdd
Tw25Qnx6d549BuHjjeLzM9RYDtZNdEEVCl6Tl55MOBJ8Fi2MQti7h4/NGDTet/gaxCqNd4i1BhkY
DrFY1/v3KY0XkiBw/oJ/9isAxne784QlCzSaoe9lDzPe26hFCm4ZHQZME6mccqV/D3OpDIRYXaW0
NNAO25pSj+/ufWDTeRUFzr26K276ZlKsYWaUJrljdwtxko1yjgxcvgdh7J7cT8yewgfaK3tFBJNH
YjYt3mfCQK1GEDN7VIzhBWc+6E+o5KIwDcCU/rOiS+AVmToRn9vAFxEeJciCscYOzlfH+v0Fjghf
gjCNSWvVJAV+gxX2eNzZ0bWCciBkRIFMUTnw5rLcik7jDZ7l0zNRKhdsPCvrk2mAVY6JZvAK9NFR
W2iDAwwLygiyj5dcLivDE65BXX+e5vPm5dINBOMNjokU2i8FIf7TxG3xey2J6RabeS7daFT5s87L
+MYbWOynJYZ0hdYURzb+orul+hBgausMO/ci0wWLEVj6eWijE0zsJPSoqDWJCl0hzEqKZqlSNmnY
6a8mZtZppGyW8U8HoPzPfLLuoUh1yGVwOdCEyMT+9bsnAxxJI0gFhu8Xy9R44lzNk2/8kCXWrRcP
nWp49YZKCTZ367MGF4fWfkupJKOKopfEk7ZAsHFk4FJGOIqwdWq3w6iEGmtS9bKEpA1Usv2Eu/cU
PKwN4kljCOTHvltnm8QAKCAsqOLlb76GUnxwIasNbkIKxhGyGyzZGgUNHOqNXTSGXYtVmFhDzeSn
DpdX3oo/u4qEAxjFoIZ3H+HcWJuk2MvQuaalq5hb/uKDG+muC4lz6uZLJx3o8fH33eMmISsevhBC
8NWU/PpI7TF0hjbOytsM6jRo7aoAZGmHrJzHtWsnyycZgWpArnpZN4agRQwlKH7ZTjPjNtpvmEkC
dY0RUb8UwjKqlJR1yvhbbTEJka5YQYE/IcjGp/FzQfbUf5mrLxrEI9PzyADrxZE8ynJO/iB+YQEp
2kwWjWB/SAPg2TRYobXzuDsisW7wGQCdN/+LOJuakF+0rFca1wRFgJZW4Q88NYaYOq7FS1PLMoX5
R61jeLarOPxsjeSRsIaw5eWpeGfV97i9cpJKTH7XRANGjjkeI/Q3V1bmiJvtSng7IULTSW+Hzbwc
3yOFfl4BbSbJ55MKM+xxI10/1tw++wwaTwk04SXoXDH7NRGVW/bu3J43plmoa0QsLQN0KFEV13Oj
HFIiOX66qSjvrydtCLtuPjKNMugDTZPiFsubEWX7Mc4d/IaJrD5Yn3hkKLhoHVBJkUwLttIPvNTk
W25q22F9W0XEpGcPzdM0vZgwpkF3lpyzPuSOmbvyeX0TNf55Yt8sbD/gUP2pP2ceY85Gk7Utu9HD
bI5qhpgtn/OUIsUiH+cda9S6pu1LQpcBFyAFYgmf+KeWcL9LhqsONr5KosqBsK+1MdYSvlLcBQp+
ygy58lMVQ0If3KyKjVZH1M2CJaJ/VQLgMFHdRUVBpZhNI0lvqOuNqvgCgCoxFrf8Vuv5DoxNb7n+
dO35tGfZR+yHGWk9z6DdcJa/tSRqjE9tQs+EMUvio2AMIpNJ9F6iyrjHcLcAW+zcsel+92gwFQyr
lpvzcAAgRm9Mw2sth+RSBZN5/mS7bClp06bL4lWF9j3zEivDLnpzY5X/q09hHKbv80WJEr6xZ47i
tdJq6M9BVsZ/LmDwyO9K83a0wppPRMI0jV3KUu8Pb+S87HUhBZ5ScH/7rZhS2o/BaxihY3qd69el
4PCBVgimDaVvmg5v5m5ObluJZzpJf0G2UQLyb6C7bc3NTgFQCpZEVZ2L+jcrqpDt7GX9W1KWbJ+j
5QS4xUbYfeyyX+wGqHglf63wMuPOLerH7DUOo+RXKI7XLRqMiYUpWU8T75765hIHqIhdGu2agF6X
ktkpdffM7pAL1pgHBlJ1MVDxhs5EbfSrVaaWk5VeXkI2bB6HW0vtW6SH9WLEEAjQnfNluo16O/DA
/dMUDhpj/XPOBdWFIXsdCi246fABRBBiLTB1xi8t17cKTPMUbUpcesnM77Ci50hDrC8ktVUPipO3
QDGc/cLePS+u0OKcQVrnf8U2Dxqw2wHPHqVsImIP6aLqFVRSyZxnmeGQDDaBNDX1SQZEVczu0oVL
T681pez+oU2ojSgwtbf/Cs2HSC68pLY5f5myz4USYIl6FNThMyo6UgnVFUdujqxjrKzoypWRSpkA
AEMXVauoQN8yDhxT02uCszi1fWbwQhgYk7hO9UyPger09nI4s4VtDjDmzFfdPftcxOG0MOa23NTz
0teLBQeMU6vU+4nlStYP8SroztLX/ZQuA3WieG5B5o+1ehzMr1mxZBzns7FpQs6h1P/NPyuMAbQK
srFOFnK0BYFL6tw7krJHeoMhH3R/AxJi1oE97UnmPtFEDuHwifufHn60qhy+x0FhhSQBnzB9WRjC
Wew80s2eqTXlpDyQav3Iqnt29RoLazJzdT3ScdILdAZcKSNfihrKeXoYHoL7LQNwk50QhESy37YO
Ese4VXHPjZK2jYkmuasv2Gt3zMC+chReNVY4yk+se7jKuHr/Tca/8G1SMb4oeL4lbKVQU1d+wqzj
p0KJ7E7ljKpFkOHazPq9khfsbrIgkJOT+MC72NcUsPp6adyRi1l/wFO69kvKbTwMJqFSW4HZdMfv
oUThdSTky/zG38WRR9lFE3Nk1TiclL01M1lavNOKR0A2alj6QS0oxHwfRCY9XSG1Ya27H06JjJV4
RikrOm8Ejjy7wlBqKTjr/T9aNA4iX3rln3jegNQYBr092c/8EPtNyuhvApC6UnorHnts2+iit0r1
wW36OAdtevCksyaxxvTbQofK2/ZZaam27bC6i7yxEs5NgqR6qLTHabd7BqksMfH4kh2jip7CmFaQ
YXOnRFizbJnNMo5yqxNoLp+DHL2JkzjGLdOQXhVRHqaaPhg/Md6pcQ33Pz/xjp9NYxSkGL0jCh8c
V/WW1YXXZwb6HOUVltXBbSeEOX1eQBo717+7Cy6iWx/3LI4NTnhUAKlNZdUixBkV4j0/d6SWyETj
KVM/PZHZIMnZVSNr/wQVBZh2jpWoMCid5BuWWOjKz8i71Z4QUqrAFDdYv0kFvrA8jeOVXHOb31i2
iSKscLErtSB3geEUhSIr/C/bST5u4vO9XVG1swrUJTwcwC8AKXGD6EGBMRJL1FraTcTiqL9CMeP+
WwA/HW7mmdGCv8AatMNKsMb4ojlf7G++4dfmgN8k2jNBlZxpB/2/7kDbrDuaF5wUbQ+jAsPSBLbB
WMsMuSZ7nb8XTmEBU5Aeik/j3NEGHhIn8BriMjNPQVJlrQzyP3zzH5GvY3xIA7/CY8j59KY0WuJ3
s0pFtSiiqoZj0sywNXOc4xkj40W2tglgXX2mvQvTFM9//ty/Hcfh7gtWtLkIPnVbVe1TNINjJJer
KaLvMaVYbpL8+eMarrUrj6aium1GIJxvug5/H1TxVRsoxFeSe7JkZ+jK/IeANjI6IG9RGHeMO4tT
RbPZzuLky3mxr35Al/UaRMErXGx6+NCt79BkOtvIJ3mmLDTnuDFZdZqMwrNjREpq0f6VSVh833ys
Bck+sI5CKhdKp+bH42WI3breOebGIgpjZ6qs8oLx1Hmq4VdtgVSJbTddVVP4jy8Kgdr3mKmH1PCb
b8nu19oKEcv8BdyaSwdcWjRT+rklFJDoyaHmtTm5o3oBpf7qJcBJjlJC8NJmtEKmBNGtXHYJBCfw
fGmwMU0jxJGqDM/GPMR5RzDx9tgZ3HOrHBrIOAxbZHYdJKW8VrEZ/DIeMsGQeQuqeFfYVWAOzlbt
s6gwsKoflA8fuR02dHdGlVoOM7RVbKT/oj5gMc6xeuizXwRMc0unsDCXCcF3nzaXQDZAnlO3CijJ
fFc8r3vfJazM9+z+Oc1NApFpwi6V+MW3OJcXvjlj1bflPof6Bc3JW3c0wVOsiLAA/9DyHZ6HKalt
FOta7BB/sg6k24AmTsjW/SIYq3iollZIH2tEEtO15jaXLYwZBNoGt4bvU5+gv2MveUVvmGGIdVyP
00OVhLkp41wU7B+DLLb0I/3bSdidAtNCSQ0awZ/KCCo7Qcr6UsxQrq2UCN+8P9ihNUXFr3wK6EAW
9EBFUuwir8sOm/TQfp5aQPd/nk1dpy2lcPpzQG2Xo1bBvNnch+yuGvaiEuCKa4IDH2hDjtdOi2Ul
aN6MvXBy+ptiZ0djdzOfy+xe+tCAyB2PcoWo0a3vkxp1oDO+zcBelg6olx/KtBPBEUeETqtlEZHr
oafWPKFujfGgNTNxI+YesRCjzZLMBNJETMK9WZc/O9wA8YnghGyK7GpKlywt8NKZEhbAgY3oLaI1
3UlMkTMyKPosK+qHC0559Gtx2DINRuPKzLdamlsBHlDh8xxxKfZZNtJjT4XGHB0g/jtf9PVkXRHN
rq2zSZwvHwJ+Ifg1otsl8hR9qLSmEOOxw1+oNRB7QqAH9x0AmFGqR4OJWwNuS5YWJXdjTkRoEaHT
M4Yh3l4DS197hOyKj30VuOYIqYXFpkSV5amRXv9ssL+s7+TXCK6tLMcxjop9gc9AIZWiWBTpAQjU
zJzSrn+lGLm2XVyyzyfbeiRmh0hY2lZ+VylluxKXHFzMVpyKp3F3qtf2D8h8QDRheQ3fu8LzMrlm
egUH2v21shRrMvA4cLDsGcHCqvdKl9RleE5ty15JNmHvw8yTeJOdmDYcj1gF+IvAbSkpdyQghUmJ
PCOrAriDnznp3jHfztcvDHoPHey1UYmNfHnbELvC5nlkUYm1J3VItmo2F/ggcBm69RbJK6gAhaud
66rvXKPARgtREGPspSUFa4x60x5n8hJXEjPja9Bn5eqAePCgkibPEEnkaaMo2pNYErBPjshi5tRq
2VOypB+v0LMAu81zP4ReQKnl4pAREyrKtazGM5s16x673dwer7vcFxviLsqzOgXZyQE4OgKKYW0j
70oGBVLrddRg5/Ps9HexZ1sC8DtDzIGBPFvTLCzbTnCQYyxOYgW0wV7f9I8WEEXCGZbc8daTJbbi
Q5Re5657Xgvyb1MO+Fck0Kf2PIknLOxcw5AFbV8UklAd4av5vNd43UeDgsat6g2+bWxjCGmaKUN9
jAObkK6jEk3dsa+Nx78VnaBFRmOgX/svftbslgDUd0WeqxziEWFeh4BnaaL4Yajs0qKfG/xG2NxG
MTL+1ydxCLMV30zE5jiV5bvDIQhbUqt+YTxweXZFvUUHcPRdYwuuUixO/pDPV/ChXnCn8uR9Z53U
tIUjM/bIxN2JBD9KO3JmjGS0Nhg9eTXWypap0RvLhXu0123NOjCSLr92oTiXS+0Cp1kfKG7JUPos
YGzFiegh5wH/yDSvANR2DofHf0NXW7sXiSl5zjuolB9WP/zn9XyIljUgEScjz53BNLO69HKr8V3L
RFPGv0TGMM+RqeYVqn3T6o2wTZeppwPSjTQf5w0LQrvZtooJAzUfxFskHcita5DdZIjzvwq5a9Pa
tClgZO3lDoY4Mkk+opZppKNQC3GBM27bNZ5Gxp3l8y0lUY8yYY/qFppso1R1PmvNk7RjN7M91iV/
PeHO+ELuH/kL+zlbSt57nex18kJwcrVhiddkppNPmYDsGktbpVOGOqP3wWzD83OAawJGsqTkEUvc
wPfXH/F0+7cPE6o6OcCvrZMwxMpH41eHIuSn7NRbdB0cpj6uAEe34656Ry/sqCqpIwUlqdr8gkJj
8dH1mt1UiwNoYB9rIwCC4rTo7tYkhB0CsLqBITE2cTdcM8zZiExP/TPMvXqnJdVpaclkYfX4nski
r94rJ5VzIIqVxQkP9t/QBHMkiHH+TJQHvXqX2xOORRS7RppYPcnbS84ztc5BmKHCCnBiz+3IVthv
vT8WezJ16krAMEhNUKAA5YZ5ZPVbyH+yLbqt1pvAM4XgddtOUG9M9nV50UcUlAMSpgIoI7q2zDiT
YDT4V5DdFVStJmpq5R5vk0sSa66LMIe+T3KlaDsIQr9e869RmYGJwLqCDeTiD8aTuzxHeNzrTZuL
Td057p9/SSQS6t3fkbE62afzgn+f19Ds//39qwOtRy7kF5F2CdowxqTVZFc1bakW8uP2eIuDFtf+
vQjNPv8f3LXO/z+nHE2Hk2kiUyNx3jZyHwhRAgwiEAT65zCPH1S3wkpogfGCg2wfrw3mlkHKpXqb
w8+Eq3j+QM7w6HKozaW6QOsnt5yGpr+HITFXSSZ+5cr43XUHOrieFZSFWW+00UCSaq4C7o9OYFJQ
OKDF+Aol4MF/5IdxeUKewu/sozuw8XC88YqO76bftokvjnQoQt2aFoWsSUgcXXwy2xI0K8HlX1w9
ccMMM28/pMC14glIE/TjKl1ZoLnm3QZWr21bQRMeNEc8KW7jZv6lXGD7uNPUwlPnXIDdM0jTLGBe
VsBNhqA60NeB1CUDee/OWpojrMxv8AZo0UYTKH9fWqNfI57/U6j9Yabrsw5tRHuTkbYmjcdBNxw1
xYUceLyi57plvBDkYeIZ6E24u2q7NIZfzrenDhxbDYtdDhzPRycaM2rmD4cR0uNVPs6D3sfAxD5g
MCURMzp+n9Ve4W6aH3rGuOAbyosixXLKb64EyRuKNmC8ZeG9PHBuGspBo/+ot2kuhromip0Ljvb0
piFzArLV1O951UVMBZyNyoBf1CguVufKGn0McX+iMm2ZDTmPIojmFzEZsN3rOuPAFgQEKgyChaut
5Ykf9xPxGcFryArYK4DfQ/tNAfOppoRlyHq1VCfDtuiRSeytJQQWWcZBBmN3if2xM9vHGixmwqJy
AweTRR9oJhA1HSbW9nKU0EO0vF+ngmVATWHK8vZXdBlELH+6jbGLJlbAdM7zcZxtIcZWPjoGQwJn
wbK3n+EddFto3zKuOM9jn2K/6QoZXIK4J9252q00ZPAwEHzs7R9RARQ9ihaT34AG5s06K+V3vgRB
/GcPRBq8z+3t+49FpKksgEsv6dYYh0MjZwdsIrbrgSt8Y1loiHyITcx5EAmQWIGCuO2W1lU5edat
0qABmo9ASAh6xBKkwV20rewF8U9Szq23N153Yb95JqgQj20NpA1n/gXsruwLvenv5GEVUFhVz9Pi
14Cvb4BYf3Hth5d9A98wO2eYfnWNJtjYrK7nTojpflzIrzVCn5hfMLE6b6K1rubEy7+jfboNZ5yp
c2zRlhv3XGM+hXVFOL0zsmoNeEodsUdBW+V3p0eGO1+wpWt6qX4I5FLPqxhWyft+bLiIYyJ2sc/0
aKmM18e0bmi4LdCz6bMqPZRaUHsbhdsNm+NNrQiEHNoVOel8I0hhI5E2XTesBgujNvVYxikV/sLh
va9xSbCO+HdHidC4SL67SHCW+7Xf3rx7LkiUJn5Xy3LuWrQkNDBjRc7u6eCVEDumecbkRDNwe3dO
w0fnNNeai/y0lwg85QTHidmbZ4WF8nG3baNhZWbY2PJT9MGlrxpxSqKgPSR0ydWk5dFagopO2+85
56cMwVqiJP0CMt3w2bcTbN6fnREyV6W1ktJ1Cx/eRdcgmsGbOnFeW1KScijImqzDAEjJHvtm4UmC
0xSbVcTVX7Jm7B/bQNPEEiFe3D4tNs2Es3yth0mtBCEIoN3XX4Vo5zJiHIzA2a8ALQZTw1ezWNrD
OPsfzpmfoR0vLCC9OT0xz5UsXmBN/xApjrXp5NAKc52efNJFCelUcZpTShoP2d9HpRxmKuCjruw2
QtCc58YEr0iFBG4xK4VM1zWY2a+Lt/Vp1bucbvW51S1PmD8nOwSseqFcSCJ9YkgSL+YlD0Lay2YF
i6GJLnWf6+MAPLkGp1N3neWrMkT5iPRyjAYTrahBGUiLnk4H4DN2tYUajVGWfwV1pMZnY7XNxian
63xNq2XmzcZDVeyIxCcklIS0+dhrlry7X2pFd69DyvR7FSQ3kyE9ABDpWSVkqCqkO8jV2uIB6AAW
5fX+KVX5Nom18Q6X2k8PECrRCPNlEVKr/lgPfHq4o917uCiPOpiDQWqiJEREQkBOKtdstmUAsdLD
iZ1zHhmOmcSnRS7NcbnCBItn5/b7QKWWA9j0EiAAQi3U6WfVFnYO3eTosMFMLgqkxtMLB39yLwTO
K2QsNIbC46K6bJbhIyshjICPa51rx5XW05isiUcUKeQgYjQo6vSctTClvNnuB17BDFof3UFgIdUj
wZIPZz+rCgxNRNj2RkV9nUjtYFB9v7swlSamo81sBZk8S3zcFp9ZjZooRbWmDN//By3JC1qjcv2d
1m3MShHC7Ictxc0BBOPAfs1OzGtEDMWEGpo9tIIL+kKCYSqGVrq6R68K3M3XxlOXmpenNISras1n
k25SPieaUycTPLb/aVN+1hnMpbSsWkc3T5/6pzDIG6BmHHGspDitywgoCryyQs06y07jFiBlX1Ky
zlF1sZHfm7pFb/a86WOAQHHnlGLTDA3yAF91f5p4TofcQmfC8TBuPXCpuKbvtGgB1H5fGq19zjXP
w+HDf5hr6bge/dz+5iB3AkozxFR6wFnwR/Rm3xabf6gEcxVSlGtmiTdBLAWAVQ46AjZbCwUJzMKu
7rG1N2bfP2VVJOCEdGYT+uz4Td/PXbGqFbH91Ifce8lg7vg4pXV/ptnIRfjF6CSZa0fTTgsdhm7w
IV8LclbvZ85C3XWHzbYRUVTWey2+8+3LCoaAbVJGdWnOgNpH57vDo9W6er+Gu0K+xuuQGZG1UyIO
P7CZK/D3doxjV2sBly49WRC8bXhr5p2CX1Kz3WmFa4fpz06jCwKKcnKwky2svZoMEBr4GGS/lpSq
Dp4I6fuWQ6/J3BvvtUGGNGKbGg3R8JjywPd8NmKIyMJLIlsGlbBIxgoFdLi8LlKo/YSsVdoF+GO7
6aGZmBnScZOowgTg4qDcSNeZ82wIizOeY9CDfn9DgmpqEfEsVd+8RspToqlh6PN/zgd22I1gBF7o
rHyPqj6DQgYPxxkc8XsipdbVCKsV6LcMFUzXyJvDTfaEV62XLSpG895cYYPYL8dZKWXH2vimxJYH
YXGdtTBpsWCd5AYa+f5ticeR6MwvjqsOhcLNfW+Tg0jtH0hpViQZqAwSoCCVz0KwJpfAYIkHvE78
A5AFAkYoZm3+zwChbThxE6xGLNNq1gPAvBNpRl928mc+4Gwr+3T97C2HfdVq/lx8qEi3XXDSVsDZ
/ofraKjE1ueq5lI7cGXysVaj+HbZ7ZewMPOByTd1b7X8GI8pIRITGr1RIVZvO3jYLRvoxVEIB8hH
AO6tj0kSng45iLLN5BQw/9lVNAOcODECiBfZh+4qGN6KnNHYNgGr6C9D++bIEV4w7gutN2CNqti4
Fp02Lg/c7vuJU/IqUk4ljVm/ksEAg6xZt6GMxfb+5AekBvlif8auUmqqr5rvSsWRJMEz474d6ITY
TXiovkioCsErS4Y6XnOWBZBvPGYqQlVae+SsQpzxOv5aAzDWKjVSzFMyyqgRvXyBTX5s0asPvakU
6aU3We6XAmE1xKjmbp2FaxfRAd+bVJ9WVZks/Px8hPm12dJqCskrW1I4MDJFsvUKNuts9IrTNi9m
QEEfiDGxHIW+CIgvKNNC8GXgyztdM0NDsUXVlOf8hTq1zBOWfGLZqbt/VTNs6HIpvdpR8IqcLJdL
lhgtq8v+fyLVSYpUKICcQuQ7H9Cgz5sMkKGccKhx29VGh5QNAJfKehcvT4OtVJUg8QG0evzaXfyG
IWX6QRmrD3POE3NJPWD74umiso4XAlIecTMlc9ZQXJrJGlrQQ6/fX9hg5phIDTpjwQ8ikyRCc7DV
ukROvJf1rLd2ZmJDIB5HS2u1IEK+b3/0oMer9JskgRBeJPsHtnES3WosOg4H4l1nP2JGJxL1FK7c
QR0t61faUe5/drWiCGDofj+j05YpgGc1qa5wMG/z3pzXnCXOnHuC2EbbuvAH4NNFM11evQNs7V2R
I9dK2NsVvUgrlwDgaHK/M+CRGAJcrVoTf7U1re+23ATQFwCuEC5uZ6Tpye4mWEfn5emdhaGheFT4
LYCPgpipKDZzjbGxdHdEiNOrprwcjoO0j/gaJFDSnNCXOss29j4pY/T7W6h0lyNFbu0ZV49NVubj
QbeCJn8nvaEYerULawT/io5nUSujJkP2UpTND5TElUtkg/5WoHZaC/rHyJ0IUnRBWXSI698oadDS
55GrnmRttP73iqnt+rXn9PmlYFQIGHwdO57xt9qEIm4/mQkSLFePvwRC+P5cOqMz+kMWkUSQNSpS
9rlBQwNg9nXOQUMpv+QUQ6QJDeOPLK9aE/MStzwQ0DmoxnWpKHJwICLfgePkTKswW2Yu8A5dbYPL
Yv83ZyyGuf/gF+qN4qahCNj2B4Qsx1IMk+e6xI4dgPr1fdkfDsCgvBscFhediMnYzVsOnypMIxPH
DOCSZMbg5we3SpjPNkmWvxyG+qPViH0Ul5LKZl2Df2E3J3+hOqGgjBBO/XBqxCCu1OjXMUow50jf
2YhICpJG5hW0iRejev6Th+TGTeqFK80pplNfkdGLdffVmVL+1sTXCYMdmY88t8KVFgGt4bL13M3Z
GkDe3HBqdoKK+DCPquMudTRe0JQ+OXW5Mqcko+mEECF8oB50O5IdhPE+PMRd8vjWlxNviJS8c7o9
JPnRltKF0MiQSoTba2g2SAmVlqvtH8FRdXgxpk8nnAzAYqpvtCb1ijhU18+a8CQX83dcN66mIcBC
Bcw7Cr+PfVO5co/z0lR7ZlTvIyHJjARwpWKP8y2ZoRc4Qi4tgPEoAyfxxXZ8uaXVzC5VTkwUWi5V
MHBLUH3L1tt+2hWGYhAtIwuwROZH1nK1bNfA6N+veufxwujS7KBaP4W6GUHg3px1lIS1j4sFBtYs
RWRd1sP7EgiqRlWUsfb4Tx62evxbVDqxz2J4xTSSJglVFWkZ/qKEgI4KUtxJ/rmJcUGNuCOhOYK8
HY32nZN8m5e1ySiZuDrTlYD19D8A26pGe3ZevpPue3spWIk5bvn38McUbazSX8w2+SdTQwsjn1nI
HL+Yd6t/ilQ/TQ9YTmbYwfRYlR+OcgLBPoAPMI6Be2M/66hsQwrc+9JchNCn13Au0x5ZTIr3KysO
dQxjrRWXWL4ZhOcgO3qJcM9S1GTT92LI1vqZ0alTc7in1UalsnX1XyZLgBNTK23SDoaBRo1BPUwM
vN9z6jepKK5CuDHdcfsEjLskXZXfRS+Z4s1XBSQ3/A9IO3Tys0myihhO2l47/iO+dj6F3uc1gVEG
f+Trvsmifz+63lE5qnEbhv+yrfiBB7hjEF6/LrLy+XQ02FukBLXjNan0pyP31zi5QqDTQmNuM03G
+jQnPg9EyUhBadef5qYyo4aCUJcLjN5+PkUF/VMnnjjPqpzPTD9lRqv/QeVhxzUqOCAgG5ARtT1C
x9uPkpgSkHcSCssmSfiz+0ex6uZEo8FpeerbhOnbQ/SBCFn2/RicyKUztFFMs7IYmQWqlAEUM1j0
wUze0qe1Odg5lxw0ikwWr1ptUjQK1GBSRtPEAVQXys2zHlP5B/aNzCGhbp8J+Vo+ThSAECJhCUOP
RgaxucfyaesE352AMuBQDcGbUua/5+4rWkrrmhNY6ZeSzmuDnZSVyMU2GZso67jS2UISkkjYqltz
FAUXAk8JWwEesRJJS2yJDhRntZBtZh/iXJguCaNGmUtWJ6riEXDl9/aWeKa4OfmrD6fnN3NM+4MM
FW5Ch3dOlJQxNtwoCOXIlg8hUhWCOIVmsuhT6wSxifb5edToA+DRVhVBwLDyPWQGxYhjLRPNcJz/
H654H9vSQWK0POnQNnF+mtH1NRvsSYSX+dotY8PHSL1LfTS2cCL3TEuIZRmWM7wjXnz5zO8OWIVg
OBLrYMRnUXx0mlrXeU9MZHYP/MbMYiM0GjcI3dSLV//cwcB0cUeotlkIYsH3Sk1GEcSoWUluMRBg
sGMiU6N27c6wpiJkcvsVwSRsP/fSZddPp4moZcKkk4/w0PZT/ddUe3y0SoEusvk/bs32Js+5d9lP
Fe8N8pFghLIZ90Q3oJlH5K1dCYc9L26KLldOl2q9waSTLFGZKCpIjps/9qLxTcc8pKWOiqcpRzX5
s1aOIAyByb6GaXNSxK04dIEieVlndsKuBuc5W8SiG1ccOac0hwsuSDFyxPfHJk36lpJkpznY1fSd
RXL9WSrV04PJyy2jSnTZD7FlJM3DbYXSbOMMui65wH8sEqpLXYAWrgtbSiqdvR9K9PEyotiOmY1B
ftH4WkOslBnAjE8qqhcimOaKIiapbWGirqw+vQ43NLNX4FWWn11nNCliub/kCeyDDGfhbmIgfKKr
ygkY3psQRSHW7cLyMPzpQwT5vkS13t/yZSKxyCVhY28YCCVbbvvYPJIoGfuMoDDRTYBiXpOdTLCf
vZn4FVSbLlXUUxG8VdvDleNy0AMlX/ljoeUFD5MuEKLPi3XbpkqRt7KgGd+XbGKBUclCx65T5bgB
nrBbI+DDTRi6vDVutriSYWokwEr5n1+J32nZhC7wT41TJ2LXx4HZfGD8JBTPHMDa8LF0kx9MsHI7
V8fhyRZtfTg14kShy08ecOdiVxQLFAbJiQBbpwl5c/qbjNsPdu1dghknq2zj4XixZAvcUujbD5aC
ye4cvxykDjo7q3fhmFj3stwm1TgO71YknbPb7CCC2/Qzkp1og0bo20ZfmuGiMJ3ULqCbd5Y3KX3/
Q6vPP6VKSJubadzFvT6ZXphyWMSJ5VwavHhMYyEC/D7Ra+vpfHTZtAFMkPsWIPDL0r/oGS/htMz+
b250VpaVz0ZXxLp1KucZzK4sKEBbVTyw5fvXTSTAqaEJ4ooR+gXR5GHwVDIxTJZcgH4Xv3gJV+49
f+/JgZches7RGP1O6qIxkDx3HhfiCysf/E9P72F1Ydp76jlHDWlgngZYc/wm85LgAJoCweFzTCVb
L1afojRSpgvbTbLgYT1OQsJIEYWgVDyqMiBUtKX0EU0s3kpirWW8OjaFc6bqHtqKrHXinhQE/4SG
HDHehYqxAgg3cut0U7vTW10/aDu/wrTaZbQqJNsShOx1qq4/gkLee2RIJyDpBj7ejvmW/nn19dTE
oDSAFaxSnK6sn9GgwMPPW2QqJthCEkKmSpH+x40QZQIKQQxnhGH6dT+6zWrZare/WIowOLc6BNn7
ApONi8c++KQL28xfqvRkrhSKvVziYvlhXxKuxdvauWhocuszWtCj8oXUgTtWoW6szK5abF9+9PsZ
aNTK+i2pjmbdr8ck9iLsmIAHoPXlgUG3duhVUCHNHVbYKVmKFtBYrMBeTetnLc8daotATlP58QsE
/TK9FTMOCrhCt6V+Xo5u1FWEp3yQPUmGYBKD4QUTcqu70h54IGlGJqAzuqda9cfxnot69hMpXvpH
q37BKhGZq3WeeS4ZNmPBkBXWc3K4tFRuh822dbeeJi0O/RU7rAM2RKZhogJ9bZSMFBLLuv/7vTfC
NMPnmDy3+UlgRAAaCCj6G2vpiej90z3NJWyA9MVDL03CzVnYAows+RxSV9bqfkC6dGAx4AnNhG0w
dG/xVmixrpU1shPM2EuRBzDMN/yno/RWrSTcGKU60R0pGCnwtVZP8HovJx/5y9tAomrEQRKz2ENs
uer4vRrIDUu/+CAYIUuzqzFGJDQTMd5bcIqN8/noH6qx8PdxeKcg5xWlFUpV4ji2B9Eip63OyNSy
S72luMBd7h5TuXwpZW4ZiOq+VSYgw/1nQbeJ1cJ2JcOZtZr0I/TrWW+DtZeTLLXjycpWOrtQZyi3
nuZ0Na/gsaZqwkL1Z/CLqGozoqvfF6Wd8hR63fewr6SmVwwf/KVYnrVei3DlntRlEn845rwI6gl5
oFw3a5xHCnLM2uxz7gLP9IEDjuByEErUKkysGKUg1UHC/Ll+QZMnINdGn7ZJcLSTSrEpVCd+danx
ZIpji3JLawbO8/KxK40axXz+qtsfeJLfKb9xWkwvsNxQco+L89yu4OqGOEitB1fk+89AAqG2dSdy
4AQBEH6w/nqnERwm7rA+gAeNfnsLCUeEdYLPR18DTQcEt38XVxR8l8EwSdAKxYaQu8F8rfXxzQtW
36iqyQ4sBwWYMzkYFUeLTjF7/G+PxYFclxdsDO3Hq8/NgQ9pNlanroNbn/C25CUj7kZW2JIxHORv
dOUmOAs8XZrQ29PGmbGowulovID0OgmDAk/8dNXgVbECWFh6wC5NF2poxbweMRzLj2VAZzoPNfWd
mbmfcYI8rzEFDVjuPXhHbK3OWMH5YXQu5uznz4jPyhBgMfIVHurebYe6LA/XTUiPRiSBMlgFEA19
nKP0cIrjQI0uDo3yRWn/6K4rdtOd0heJUWm7/q7Wv/ZiGtLDZdPHw4QEpIOsRYCh+h3RSkiXtFqp
VFbx0uDkOOllvSmAUseXy2JYd4OwYCDHA7IUQpAp6slKmzj1y4duiyxI0mE/2oXipwJWW7u8ml1W
Kfh/BNLj3AboLXqlu8Fyl8NH+aZcPKAKOjj3eYH6Qm7J56q1S8CChkWaW25Du7OhXNl+JG2l+Uid
5f56A02/n49bR/zgrg1QfB5CXseZ9lrIgxHePiUWUozNnHswHJWKDNa6nHafeogdmBYdwbUGY3kI
72lPAYxDlKCPZ8XZPODomosvIIv4rZFSBkruUAO0NrlFSm7LsAalLvOoO5pvstvUaAuEQYcvHvI5
x4CY0ru+JCHUapQ/SVChrmp2DOleBgGdD184/nxvivjKgYOTlfxlxxLwdj5Y/4F/xxwSeLPbpTkH
UeF1NNMAsz0Jvag2zfh6HCZZ6xOMFYWMiFu+JxuKWTxxl1emQa25yJkJDefZlpdLsWf1rkGmNA+p
8pQUSfWVbQwn02yvUSTwDIP2w1VrjFTg+nlPMEU7HmYDMLmZdxz17X79ae4Ss84oYg5YjDULpTiT
Ok74WCNFM5MKdRU8Rr83K1Yvr8G0E3P3e49TFqY9dfc0fDWBq0/41WsZdEC5jxGkWTBILlQq0Nr7
fN9CwRMgEZ38DGIth/yhwh73g+X/FbeYZ1qPgNDMqvL6QWem9Yd4FRllIMlzosuxldhG2XAetrFd
BOcH8v1+kN6+I2Yo/AhKbu8Vc3uUoh928gK46DjLgthNfIc2b6aC8GbwNVO5xjK0J/xFqF9nbRrB
dnlISZMuAp5B/HAAnc9On7u34BGVjJ8tw/aMFi7k2h8IF0Vc8ioYOmcJEpGhEjB1zb3TVdqfzdCh
ACqx/s+MAC9s9otRRvGZ6eLncen92ndBFziHIfAGv0jdndzr+PnzCYauxqiFipivLAN8YXpQURPo
PQzJ2ntNObuQjV+1RMxehNa40axg2aP2V/FsyMWChBqaJcGFZ4xq8LlXn/MrKtQXeshJSdXOt2TD
/OhE3Vy54sO6ZvFclz6VDj62CJ0sX35Awh4YOSoF16axrv1sZLD+MxcO2O1fxCUHLmpfWGRirUZW
2IECCEIS60zRX2OAOzAyGazKJmtYEJkdu58+oCWVHiC3WXPscFOcglZzqopiwBm7730vMmM2TkAb
NKX0y0sKrFu/YcJyBmB1IX8Pi3cmM5rhw0Jcc3hdYHZTk5cqHpZ2vTUz+lKIbCOCmGteXs7nQnFk
O/tTCsqRKAVRoYJsCUqupep/II+QrlP7dhBaMhVXJpvilA4tPL1CyhGYECve/7Optrk2J0O/Gh+e
RsPTxLW/RlkIejOM1r6fzjxpueIOJ2iCD+tmooh0prGkEX81tnmOq3yil4DVFESbUoGdzRhV7v43
/oWiQMIAgl34e2qb0OefFHFRtHvZY8mgoIduMOYTyNJFsUU7bRODhgaDYsYyo0XlidoS2EiSpV00
//tQ7bUeQvl6Cr7Pa8MsVT63oHrKbHiJdwWl82RJsymzPvKgWemkgoeZkHA6tnw7bIuOvN0BSyH8
0Q4BACGFX0NYDOIQFUPTKTo4kGvuBvskMkyjJjNMUPEge57zPr49qZSlD/k/WS8DYuAmIGUOvLa0
2A4q3u3trOevgaHIMAQqB7EsT1pnUBPmDfk9PuEBKow2qtifjj0win9hv+HuedIeGXBXI0fA5F1R
ym6xVn74/amWZObL0xq0EXaln6X2GKnX7Uu6DHco3+zIXaF5mmtN24y1hRV2lOPEtZQ8S/39rQMC
oKcZR90MBwlUB8BMEHpCqAJNcHat+nZTq7zF4B8Gn9WN29EFCVGn6GwJTJRPWVzMSvr2hS3Jgpn4
A3CEV2HC6BfBG29cPbPya3YRbuVIKWQzdV6fFSiX4WZwdjcuvfX0HIeKobgC70guptOATLckOTSc
R301fS7q/GgqsI0iBiCBcbUJxRDcL2ZgDC1yb1yBx3F/QV4cWG4ksyK6Ag+ptvC8Kwy84M5qb6mc
8RrhkMCuKpN8eNbR7LqIBlAKW8oTRHyF9USKeHU0nwFPwiM3cy+dEU+UvMiO93pcTSi2Yhrz3CZO
jRui/7gc48mpNRmLRtEF1r9ZKTAlJoH3BLk4DAxBLUYR6IMfj0avLIgxSnWSck0u/Y2mxHohv5Su
blyhedPHEDjhffeEPH0uM6ROl5/ShH9on2NOQLKi9GUXEkx94z5WXGCFj9z57HMbBIyo6lvmqGup
rbliRE0+1F+JcUvfqurR9NEUL+aB3JuYF0Ur0pKLmTo/SuRIMyhdKKV9mpO2a5CI8obdIHJpYTJi
7+tqjUehlAwtCDLwZUO/+mq1wYwglwx0UAthKgB7J2Cn1fvA7wrn4nDoanp0/wUltOSG/3gaadlL
9GU9R1N0n+UYjg75vk5YlEU8Z7Ytn9YH1b6mlsc+7j4Ai+ltR2/OrKvFs0U+yaoC24tSRlqDTp4g
p1iH1KT7hYORP5jeLocpVEdI/3AjboCD+7BsAWAbDlLoxnXUU2uIbmhxAjy4H1Z29eGsQgZqdk4Q
s5luPau414kyhLr6IpFzX7hPdG5nx0FnuRtRdv7aefKYJLqeyhQSb/6CE/Xevq2cFlC7/1v+WK3F
JmmEu34S7/74ukRNGXT+iKtZazew1jpkiA+SnfILlqtxLxgP1wcnWvLatHkqt/8JRkTrDGNuVQkG
4fXEOMLl7cdztkDaLaXfPv6Nby9LzE3bfVOOIekPgXpixZj8/MN6eSXTkU8Ewnrgi9B6lkNCGtwD
6O7U5q3GjhcLukFOYjyC9HmYvPmXMibMs4VPHrkAQiQaILh4q1yl5Qu2pClijwraJopjn+Nl0cty
JjhbYqF7/qU8nmg0O0jg2BIFU/5QrmMzuqQNek9dy21U1+7mIIm4evQUy92kY8RqCL1Mt9H/GV+I
f1+mKqupOnrEg5XomvuAmSSa/mq3AAjzr0c3TthqLgt5sWT7rIEnyfJRXPYMwuu9b9mS6mq55BGP
DIDW8kx5JPpXPxdjtRPH0yGQWw9FsZLVVwSIHUnr5KHMcep6nscbT8ShIy+cSny72WIswichITMi
5C4KGZ/LRMFPZWTa8EoksgcgJNGrfzX9UghrleiGBWJeF6RwC67QdLuQXdsup2qwiBPkqW2nxlVN
6mSDfFjXIMUz+BvPlLEfnJFzO2a5LA6eZFnChrnc1ELLyogLMLF3Ne81I28wJNKb/dY1YuImo/mC
WEacJbKShiBkskAm0/581JyiCJFuv/4qnsmzEokgkyOYcxOTC6wfQp4Fe2GoYr4R8sapuYmDO0+B
+Q5qyJ+uLIEa7m+BH8ydYR0+W1yBwrJVwfkdj0gF9tyv8YWqWJgWGp0xb0eZdX1qmgKYMhsAaweI
PYKSYMWa5WkMS5/GX33xOU83BfSexGEONL3GT0o0Yio0pyqh6t9gysWcSDl4iWiDYmcP6YGJlAIU
CScVXJm4HxYDk7QiaCwGaKE/Gr9fSudALpR5RXLbKGdPMkL2AezaN0GM9NRlNtRa/Nd+SOgUJKip
X1/hPC9Z1g7OqPBGfGhsVrPdNRAnjYcXAFA/P2LUbXpO4gSByvhXWFKzn8zlVGWvDSMupb37yBzS
Hq0ZcNRVRYYOIvYY87+EJujHcuXTxAB15x3RlD1dKTOKQLHQXfyUc4w2XxY4OH46viOmVnXQJ1O0
h0DDKmgyluIn1Ft+KCml/XBpF6/aER8h92vFX7mzr03Ii3V9Si75BESH8FSgFT+NQ6h75xcqZ0NL
CgqjnHN7LZd7vP6kBBQPZPfRdCzWz0PYQDaGes4pFCDnCooove0BfsVNFnZGm750HkM/rQ6PYbJ2
yxbCtwvbKAeiC49SzJVjFNHW6Ol2OYqNhzVpNz6YdVv8yt6h0DfwLTWNjvlVb8WMhX6TKqNtCnB0
OVMjM4n+ldPYJYbfOHjC7qDVpeaInvVrBCeRvH9GWAo8BiLhq1MiXAN8l68JP/B4DgCVdLtqYtyY
mrXNcVkqoL7eHTakyIgDU0/1ASyDJNgg9ItU6I3on46M+dAf9VMNHPpmqz0deC6plJDX8ZsCbzqi
3FQYp7zJNccmvmbGTMMs6D3sGWA6zbGFwOEl1cuEjJ9H8UXlLvJFYrcwBi7d1HUI6w5ZkzMZufsX
ZMPVfn6CP5CDKuT5xOx4VhQ3LPeUphm5S0MhK4KQC1n4fsk3rx0jnQlRW6+RwaSlgqmAJAIlUioo
jLCmplSqMdsySKJzCz5FfPP4FOTtBf8YX6l96sUniANArzqyZB2D+6I1vrW+6w7oDe8hGWcUtvFL
78YZe9pp5cNAoQwRMZeJjocoQ6jbJ16ASo9h8VZu7oplpiEodiMBETAII6ontnsDH8tdcY1NVIot
4KzBo2mv/HgE89neNKQ3WjciFtKsePbuaLFTWK0GWv2k2TAi4tb00Indqg4xktL46L0lIJgo3ALe
IYYXqB7ZG0S0lcMovat4t5RTOxh1eh1lyEFUet7/9ljgWXtRMIFqL+jdvF99WCFHFOp1IZSF+Cqw
+SIodR+GIC0zDQ0jJKTpbKolFh2RoBD1+Kp3D2CWZ7yAVa6qYKlqsSvkshvWfVu8WFLNFRytfAHZ
2rzCqW1dFElyW35CGKGythD0SXo/cD12U5pXJu0yEZVmZ2oNhUEM9Sv4YEB7o/bQoOgHA0UErJVk
RoutHW1e4Dfl3A/PAkJGNX1IO0/fQT7hjrHHq6I+0ulVC6HphqJ1zlGqAXlZNR+AwsryO5UsavRO
z+BvLo1ahjHuH9TGtjSN+DD13TPdHIsoZkGGrGKMd+AlLfU5jr9t4tr3ZJkeRQq1LWl//bFSNe8H
Hi4hV2ismbOa0gkgp733TASrV4KQyILrGMO0lYOZozrnK3KOAO+qLwhv+pBMyGIjNLpYWlv3rb7o
xtG/ie7MaCrbTJQ5zqEOk6CzbXEtV4mCtCCqiipZFiBYH9S6g7Ub0h06+qqn8LrApA+KaVDLm2bK
NKkbn3+FVUFVdODRnbumMtcpsvT0TllGGS+1/BS5c/SICWmbPgOhYP8J51xLv9AFuPgkpYSyXFMW
/yjKNx10aWa3Al0m2XvsLBUT+VZDsiHPS/9lEhU0GzzEVrtg5tkP+TNrXsqz27h76ACrQFNofK8+
w6+NoB1dXc1SH6wuffhJ7tHMOMDD7liQwcTpxOcwpVKoCjxgIKnXa6tKe4TZSX9VavEFzWTFzpBy
t/ONsL7YWWlchoJL166xEkZWsdV8JizLJjoS061tSSmchQtkMw/mtIfBSt+/kFfo9kqBJatY+iU3
gxbvB4vxpPcTVHorPNckWIKJmVWwx3GXJLTJYMS/yCXrME4OafasMwpgWlmjq3bzF0lWmsZXEWmU
uG5IUf9KUYL1VoytiwxcMJu6bwXRRn5Yjm6gNuI+W+yY8hLc4SrEHmNNtrahNRiJS02JNEO/72Fm
601kWhWdjJ1CYZ/sf4xrX7/GV+zvbRZKxAldHodVk10q3Q7WFCCUmaFOZbBWZFQL8jaDGNZEKlkc
vgaG8AOT7NrVwG7hRI7WJ5DbR5WNW7KMjDuEcVcwxtKvQUmlS3qHp03txMpViEzik8CIsJvqA3nL
Z390acOqRRuTIzeocj2p55iat8t2PIlH1SwAkrAPKbv94iYjdUwaMTQrKoFCC01roaL54iAd6XPK
cuQXTKPf5qqjsZNb9klPt35yIberUmk0CcaGLUJfitpN/1QrrI1+ewwLKLU/qF1/edR61rHHjqVV
ZUKWYqBB2zaJ0UAKrAG5FCJXkVnh4sIWHb92TDWr6N8Ljtg66I22el1wV0PR+JAkOnL8270X1sNC
3x5mALG92O1dLIiyI7KspbB5/93cdfGDVH3z5u+knnQY97Sfy8mF40Z8PZxTGHTf2wBsjZHhsXJV
of6Thw50qLpC97gLT1mE+MXthoAXJSHgLWPd1noCheWsLq8xn3CkfmJ36G3yvMJsqoCdu0h6Aajp
gyrwhr4KdkLgxf86/BFu14ZOdxqgJT7ZmNzNoV/1ya2M8QxbeZXOtCyLKvoJN93+xY6zq4Oc1NY5
W37/9oLDJcvX+hD7CyBCVLkUET9bR/VpxsyRV0hJ/+zCTvR3shshAhfPA8/n8N93188z77ea23W9
YwEeCL+HZr9KAcq/A0aVlHFl+AnKANFDA2gq5w6bbIxWY5WEjY3UTK4B6s6FaIm8xY2WSEoj1n/0
ReiR7XuIsfoEaGCHBt2/EeVRMSPjj6GurMvUIJOXpD6lLypp5+07162Gyl72r7n96Ym1NiUm8Ld8
Sdwh1D3DhyRu9r5HD26IDJ75zDUr/28EBouKpoKWFTqloMYcwQlkOHzepKzuKt1TGERld46OcT6z
Cry4PNT/TYDwN50K43JhRim9mDTguZ3ViHu1hMJ+uTInt6JrnWxicVZolKeFYW5WybRZlR08ZYoI
2rwtT0fMxPXBsdhewwfKTN8FSqczCScN179FlR4u6qTJA5tymwf6LJ6mpbSNi3Jam2+WwpwhIGWg
74ZOo+T68ceIJvsXI3dtwXp7HJ8agGaqaBF577dAsvs+tZyCfj6VyqMpyXj+ug2pQ8TJJBw0vcyE
l6Puwnkc6GvvzBuKEYCnMWupzWP69GSLjDy30EIe1MZRzQvmUtaWbUS3ZFy1LMQaJDi3dHg/fk0r
937uWvxPZFFk44cJXJ9xzB6saiMQxmBtoShDmUYO0htxuzIBk5a67QCTPe5bjmQFXA/KUMYVddax
Pp/s8VBOlNkt+UDrtVkwjD474T91ATbYcTlveLiYGuqzvn1Amg7olOp2RJn7/N/akUaqV1o+x2UH
h31mqIP/YkjIV3XXsZUiJroPAsKd5bReigW0WN1oT/7Fy3FeFPVywu0VYVzb/GUgggvI60ivBTjW
OtIJTEpNHiqQrsaFe+4TE6iZ4J53SomkHZHswqmWHlw0BEzOHtcO+LDHIUDV9sAZL/yUQZ5WTcPR
S+jByWVbSdmXFRC0rRZmu+92uDPT8FZ13dDSEm+42E2br4eiAiiB9XzsIHLBG8v4FGmHklI+GV1b
e12DTTkfafr9yW8Mljdit7w7DERaISMq+gJN5pflB3ZE49054S09k/lrR9sLYC11xPOPDMssquFc
q+ijViVnAtRWVmDG79APKqUKoogc0DA6lGVbf+p9LjrBt0pAP2SzC32KtwoLYXTqC1Ow8xhh3xsf
HLhQ6zyX+F7+vPz306iXpoWkSID2YW8DMPiihHh7tk1sy1cIlSjWCJ99R/lg7cWK4zVKpwjvNo/4
PJ3+ClF6npQSOJ+gW1ff9UMSPt+Qz32vL6YBkOzOpIbf14d27AfCPek3p3wpa51PU8FRin4t6IrH
Ei+R51vUhwTy9TSiEQhCM9ObGxOcnkoHlGyRnfcR+WBGEJ47jBpdwpY/GgfI7V9OGnVp/TBYL2PA
RwFv13MRQ6p3TCdFQlroZtZK6GBMhwtxKmtv3zGi61JNT0Y4QucIbObvgj93I/aGs+iACZLXHcx7
9eHbzb4bjkTwUZgSZ44fof+6YOQ+lYW9Ku7BC/qNNsEwDbArbCRtGj17zH95jL63ipfsJberZkAq
k2rfWWcQiu9N0r8gbFov5UjgVKS6Lx4torZfh0VrO3aF0t8EW0z0yWeo73yrbXdkXPm1cnJBV385
F6y2y2SMngVhaMGVLd6QUTPuuHE4c6kNNVl5udWz+Dq3q56DrQ6SLnvoOquX7TvJEXpJU/bsi6z3
cRcS9rUPG9L4yGRgw+8Gk4IgZk7gIMELeRLvVHEVcTXMzd6l+/GGP5rbSVrIVlxHB0JHUiuNyath
JAra+KWGSDhe542ecZbQ4dExw9zs7G+d3Gdl7SlIXso5UQdGsWyE/X03yD/SOhcepYJFlvOD0nku
Ttd7HH0ZUgSFxgpwTsI3FRTNDNi9ZBMUfNSrKvP0Ykh0iJHuFaXVI9JonWWTx4A9/PfGgDWElcnP
HIKMRT/uBynwV5otlW28CvheZvLJODgndggnW1FX9zpqdURXmu2chwmgXvQOwYlu0tlx2nTLMvHn
UKBLGDo+Y5P79vlOolgzRTfxuzj089ROHxw6fMYuLSc4bm3d/guC91B6r522c41K59KsLN4LS4Kk
y+BmNyavz+HbFgfTYsgaxPj9sQmeFQHRtZlugdSW9WTusT16nhO8o6kJekhdYqQzzQfg23ABEBIi
NpNKAWvPzuEoCsoTfjAo3fRi0kPCiSXFbMkyHbU5P8qBxuP8YPpmKZPFpVFgLJzz++EPZDhNBoQP
XPQXmTtQUMhWUbNz4YZTHCIFWZMGaOpOnii02Rtr9I6zqsK7KeUbT9KnM4NA+J0w5iXSRGt5pBh/
i125eiC7UhCWIzFE03f0Tk7lYeXpan4ROvY5AQKobfvPQHT+egiHssLPOz4TeBGy3QB8oboWjqF7
7z3rldxfGYRsXLOv9VuvGOAouiNkiDZapYUMo8aaV24NyodYVDHWjmFSPMNORiif34lxsHPwYx0/
w4BDKjYmGonqnWkGqdG7TwctNddgkP2N0dodDLMyJXh0clvOt171ff0FFw0z19TNniZinNOFQGxQ
AQh3bgE/CGWcJJvGgI3bpqBdTa4qNw3IOnzsj10srUlpl0HNb2sBy34/bGK5ezi+qqE8JniRsrlt
BwqzGwG5sK0ffcsQhj/6cm6RxtLh1P1FAPSbAEcPLdFww7WW39dQTUPYQVEDYaJk9djpcqt/dIuy
JA0A7+hhD//y1XeQBTk2BefQGTGAwQLrH1DFdKTE7ZzYwIaGyy30VrJBuV6HiAQJ/rycHZNUq5rR
2+FgU5xq4fb2qLnOTjZtQ2q/JnWPibg1hYpZW4fEz7FqMviRZEHyrfi+gPi1lahkC/e64dNhNNIL
aqmIXx2LPUVN3kiyBcANhR1VhBvIGzWIrxn0J8kKVu5dHvR1pMSzRweQFIsSIn5vTP2jZhvDNeOq
fPLYoebkdI9Ri7AQfdJU5+IR/5rp6ct2kkoU2RbaFrRrrXmpEmBc1soc5U7+FKWbX3wABgxLxEvN
JYTIyzQYo6mV9rwqw3hDHypWQIrbJCCjWKcghf2gIOvrNevt0OKx/goW3h1yWWw1c+7ZaYmaRxHW
WqQkYv5/XI3t4KdSG0zrf4dBVxni6pIpeeCzyF2R4T6EOfePo9bAfDfmzEnkNPwk1yKY7/9hRGLm
leRznFC1Tig1sb2gTttCZMmoav+xgjp88RAL/35BGthxJ8LhLAHgagzdqo9nNVZtpmy27GbqRaYO
daCNGm9RJWY87mwyrQS3vSJUG1VUlmMFM7J2dcgBrCag/+4jmHDJWZpPH7Ttx7G9l3nvDLDhwnvd
TQD+zW7QudBOj//eShRFqecJen9/ic6+ydg82zjFgRfHLEtIR2WUzofqFLrSG9Bm8coa2Ys3k3td
v+jgT+xQpvJE1M6dgEn2R8A3lvCl6R4F04QZFGPs4d1geUXIB9kMWu2Zf5CvM7tF/YqJKhy9tUrw
P5GbjsG6QJXnyK/O3oTKTQ9BdHgo1J3gElx5E+nSm8Qhli2cP/4VwoiI5Ictvl32cjPtUqzvv+mE
ItzNrNRb7xxPZA6Lf1H9+9NgZCi77e6nLzr+ErqeZqkEReYMb9snLVahyyCRu/NoMnQa8ktv4sgM
4PqTw/aoMLGXAuh08MJ1DlE/S4NYDqfmIZCY7bN/XFUUdjWCBraBKPDdnzsdCJhwxFUKdiaX4Qlv
BY182McMLWNXmBrLRpPs+WeeCpkpSClhX03lReZq/cJ0sOYaWV3aDx50x5lJTo734gbKMk3YlKN7
X+ikwDEAtZHyOzim8r4/ZpZhNAbvSvdWrB+CUXOWRvQdAuS0uVTnJdgQAD7VQrzn/2kp0HPxbgJu
CYLR9e3qWA5ZxW1YOwxXvoJDpT5sQJ6b/ei5daa44fE9I3OsfIN+ZhgvZYOZItYJqT/rRcbKQEpV
ltpYCOFQYg8n+tJr+Fd2u8n12g7TI6xwADSn/U8YmnnjcJzlqryn21TSz0o9mHExvZfI+6Cua7Zd
/wW2j6Onq/TMfb6CBt8y/kfqObX+Owz4rPNDPFK/SmuGmrjdiHbY28YWRu6ir9XSGwR5sd+BA82n
GhfT8tgKBDKYPMfZyg2toWmIiSFucZ/tZrQhJjaugQvlOqFgusED05zlPlePZVxauqFG1MLlLJL4
byqjpeUj6aYzpnt2sjLzYM0e/mYx62pTvFlSvzjCt43vnSfdqk9n59MbLvK+sGnoU+Eh9RqoZUhr
R4aA7T/iaFH0NxdnnzZkLwW8nK2vpDoZgNYb5i7QBChOiC6CaUEcSQUjaKiIPO8xuJJxJK1uuL1D
ykHfSnx8ZYOTb5bCG9sdCLMYsGJFLSv128HVXEEV5ICGC9nyRwQwA8fOcL1b5g9a1gkwVooskV0k
yXuLkT4QU8Y+MzHjeHCcKMkbOJ77yr1fpOcaJQTWWXo2HOiwcgzwc+XLOSXj/nX8r2wDt9vgvI/z
1sG8rqjSsj5ea12XU5K0lS1JjKNsYYxniSXtzpNbbhsTdSjNEumxeuPPc2gQQ5LWIdPvc41qauV+
Rbt1SOkbR0AOIqtoUSMkOJfnmdqigLid3B7CZhsHc3mLVc+XMzffQUJ5ttaD5pBwA/9Wyk6tpHfM
FXMqQFCnbl1WiA4+zqL2zvI9xNCtRmIEZaenNxkDRn6YVOlTHdJ/YAAeGrfUfRILDE+1idQk0J2A
dO7xj1jihy7dPQRbQdpCon5gzf7opJv/LtFEcZfOziq28NvoiyW+dGM6dcz8pRaeQTGRH1BN9dRe
i8PdBlBUkkV2gD/zv31nbGb4QC6sr7AFSd6pNj6zrIM+8uwxuXi8C8SpT4pSwOytVR99IDbw14jd
JB5SRSaFk2oN4P1LZscdYpDE9jLy/XaSTmV2g2bnIJFAcqgrZitsuuRtapAWkeG/DpEDTydMHPBw
z3+WUJFxKnHN37YC8e4PKP1zxrdtOvYfkNFiZkhh+YPYlgD8HwxQePiN4/vudhIHFYxcfA3c5Mrf
ViUR0c/qxPrRE8lxF7TqP7v8mBokWMptlOgW51ITbqnDqNCJIVKDXS88xJy1NBaE+s+DcbekjDhx
0SzZMI5LnVYG3M/G18vp8EPI18tWqv0KCaMgCuBAZqioAmh+oBPU2STyucQsHE3lqivaPTThueEm
w9cq8FwdmtftpDZyonTnhuynbu21O05Ufa8t5rZcNf1KfBD1uKcPEJVFpuOTzQBFcrumkcmj8Kku
SEygtGCxu23OMx0hL4+/Y4A9GwBagfYqMqm468O74mmQeWeQgvFwxoL8qAUYrzzcx9P754FO+Zic
ZoQUUWqm1hLlBjPonX8zbotAQH5GE17qQh93y/EqbixErbQt9ghazaAM2gVn5j/Na/dd8120WUpQ
VetApanyqqZoBeVUyxkPa0EuIXHm/yaOkkdDGyU/3I6uyiRI/SXjzZjryODRPMUXtzbbAXItqzUV
54c/iqsgYMOqQWODENDTTKaC99v4pEeKQDVPpvE1XOelmgkoCiooH0nyhBXUzba+E9tmBBO33xcs
T/Jcu1EZ23XKwMnugOykllgesL5d95NVwosSAAwiwu+AQs6ZM6Kk/yJOvrQS4++seMO7gH7w3voq
a58ooXPyWR2icdvAG5cfM1IZlw6D7iazBEXfAG5OotzJRRmQT0j//07A0am6+yT4Otv81L497DgE
VHhNyxDQ7h15WbW31VEjv4p26uBRQSXLOUP10HDmG5wcDPXzBgPCpYQ1pOflG+dfxf5TIzpFrGZm
A6Erd7T5SBgQQ4wP0+AdkS3IOk7fL6AECZj62G3OmF/Si2oxWx3Nb6e/1dFU3HMADR9gkJuzHq38
p/tAd98QWw59OULaL7yrdrHJBaZ8aqiroaXphsXI7b90rl/e1al3SwIW8zqk7wOrgFCWXl2eulnW
sXUNML9EnYoM2IZOWaz4ch+Cme1KC/ZOCmGzXzjTKfKAM46ZTw+FZv4jJyTMUivtOPhgsDhO5yLW
8/XqQPV4TiX4PUocTb4WXNt61iAhFD5QnmQrt0W8gaSvP/yrhvxdNeLaXdc0WrjkRqGrqKIA9eak
PDJJPHbc3Rpwck/EuYuxE/PuWKkjo0WSRA9DkpJM+MzOMotGsp2i/AUZgrw+lkQmCefR54kW6Wi9
EnqQORDbU9jjcAoOMyI3JZkmy45TItOQTQ2oLrXINTs9LPRx5vxU69NBghi+KGa7u+88SNku+HHr
k66Fdg8sLiN/iakBLofyk39J7rwj5BoNHbxN2sCl1L7Edpk5UIAZmIBaR6vLtsEu9Syy6BA6HtCx
B1KwslrYSw8UjWIAp6JmrOYWKyFQYRRspzxiP3OdBKblwwZ8JyVm+DyaUxfEffW0srwNrQckvlZV
YHXsPa3qNhR3CYtZXw6m60g+p5DmjmnACgX+ZD2wO8zJ99RffHjgS/WREnQYaENRCfP44S/k5jG9
s/2T8JlxC0Jlg85HDBCswtA0OMXFS4XgOMc2B83o/rglyn8gSBINx2Wc2YRgBaKGnSzMNm67lmBm
NKcA4+GcUt8CBaNvq0ZtrsVQq0akTC6HWzj07geqmvl27Wd8dP+3dENw7Odt3FEuu+7axsXFrzEM
7Q9MJwTY9C1k70usifRY5csewtD/gmMiVM/Nxp76JzaCVX+99gNnPuX1ae4TrLkDykP2+PhNTfkl
ccd7gU/e+uRujn+GpPk+AhklsdiJVtyIWXl9P7Gbb8otlXPom/PHP5y10EYjSmu0UD1yVAuwf9FQ
lez5VdKZdY61aaYiYoPgFV7CNF2eieC1xSrss+S7n1Ny4XTWjKnBnS18YZyYvLEGPVZzLPyfPb3U
Kc7DvBY0QlO+3GNxTBakRw/Wn8PtdcUD5fiER6hAWSkbd7RWNMLVBR84xWdKI5FyRk10hjP6bZNG
rqQKO8pzUPo35eTt1BwMRIbD7+MlRSxgFiC0lWQezp9P5V6uiud3mjYx4/rqQD5kMjbafGClbFK1
xOTNk/sk7qdp6IpqcoyNDB9e8GSK3TlBSgZ+1L1OLZFYEKVrbUkB+NtYhBfvuuHpV0dwQmCxRQbA
qVmSVvDgNIJOFZ1s+zmzgcARhi+QnyT9maTv4G1827JNjJK1gK/zAy8wiU5Yp9UlJS9RibmH52yO
hl1mWt79LYRcHr4gMndtzyDO0N1LP2XBuNWinwnfviX6CfCUHGav8gHooS1Rys+aiG2jgqlKpBy5
BkczXmzQA1Wp+yf5ObrVFkVSt0mnL6zgrCfI4g/Ojdkng946Xv2u2oHgNFi9attGcnEnw385EMp3
RDFTMFpoCgLlE3HLCpb08+f8zDDgbbJVL9OMJkMzZUmYycVxPgxrQSS96OOH9aZkRU5A81GWIcan
ELf465hDOHzxEYBUYZeoi+MRuLzuTz1XSv403xIczTmvmOBHIyNyOZ9L9qEjF0UWJefxWPFhrHLB
ZZ14qBNBQtuRuIWQF41/zWAV0Yc36Lu+r2vkHh9UUYrqYHK7QUok1NB+oPGUyt3gnsjYa/8dqnDi
XUSxC3q5Pd0JkiohJvHT2YOncazAiRXaQdiIBpsh42t5CZaEJpPldzapbnd8zmq4yVOSsHfADehg
rRQf8s7C+Oq2tJ8CnNc1Dt9mD96LcJLpQD6Z7paBTvnJsbJOSyJU8z1IbKekObyAGWUhnH8jG0CO
UF7ZVRJrY8Xai/8PiGrFv5x7ZG7Q5EDiRrPeTw2jQ57BICBDv9F46egjUpCqFl0jG1SI8OKXhpBM
iFcaPQ68vByIh1+0zv+gKWEcAAPefuORwj8gIcQnGLUsG2iD5EgMUIzPm9PIMqGVrvZEw1523rrZ
rBmThMKk3YgjP0T1K7zYXeSq0ESr04YAFn/+Ekk9KSFf/T5w6hM25gfhKhaKaxhU0ExqHUKLlXOS
HaBKm+Pef0+uZESg6QaeYJOkv5LpN5ovse2e0Cnq+BfaF2B8mC47yPKILVOkKZJdxoFVXcY5e7IK
mYnW17whz0ZcXaQNfOWL2uTZrVf3ckgtlKqc+SYw0+bRAur4j07S3/x8qDC3I8xGGVXiSRWzyG1l
ASXjQWjU6rNXARKDL7lxL8qcEjNTHkmGI0h2UMPlvSgD43KKQdDCW0pzTgx0Hi12aoe962FIcoFz
99G+kxNh2X4YmETI5bJmaEdYZ7xY6TeF2TkZS/ujsmJlC+r0/VQxKbVCn3SHaNp7cfa7X2lTBqNy
iyrb7Z4nI6l4EhKgcI7uurnDGmc6FKQqSiTmpHyxFUZbUsGyeQrfGChWNkbb50nkiv7cG60MIE+K
Ibl3m7L1xWnA85c+a5XJEhuBf+b9IkwJ/7OQJPfNw3cfUY5hTnZeogsFTXp4N8HiZA4rfqqYIV7Q
PtCSlFLux04rShOeMi12UHdVtUXhZ2CmN8UC40Bp4RJLhRREqnVLK7QqaIfrBeZCmFIPrAQYh6+/
SJRqXTmvYTZHLHB905C6jKCUfeBs2t6AcVYN1rMIp7tZO9bBs1glA7f6HnODGLz+0o0N9H0UkKPd
6RhODGrMkOnhHFc99EiUKgTtFtfo0OJNaMajZsPS0dw1v7a8Sm6rm92nT6c/bdmkbfCseJ5vpD4Z
Zpo9YD6kWp8PfwxI8RzQRtGWHQwq299fZ/i/qK3r57VvQi60N7Z5NA2YvH/wMoeGhp1xo+Z7XaTa
RD+7BCYPbiTfGtQHjFO4YwsQIS57X3XMcJCib9pE+d7IRfHSMJMQpLA4nxZbMRSw7UIu+eLzBZum
jUYhJcNJlM97LKAr/K/gyjs4sD3JugsLjqlvGERrx8TlAea5YWw3d1/O+yKuhvEqNBCbnCzdm3jk
az7GXHjlD0HnwAUS43gcjCWUMGG5apwVhbZLRSdwYUDR9zSJMQb30tMeVvw/+3vN82V5xccSftKB
CMiZvOipWBO1ZU6ByvoBf18tNy9WeQZNSe0tnBxdpipPQbD8X9a5do/HSrn4ei11nWYq+GTxp3rB
GKrp/BAAxVl+G1cz7fhhgj5peOwTwaupn/4RZsZ+T2AovbHxTaKi9hAVWkDzDDdZwN2z7wvDAUvP
ExFpNvq3gIJzWNpssx/tyl3uRewSz9lGW3ARVN/2+eZOy7S36XWYLjbHQOc3MocKBqdPieVd0gtZ
yVMd+U426S9TsA1eAmm59UuToBpxgsmZgcLol7o4Iw41/0v8meo53QqUh/0VKhrfGyzL3iHTAhZy
Svc4ugiAruDwLojEwMCzlv5WkDrSftfGHBLO7NkFFIwcZxPxQR+Eu3AtLbyw6/25TLfPvZ6BNn7p
awNHZX8HKu36xJ42ksCjsBgcUCpFlINzZdpRhWml+ZzW8Q0Wtw4u1gp/O0lLR3ukBCU4uM2iyWQh
EvvSNNHi4jOYk3CcHOIk/ZEGT2oWc05aONEPCHYsA8xxdyDI5DmB9ue600LY5oZdO7SuuPfNfPvG
fjKtpsG7lZg8Y2cst8UsgFLGjfASWOSv6nWotJ/RW0BosKgZsCTkrXcJzppymyadsztigGtDGShG
jjrt/VzM7ISp1j5MjEEgx5DlsRT0REcO6qcS1xjvdqsJJj9eEuBs7L9wDgRj2MhsYzOPlEve+u7/
33Jg4K1BCQzASn5Qv/ALm9ktdX9Otlwq8Khlnxw8gceEwvbX4+cXobUXZmNoSOJOMMffYTNL0WvV
LcVB2pfVi8QTRspmBNy8Jgh/Hn7HKQhWZPFWoqXNKVcI2qH3/90PLUFfgc8xCT1jBBF3dOOjg8Wi
kbm+3ylKz/Hzaf3JMfl3Pl+IJNG6NsxqWyS0eQpsQ8lokGv/gudED5+cT+FY2QGCUKrEJo8r2XYJ
3USbMfniaRQDdDjXKnGP3SOa8V/PTMOxJTvJhRNAddXIzcQSeRMHuXU/4m9YmQd36yBjEyPOOAzc
lw8LUqo3Y77VqxOGznqIXjtKJHrbgog5ItrIeUG1dWU1GRH4QUBE0aoFQ5ryyYhX/Z8jtCmPs5Ay
Xhw4tHJU8Hpwc/+rTn3TyC398Dm7cxpRA1OuaZJVVuxDa92yZ+XLU4ABIywpMWro+YMB0V9OWxv3
0kC8fdTVw0YjVZg5CoYZbxZKj6ZGZ1r0CPTdTYSHCuhDG5vs/lPE5PN8n19+EdpEgvmqSCF34zhA
aLI4v79Py6h8R5feLvfsQDaa8/uZD93Y00aOEW5StUis54xj7cNOCN8fPQ89W8hxgNo0jwpcdBFc
SOMmfwW6K9+GsS8jREKGBL2Mjh/PkhIEN4bZfTYJmSD4IQQM3ccASJZ60+0KBoTZ8FKQlj9V6kSb
Z7ddql6CklmLQrCZeCcEUnMMCqyO2W2q8SEV7AjGkgWvbPxBoQjBJ9ubGCNDYikBJwGqLHQbr0NG
ePdAk+mLzVVyQmq9POr323D0CRCRKTQZWfhrQCiJZEay19UWoNNuojT05z3Tf7xwVYdYq6VpjxjA
4IvC8j5z5cnoThViQG58oLfvno2Pm4Ui9gFZ9A7txnllquyozJmjZJQ8hphY2qBsScZhIorxrTrX
O2JxcY1yLoWVTQY9OOeTy9lqtB3+w6fTxxucyCjlnl72fjyAIBRr0bCN6gtpEVHfIQbAqbAijx0Q
nLFO4Iczbtl7WrAsYbsz1TuaEKaYV/TNR3PWC2K8iltfQnwkAFim7FaWHrzdAfrxc3zl1zLPidPa
LjrT3udCASG8vZmgUgWIjb7cQ5C0kAdWBaRTLglZ5vcULA73GQ2waCqHjWG78NLvfdw0TIPs/Z86
PJ8f/YHWVAHxhJUORtfwNoTm4yWT/tW3cYQLpUIRLKnQWBmJIYEDInv/yK09jej+Oq6b94Dwy5g3
3H5tqlvkQ9ZXEZq/wNAccNvyF2xviSmJCbithqLoQeWeEGPbyHPE+oa4gIOjHkIHy5NlguNO1b2o
lXxeeubUIo/Y1oRWJTcbz85zAQcBur1GDdbdgm2AShdzPR3sNjbPnb4KP+GiXoyoWWj5HE7oWMaS
Mo1ic36xC2Z/OD0gt8GxYwvju2m9qAfolUiV3odjkyPstzQpqgHRlIjhGTThvDItA0bnSiHn6b2E
Zm9RyHoGfk1p3XduxW9qPv8QA4zWTwKU9nEzFBQuGYXQDwDDt6D334AzmD4Q31zAeStpTjtmte6H
8clUOfC0uPHnGU2hhGZZXsIjoTVYGM8PeWqMbeu00NntMusWizTTYRbv+CVEbclRdlZqA3KJQQTk
wqcJiYGbjOA6pMXsCif7Fn6SYi0nzxI7qW/PrZljnvXRCNouiAdsG6gePBdzYmFCQN1AwNSrrPBN
LcxmLyvpko0E4CIf+sGxEzZ4D8ASHUsIrVXLu29Ew+oO12vEVPcr3CeKLbMexsCiFcO3XIpIZtz4
sYnJvMimpBPsUGaKzJXpN1uu10tVohsfaSCHZdsnKPLLQxUkXusJaEdrFGqWwXlVw0ar+lQkzK1Y
5Gc6FVW0ciFPM2+S26934ZQUFl9oXnnZamu62u7gX95iqNQkUXO21ju5dse63aJfaUmDIOC38WG/
QAkrTn+DpLR34Rxob/Ze0VDj1SJsz6ZaQeo7ZJXwfXa+vESl63LYt1AUx/ijnldVXcFd6/2PtKsH
cTIURxB7IDthov+gPrKi1jTNSaHexNOXVblg1UjTTMx0qOc79B4RkF2RAqBTYglUDaj4ZjZoZIdZ
cYPMtysz52pMlMuAjpJ2zzVdTXamqE8zAf5CAKTLLHHsqr0cFcEjYg/1XARpfa0mFIZCAfRQBZAm
fe8T+Km1Z9aUQjlH73g4Ba/RD8KNsjtLDTgsME6LsX8sw/GQA8gQmbg+0Ke2ebSycu1bSMp1QmNh
f7ms1zwdSAnPj+JXNRSPAu0zpx1iLQxyfZLZxJ8eiGXU0/jDz00j/iZUsNytk4tqGEVRKkOkrH4B
Xcl0S+t72wtHIsPu0dupvawhSeeP0PV52F4Ms5EULJhwpsfO54Na28yej9JpCNqoVs40anIbqTf4
nDi0TORQeqRBw3Mu8WhUO0ecNetIpH6+Ee1BuA9DRmlyAgZImvU7aREt+uDZsRgCcY5hIoicht0r
2y2QfP9fzgYXeIP3wkjuZHXdcg101pppYxBPp0opf/QeR8CFDoNRBUiXQ4qQGg0CH66Ix6GaCPwN
QZa/y4RP2XLGrjdBKl4sjkOJsNFEmC5tAWdIF7uGLNMyn40e0waSG7/g/5tPho4eBe/pxgZD5Xdp
kFg37aMvf3gIHmBBFBUIn7+vy4LYmDbSpAPE5jAGI4FDfe1DLpFtUERC9qrmqirB24TLck70m/bV
s/vAhPt6Vogc1Fm0jyrfwycMBOppfPPdYvZ5Pm7T8LPVcnKD2BEqW0Ub0VlvYixMSm5OtjkjLv1N
44c2MWDiW8wb5wb0XeSv3l5ZYY938tQc8KAFusMKr8st8oOY55q1NEXlDPQKOKZEy6E1u0HqfwHw
jsvoEbY1xyPilz5JaUqaR9Zt72Te6GRc1ZKD8UgGJ0cGYZZGCUAIqT3VarvB9O/Yos5dhbNbQtjv
/uXLObfIOmFangdWLjdduTUE+f1phe11qA9rBOdl8311RH+3s5JBnhpNVyGj5G/dWu0cdX9X13i/
FEexrunGtSQkcqlaGJ+O94FIzRJsO/X/kSXEINvqj9RRRxG107zjxH/C84ewn2SLRF0ZzA4uJ7CM
pp2/R4YDTfsFnL+5cK9CwtxfhHiaxZzb6smJIVWe7Yq9Tb1T7VemAJSiIaazONk+zjf8ACVAO1E3
qZblyOf4UXZBHMp/K+SS1B6qKqFfbOji9Tcp2rvurmmgY6s1xB8wtZ0GijUyth38rqqdlhIVlKB/
R3O4JfEhJ80jy/ONNzWzbGBJYbxjYHze22TDE5avvUy2Eg/vmX2Jkj8T3VGZ7s6/uZez9bo7Q5NL
yp/Z+bRBgr1lnld+cF6hCWmroXTAFKLRcCxclpJC0qfAyfWt8wY0YtARUW6uscQufnfAzzC9eOv1
Fen2sMInC+bWN2UrX4D/tfkUrJ0SuH7w73rBFWU5jvZ1dWPfoBPqa1yUByN8v9LT9aZ6uTaV4ISQ
FXpzlSQO1lZE04lu/sQl3hMXUmdppKE2wwCoSn/lYtXsAuSM+S0RhhPN9GeqTODUiCHLlatgF0ET
3sFoMC3eeiHYwkHo3o2mnMcaoWTfIF6b7e9NcKF84Dsr6qbzirUGqUOpZ4yy9Dul5G5iL+C/ATqC
lW1hDFhY23824EbCGgmedYo5f6pQ3eaBXcJZ3hhmo8DoqWpn7tDSwQf2tyzcU3293hgl9BopUFEO
cRRZIQt9payvS/YaFRSAPbYz6fDGvdwU/vDLEW+/n0TzC9ne3m+woCbe9SoxpLVgYsF1B8tFuIn8
lhFTqvFBEam1d4EhL983QI4UOpomm82FTxmF9GaQH9D2OVsAJR8lDBB0mIBKo8ThSTNATsuK40Bv
/M08g9yhn8h16izTWqkcbl5RrLUL9QjGLSB/YdrGdEyhH7YnmObX8gLu326g8WD/3Wb0i6cz23DV
ERS8pWMJBzNO3joMNFCsLzzVs1dDvjDo2TWFcji5gTU0wNIPpGZsU+9DSKe05Rb6vJuiV4AmXUzB
k7GqZAkY335Me6xnkqZYce0ku1TB5iJIiXWGZSNEjiJP3CEr+eO37mMTqNF+Q9t34TzQEcS3bS6B
zZpblIC0eDMU073+7WnmT8cFxI3scJUvPUR+rKnDDTeFlTkBD0jxXa6R45zM0my41Z3vj4lyhts3
oi8cEu1JQGo40GcqQQCnMXaR+yXKS7v3purUacEmv+6nWHTel5de70ZPEdHM+G76VSdyOFaCFTsc
mFlks1jAKmGFJC51NDMGbDDMBkVAJVAcriRtQNDueWKyfqR4LpTQnsiVjUUGPAFUOqdhot3P6h07
g9xgd4L1/12OuK7Ayjd97l3e9cpsj1AWVUnugiM7cWPASj9fIF+n5ErTXxZoxJ63IPHRKg7t3ksW
+KbdaHtZ900RK9HTK+kAVcNQ9aoiPOEMq3/Q/adLMzDXuEh89G/0SKL8I0hOz1co5HkMViZNiObx
rzTvIVV0ngviQ+nVehXic4IzFqLglpCKx5/yY1IhEA/xqpvi4t3D0bFdCvrcQmeOG8ae6vzMebF1
l7RezG430ETIxTPoSbc8DkdIY6x6XPWrlG6F0zwuuJMWnBWl5gPm5bsdsqEsBd5nMYfPTOA4V0Wt
NZjiyXUw6LE+WThioLbEy2u7WSSdKvGeCJGom382WzWGx/GLkuJygxTYd9VrBnbUKcj5rxuxU3Zb
/LexlPmZDFBlxQFW88KPsI4rKEIHrtr1fTdBoewpxZwld5U/exZmxDuH74cJC+HbzXZPZq1OSMPz
brEAz4tkp6vRb8KHr6aKmR7S+iPtaU78PGEz8MnZDV7iAqBxstcf7DH75Ec9+F6a0Pf22t7novl6
5LW9xxX8VxPS4zrrs0q7S6RPMAXyaQlL9cVYxD1yTLsfMwdS12G2AnxB8z8Q8TwFPOK89+4AcSTl
iJbScWghabzprB72PbOq6NkZOhCbJ9iQ+e/vVES9GwbJTsyRC4sd302QvmU3BWiFhkrLkOKndV8M
bZK3tIxv36c77IZazzREyNlMsN+bw4LIfnDpXLAoTBI3JDfAEy+yenNyreVrRky/R3N8ChPMytWE
6SJM7ELlhDIbav7RnMwuD7G+oc2YVVyvgZ3Gq5gQbb5O74uxQg/DExnsc8ifG9zWuUC/iLqDlOQe
oKLSfv86kswdbd1xltAXUuTOeenleXWnDkZGwqxv23jya9q68hO6ZzQkeAhVW/RMKLcGvQQVCjot
ntocp6fJrBEoI2XL2xeQbFNDbg6rxlDtRG0wOGm/H9Rm2nT2eNkUEDzq6MN6aBGFSTnF+OF4AZ9P
T3SybGmM5vqqWryS7SfBYAVGA6MuXRgpyEYyP2EeZZfXMwarBBxnWdJ68sT5dyg8k6lhCH58/z0W
E5o4BjmhshprYihv2kQD8MOuHQg0A6HokZwj/9KqypzGBDlfv20Stu8dLR7S27oCjKxABDVmAVF5
IOimn7qCfvJfMWU5vd6byrQa5GF4q5zr0do8X10aKl0wVmO75qY89f63ekZP/8kYkkanGK5sDrLq
jMI6s6VaCy3DHxKERdhMALX7cDlw8xsTH2mTwpWuODf5DAa783dSwgR2kYzJdLR9tVqH5T1I4ACb
uRMEx8Ud0RJxslBAQ7Nn1kNJmF5pteefu3N7asPXUrnu3hZrpfA20lnrZ32hD2zqv651dAvNRulE
BJI4HM01VgIueCFLSc411RVfiYa6yAs3fN0uZIAk04Oas0N+mcSzFokvWEIcwerOfxX28YsNl47g
U57X4W62wpZ0Di028h73hBlOjdM1E3mthDkySErjJ5rPSpoo1C2Zbpixkj67UYQnEaPBtNVUnCO2
ZqZ12UpeFMvtYGbmPpWQ15xYmnR5c8qFD3nUKILXQGdCGrYH/virwA0qiBF06iszqy98IFv+VMN+
ij9e/fQ8l9twlDDAJp0OdoHKvc2h+GmaQow6C0M2zXVnYD4kxxozXZfFfJD00lawj25JvEgNsBer
pPxtB9vpu+AOkeDKaXvDujkjAr516fwgnnOYAaLUQNm6Q4JayFV6Zahz8bw+31QMtl0QM76B6/dQ
7k38KzNonpEwDfEMe58kbVQDeS0gFwkvqlqIr56ddLOA5wNhJAemWPcttG75ZhQsw/gh+rD6xYMB
T/hehFnoGnU4+ySQLRWiP8+fyrs48ZBueQEAyh26hS8IcZYZdWrV7uNSD1Y4j7yfOtG02FBJY0IN
xJa0Z0TULcWeQul7NEmTDtXOlQ5uzJnhiZAayQlVATRfZTr9KcvXf1o9XyikKpk4W4l5T3fw8uC5
ouQFn4sBuJmHRO7nz4tS9YA8vIWGUnUoa4I/ka/stFYxjkBzdMyeQwOFj2v1vniys7pg4yrEtS64
gAbFCW0EXVoyxT0qhta0uchR0q/bOJLlNvP0EXGq8b8zYDGOtnOzaYYcBljNX+mmsu90S/xzz2fX
xNh6Lm7QrMUO5ugQdP2CcRY0LmO49zQnuh2ABKsMEt5meeBJCComgmBPNMd43U8ikO4lF2EVlX7Z
7gMeHvtTJIszi7iBHY1tSwep/SNxJh/p40w2B7cdPRxEzJ5240vTaZuBm4Qd5ISoJi+skpXRsOch
sdIcfc1eZn0yUUKn+8QZMS2XyBCeSVFvkQnoSdiNWxDPzKu/gYwggDtG6/y3LPDkWeHyAX1qBrgI
71tFSzC3/WvM3OaHX01dwvK5QVYsNotKW6TfGfhPd/zh2O5nm9JA9f8/VhXQWdbpG2SMK0cMC1Ei
aKXxIpcLm1m00cfNtDHZ7SzAXv8rI6QY8rbxOQ9DwHQiyW+3GLc3jjs/Thqx26WhE+nzhwbLfLmo
caXUODsMOqvulswrdSwnZVnUFiokiutMFJuLowx8RR3QLynKrS9aTOPZWk37POMvOAG1UKXbNnr7
ux2VErLGRlKCof/Yks1wB8ye0uIEuNW9I+kH+c5/2t4cmNIblDMYdLnmYiSUZpV18J14bTCy8uVN
fPZ+7H+XdHZFMgLiKg59wfsl+nL6j5RzIus3GIBaEiKGnCPXJPB/8OhqPO1sSAHjQkWrOHBke92y
H4M3dHe9Ign3KytWuIboIpGCHhM4IRzbKK46LpsDf413MnYRaonrEp9qmA6MfML5GSKgnkvWgOaz
o7pp6zlesN1nSGRQqvA9yMSsTMUjKxcL5uULH1XCsS6rgSM1811BL+NjWDsTLXfgAEbdHUSV54cN
qx2puqe+B8/XOPwJ5XGD3vIJALNuwgL9aKx+N0PajNgGAXKyTIuKgBYvuwEAkTBbYHeGWjpMlQiU
EMcsYaDvxIU7ujypxSJJx4W5sOwJqwgO3M+1V5SrzoGbijQX84k/m5YaEyPR/AmeUUT6+Kv5i/q0
pG59k6Y/LBu0F5O38EHSNPSj6UYLteY5r6F6J0gVNAZvwEisSa6JBFAmMXtxNn57TAyjVV5EgKpT
PFSVRDYep9DcW0gjXvlEjGfPEY3msmNFDZmW/IzhMc+PLb2kLF/2m5CRHUUrpbPKHBUbt36ccikM
h5KdL3bLFizh6wlc50SQsYC6sqn9ONiGWvmwVTNBtzTZkvD5BsciMWJmm+GLE6MQSM4f/xnZk4Of
L7MUbKlVg3+XQqu12whl7+J4MSjaSih42AoXAyVsYd9eE0DeIcAxcnvgzkP0rfuiG7vnLqiWWnIz
VWcp0mi0NngSi0wIfpmkBdXaFRTERPE67zuSUqNxjgbYUoemy7cvQ3C0TFy6YT/EpY8F4hShlAcE
rIJl9DYdWB8IT3lkTQ/fJARCbk78uMi6Xf7EmtIU5TZBypI5/HFRFRu4pgHNj5RB/yk5v0mzfS2x
584jBbldwglsV28j5vvK7g2fG9ZF3oyIlNHS7xJuFWmrKF5fpqcSDk+BDOkHNL+fNUY929g4Jbuv
VahGJkjiOEJeqwqgcYN0pbKKPQ5yBXZ3qEMbkFAbcrkeABvRqAkMiA5N4gFhJpMoiSN6kImcz+m3
MZJ+W4wowCQPUkDo1C6IoUkQmiTchcKwcpuLMlXKoV1UbEn0bQa1Jo7RtemgUgSxrkTFHOY/HTKw
DfZAH9wcO3jBODHEm8CqjvqFAD19vG03647EkpcR9dWXbaWcvDRcF7p0EpybqCmtlfqRKdp0+zta
8dSZM8PTwt22LojenjH+Qg5f+hmNDMWee+DncE1S08ESBXVKd7zd2zwz8cdtCqYRd/Km/U11kPuk
/B20K2t5GhsbRzSogGhAOyaXcAK/DgMfrBmq6BIAReX3lxqus2xq+nNBcoC6hPpxJl/s0lOvnJcx
jS//EJel30hAVKpJNnv8vN2s5B55WFo4wMtqk1S3/CvypdT4VYZa3GZr8aIswRFtPsZugeuad6Lj
kJlNI9ADydhso5Ax2nk94B/oA8iTINCzRSiyVkofxShix+Lu9qlTeK73V/9DpJMFstbcNrWxWF+D
FU+O7em1+Fq6rQNRYjL3Vy9oQR4CUZ33QPnGyxM7I+m4kqu+NO9LCkVPJTIH8h1LQj4UM77sDSZR
xMvtO4ixELm4RE/JmbivcaDHFnKApYJzsyycNzj4qYzt4F2u2RIGRwuCi/8jIoHdfsWlGlRUSzN2
zDMI7zz2cXH9KvQPmwfmslfvjpWZ5NSyAiIlvD/Wsz/cMkQsZczSOsq5ttaLO0ImGpVaMXx3/bif
pXtyRR51sBMiR+k+ipLDEoHoklFO7XD1xePN2yoZaz7Lq7E4YrbfbWDZ1H3jg7U2gzbjEsX4pXkb
QXDqmqDJG0KqRQURPaxdlgVBfPKq0lzAM7wUSpPySCaRKs2xbDsTyGGlwosmaxEmJIKt4ylPrgkZ
BPYSoZr3SgdlIJlvxJrXNJAjIFHLNHDhNqK6m7bvxCEkYkoEG/0oZFg5w/mMHwVtiMk/zT41+rm0
Uz81j9WFFEBn1+Lp/2NyNu/ZLOcIWwdC4J2QB8JRhkFrJRj6njkZIVrtxmiI1RQCmf4yR42294I2
SBTMgvywvEGuUQQt3uDGlJaj0K0cFMDVMJJRUXskRynYAcwwgCB1PU4yX3d84gFN7Km5JHiDnfU7
k5HsO1qDMlfPkIIko/xnb6OvQ8n6uB+W338sbivxgORueugJDCXsyGCoBRj6agIWwlItNYzW5ljK
UZ6Kwmca0IAGe4kvyisouHWu4NNqvXYPMZai/AGnbusMGTUmQc4TBi1HkxotelLvfyvkFU/0uHqC
dO7fFSNvfNj7cjIPdc0LogNoL9TFTxTAaLYrbBhyzxBSYkP+hQcEZveMlRlSHfXcdOSualznjIka
UHdfKMal2T2XD9p+FRKtr3u5f1sM5pSaSaUEtr3kXfXNZFe2mGTmAllnUP30B5RbcVq8SD1iNyUY
0Kjr5yaOG6gEWvsg/Xoy4sAIzj7gtfxrdH2scRAaraQQTrhuXV65zi22MlvlGIkFb8QhFs2jEvC7
BRaevlPoCtUnDjdxslDf5DpSaCL0zLu+rqyQ45PtglxNPJ2VE8w38xit8XkBTYLvOBvDlXltUeGm
lII+O04wmcuV4+MCuxFZ5WhNyTOfgMadaoorCOaELu3e3aoB8/QFMC0/amEbItB9OxI7zoN8i5ek
tcKDgRNCJaJx/G4oY6KZQAtHvlNOmT9uvtbVcTkUF+4qADH9NeJ4cS2EqYYNVBJf30Mas2VZE32m
5c/1uLLUVszef1Y/fvcReln9W2U33UdU27CzX53TuJBKKZ8m9RFzraAhx8ivhblVJsxQNKbhAn7m
B97/ccceAEx2blXYnu6PSbBaXm1HBjOKMrh3rdOlbZVylFEZ/H1zrIhZPrTMtdsnYIFlPhFwytK9
ckGiJ7HGD64DHjXk3slpNFVsKIWQgUOO2I5k/rym5bBO2qfuEJ3GQtABYB32Werx97MxSaycTRDD
YmmQyQuG5PDSXP4UetEkIFi8RLyB1xShTJxEoZr1BFU5QDHMhnutad2iPkzTE4HLiG/FWwAawZQn
A+foZF335MIB99Sk7pIYne2KlfbWupY50GzaIflPl26xWtjyV3MhfDaZNJ7hWMSCXj/aAkrAmzoR
iIl96zvK2vWu5z81QxZS18L4bHiQT5VC2YQIlCn0uNlpXP6ksT66C1eW5ie9G0czQ1HhX8D8oThs
pdJo7O21O0zIkvMkvoqzUiLAoLYqVTUS7sQPLAhmkB+w0DxB6aWE2ISr1VJFxQyoMKm4+dnMxSS8
+8M+8JhJ7Ss3mQX+p3hWTo7XVP7/1SqtumQAlHyFv+t8zdl8ZbN6LJEgavyc7SSo+5W+EyNJfDuY
xWfHkJ7+iEyMHg9bYhhEf2ah0FlfsNjTXLCcibgzICCPdTgSPW8NsT2oT3E8jl2GQPyt8HluBlI8
eWI5XhLIfwzz7JZiiyMYYSYgqMUwnDkFQp11X2cNs1Odo9EsSxpyb8iFVOFSpqyKXNCjjAox+DE1
o1DBEPGp7wP+3EZQxUUaAd95Z2n7+qaD3VFyV99J1U8cENc3Ar8ayriBHlL2ER+ooZjR8XHA6b1t
l+GPtJ9/+9aQRuT2mZXtGTR1H0Fc3WjTPLKB5owhMckb+1B1bj1Q+Ib4Ro+oBW/HeIg6R9Bf7v3T
WiIII0VqI0XIWOgQ29sLhvfa1tWwRtw4Hu0/pvrkPq9qhryqjC6viIieTj7jyBk9p06Ocqoac08k
96jelK+93WzgWkJjyx+Rxqx4LMt9pzsFmaM0L2OJKJ4AFApyl5EVF/k2YCr7YhnVcBJMYcTIPn7a
cQYpNIrNorylLUs2L46QSHDpT30d9k6uy2BRrjXNdxj7fZgD9rvAl1E1OnEOUZuBlkozn+ymIGC/
RtMiRz3dg2PrhOFFBh75wBFfQyE/FAFT5ro6xJsM2fQhYYBl27+LdZZ4Ou/vKI79EwDMIPR6JbPS
Ujs8JWZ5iac7iuvLICpQy6n85lt3HaBBOr1HHGDcHra+WLSebKZSRT7KttUBqUGA6caKiDU/llys
mQopv2pmIjZy10gSaSRCSLdiD0CXQW814YPPYvLvUoNoNLkEO9XduzIM+es/GGTNgCLnCDKt5kIQ
RTkZpPHEZ4rKNQmT8NUqM7j65ASqSwto8SkDAgRJf7XZCR5q1nRBh4EE3KwkdQkF+GfDvwav2OwH
SMtJtdWLtTz8KC3/DfeWgR2ZQltZFV+O53YWLSyv7UYiIXJhKhWXAgS/zH2Md9fuq3+DBdOzKkcQ
DUlNYXhNs08hK6yo5+ASlS/d7UMmSe+OTHkH64mOU26nk1RDp0vAAfhLKhgHn8O/hrAP6G2S8W+b
x9TTjyM6f1q8XD87ivvsS68+tN4l2HB6JYm1UxTxf9uT3ZRSsdu1qQtnHqfccss9N+Xl8ilOZYH6
TRnVUK+cjksWrPfSQcK7xe5Z9v/vIZRy8CQzG9KGAB6UHTvAtKSRM7BUqOQGqBb6hBl5GGLrITcz
ndKcklYLsm1as8ABLdOfqhva176ZNPXV25Q6oVJ4fi9aeqTaRoIJWJyytDyYRSYhutNyXUdluVap
/QKOBqpaw9O9NNTjjeZ2+AvCNiRQl0CVePdkhUkEi6vB7/mlveseT170K6HL1O9Qs19NwmQ9/AGU
P7MF2QYcI2fRPe2DmvW5R6w6rF3eEVQolqvzlsxi1iWFUV96qbQvkqVyeodFexNCEpao6+H/R2tk
P+DyTHGO4jGAKlgYmBi3eNtPbnHHljiCwBanZOKjkGiz9UO7sj4aL+6WoP4Bn+6+3cl/tTyF5+c0
SKZSi8VgjcQGavbwilu/MhfqOk9ALWQ4MBMipgwrZQ/1fTnueB+XTWZGlNbV7ctQ1alUZYUFkS2d
CkXhduB6Gy8wW6/aO93sNxW6AG2TZomHh2ZqmHlJQFFrjriI6YOrcInXJV8GCM871ZYoy4A7vg4J
lvtbP/V79EQy1g6LhKyqjEpV8Si74/yM3wwbumwmsaAtf98KrShQG2L6BIbKSEBUANZuJIjEnZIu
gnCYuegVY+pyjdGrK44ps8hi31rNs3aCqMGTRFiFnjaOU7JeJ095kFTluSgYorwzFdzDQtLusPXO
RcoJX80zJczwNclr54MP0/ykVKmN8zfRe6d1MxRlY7oh6RgTvcF2gObiipSZyW11+EcY0r6buHaR
lcWyAvlVL+2oqrMhS3ogfsjkJ4XL5uluwx5dFyzdpBCmDcpSBJdqb2lDqNKO5/gMtGEOB2o+bQhR
0NGZhrmUW8usGGaRWnHJZU3WSar7B7CeuHYL0WGl7oR6DBgvswOKYIeLaH9ltxYnVQ0Y4xVPLFaS
wFq38bhwyYKq6WFOTY6/JgcMG0iVR6ZNq1SSmwsrE8wZLqJO/5KYjjQ0GwiAFsILBKz976AS+ibb
TXGlvm4/VxV7dZ9X/SbeVrHFyJ58mQaewGz8TiB0hzwD0AtymozHxoRwhzq375I5GGPt8PE1Xuag
AP21ycVEyycr/kobjUAwkVk82b5QsS2a0lSBmlRduAaZTBWUMNH8HhEVYyGiF80+pvKPLR4+rDWT
8p5gJ+k29Y+jRLthGsqy5Ld3apdPvVor2sqxfldhNlVQRyw/7KdYb6QsmkcEDDokBnZwE1vhh9zY
WeSGLu9IA1lanrydfH7fT9RLIw3uVN04i6r53Kdh5Mlo/AYp+Ikm4FDC+dj04y3C36X2J8fVxYXK
pMLu1KGtayb+jyZDD+Ilbl/I/Uy3sHOhPBfXiMFmBupotZilFSf+Jh6kOEbYp8iH7RmKI97Xeb55
+RVXrD5xj3Z0GEwtDNRkbKhWq36v5ghLzCxiudlRAMNMOGZYaL+H0QVzO+DC4MaW9ooQX48lhdNw
3b1/szeF8k7dUtzLVlecPn1FWD7U5RVeY7ODpion1QZb0tqDvOXi5Loppk+f9ZFZXX0hoMDiDoAP
K4KSO3JY+lUOTJVyHRFiuHUfN+Iv30qzPDsNUquc658enZzUVtr/wJZ3YfdvHKsdnV5FusoLeUNf
ghRHJ/6fSnO6/J4L0WH4+ZEN0mheNKo+N/Dtj+Xo+yklDb2/bKdAuNFbmsdY39Da3hwmqacMdC0U
2CC9+r1DXn5w7ThHDxKoHePVH3xf9OpM0ID+tLhbwIwFdPOXvMIgJDXikcC4aOv6Q6+WaKEtO8Ae
AltwxrbVIFirSCwj8bbDrUnJ0N/DP3Y3t0kNZ0wSV5AtWafjwIvavcxHLPpXfCv2Z9RdtYkmTUFk
v77IlVJfmpt8Ylx0STPDMGkCFlxVccnx5xSXPrIR5kQr9mltkZl91/W6BFOTyd3zT7hC7aAFOeiz
ACVeIymhLNa3sVfmykc/ExoHHaeavf/jN9pkAHOF8I51IvYS6flJGdBdEbMUOpJu5qBjoDgWPTUE
q36nEnpwRWGm12Jwlk8dwTrdiUD861ZnDKwybL6BKh91Wo/YeG8X3Qffb4kmqeNqal1YWstY2fDA
lhA5FQyWY7sY3wDtot9xIeN8OzocYwH8MdcCB9OsMVtlGYONLBILarVHHXA/tpIIncyBlk//6hrO
/o6BCa9f6Kkuazrt61cSR/my/R706y1c66WTlpZmmq2oFvloJf3cTmSC/Fx6CLFb1c6x/eJFkYVp
2SsnbW0/VDd9Z3QXoEts05PiPM/v8uuEYj74jxLsw5vy8yM3iNhSqjITr6WehHFC4JEm1tLoUoeS
hDnOHGSmaXbked4BbZsE40qtRKfKn2NtXW2d758EoWCx9B7oyFEZoF1QIzmvEQFc9XP6jzUqfEPj
IuNhVESmivubvsSMKClAJDw/CzCZiN3CVHgOZBIjgfrK5/5u8BnUL3/lp6p2QG+HxtavLiWxwdjz
N8SHtEGAe2QkceMXqC8IoceLLq1XOgyyGWAcLPQZrd81+Pfb0QPqWgIgVnpyl8dkcPVD7OUKp1KN
b6i42fNn0xn/8im1SvXLN4uxm+YS0f0s4P9AtTAPbbVRdVh0JQgrmTbn4soSwAOKgXPxvSs3VZu0
AyV9dPkKbgH3IvW58YZAM1RuN5ZIOKZDWHu3JG7TQmyA5vWLQ7xKZ2YeKlkW2ZRDLmIDBdrZ9ps2
PC/ARCDsu9GjxwvpCCGe8yTJu3yasgVMzrR+aSaHudCshbKa6nyPskBU2g+2rBqhDmuhjF9nyPIv
2C2N34qyJEmc2B37wrDyOxZzPrF5jc8+QePH+mBcn4X4hjWQ4ej0ePyBpirSNsAlxfB2OWwctrtN
7Kk9vo3jROVsbiLqtBKXycIhpSaN7p9dskdTjfw6dovkAxYWWS8Ftggt5TTKesy7L+JdudIufiAc
hENc1mXuKVR4f3OcsnPvO1A81QNOoN81/Oxkkiax6c4r7hudrH5SMSGzeWldAxUKb83C3h0LJORJ
eI1iK1XEYDr7/4B3d0yjN3Pu9Rt7aHEZ4mBS3/++ZnR6B1LkYJEtGRzask4MgZLP73UNVQGO3Xpo
KZFY4Z/WM0q1YUwh0oIp1Tc1LONB9cW84jcaPrbLlkoiEuiF9hglNwyCw0CA9JTAroP/r/vagvSk
dE8/5kRnCU/YgYQ6UsDQq/y+4Xqt6LdInlEP7c9Yfqbs4eFTtn7xq7AtLfbEofwZuCG2GYQOpKGT
fNU6oltpobZSsmYvJRqWsQZn4R9Gx1hTmuBblDg24JxMFWnQ3d9TybjyF9l/bIFOi6MUQZZr/TGU
WTfZBsJAcpCgDSS3qPiZXZPj9UVPWiA7M8VkZiFwLQ1QiDu0v/jncC4mrm1jEVYIYl4IrpoBxBw3
MxtUKZKW6+vK+ismBlNSDOZmONZbtHzBGQDaQkPZpDQ2XMCsaZI9cXtps0IuvrooeUr/jci6b7OM
CoNYU1bPaedGCCCulmts1KhFXFt55poU4BtL2pbzRtLMxD1PKoYUvj1fkOi4nsrg8luZqk3HfDU5
fYk6ktzQQJGpIAKIg8darcmfNE/HaMoQGTlk4WvCZAYXXlCLXgCqwMtTF9Vc7NBrD0TLaeSeYCHc
gbMljm6yXkRfbTiFGG9vUuE9XfqiwYMLK2J/SjYKlZfuTwfNDTdXOZiAl2WjvFtzYEpGuCwv920Y
4fCu4Lc6+4P3c2Oq9fhqV5RY1HA48O3Ty9BmYolxA6Hs54/zyKP+3s3T8Ds0TBZ+CyKA4G4VvRTf
jH1NAUSg4VxFCUHal0J0HZbGlRenWoC8fmAExf3fuXrqKt/YPfhxUvikijZnYAYL2caPwb+KzutC
vPo0QJgBwD9JXyoNc7UHTQL5jQ9a9+ZVidgUPo25EWIAoxaV0Ca5mbfHKU0x7QUD42hNxsTwiWho
RLeL6FkNfOgK5ZjW6j33Y5ZJI+2WN1D1miJmgQ6CEYan6cMnBitD/NtfR1PYZhTiPNn1UgWDJTzz
ptYQgqu8Dv9pa/ymlyVNdmSWD4jD5m2Qh5SZyc+EeeT5xxuveN+HIvVYJ6vKAEGOokftVGlaE4yc
JdnrVSQRyYHzYKIx3MiBh1Pd/I4BDsLsDOSjE0LHUbhRtPxG6QTM04eLn0NNVb+mf9oxH1+RDFx5
XCBaEOJ7bwCRegTtT9EWj97w+IRw3JHYlA3UBCJu72+IPNcnKs6QGEK0GhRGJZ6x/tAFqhY5RpiX
YOeMBZhcpSf+AvR6itOoWSAF2Ed8l1ufhEVBgIfOKSyyBBVYdavsKXOy8pfunEC7AtQTiiRMHC1+
AkYXTka1q64cgTV4X5J7ZDW6PUzKfuSqEghqaDjLSEtJn+5YjXT6Yry7udNJwEuIg7Ce/VH89tzl
rIRyxcFrzMvKQPmSM1hxNlxHeMBQ30ulCNWq0Ms9z8NWelkW3LW26qHrPyhE5QA35lA7CIo8tAAt
JTk6QmF9/Jd63im5GLSbJgtlw4k5KkIwt1Zt5glSz25pDrX0GZ+mODWj4eX25dguBWWLL9lqTct0
qIXhHnLxMxINlVTD1m2vZGLY9FDXYhm+NyTe9MkSCS9mVUwQeL9QP67m8dUaqLloCClw+bR5NwGm
r9ofppoW0gFTF9k/Iuom8rvTgO1ceoe3ZAB0t0uoEO6hPjurIxT3e5GSoerXOtzujPS/31VlGp5q
aUTqGlMFB0ICZSgLy+Qutg572B2+dnKmoSq0JbdO5bQIZDRQmQrJVxujG6Tz8WIZgRhr7+eBIIou
CUwX3dhkp1Q16RQx2y95/q8B1sON+mR97oFhAh5arS2emz0S7wrwdvGcjfgxqjTqjsWENS2EKdMZ
w6zoI0q9VAtXVGixswbOb1MAZreruki0yrdUjt/tbEKh/KGCKCFFk+ONXy2rXZ08ckXpXdN84XLJ
qPqh2esUCevNvZTR2Cb9DMkqyinmX47KwDCGHvJyDK8L3ENU2thnPoINNHZ0FD15xUva2YqAIax3
lBxj9U7+46wYFmYvWgkvpmQFohLa9KRn2mHTlmoloHnQ9ylRl583DFmlOxFWjrb5Jrc1IFv5cIL/
IRqG3eY9Iw8MEBqmxeE4o2/JH6gqvpc3ciCu7bh9xGFo7oawsfmjRawmLNF91KVYrarRmT+mIl59
T9W/0nqqEC3mPqFM528asGcAcixUI9C77DvlK/FJtE0bXA/Rb3LNg7SQEMJIa/R012nXqV4+FoIN
pSUu8Vbnnf8f1jTOgWasv12VnjS/HqEMPUATjwmknAxkWRV+OiRK+B6F8jAy1cO7OKF7sOvjhXKc
tLD6Tg/mFE0fevP2kBAmPoQ+MelIky04SzlUTbLWBVh4NgypjKmGV85QBiDMmG2yDvglCoGZ5k4t
YDfo3OOn5k9apbBT6TFBofq5lN0PR/spE3Em/trBomcNd3C9zYoyTq43UcXnEVDe8xUJam4opgfF
gfUsUv2WU7NOc2g0dCmEyGcn/RVG+e0MgPof1jDndsHXK1Rq8tDwmuDX4N5b0Fxyx/aIMWmLmfCZ
0/mHZ/W731e29jGRVip3N6heo32AptTwRriiY4Ld3BEEm1pY0gTJz1cgxrvDyY3Re493/XBDC0nM
2xY4aEHokbOeiqqZKURtANhSzr1LL/8UnX1mfwZ8eHxYsxbJLLaQR8OipELt4XLobnJkxh02srfD
e4fe0e0x/RVzpkyCPSddBLXUaLjK+JuDZdFRN6QaPO04VBFN1u7Pi9SoryZMfTqMeOHiTOpth7NH
MLnMKm7LpXN/WrraIgDkMW+AGiEx0/fCD/xxsn2c3eg9fiiXbDh/65bBiVVJNjcrD16MwREcbmrB
ASMPGQhBS8Sv9lcADF1UE1I19QuE5JYvlWS1ONAUWfjB5f/AF7TmPSXplW8psFSFSg4gqEAihTFr
gLN626mBBpOqpIyhFy7JJgIH647YsDy/tmVkdR3J/vcva/KVO2ZPxZYRW8gvLfOFbBNA+OPn+iJO
mCdF0E5t9QTZ8ISYXM59CbqineMLhF76hSjwra3QuBwC2R0G5zjVOLaWF2PSiknlRGAEI5Et92Q8
9wrvSugz0ybbQipo3Ikpm/sCvOn+1O3iI9OY+xwAQUo6D6/IjQonL6SZ2nVZQrHU3mmC/45VmlcF
9THLm3FDC+EpMV6m0hbY5lb2iDYOJITd5167JYcg0mK4rEWAMLB1NYLO/T+AdnrUSx2Xr5tiesB7
27NE3adnqYeTnrHDUd/bjm//wAdM4RQL73WZ0zdWYy9+j3XpdNl2DpRqxDTIHqLaCofEiJe0DO5n
guronI86BV7dIvBHdYnYv5P+1p8UCTBSqP8WvsDGVPWfOE7H8ljdYM4fGS2OJTdk77eg2k0Cjca5
ykSmH1Hmov0ByjgDkCEzMq72eeizSBBZXFS+A6nerOYNCgxgdChSddqdqppySnE62/zKIZZXqLZ2
1EOYPhCxR7FINfXpsufFM/L3qXSrpoe6HZAeoa5M+yZbStpMd+V86SXDjnCz1Sqmf2+4gFIknh8e
E2WSVJvVTCe5icpo/KIKvCXcpoIsI09mOcVJ2G1XRvIyAyDPgdigx2ew6J9FSbq/e2PIrLEIP1Nr
MAbYwltOFLBetR0VApdW0bRsPlfdLiIv49DIW4oispZiZrpJJ79jFGVrI/bFANzq6SAe8DlAi3n5
UdLTrpKoyL2g3udBGeHaoHOzMV0LYfrIEJufnXIk/wa5UJMWYDLFX1trv789xJ1zOysN26lVsgeg
H9Q1jRHu+jNvy670MTEI3qgpEjBA110NzYh7NzhKkym+jtqp8X39S7EM+kqU7ySAqeQJqUioDqnl
fBtI/09bcXKgkjELVDBEnmJWAom3BqvHsB4ByXVOPRt2a98tiwVjwlCHPG3gD2vMVOp+q5MqPsfn
syXYbFHeU61z55DrBr92qlGNDzSsXY82kmmXDeM2oh+fedQjySwJQnvCj6BL2IR8GV9m69Wlnpeo
86VlQ9qEtlGTX0w8TA2IeYO+EG17a6+AHTKnXTo3GjEpJsXJPqbe5uha8kZYc3zuNPRFuqmDZgOh
WSN7/XFuMZ29OeB3qjym1xxCSh7ZG2hgkjxep0GbVnPFAPjVVcGtWBXgydAbs/Qc9blJoMSQ2wSz
Pcv2WRPC5Vux3eE2Xytb5SoakCy3fxGvaUWfb38HC+7xv+kowLsMnFMviUlI5W13PgIc6N+83yt9
8rS79peU+bcRSBKfjxkHCH/txuh/I4Ax8sCr4mIt75A/evSogcDOUlcmO5fU2zahmtqpNGmH6X2p
+5tBnxREMSakLoR+tvBZTqnlah9eZ2ZqL0joTO7u+wemVf4A94iNcmy4jlieRJZPj4sbVhTAf20e
vHkBASq1++uqX7oHP2Cx6rpxQDV6lV1kvgPd/mLyTHIzXJzyiKDq6cYj3JPdoe5iy3l6anOIewSh
fpDYk121o6QnIZtyxz7vCwByAKP1JWTDzva9KAtcciS7sY7QkKjCpFhyD2GFTrCVkCthywo19snE
StTxBOsfDDPTKXzP6Zg1IvgL6Jd7cNp0GHIsRIQLY2f9Y8jjTw171S/G5RNlFxBuJrsDLxs8x89w
AiH/jmaANWxu0ErRFVCzKc+gbmQFQaK0RNmoBlJSp2hk77u6CVH1gZdK4rvSGksAd0T4KwL7H/lb
RhknvzJQ4fiyrTiSmVnxWf2/0yW4MJDgE0Y6UhAQnDDPGk39duREjtbt4lfcMWkpKnrgcYYqamNS
WrSS3nZ2lSEG3MuiisktNSzRVZp3nudmz+4X20yHYc2vuef0k4uh1OaHQ7jPjD+etkqTIf7u5JDw
Ep3noGCEjnZx3+mFZ598bDT3/UUjcIeuhUeNoGSiNyP9NoCFItBL+p+rg8MmDsvj7o/xpWNT4ClG
oK99Gn/UO2lnMYQJSIWbcGeQYlD+nUxX4cP6eWdSvrCTmLar7twVvYLy1VlrQJy6qn3K8rGVN9QS
wYjhnHmzPFSbyPEXTViqkIzWSSWuC2eQhfFQCp/qakvG6WywffyGojps6r1IzqCV2ABeVDuBjQ7l
vGaylV0yWnbwcGV7RdgNHhkS82KuVEEvHl0VthSEPpBPnavPtr6J2Tn4lNzpXZhT0mwLUeYLWlxE
D+Ga3KnmcXYSWyl+MrmHp3Oio/AaLvXo4uZJaTv3SNOIt0WaWFh6oPXrfLBF7CSwpzj+a78dtNLr
UlSAxGJ3cUWiYJ0HAkiSagpu+op/C+dlHnBZj8PCTYjj7AHqaEe+BmPlrWnOZPSfKkwRcJT/haSc
0ErC2/QAMNWJYypzEAB+HnQtCpZdCGXE7b2lc70/mZlR95Y4Zt9NgM+EWgaN/yUugct/mFjkh8pB
QpfiJKOm9j95B0joNcUD1Nbh5OdeyOTMSNJpnwuiB1HYoK6KhxitSdVk70/tJVCPZU/6+C6UHmlo
7eVSODxm7tpREdpU8M1KN/NO7bWUfxAIsPsyXIOocaP6zalHGIPzvS4gU3kKcKpBT8KFYB8Y0bSR
gku6x+PVWsxUmHbG8+9F6uKJcI7zOsDafASvptO7ao4oMgao+aKKB0tqkipwV3EXO4knk93WY/4b
FeuVwSluw7PBB/U1qBNtD/0qyNlb64W6ikQxJ2KHqHaAIi/6+OxHDVB9Pe8jcOTOztlxrxbunw5h
OQFm9S1O2QbDT7I995FKCdsJa7XBuevrKektrezQMs3F2ev7FUFgRN8o8IfZKXikldOih9dnMG8z
wPY/n3aucnvdcOcq7mB9t1Nqj0bwijqYMbUdappuso+/vBC/oVK681Gq014F6XitgASqYLWv3KrI
O2vLX7IH7psJv+0t//WeP62ugwpGA8ZNkWGVdhsfUdQ5i4D9TFPU19B3SbmrIimm5CqKfdA3W8Qa
RPa3maiOZTHSgZ0wVQl4xokxmfqW93lG7lX1McgsTO/NnvHiSXPUMaYbNrGpu3axS3h5fHEyPYw7
f3nMInGfyl/ISN6iqOevrJOmz3ZRqL4bMjXQIv0Cd7zvNujA4A0Yd7KMDkQSZ6MWJKjxcZ2GdGh/
LPQT7cL/ymURpjDYJexVvPY6wSN29mvzvKBVDUP2pf5JEabpz8ttpyi4eIDL8rkZvctCwk1u4xQ+
AanBXNlDxM+NLOC0CnuK4CVB16YBvG3lZ6ZEiKHGcaRS2T4f0kPLWd0TrvF3jk7E1yqilo2Jehzo
ixF1CEu2mQPMSO/cqtpX8vTjRdRKe/fyQFF6s5thnLGrtO76xlTQIfRQcsK+xp4Yxeq/Sdy26MDt
36SZGS825/oZjzwM1/2tH7p3pMHS9VYFVfp2dNcTRCOV98Add9bOxNEq2c5J/pC7NomemuQG0n1G
4Sk96+V2pdjdjtAUcJU3uv4mmPMepz5G7s4UcZ3/U7PGfq0ehQZXGuTPO75R+bKgc1OttYzoyrsb
2Wd/7HTiw/1xC4OKG0bCYyJUjCzHQmguycZIEniK5RhRzEKYckovpeX7FpEGtI4SPIhy9CO/8x1q
ql339xGxH/gqqUYUrX2vn3anWnUg4zJSdzU3fFKF7QDiqRVJWUv1xbKzr7SVIEtqfbreYkw/6CIr
V6emQ5b6kECzhOYS2bR1F8HDdE1WUcGfBvvzilciemQ5TMP7e+3HBDpINy3iCKy6Ysu6mRdReeF6
oyyMNUkd3rpyL+5imQ5+zHV4Ged3/ewDKfg6whXNL7e9SRBvXY0zi/54InS54o7gkExBDClH71YY
ytcDYS96A0YuUakcDqCdryUpbGCI/PnN3Dp2sgKWIMsfHL0Bz21R3C8NzCG0IkFeEQNtUuWHmaUG
8DkeLjIbU0NNbLaWt1rmYj1WZVG3tSxrT23qsb3EJEM01XUuo8N+1MxHyANXwFhOApJ66tn/cU9N
LZFFBoO+fow9cRPuamkEzhFAiHpzGrxirxUK9qirGoN/ap2uNw5rNgiz8bL/BBdhd3RYt4u3nFZN
nZXtSERkQaXjjjqukDNUZCqqg7FTVbWtySTjpPYQ35Bkvcw8cPOpXPdIY26eeprWS/MD4aBuxFtz
ngDv/3c/fvHb7+TO+eCnrrDKWKKQrebCZLR9m7A4ZeF2skG/UJcxGP0zrR9MagltGLYj8xt7urdg
LrSa4/ZIpK8tkTcCezyF8xDRHO2xrmjyzq6aBJnBveNbfqEtK5MLRp1d9Gxudot5ORb04jPgI9bC
IILkmAkBWwIE2ALC7U07A9AYORt6hjJzVgu9hYwYkMbNZ8QK1Phue/GJCwbJ+Q7QFqV6fVZflBST
/mxs5x08ZYh1yMrxldbaZTiiAQoVpfrefVOeY24sXrpQBGSQ5Kb002hO+SPnIaPEFmVdC7ujAj6A
EsuB+jg7DDGxBk28e5cXIL28lMo2RFcAGE8SkgeLbnNdv1Po97pnTbLtbz1lrg9XGC8excV7UQ29
6MYaicgowN+rEkdA5OK6pTPAlgIZf/2SJBsdaHG1TYYbPCMdWLmtS0KB3LBE1r10/8zqaDiotPc9
OZvzfey353KGREnHvzbBVmb1CfMS76Drq+COUhYL9PxVUJ6HQh5q9gDANhXND0ZozGabscpffIWP
7ftnmG2tSKT1aYrqxsXaZT2xMmTn7vCWvty8v8UFJb6NzNHqAj6fY1rzRKTX0PvggyZ8SFTpvbz/
yuKI4wvWoA3ULLyWrVTdK+oWB0i1i4QWYJP1SS8Omy3hfeZXEkBXDcvJUcsJV+1l6Z85kHywkMvV
W7yDvVL19Zr7Yid6zI+KpTyloUnwZPcXcvVaiEFC4Xh+cN7IfR8e7vSJOtjTnRG3YwAFDlhE8pV+
29c/b5v/wukitiz1oFoxG5nZc++Md0gQcn3VB21zJzaUkjOY94puiwABIvnaWWyGdZfvm+rzOCCr
kq4rNhvJLpnsi5Kb7Ah6BS+gF+EWnnlNOCCWZQZK8zAam7cQFR45jvs/qi8rulk7wqpyeSq+tdSc
XY0G/SACn6NC0jldfiMPKZvpG4bE7pdczn7/Lg/ucMsndnT9i08rB6FUa60hGlPX9Q1+Q0vJOQah
FxNbz4D9mGv6OXjP3CQIwfdR6yC8mFsFyX2lIRbrQuugP8CkFyDgMouK1j1FL2YzIeHO13gZAKOH
3EoAsrVP0rKLpSNU9rEBr7+uyxmCdqclnsQoANCDeJoI6yTYo7AI6dyyvHgsKwaEr2CC/UA/vlOr
iAMPg9lawXxojy2oTfd58DHoDO+lWUzr31iSHH+J5JMrJBPyV+58smoIrY3W+/+BgXGRaRi4Ojuw
ztVHIY3PTolPB8XCRH73TZYAhE+vYf96BZlkjigZOq63suJr/v/ty8P6Of+pWD3Bhl9PKa2Ag4pX
Ea+N3zvFnvz+Y/KKiWYVmgaoX2utXDhjjGIJXgN3RvsYJ+omKZaB7xyjkSyCW2jhVQTRmNSKO3r+
O+5ZL3YoXiTisUcXMqcIc2F+c61Si7Pl4m7AdWNEMAqabbrjGOk+8YRh/fejIMD7O7npU7K8hO2x
UMaokQjnTKtgg2WoCQNxphfBub10egLBUsvcLgaKSPA5hilmF1fmuPJiI4f0CUPbxrh79ZZ7wfeJ
8J+ExDNv+voR2fCjhD0ToQQRiILGpx1sipNI9Svrkef3tTstlQ1KFqZw57wtnc6pBgxXzhnhU+gw
K53gU0Rnkhz75vJrVR/9rS20778T7cMVqVsdt49jlIoZPYfuwieKLLvHnlsTLmbkxkq0hQCN8eMJ
KOXyc3MRBxtGL4i3gf8kAdQptMBf6LXQ4ASft0oki7aM8uiixNFNTqFTLQhxhLyUaiHIxwI5UaGq
YwiyIwn2ubPK/Raqp+8Nlg8C62jr8NiNlLPniB9xsL/PIHlRQpf9oMyo4zH+Gp/b8NJ3vLgaVu1E
0MmlOsK4FC6AJTTHUnNQLiIGmMAgx2iiq+Go/ph+ZeBJXDJRtsxKN5h3lc1MNGYF5VfFKg1g8dzq
aAdJYZg/md9AbxwODv1GyCvha7+wJWUenVPC/nYDxtuVim9rrkgoQyunuOkjez8niId7AJsW4nTn
XiEcjFYFL+9+3EoVA0GnkQwgNJ1kqXFBCnSgZPuCJ3+n6bMpPf4FjUT8SKpwxbQDbort5Q1lwB5f
/c5+hbBmV9plquHdQp7lr6YgDD/WqOunN1tywFbGubx3n0plNhPO9MwhdOy1D+Xmupoc+b2Z4qVj
x9S6GkXT2biBcEgXu6bCUOMeILg31+JjyLkyi5IaZ42w0nw8WGFWc5GsNrLa/E+jsJYAL5wuz08o
f+jXOZ8RdY0pSBAuFvj7izzKKDFRNsyOT+zmcGkmyBGhUjpFMLK2RAb3gTZd8NuNgvBhB6acvXhT
RAVMSH+2a/4bKT05acuJKzih952PXJYTMKGBKbY/o80HZXVdaOB7HHT7u2zIv26qkDnO/s/K7qy6
XuR33rPryf+fU5XjkyBi27EavoI9DOTPep8HNMEQgjMKx4sXFaDwgKC6uVI48vNRc6YbboVz+e8o
eO8IBt/g9Op+gkg5i1M8rAyAXi2YOr+nTEEK6WQAT+cSmNhPfcgFSBGz3cUvJaXXQRnBUUqEch0U
PPP5q8tEO1hy4uaMhgx5t2LyfJQ8PV+M+LIcezYXMgQ89cOdc/i5cyMMER7nyeOGN7C83jYlD9T7
hmpisa9XCCpeD0FM+LIw/pP3/LtcNBsfbYY4Phr16FOAnvvbOCe6wg+ojAL2BLcUHvOH1nqqSoPc
PGgaQ61QnOcHCQbAkVf61v217KhHL+zDMRJZC4jQq3PNitrAAMgmJjYBSDmr1E45MHRGuCmVsmv/
zrjdVf9c9UkrhWPyypcf2zy2ICyXgs+kK78+B9t58UbpWKuRjBD7Wzw4mx0GNtJ/wM7NesyAgLTP
guSvcCvdS3TXZkfX6G/rxKCwO44MY0SStSNdxCk5Ecei57amkzYXCkZJyu+usK7uxWAtS3OGWCJy
ib4kP5QgCiUDksur6MFXtSga6CwqpMF1EFNG+7zooKE8MreA81hLnI+DI6mj9zRQEJgKi/i3jT67
xfQxzrgBQ+WGG2k9gq8DYN765E4DZxu1kNwSuhUjzpX7SGay3J9WJcHygPnV6FwwEw29zCdKNzw3
EHIifKHHWqKjlPcLZAhNlsp9TJ/+DK69B9aEeTGgPgIjCvYKX8BNBAnEO+WlwhGKxU4v6c8605b5
LxAVaCom+4PbxU6DvSi7Er4g7I7EyJ2kHxZFEfgtMYGRCj/RoGkcsb9NEQqz2RNWQSEtA19pqmLV
NyGPezNVKsdABVm++WAynpQZkoPFGQt7zt/Ze/FXPmYY6yj4h2aUs9tGGzcMB2r9E6zKbCdgmbXY
vYeXwIhE0TXpDq4p6SGmgRYrKM+AHckcdREhumFtgDkZyAIttvsehnvRS3u6MBuKlZFOTjwnJO6A
56jB76FP8uHDWOaFKrGejRIS6gUd4dn93WucC81zpBKccwJSUCMKFyXmQ76tuUTGl+tqkCJ1USKH
l9gaDMBBiFBvfHNQ9a7nn7RWy5biGwN25DcGR8FfnpiKY1ovkysCW5CFDPs2JZtgfaSKoWuZ1tFj
mumIQXcz1yZjhrTljnyf05oTZ4vnzHpK6qSQ3svvOlfa57J2TN2zXDP3lsPP5TB5G442PMrbRyyJ
SJO4wR2Tknd/tD1xWx6h31bBVDsbDDBZB5peD9/KYjk7jwZLkGekXDKARzEq3XGvVR2XgWU/rDaa
FVZlEucpt9SByD3Uh9ojN734e0Ny0+UaOpCjZdKGgWzGejdaGk6HEbMGKoyHIFNNkYFYHaQ/0cNg
xjsxTuqg92n9He1wt+Ath1PiHPBACBeezxN4vkGZZY7HJ3ZtZ5kFxnDZ/MtWd4w4n2lEienYn3EN
HSVhCLdaM6CeeAqJ/709+7mR4G0oIDhV1JWjXRmYO1RlKz13S+WymaX0hyzmYjnbGa+rLpY4p5xM
c/jLx5w85sIbYynZYuKjDD03p0HtQzUOU1Mq6TBGY8x+DWzSjOfLQz/39vpMC+kwekIMg+R8Q04m
tG3rcvCA+ZuXFJdMLpFwcQ3fXuJGvZZMdAKogECccoFkmtLIhkoq6A7scscHNZJt0Q3U+zIQAs6e
o4lwsPoVK6xf/JmOH4fmw6/eTc0u2h91VwLkrarxAjJc3+zLmCi75bl/Yi8lxtrBOwK5jyH8YtR8
gr0t9Naq39SkppBU24UcEARfVEnqGhRpHSVqmNTF9lP/WVmOCwX7E8DFADK1YGu5qG6uw6dJnGDu
ZWQJ5WEdEoRrs4Vv+gK1KSyzP/XzssQ3UEYFbp+yCEWk7Cpp+/3Qk0XzL7Q1fXJ4gfgxXb5XKaZR
oPYOx1aRB5bOOohCPiYcaHoWZWvX6H2iS+HSvWXDaDjhEA+Z9sY9KwkUTxnN3arN8zt82j1qNzj4
iS9wWgtoF8edvo0xNwvREC2oBOG631LD5vKIhJv/qKoU4IBmt6a9rS7Rt3R3nFrHWaQlT2NRD3nK
sjHTePG+fcH+PuZ+xhL8OhK1t/FmNpX9T5UozGp/H5kOapSrkymlGmOljR1AjdtLII6ikZFwJIgm
15rbv6D5x2wvTWa2XDVXE18BkUL+M2gKvkEIMTiHjJgo/q+4h44kauamiUDXPsOx2N1FTHEDqUpF
WMQOkQvDcKTGa+Yt4RRdUsFLdYcJGxAOvDazaITmAwurJ41sNRk1AEh8R+WvSLD+TQrfnH0h7wfN
9ECZX5E249fY+1qEcFiN+qZv93gHwFv0LcJk+Yf+n3j8Ibj1a1QPb4xgW4CgOG3b0tO5v22NTFAS
/6fZJOmquDRLPEIRS1n/CRIJSNMG5i4ceg0ottsO8rCLkfQpHlJ+u+heFsyr/A/HCfE9NYiDBKlP
Ag5nJHz29AxbJkhMjOk5cWoaFajCefpPS4w+8QczCTeNj0GDnVMSBf72XPQCJ+csDrYFULcA5lH7
y06ND+YuXUqo5ReDxyTOb8D/XnEo5ixsxB278m/0rfTXoGqohEYOtugpzyAQ5XMcvuD0BcDfGWDc
0z6ZJYlZc8KESQvvrt3Ei2Xm7xiioiTXe/dfFNG+PrQJ7v5FIStMwmk5T3SE4kZeK17viMyU7hlh
vD8oj+NzYXAUv3cbsmbbX/BiS1rkM+yzj3ih4tUyjGO16pHd27YtQy+Ykx+j9IXQ9C/Y0B1MutpP
c6kURV/+RHf+YTk+czPzgPlxisYT/ohxZ67EyyPiwSD8hFuhbfB5QehTwwi5nOeVfne4E4r6i2ZQ
3JSIsEbTDVQgFt1pnQId63zBU4hxb4NjiwvaIsH1az9doq+YTlijn7VapXCwfowm2DFNt0piXYjA
DJK55LB1HfWAmeJv39UnZtAzIyR9FTBB7KM6rsgpc2BGAAgtiKv6NPv6oxuculs1expjsa98bFOC
GisODpAx0DcYA+BqbO6wS3RgzHFt6CkkcWrWo4Hrl1SPH4uzqux5N1ZXUUOWvPH1Umkx0grsO+a+
qq7+nTkCeXI2esiKwOSJRvxdA2e+u+v/41UGnoaK+fpidcd9PTri8aG2N7i1zKEge7CQHYRlkXRb
0D6T3LIEzjJLzm0cNju28hDfhXjEMjmR4iCeLggrWURdxS8k3rH4DqlEaeLppAPK05MtJQe5dDrq
9TZQS7UmNWsFNKS72I44qHydXjNWzzfNdM99fuZMWf0pSScdm3OrgaRXuf7LX1YaOHzYIHiqMjUY
MtjxXHb9FdU5b07m/lUGVLS8N4UN+SKj0AoZt+HMFuqw3Ngt94Cy1GnLjfabVeVncqujbbxVYDA9
fEXvPB8jgwt3FxwUJhkDg+9f4WtXVSzbE5NDMEoToOUkMKBPnKXx211+L/TABcZ3fyTcXJyLD60l
BPqp6aRCnu53tMOIrH4cfxJIqAktd6Yu7OcMxPbrhiL0XWlGZAi6L/WQUxaaCgxyrBSqbjy1IWzZ
gxt5oL7LzKB2Gi1c8a9NI7BPNNsxkQvlx8qdXjPeOynw09kncLFPuunUfG6OQJ1h/eEWS3zuB3g+
w4y3VgvfstItultx7EHydvnfOI78rJJb/6n2GnqelFU92M2vfNiFMvNCUbzgBAwBvgIHaFTABe5g
e8RxvKImOVFkgN7jAbViOjBu2xmLjXuvQeBDH+32cSX+KkySJugdXkL9yOeiu0UmN2hirtul49iO
rVzqM9NtsWwBE9vZk3DB/HM4zmKlx7meS9mhAC0w1oDNyWIu2rbNULP7tvKm/NFFwuOWUL9zp2uE
VgUoxrDglATraohNnBrOE2wEJ6z+sLESnN96W/DAjaasZPOrRoPEfUGFNSt550PJ0NMFOb4dM1jy
EwkA+cOf30u9V6azU3YyPX5iATs7IKTCc+rx7Ts7KEAga0dQ6N1nHTxlZNeHc7t11UcsEn500VCB
GmOL2VHxQgfGFYXTvt6myGRcTjmXBTT+OUFCay4vnbNyrQ6t6gf20BxTZgoZlJ+YluMYm2vbjSDK
wzccuKKNzCDbsHu4Aax7hSxB9M0+RF6TNvgBQYn/3NsG422EOO6dAZ1x9bXS6ONXXC6lYnBsLE6y
zVnmcyhwhopfP+WfX98/PMr67B6eZhglqOL0LAFynnWzoGRcXcIhE2NRAL0mCOb66G39YVVIsXW4
VgieeVXFjj3tii+wqNyW4Dj3w9vHzfEVPjV0I0aXJgmzbKNZtv0uKOnih97rqHaHUDw5zqrvNyT3
uMkoCaM3A37EG/a7qPerK349ahKzR6dWEnbPazbKbkB2+zHl8R3NWcAxr+zdlPRgxkpmte8S6rdD
gr7idzAw2cDhj16oUJq8duAdkovsUYj5jGrADOdyn4baGu0o2/x9uEBZGPlyAj31TmAewmzlFOJz
/aDR4u9FRj7+4LBD9IzckAZLJrzUUhTA3oC+vOgknT0ZRvpPjQICgM1hKmUyonu0iJGN/HiiyrAc
RhdLQ3eNPKjXQnNlaOovGyBV4DpvJHMKIUFffoV6or6RELzLoFWzHHTuRo13+VKJglgDXcyS35E6
HOgNZgoN8V40UEeAcFWVcKbUHeWC/S1hAVFt99qRJeO8EB3ukbYURpFyA3beNFnsIvLfyUX2xrIC
najcRKixja/jxYBXHQPQZYTjpobLLG4QfHdFAYV0uXuAOu1kj7PAT5ABCN5+rPTw5XpmPyTjnjoN
q6yYGSya0GOA6Ixb0Pk/rROiNnLfnibHFcJVYTc4YPpqgTuJ6YCNC16bFasy7qM8fBYqV9HofyWR
y+hgdNrlWREO/WnV5RhbjBnyPm5eUlAwhEq8ty18iQP+O+6l1rVqwXYNfQNNAa/FzGlE6NL3BgKP
CyfcZ3WyQgSU9BtRJVDyCAl6k/1QYpSK2otjfXNHUagVZ0P1aDbEn3MA7OHWDyvejCwaieqOAfge
Xbn752voCkieXR4YOa0QCjk0NGMRCMgvnjRQMypvB0c0bKFkcYbhLmum5XPDa0c6ox0uWoB4E3wZ
BppG9mP5+cuZzPrY4dLD5HQgzDvJKeZuVdxciKBQ28QTU/TrlIDv7EeykgpbR7K0Ou/V/MS3VZ0R
7//80CYOC37RnaiodLziCBYjlJNHfo2H9dyeskDo2hH74uixCy1x1nHVMzb9I3y7zacL4mcWCAVI
wEjGKLEtjcUjF1SuV9GXDtqJdkwcdKN5CAG6MMp4M2DaPneyiY4RqGPpTQyjFnQCOjrpszbnAYm4
BOfH86PIcJVM98gf53KHzM+RMBNHAr5dl9iGq4rRtav/XzoFGobBp7JgAhdzYA0k5xR97M9B6LrU
3fVzTHuAueLzqQKsWGVYKMbEmHGNioiJ6TwWmZYGgIHemnqvZOJ1Oh9l+jxruURiuy6rAx8xotak
3dx/i8+M4EW5Meb/pTI09JkfwD3ZIlX1k6k5zq2Tnzrbef09Keq7JU3royuHuRyXJqk4xzBB5uEJ
I1zUSvIYaes4ydP98PpdkWZhYGAO8iHqagEO2MHONcJjOSngFWJMu10v1mfq7vcW/ajQK1ZuKCyO
kPHqpdLLUkxVhhG1VYI97dkDPf2w8JGC0+WvwMJhX2bFA/JTZo1GyZu6vj25f6UQhtdpUVBDrv0c
49csazrGWWe99qNjPZhvvWl10jH3nQ1HDAZwg5kEfc/FTCo22pKYZEUbYbX4CML409Buuf1iKvx/
wPa3/vhC04jHo6jGz48kCcETqx5Ex6g8WK98OqO99Q2nVDdWfuU+yQJ1wEjgAcIGVAk3NuZmACfP
saV2UCyXWJ1eOX62jO6tYht79wqu/ap1lsoA4VSaSvdNVe35VS2mGyn9/ppHzaX6Nd/ESm4GKClU
YVaBNh25pzP+0j91IOAjdWoSkhZuToFHZH7mXYqLelUUFvjePz+O4abslnB3QRWH5cxazdVsKfdI
BXLQdJhDaPVfczaLl/Cxcm43h3jjdOR9027xYKAbwKR7emBZvRPZRQ50qcDcW4q7ObXpEn92HpAd
WApdh6SGt8KpciSPegCgn4fLFuXIZ0BlEKp+sYXOFwISxIrpGAKaOz+tOmLa0xtw5YlWxtTDIfz+
Imh7Mtk8VB8GInnc/ifEJspSscJSXRkX2+lQTnsEGvvJPw0Y3yB4lTMbsjpALSS04KLp3v0qrcii
au5lkyNXkRgvEEi2EAkcvv4PtnS5bxB8HpDBINIBjnRdaQsXH4Q+y9bE50T3fNZK1+TcQtfPCS1a
2xL07XMhKuf15LzxyYDI0bqnSPm71otB0Cekva597ajgnP6UMvpQndwISiaIrKen5+mYz7llk1zb
9dI48X3PR6B5027fZg31MPcKdhIqf0cv7s57Xauhm5SAr4JSz8DbgfaRyRHSOiXsHlwgspQGr0tW
WEmhX23POPYJ2JyiXE1XxWFzuGBU0uEiptV03jnrI4spaH+hYGEcBdgcp5RMQG+yKFJsECb6oNEt
c2VYF4sVWYIuyPzh+RL1rXgdQqCv1FhEs81gTd5D7lIiTCnWnkCx2hzDB9wE60moUzJP1p6MCo+K
uZg8HeQGwBIKLAf5kfWDcUQ3DKuA5IYVzmEDZePBU3bLzRke2gmn3p285IAD2qNqzpw+yfwftfo8
kyzYoVeeKeiVZUMDkXIlYaYKGKNuRs6w4xSfjyrydpVuv4NHkLMYIDWfRfOSMDuwbEaL2BT9mqY/
zLUya7r4sfRa+sy+5MJ6K3DEuJFbqm/K9KE4Mm+XutuG0V8MMMVPhesiT9urgeAoRxIEEM6L1SAx
8VtKz4nFjUu/hFBwXnb07kbA4a2X5mxvv1310qLZyIp4M/knBpFWe+TcCvw7qkpgh/aCUlnOkFU3
wjegnLCRPJlH35nB3P0I1S5LPJ1BqOL6WpEj469C7eHCqmLdIVeze3j4rTSgvKxbseFj8ztwFBpX
Pzqe2UU9poqVIE3fSHS55Tod/IPnsOjIH8LBO9Z5UOHySM+pU17LWLo2UWKqrk3PhNJwtLwt3pUY
sBBirqBYl4MAjXN8JLc9RWACbnePGb3YV6dkCIQjn5Y7xXxmTQ//rRZK80D3GJ19z6wyFdYCUq/h
8/PBxa9VXejkOArSasZkbAO8ls3ynCUVK3W3Hj1CIRVZ2g/N15uWMSNJ9XalCmORiySc/PMzeJ5y
xaI/w8sKeyk2dnTxnd/Xk7srBDKYchp73MnjePjr1I3NOQeWd6QxYkRUIyDQRrHkV+4nzBe3uHCE
PlZ771ZMGM2lMiYuLiEYKrZeNFz0aeJQiJbUiOtLwJhda4pieINmyM6ZcsGPx3Z809EdEl57n8yJ
vMLwmKQGiANOkj1rZ/ZZm2D8x5UMpBN9uiDEW83fQqFgU5DgVbgPk+NIV89PhkrD6QvChfDEcWaL
DN0lab83Jvj+nB1tQCWMst9Lt2PN+QzVyzR7X/wlIPR7xMIncSurI4H8b9jc24hs04H6FpvDShS2
9Hu5bdgDXR6mXj50+OSRdd6pw8BwLG+82/HcsZ12lVsnAUB3yo5s0uQAa+o6nfJWDW8fRgxEJkfa
ojyx8qPrzvyesz7i7X3hcWyUGmzmigg2gZkCD7rAIPVWC+7av/XEhdC7v2947ST8Jr1nCHCWq0rl
alPeMyQfEerb894Xcem5qpSknLM2PX2L7B5pErEOdVYa4K8LDqmzqJT9coUlQA42fFARxSwZU8HT
RhneQVXF2nbDPu8JtroHiGIK6pR405A9SgUwk7al9E3iDelIPSPy7+v65lv/ADmK7LAkcuKoGLly
EnqGCn1WXFmCS1AxSIWAuhnPXf55Gmp8nyoLvrBtyqdOQIvazO/0QpjvRXzM88Iq8rL0dIj2VDoc
5y7JWN1WEz9ly6wizU39vfFHyljSINGOIi9rPNK7I9v949fKku2twyr2El0tlkGyckB1/rnVMdwF
/TznwzQZtDD9VK5iZ0FuxpUUH8vCQH5bravbclfPNw9O5wpln3u/45ds2rthP0IQfMyswP/Z7v7L
Sq+k8SmvDN+knLvc2QQRv3EA9rnTbu5NiDS5iOwkiYsTzg3x1NOPmSJHMSmfneUTkRUIfrV5OHbO
mWUyGTDyWwDPzEh7NWiuKBtHu2JH6T0XNtxUR5x4Di1IkAQAg8jQphbd3IgI6ZShYEbPOhVVDoql
GxoC/nhlrCZF2WVxEUPZcscqH/ogGQCtV8xPgSoHmO70d11zg8DAa03dkejiUENfMDvV/QM+hQ54
0csHOUrryG3JTpdvvRWoEgYwu0OpQbtsrnM02yAse85fYxFaYuhvax0O7rGBK2gcUEwta48sZ+5E
MKvYrLo3swoZilsXogVxrQKkEKytItw2Py6uHL+XwnlouSr7mFbtJyvfLTzb/dcqHtdzscNZGB9R
88tGlobRR08lENt/MhR0zLPhVqkO+yBQYFW2Jm8H6KZE4uYKned0Zw75/cwGm0+BAt4NFh+hu8zV
9CgbcXrO0P+1xn62Di4LXhzxBydN2/AyxvQItxyFHHJx0jMgFfgBo5XuNUmp24eCaaolzHLpyUAR
itRlCwChSi4DXEJiVmmKjGkgiCeoYAAlf0NBCZwqj5sne76j/EDXBxnRU6VEujPV2SWNuHP//LCM
jUArCtpK6JF1+6ijjmCoOhwgnPHRinO70vZ5tJMjNKmbPDhdWFAZ5qpi0rldOVXkbUgLFaZ+jRvX
ZSyyH1Ynf4TSPuUggaRPeThSS1yOfxZf7SEFEysis/rcwStNVl3IYcBoMorWm2W0fzGVI6wn90X5
OSZgr7kiTJEWqW5/bB7SdINSXwzJgOjUhuYNk3cr+Y60uHdROuMV6bnpvkmJ/4pJvXvbgouq9cyJ
b96/7PccrTUG/F3eQeB+0fFPFr0S1r4mGcnVsALcQlIOsBD1mrpHFlRM+WvPvIgArIW6zyqYttIC
5mN/WJVLI3Hp6McNgRWyI4nHb0FvWofS5OWaTzCJxiWdxw73BBLnEYWzfMxIyzHaqQf7flOjg7mY
gr8uCH2PEw3uOkOO+VRarIDU83OWCiz67jwD5HeS+wNS1Sb57o5yZJjJhFTNVzMoFBbQAP2tXD5Y
/Fvk3i0dtpq6jMMYZFgoLBxz3DZtT02PhiWniOyEobntKyXR1Lr3VWc4Lv5ZpnW1zL2+3Pz1fEG7
bBhoPLBYgh/umz4vTzAFNBHl5YcOQ/2hn2jVim8nGOCCaB/oT5G7GpUmWE8XhoDfSCSIOrc3kcUg
iB6xYOEXw5quUTZqTOeFTkskfV+pDKFrUyvnhDvtQ9NHcQvBEyEWF/62jGG6gcvLFcvVcgy092Em
P7BzCl6/RCUAZ4AzCKxdPdgjF5/YN1jZyEosczX+N/iUDbOvwXzdVrO9sGOW8Hr8zQC51nxSD3+Z
/G2FLkJ7wlIyAoMCtmFk51k9yNrNA+HSPFHkoxp6ZovLQ58rr+0xgDDNT2GLuQxZVIytpI/Nfbw5
L9wf/Gesqv0WFO29cPZe73uTyOKb8QSd62MRw4nnv3CoydVdDC3N9mCOfeOqha9uBwzMm245/n5v
vrlRbSZf0eGEr5P9GG1UZ7WFH8V1rj5o4eqG60dbV3WaSHl8pFWH0GDefqiDGedh8vpjJ5BbHTTY
gCDIbV+yKmy7R5JMJm7Deu9FYZQDGERQLEIswZ0UyVdQlLVCcYNI0wnO4xJ1DYyTstbPvT+lKHsH
JzBGFxt2PYpSRnwt+CcSOn0ZkNeiOg2EA8AR4CLil6wb38x5lDTIc+NN8ASLzD+NAtW7ogUtu7VX
f90eIApd4/gE6M5jbE6nk+jEXh7HLlK38+OqVTsDZob79BbGD1zLa5kR4KftpStQkyT5TcE/7C+h
PMWeqG40FYqD7IueIko8VJBHj6Q+6bjeNhvo8Stuo03NdBCLh0SBBRSWxHtD5qtUnRdU3pf/vMfi
Xg3lNFFdxUbnf3hNRK5N6l7mOKrm6FajTcXCZ4HhMJbLrvBkY6F7j+eVRV1OUkpOdab+udjHQGJJ
b6ADhbcbIhnSOTyOZEfWFfkwlx0n3MR++1RPQoFlNytK1VRHi0nJSBg0xU34c+gJA/wnNLU4W7GO
lYDZNZR+P7JY5szLZEd1jAjKWkQl0d68ZHCIAt2NRGSn8n+OoVxnL+xbTFxpilzQe4LqUnGhOlCF
Y/emon6/1/4hdq4oCJvY+akC3K6c5e9zU7GFgDl/kNJ6Mxkyru+QQWo2c5F9aSVlL98YnUmWW3r3
gDXHy1/0xNLeF/qTxz1uhaiLVhJRFemKwaEsX6SQQRn9o3gMXa6ImMVGCg96O1Pw+jRty5o07gRP
SgIEopWcU8/meSMPhWXB/1oo7f4S+93l2hmHdnPbqzUCQGGgY1kIznpSuFjbrqzNGJwugXYci8ZU
s6WOCgihyZMAdgKUM0vnFvKr0BTWo+trw5kFaQyIajaGsnkRvBzEbzBC7dXSwK6p0Pb8sSsi7FBG
tuTwS/4oIiO90pfzQn+yrXzVRToFRkUUDknwqRg8ot7UpoAUL0rCBra6suztn3PFjAm8gKPwB+Hm
6XrQvEfbwUA2y6CqwEs8xhB0DbYHY7N0IBemM5H1E5OKitt9BS6wFAkNGvOnqWCr0EB/P+a8W2hk
LedDWaj2ysEr989xkOApYHoF/U4EoGN6yhGpZklbqeYKWpBKHAZLn3AEkmvRXIuN+P5tqW32h/Pg
Yeinfk6wWjXiB+aaTGuirGZ6SAGhe34mzfJ+yMPau4f+pKPxf6arg4XxIZrNZ4w0KXr20xTatHRE
rqDddkvwgjVItvrCIG0AWF9mwjzHuOCzuW6Ac8wS1NzAxzNcpcww41AtZzPBj3xr7U+JsJTMKKaU
VcumAhoWeBZWL+r2y+jFcO6izVy/BrgB9lerp5d/5aWO3J5b21x1LRC+bd8ThwojaDh360dUFOzH
qizG0qLbqkB8S/WqcRmq8r5+5Egj6iovpucvx00WzZaItv6SbZDMaK9srSyAorQps11BL4Otwf9u
/8GYfTcIjAGpOZu6qUT5ddCdHw5stc4FLzVg/ZGT2ExFTeH/UKc1Vny97zQIqv6Uo0BgtO3TuX7N
srjqVJ7BicMNWiDYj5vSMSoStSFLFfFVfHYyRI7XN99jRt8/+trNlKsEECA4/cvJhlNLrDaYMqFN
4Lu4/MxEP1y22o4mXLMw4W9ehvv4PuTnAsPmzmpzmWwDGw8Q0yXqpC7y7z5wRGpukuKwtnjSiKNU
pRV6TB61I4XmXFomoQCgrOGegj1s4gLAysjDn1Vu8fydMhJBCFQlsirca22sYgBUgN4CtymKZEZR
yxx49QVqG+RYAPqqKz1iVeS75zngqCwr7BLt/Xul86aGW/HrJLxTYstydTsDGgh4HiMWZyqNVqnx
MOt710ilQPqoC/7UpcibU2xt4tuzpW3N3lEe++gi+H8PcTZFqSHZP1+MBFK9Zql1mpyERbxWwB6e
Py6ahqMcGlebr1OfBvpdIkQl/51OWY+Y4BB+w6BnyyFqcaECh8QLNyh/t/lF2pjD4MYF6AMZEekW
FgggvjIXIq8zQL6NfpNm+A5fES6qH6zdy576eLlkEh31YqE6k8xLsCE05ySB/llJmZveFNB9G/oC
O9aUnR8Z7QrcffncMgc4S/DhyJpb/kEbCZ9r03pVs90VRemUn0ZwkcpuF7N+LI1xgCefV4aYvxap
WV3UXNqY/a4eU87erf+cLKW1cR+6XiLe8btE8lzAMgyPUsO8d+LSGH50UJ0zIvdHnrh8y3+MgE9r
en3WMZBr0jX7sqOIOG29z4HUpeoB5iELvcTpDqjR/NWlPcWM9HoMl4wvVQSxshQuHGy8a6UcHnMM
cwbNeRaNvMsLYLZxMTKldPP1j7p3bvX6OdrivOG6oRJPtTU1KGHGxDZGjHRKjXeMWLGQnO0J1hjh
w3amRRDhMdXsgt4q9eQYGaF/bh6AVkypCCLuCExkBOlXNYrj5yJTNbc6wPGeS//ILvgAcwpHUhwM
UGOEMtu3z7q9JLYN5uB6baUeFPAMkj0/y2HW3KePGQh0FjqhXnvAZjyonDs0NYrMx/084h9Qo/jh
ctZKJJLGpvUeYhLAHJodoJXIMJpRCR3xjG167np+MBgLzK2XSQqhp+ev1DbEpXhx+szPqTWsVRFY
WZvHgObUa40WFpcSm0OB4S+MeUAe9w8IhIxefpmNW0yGCqyTOAMZEb0NkvAuUjFylTnjnfbtjA9X
rAUB9U/OV5Abp5b2ZICsSoCcAaGJkZvyIZOiBrgzutR9c7ZVtz8Z9LjGWgaumNUSOdAEV9Fxr674
2V+5lNNNGlen8Jz5bAKrDaZr5jS2az9+pvCBSw9Hq/S+Cw4W/QBTko7uJqgPhbbaGhTqcozqAWCF
Ys/qLQbL0eK5hgSznMSNIpVPRvLeLUSP5LBiQ5Ih94KQ4PWh2R8fe+7M/hEM61TY1ybJJ5L7AYZ7
564/unnT0YObj6GO9YOFYEwQmgeSK5N6TI34v0cFssxQagObIq+ttSMjOA8gFyvEi7ctpiDioPDA
SNLQ5BsLOZBB1Nb8rlGM9ORRYMY+A1r/oPmr5MYB9OlrKzdZ8mrXezEE5rloW58p0W9uTWGuHQux
bCWQTxeiMc4t9sdeQRmvF231QXfGOwbnWs7AV0uI+di43BCdsi7/3JJUohN0z4KaHRZ74Hvst32+
pFTn7wWjtfMiHf7OQMANYUhaGYGwed6C30JdipdiDsRFkWkoI3G2I9UPdOYPtJ7HNEqe7x5gquYC
moqnN8eT4l3U3JR2LopyUgLPv7BL0opM++WTQFBaaV8+VA19DfGh9BMnNOtr2vq+oltTZLXQLGaW
vCJ9SvbDRKA2CL1IOgfOz1v4SVdb2+pKov7lkMu9LfqM+CQRYDLSme9pDBpdqWbDGumqEA0WDZ6W
keoIcUJI9zAOrThkaBefvPjD4CJlZwyrs7hSVCqMZVYedCAo0hmmVL/d3Pl3T1cC7iS5yZ/q6lO3
IqM81ynsiMLoKlE50/+GnUvOy2Z9KaVc1GVruCaOTj53OxsV+jEptsPz/TH1nflv9lYZzsBsrCtB
HOuj0TFpo1DAGSkt7qb5Kg2k8/yeoiRbZj6psATKsIM+1wL0jgrDBtWyJWeZXbek2Y3ExbPBOqTG
RAWUzSycNuCq+QQoc18fVnt70IeFGr/NIPLXeMVMwXgx+f4E1GkKYmYk/i4xg+PB33Ld2Wq5GVWl
lM3cT5A34AoNAn9RgZPfmJKsv1yTuvd6+vFGZCrYTFTkFvVEvKmVw/BxCdaAbyrXfgAuD69u93zU
R8gdgTNtNuTaq+kgpuCm+1UH2GxIOUk4NUw8Cnvfd3yx+6C8IdMUhQ25hpS9w+E3TROPflYvGnRl
9Xyh/3P3kYb0XIOod0H57OF8mYgg/7/DGeC3DCnlHow/DDfhL6mPqcsz8/NuUvFIfYgBbqnn27IU
7gIccVvng+oW+TpFua+EgVAZv8QRRC/Aev/cmzC+7QMrMVoP9CsiUM3z0UZecJufIPHuXxCkT5F+
YkkY9d+18X0pqCCqjO8ZdCtPmMOJuAOp+EgwFsbTkGeCgBBXfB4WtrJE+xbWKo/V4CqNjFdvYA70
WkHPYDmykKN1g2gdk4vaNKfzg4jEad/vNnDh8Ff4u9kP7cbqle+8ciLM8xV8uDNZk2O0AKKi7Gc4
3HnxcO9yjLykq9IHAEazxa4QJkRoggk90hagxwrQcxysU6m5VRoJup9TC8XYbQenC+4jHhwxJm4c
XqalDlla8LrHp0APAQt+rJbPxFqR9zJmrkajsSAsF/uO+HsnQ9yAqCCW3NtX88tzNCaLrtllzFxZ
jgd0SZBbUHKgZshfpTVkOrarkcd4UsQh1d5Ta44qKqoEvyGvrEJviiSa7KufIAH6GbXyvlh2Yma7
fT1qfuxt7yHKXw58XJtmhduQXfGv+pFpWlVZXJc/P+pBoquiLRTLyqLT5c2dTuBNKiTOSCTNzkb6
eToJaJAeEYlJt6ZNs1siEARsNFQDJ80Jx1M8QLb9BDcCQ4vhhRV+AnOG8mulL61dC6mH0hsu7Wv2
2aQDHr/A0IBVhg5HNOBDmL99mk2P8oNub4ghbZU5DibxjsNFmujI+OwT5XfOWqb3FhWStCYlLZue
33Hyw58DRcSA7LItQq1KgnCSmDOEPJrItesHpJbc6N5LfXbtpJQZr3m8NI5xF8JWEAb6Av9rB9U/
KGWh4UxuLvz1Mst2oEc34XkIzVHllcXSv0CCiJxtoM0LfUsf6v3NZeT/pvOAtmDP3H9XGCXInudE
cXKPbHhgGVIF/0nfBZ0xDRV4HyYsYfhAYU2m4eKvuATskONttIoGhNaYLBhyhdNsZ/Ac12Ah+Xze
AZBKE9xp6go5/+artPdQgq67hDYdSzG+VrI+WN0hXT01NGMxdW7IkcKXihnrya9Md8jIVYryUqYp
EERcJbhNcmPV1dGM42C0HVrUO5SevUSLN0FBXL2/bMqvGi4LSxa7tLSloEOz+zG+FbEFBidWoe2b
QBU5x9vCcm1gMkbpdCFNrK8Pi2fJ7InJn0q71uf/a9DB/X1IJfnYopVFu23unI6SWmZXiMteeeld
HsdWPeD2ZrhhF1yo6516PJFRs1hlnsZU2wlaH4HHt9gbjlCCK3suRm6tMWSeW23ejlHX+6WiIHSn
Fr6snO4yG1Ln88T94A+VQSygmvWtgi+iUUqNIMjJ4/J8qGuxc/fN2AvkIIe1va4M3GA9d2oenH4o
xqDClk/yccgCdWM0qK6B0CE0yaX+7AX2q27cYOkBs1JF6cfcUclemDBZxeWF6uC4vBNBKU5zoPTK
oO0/Uo23YCb2beqduy2gVxupSkDl1biavobIczCgDBj/7kboyfdIgSN9tE/mRVnXzVFUfsSJdIUx
Zxhz0WAWrvGq/Hg9T4n/RjTQcTXbakVv+UlLECfRq8ESh9zc3KASVVOlu55TgP1ovuaj8AXrNsSm
JHX4DOB9Tl9KYo3+1gP0tBmfTKXZDy0GUhAp7bzLuJKVoaCnAg32A528rlDFjP1vORRBP4gjaMof
yZYm6EW7puCJQN20OqGav+m4YgOzi6zyWvxbW4n8OBrwoSL2hofNOa3z8Kwbg6G+kIcpNXjkRTZq
lb+CsmiHd3jsG+7aNuWhGLoy1eQUl5JY2gYXu4rrnZBp9xmGs94Cby49ApQbvC9DgjJTVtUW5iPV
gvJAapPzKMvRzVn6WvnHX8hs/8W2+PHnw8ikJLiA2s0dc75Mk3YWNCFTbvMn79AIZDcLtM4yfN2/
s/RozI7o0YsNlTjdu0yX8n0gydEZe0uHwXvrKN9dL3MnttVlZ4nIPbQS1p8j1W3zs6uuya6kFbHJ
RjezzdeCnb8Y7/Zfq+XX2hGL6XUy4Gagf1qqIrUkbanElvII/Zqd+QMdMV1EqKir/t7K8738x7DX
l0oEN/3kJBHcu3+TVw5F+9NnvuFdXiROCxwOPuI3NRdue9UGr1Oyg6cY/RW/XCejWML/EEX4QdAR
+s585/IgWuLgg4JKOF3oGOlEwOpzUlZQdkXfFapSjdbDJiuWU+lMIbjXKxHabYpv6ZAy/PsFXKvj
5tXAA9622H4VMTerzmKK36gVST0ri3uKWODTVsLJFMUDu6DTMvbcnt5ShiBv6buC6EKCugE1UPE9
h1wCcJZahH2ALm7uoMEnp84V6uOj9096Yj76gKv7F+3veWFmWbPvjFg79SpGhkxpbLau//FyoHJC
auu1bSyO1591kgIj7eEGztfJJA6aKzLktjr8dkjrNlTn25zY/ptRA1Hwt1dt2Z/TVOBzvWk2wJx+
T5f76AeJENUB+KgvWEpopfZWhdZhLwN3K3eqX5fRIT0IObjjvVh8iWDxe+fvq/17WQVuN0TITWjy
3E8Y29zRQaZfkvN4+fn07wJvuzJVqbLiT+dBgEEnHXdE8IK9r+FKeexbDKWEhY7+TAzDtTSzl4sc
rExIYvg7KPpomjx/BN8JffhRAmkh77mE/dM074B3qXmVmKpjSCGD6qiFV4f09mAP2zi2Y01oZXXE
g41Ih77Sa0LpWfBeoAcSFN2rcnGjZ4/1gXKcgnZbXlNyoKlb1mJHKfdHD6iOPaqS4TQTFHssM1uR
pMJctBZdJsmkYCfgTsfPkdJ5ktxVoeW2ugV8aZ5vMGObh6+m+F7PnSdMrqzaG/66Ncs7SNsKjeNY
0GA7PWJwrlgXw8MW74G1iowy94qvjX/6P2hllUwbHLtST0ZzSc7PGn2a2kKwSb2r1iHlKnuGzNTI
u45DLHf9hhlano5oKm5dwyT36RV917SBTGc63fG5ZE8XDTm5nTxvT1v+GwX24KfSRVhUmPXUOhNe
mwUAgD3noniOcLLE7pZyV/DpQ1JO+Jlrkq1eInfFigHHuERBceaxMfeGZ0aN9cLs27ZW2ZsY007l
XXYKWMXHHbnFfYYv8uUhFARJALdKVDHt+jTFyt9rGG2izQRSbBNYiap3f3qpJq3mIxkZDc48eMsR
nJAXQ3UL2ammRm5KUIuhPTR/fDSxBEzFCEK3V3UG1qTCuBHvWJnY8a/gWalKhA8p/E1pGuDrlXTz
ZbQS8742GrwHICS369SnZBx6gvEhUEfZgT1bI9i67tn2qUiZSNEOjRbUczjH8a4IIGAk/mZZv4eN
HpTGDqsjc46XY1a+dZG5WqQ3Kp55Th+qiJjX0jLAjp34VRuZKhbjXOfQZ6TUKMmB9O9TkcGQhKlP
+Lzsg7/DH7i0geQne/c6ThmkIjFwCvcdPwz4q19wHY0aGRghiu+oz5FwxYB+5S25WoVyfmHlLlWf
LZ6kQP9kQVSRgNKgXxBBeJ1p83PrwGuVT3Xgm33ytki72JNJMfiQgUrO+084EwsYWdMNoTq8OgdT
QV1ecxqIR5FFwW3isp+JtnuA9d5aeEGAWcVXBiWwjOnmZce/RxKMtAUGHWIMI8/2m3/hXS1zoYf0
YRjcDLr7eK8HKLxZgkMKgXfCaJScLzURKOFdHnTJuZ0Ei0H9dobFb7cDu8tzbaLxhxFtxfdUk7C0
t0FWsQibcPnzHD7NObbz9ETlt6lXAKebF+aw32yDicVvZsMUFYgeFyQxMqqtTaEBHn1wB97F8oqr
0F9YQvUN28+kqs+6MwP7zNf5Y5XAZYZtBfc90ZlAp65X+vRSxiZupdd8zj66fj1fu6N7hPDVoj59
gmsSIduFbzN9ZFoswnxouCB/kMVpO/z1ExsS/41+/7N8mYJFZigIjGbi35Pon1MJhwMZlYKOAPPq
ldU2pY9l/yMV8i6iqjPfPThRc0Zz+w+qhtj33jdM+zabcUrSlS6GlUHbzAYpon9mchyWKEOec8jq
nq3LGF4Z7eIjMsDBTONXpAcLQnGujbuqoUzw/jMhP7rTMZ6KPF1IIy/uoOPZFy0MnwKO5Xb5GcaK
qeTw32apA15XZmPPhfdNq5TaUkDuaCbl/sEmf0aWHrkLY7SUFPMKipDa2YcNNkYhbHXFDdRhcaIz
rherfAnNePEqvKEPqZ3y76yr4sR3h0E84aPJ8qDD4zTpCdgg+1inmzOoRwYMpbDsuZD5d3XtJ3Yc
xGBfHI4qYirCqFnVrQ781lQemcmuHNuDx37JnPRQv+4I1qHdPbR4z1O+mWNgAizUJQs6O6cz5kq6
0wQpvN7lkhvpDkSRGsRZ363GqrHHlB3Z0U6FGPTDaYH7p6Ilt7OjBvOtjBTn9ZnrrpyymDJq/57k
D8GtVU8qcTEsniDvWXzbtXSzUuYALJ7hL+dU/8+0e3i+UBJPSe5+BzVUwwL+A3UOmSbq7UuBaajg
P4vG82Dv74SSmA3v7qO/J35HPSQyexvlmqzqjn/pYxhEgqoQssnZDSTXnzfSF3OypLwYp8W/3PP7
hFn2YSVg8sTeKL8WKdVcUVOlSObyZTf7j5Y5fZc5Ycjs0WwYrAXURmjCDsF30EN/VJ+SRVnqucaT
zrOW8oBdRL+L3jgJTqVCLW8WQWsIFL9mUhRlhYykUTmzsqAXT5hyvpBj8lWP0DHclEhDCQhIiR4U
aEyM5ZQBwDbKMB0x5sNda/G5NS154XrzYafDvx2U4h//gZrhjs76+oFxkCrSldBHyhrSgJddXt1R
Vm2ULoFh2chn5UvNfYH6PaZEIIN2CjkYv+1mxR4IGAd3vEqafl+DosbPJpBBg/p7xsFofEUD8rVF
8zZQsc04TKfoSyaH4tEAJT7HqldokkzFb7bQK9tP3uzO5FBUfoS9TCxDs5MQ+MLODouSEkoTFlmU
Wg+9jCvWtdL2/UEGcxQyD7C5hPHrIcVpSzRwTx6oQy0NgqzDgMsq9Vwe+xRlcQjmFXw4PPS4sGjP
JwTy6ymU2K9tMGQwFuZB1wpau7X5lZA4FjAJMiLCVJgnV6VSaPsUeEwz+UF9MbhLkcBvdCyLPPAu
D6kOgakDcESngaCbTc+lGk5LW67k3niuU080g5+jbbwy20rS4EmTFAb2hk6etsTDsaBtIndmMnt1
cR2XXcs4blicdXdFjc4b7mrxbjKtlp23XCbXwFfnjZQ6k9+OX6q0rN5xG/BGL4lUF34pD5KErwng
77fxnFi5lC5baEDw7bxhfnyhQ37IRow7f/xvRdDmyrK23UcC/Vd/mFen7JgQO9AeGI8Cpy6/o0yp
pz+3vFXyxRnGXTx/NXMNL0wElRcNEwIRMMTNcnO743WoWeGhW0ZLoHZplZDiRBdq1SVFmqAPcwNN
8IaIy82U4c5clhAEAlFF7Uh2nFxxrSRyahfZ3ZfsaCH2xGL+uC2qAG8kuNp+9gluFWFjJ2oedWgN
3AqR5xu1A5/JAyjrXbeIPd7V3oAct+Yn0uw6U2bs3t1m4LG437mlm6hs4p82MW7384KFqcGdwPpM
txXDhH0hqBuu1dcShNHZwJf1sN7SV1p1PTYE5OcIGZRoH1dgHe9GKnfdHCyjU/TAv1AfSWRgxSYi
NanS/MWzVOPxUuv/yPIiHsZD7+xTSw5jl/fdlNRqWHyQK9sCqYYCyS54IONPI5x3cTzNrZz7UFC5
uQkpxISoMBm+/wvJjENIqxks6OKzkmDGOSUOOucWg+fN7Grqv7lg0hcJz9EfJcQ+BuY6V0NbHdUO
PY9koPfj3njoGY3b/9d98YeMqZWnkX9dTO6wzo88YBiLzzytAlm/bnPlc/PSNdugkganI1Wx/FTm
JrjssnfyUrU3ysRlOqxXBXjjpfQpe4do7xlxFDRudGZrEV2T84hdXZ/YMgs+aOCqty2NmjWkVmvN
NWM3VF5GuMsQJQRAxn9hXbMyySIpiEomwYUyC4kEEiUswIwbwQ9FUhnwA1R2HTZ2j7lTjecI69Qf
/iFuLmrgn18zC9LN5JyRMIoNwNFwEvx0qauC/ntDZJOFaQSlWSizpmKLMihTOAdfv9HL/2AVOR7C
MDbZbyh/wq4nVnMapx43sDJR9r2J9uxxcQ3iCN5cd/s6ojvpeW1B0izXRzRLD10bRIQnB7WHdcss
nmv3nzlaV+dyvHT23PiNV1Nx1mYffa3CgTfXO33mxl82poN0tW0w9YxBYIYuj5zbIxd94bFJ+kAx
dgCCj+ep+5cGV61dsK+KP6YCs9YpDWciC8Dx5O7XTQCTnk/zylSttnpaBaEl9BYiNNs0DCmLUsxv
XRu702m+SYoRrWHDFKfeeOMt2jzL1a+B85Ep+1AKcxTqPBTIOEwG59+emdhRQmW/DdVOCbqtyYWn
sX2B89WydW+yeTx0qxcyit7PHBw30yZyxaujxUxDFPkjq45CF0Pdo8t9TCKtkcVD97OKKWCXXjQO
wYWWa4vD5cO71l4DVCBuI7hlxxPLiYv61pyhBETGAhb0envV8NzUW4Sne17Ohrq7Gj7H48kzxGbz
q1uqpVlUeN1w2qiAzOxvnxTW2mQA8W/U+DJVscMmsXBWlXO4JkEHLmYEZiFABLQ1Sy1qmx43gVqX
LRxPhjbgt9HS+STLY4vZm9lRoHtlPd8EXgz+m/zFXMvC3LgAaJX/pbdVTkuAno3SMJqMbXUT364y
dARYawNNAf/tMf41JXDMLigFQIDb7mResgPce7GQW/mxC3gI3CyYPLOKtRTF2/ASKTIcW42cb0Gj
nzHdbZha9f9rp+CXcd/zmQG73z3UVbNwkuYBPyUGKP7KM1Cke0hHLXn69WnrarPRPI5p6OylVjQ1
fonr+R0Jlmdvc+rreyFajRh5PmEnDP9bt4pyFaFC/OSfdFbdvnu8cOkcUesPO5NM58KNJwO+jchQ
G+4hYSS+1gA92r4W7Xy9HM28o5YdZAwMKEvOwn1ptIHAf35sTMS4PY+xiZu/WyfocKbHMCDOq3kA
L6bBKcJMGhSuZ4EQJ1NqPHmbyXUjzF0Rfyi810IdIY182htBndOyNGOIJTOtvUXqyAyoPHSu64Uf
UJbgaXq6O9q5td9ywgGC8udPWRpZu8nFfdyiQlpKD6salj/z9Va2oHnJwpY7K1tqYf+KHHl4bnGa
CWqxp0b5GD7ui9t0B1dYUcoCllVTUSGlDxk9/sKUzNWk2OWxh4gyIvp56xlXvIc8hHDu7Aj/tB2K
OAJrgSeNOW1dcpAcKztRB5YRUqkxd1s07mogELLSLHokKZnTBmnTDwmEdiCmd0QEjVVY1gYRnl1m
9Lr/b7n5BhpesL8ljzwd6xRfig2IFPWLFeh4cej5pei462leMPO4SMLEukJ2xKZVVQnRC7qyaObl
mfanN4QVioB4O3ZdacnvNjpohG9Cdf+AUV3kZfYFBPpPjzVcSQ2OlczYo8+OmJmt3J887mbmNXrb
S5Q93b5WBe6Jf9C9/K9hsrU5Kp6h46epgGGYoVOYRmnZeEv33MlZGTBAKTox+iujbNvtmYZHB6/r
C8snWVow9+zT1XKnkZk/WeeKwkasC2fh+TgSKGvgPfNGtnBl9IUv5WyVG3BxayfL+9UOYeVitiib
tNjtPcVfgrURFTxYcf/l6iZ5JKdWadxiROVr0paWgl2zmXKdkXWipV3X5VwfCRqlvGD35hZxogs5
1vooLNezpvBvI93aabG0xHit2bS5RidP2vfRZo5odoJsXk5O4PjZ7GlY9THqwKmZiuviuXldgfbY
YFusl8WYrpmlKXxg53DCkOWdlhiE+fTCzTjvV9D6ICCYK2agkrIiYPNC/bR/s9V+yeWZgdkFeqEq
/BDgQlN5BefRbigNfdxVbSNqJXhwxmy1qZBEc+c3djVZJ6kovLIfa2c/+0P7eCziqQKwVrohCYdn
G692hvNNgPXRA2wW8f10u0M9gRBMTKIvjfRAu2iespmVOEt2eUeTWi1ca6T2N/KQYBkdBAPRSO4S
mJv4S8QzYG9j5r6/tK7sHs/XSVOH9fkBIjQ/7oU19vJ+5aF91Nj/Cg0GVosScseP86ZaKmMvPKgF
aQtYqXBLuFjC9UNiOoR+zo60+Il97p8SaOGzsgsgdaBJ3V2Sx3tn2RFoBGOW9EweMlmSiIYoKa2m
3VKfS0GC3q6nxoR3bKf81R8fOSVMuD1GZwEuSacvLiNEpMm2IRAeu8VYnYBCg6yHkq2R2chl8cej
10zClEwWtlb/3xiCf4EQe+mhvFFw3bZVAnXBVfZ9I8hZ+VZYpc2JdXyUj2il2sSQZm8TtOCerL2o
/eitGUXSUW4Q9KUOEwkKXPM0P0+eTiAEaReseBRwhsCw5dgR2ImSu77WPlUCEutaF0CEPQWLvBO7
2vzx2E7MXRh/He05pSeFKYkkVyvIy4iHocajIo0pEWJIIM/zdy+jaQX7PkwKfvpiZlRt+RIJigMd
Qb4WzyWERdooNWPzbyRfTX1koMXhrIeCQhYU70utN7PwzGdYsP2UU2nQukisBVp4JfH301Zz8+7r
t8krx+8Zdtt8VYgVy09aqd1Cdgrn90xYMLOj9ec5/AiXodn9O2veR/6X+G7XTFHxkfi0G/kGseVf
nPZqtF/6pYIRp/Ln/5DrrYKMEZmZsSBqRgfcULVDXf0o4y2AavaAuDilvarWcOn9w8wNVv26TjlN
LxIc2XwapMPluwTIbKAEfepWi6hx992xQphmkMI3ty4OOQDYJKJDCxuGZZRkZi3+yRG1qL28ixbD
O1sO5qx/z8psq6vABj2LqeLkSJ9QlC7R2X6H0QFxdozEnyRDgDjO+fNjE7QoLss5kAlrZVn2vv01
h1i0Eih45ygFGbiGtoeqFFSEGYSE0UyeQR4q2CEQD0iYGpfaWjWO8K96Cw58tSp9+mYshHUogVjr
GBe3KRhuPEIiZzJ8JkYO7bnwgc9mY+Slfmbwtdm5h055MMlllneh3iYgAX+dp9HzW6fE35dsBZVq
WQzpAP/1MXFyIRKHjJETVNbb8W6Umu7FopCpFfTnfXWQ8Kvph0ibjg+f5vSXYtyMf2ROP3CLYoQ2
2gAR1q/YFS6gTFY9mMBuFM33llb+0DL2FEQrOkYlfxxaU2vIV9kpOQ6/bUY9z1femoI0T5zkUApR
SdgIW1R6HCcFkJxAw/rTJUc8UF2pGSyteCrtsX0iGJkdv1n3ezCnws1SaJlCKMj9+K60WgraAwH7
98uDPGbep+obF6oxUoL3Sv3E3iDgMmovqKWC8emjxO/RAUiwX7VLNzbsWLFPJM9ceW3/N5kjBtzs
jdGOh2+wCL9Uv1x4FeNJx8hWUQKYSN2twbDjeFLBaW5FxPZ1ZtUqBfoYhWgTm5HV/KQx8yao/+am
nnFnLX/2G7jzJTMXI+F008RvXr4N8MR95L98t34GLRZwbpPe3jUNkjKyuHoxcQeaRcktY1ojCgwo
9j+QRZWabNYKllfOVhWTEFnj/2O7vXzCkBvY4EO2a8ybLB96IcY9TTp90Qo6B02t9BGdZF0qEyXC
4rc8kCC3WUm9BgWAydtuYUWn1Rd5cRXSVEAmvkqhkCH2xnOjGJKdzP3ueMGTv97jbUEVvcIqGXpZ
Anrinqm3GZ+WseiMaldJXbaXpnb/+Whi2MDwIs7iDkMrZKVDAxy0V5kVsoaQ5O8BQcoHMc7j2vF4
AWl7FkuDvPiBUPDrT4PFtqoMriicO3A/RztNpkEWxdiOdbS6xG2t+l98gR2/rF5zzzQrhrNqo0yM
AIvQdERm2KHx7awjsJGiIVqLYCJ+DTnsk9eeHZdHcrhcv5dUHq3WckKlHdbsVlHE4EzwNcOd23AR
T8kGbLoOCInmGnvhXYEkxc8A93WKIqRI0QS6x6pfgX70o16kP1dwhvL+L1h73k5f0nd0n4F2lyvg
1oQi6MA49uPTgMLw9z1WXSUUQ2WjUtfNeyjN20unFcJxc7A00NT/jCnnGTndXFfKu6EiT8rRpMX0
yoeyDq9thCF1rFE6EDPHS1km45+js1ePHOyUj47znom6/4VpeW6WHcSzL0iavWgROldgm7ulpopN
8IdtoDalu/6zYFxPvek1ie0Un+5TLuktdbXyrqxVWk4IMr8u9NWOSfA99e+UIDDjXh+36/gEzCxL
NxCOW+Q38fT92+GcyEUvNfEW3zkVe9ZvrcRe11fs6Qb6cPZnm/qhVnLCRBCJ9Hu6IxJZTQidRs5E
S3rY8fyHDY33XUePoI5jyUmA8CuAya3/MU9hVqv4JNX2WQdoAQbe2ld8JOntu0EXqOHVMcH7V3dK
eg92K6Kle0MTcVWe50xfE/u1ZLG4iTUmoyscLBnISnm6tpZCQ9iDZNfybcZpE9OHlbnWsMZazLKu
BYns3L8arYbn2oXldVwQeA4BeaDx/XbuiYeNAk2QZ6na8yb8nDmnN6aXZHtQQos0MBRWtWZvWyG5
/yuRZfijkaXvLEUO7WlWDfcnldFjlIyohx4jdaf2Xvv/4NWgi/xnDUlXU+nKveXjL17L+tUdF/Z8
wxV0zpl+mICAHu4jRAee1qNYxk9Nad/as27vdyAKbh1lFCfHkAOdc3eT4Zy3IK6dUB8W1JBX7ZPS
Y9jKqvWeHepp//bF4UpriOHqXM0sH/hm7D6sa4IhkahXAKtsPWZrnvod3/D0fUhniMYFO2LV9OfP
h/1Bjzfm/pqOSgrMzQ6pRWtey6ATAbcSs1nLqKF+aMK4v1rDBewnSvnS1rBjagY6cgLhD+HgQrVO
yAWHZBqfJcH0mcKe7TQNHCgVL5q8fmSptswL66yEyEVINWPq0O2tOz5w8jLdFZhrD23q48V2MGB8
bDgYTqA5nt2jK1LMIS/QQqZsp5yXVksy/lLcHln6TDiG00Lb7OhTtjXvYVzi8rJojga4ta8MHz6Q
jkxy5Gx1dzw0GUWKHlVyUZzQNmnRgs8Jsph2JcdIEBhuk9bFjpCYFuYwEuorUhbmp1Ql/xel7Q3b
QdmWg2lZVA3+CDbJwSPnsQsoNodPfGQizSD2glbI0Rzd//Z12VmeOm8U9FG9qGyPy7ZRHKegikQC
8ZCC84ij7x8bvMtjgRBFzF3VccWirQm1MffGYLy0oq74a2wKx1Q2WWVmtJA9kxCTAEJ1YIdw8e3b
kgG2UmbjzYxJ520RpaznrIoourL9j58qlFZREXtPOC3opIUlxp3Nz1pgwc9lqH8QiY80nxjrP0wL
HYe124GfLqLnFTu14mBW1KHmCvNPgt9WAR5H6C8RLMTkquiKol3XlZwmAw+jsvpBATl8AsTQyxKD
ychGtintxtx7lJOHFtRY6lkcgmU4H0cCveXKExY7tjBa6mWrjZC/IhLHP4bLELpopApQRsjb0kUr
NkMU77slI0ibRZ1eufwppgM3Ky2wV6u57TZ4Son5F1rpRVP/JXA0eSZaIcu9Bg8fR0Fz5afIkLT/
rp0rdOyt6lITMRmDRk+Ykf1Ivs5oJxIekKOIfNsEMqWcq5BDrIyJ+3ir/jZyqo6R4D4qZGiWoapv
qSwhhLQGHgDp7ZtSVdBEgbIBV9VW76oIZvUKggLkzlJZCboSwd2MU0+ZJaSfX2bP+Mk5yCLMc4W4
5n4EmYPLP8gdA4t+he5pH+WIi/vQyDMhcFltBix1kkk2K8BgB88r8triatF4laz4vRrF4oYCu5ko
gxBQVblca8m5xU4QQNaPpJaSeHQA0wsCJGo/RK1vRlOnbk9ybzLW/LKLKWdA5iPNMPryT+PtYwKe
Oss+rfqEC7hSkjWFDrLho5Jr6q4TXJh0qTEYmU66KzXNr/VDILMQgw011SiWjoi+6JcxglgjvSdm
kQLx0nV5d+DaSIUqElHEcLR9MygDw2T6L5vSZGaR9jfZwO51139hhFIDxx7TfQMUxTTi3EDAI45n
IyU0HUPbS6/WEEAcfOa+g2EdwIMQx4KVhNVod1R/QyvhanqST5Owl2JE3vwORKxYgyu2ZOKAuPQV
ucElnU5qLVIRRmjsyAlfUT7jGucIoI6zmk7E7UXPJ/KU2ctB320WBJ9/nyWFPGa+stFvtTLWgdeZ
hGXJ3j6/RCxzjdI2UeBmUd1jLLQ0OX4/NBjkCksEcVwwOtKqqd5vPUs/wJ7kfj5CXw4fF/4iif67
n1P8GyQPMUz2s2t8AedW96DWAFjzjBmkHtdbHfkOpp4ADpUFU7QI4KeM2Y9shxZ4IbKLbTInndom
SUc5qWCfzr5YVK8QGiMp2zgRJsY7Pgzr6OI4Bi4js/djLGKg6I20A+E4J0WLU8bf4S0LusuykFpG
V/XWMfYVxaU+xPJemzaeF7zt6dEIpyvvt4bpkxdHjNC4ya3CeF7lftt7pnM0eFLmn25hhT6SnBBU
E1Xa8rAHqAlrTqj9cXzZ19FJE7tuy89rJIjTgV7ZJ+A2D/EdI0P1P7mJ4+cVmnhMocR5mCYj0XpR
i4rUPUtGLcPqSN6O0wUoD6eGgQr7zc/+WCMawPzVVHg6eagGJ2Td7nrz6zUBn3w977tMG382Ego2
kw3SUlHJlfmy2dpLGt+Ogh4nJH8REdL94Y7/7BIXoGxaKRqYwuzIOwaaCjSzTNyss4xmlWD+rklV
O3+LuBErdc6uOPoKUefCOx5MGDbdTXHR6MMU+Nyj7ow53Qtiew4uTfsC7KNDgeCvaHM3rB/jeOH2
5J/KoIO7GBd00kM4guwasg/cN0B13DKGxU/xF0Sz4xkXRnPkJ7SHEmBF4OXyqLKp2OYDb3tEsMnw
4LPL88Vih0Uz0YPgWgR1vODpEq28kZsTRDgMFhsVN/8tVtkFJXVdo/mIr3HreSyti/4ts8uh8HIr
u5+8Eyj4sX4YbycaomUPXk55Z1ayrUO8BsR2nyDTjykXDJIcWgmv0zqEE/cCfVIs9zZ9moTOGHUR
UEAGbrA7+yqx8gATGipU39aHi5K/YxTR8sLet98bKL9l2Wl7Qvomk9uAxVQnv95wbG1psGZhhPjs
BN20PwzMwmcIZvNZTBMXY7fTnQL3wnED6MtVMdyGFnIQqMClBiphCfLbrM/8lxD28SKgZD/biv7F
c06B7rAgsP8QJddQhVCowTM5SLJ72XS7xnYxzRHuccbnQBNsXZ4RM/RIKSlKRxpLtApT7RtQ4BRA
bFKlvrYTXXm+LF/uahZLrI00A+vKjh8CmSaHKzLSRGry8O/7ZhPJuIP5XPbPVnDlEKjWDGdlxgyi
SBcV1X/XuYxS+59CXICBkW8ba2eJ4vxtnF+pTsEVYorf0pRKT4Okm9e165mwXyiY5BfpqdmKl1Wz
FTxuhiwSZNWpgzdMCi2n1z0K6mQMKwRBJ6OYwDS6y4iinY3ykZv0axTxeKV8mliApDcaHvrCUmXJ
jbSP/0fThIAHyezwj+PDRC01L+0TZMvz1IH/uvSDk+bxp8d3g3DqbFlh9y3cvv6Mb2enlYPYqJIA
cax/LFRrVZquc3Q4z8SjkGy4j93R7Z1F5HpSvOzIg9270c5bXP/6m/9ldR3aZriT7B937gdx11Y4
eTzd7QMn7gFYLtXX+N9TdpthwLay/IA1FaQ7qLEEpqvMgCD5/2AE0ILQzc1lqoYQco8vekmS2xc+
FrPe/3lMB4D99f9ok8qwKuyNKpGkCg0vosDFP+7SztpHaSq7zdTo48Y96ZYBfpixWwOmAq52THJf
HpDCRznE61G/OfRa87A/RpsgzEIA1OM7fvP8ZFIPtJP71yyGhzVNJc5+GgBUP6DOFM84EICm6Sw6
LYJRjWUFslupvZiQ3hVeSQ9NmJDJd0WseH2VnWVf6z33z1u3vKgy00zUUK2BLji8fZFCNZyilEqj
NlYclElSUjRYFZdiGjF9SfDoKrFaQT390cjxnjz7eRRSWq4rodLCXvkEEkobHIINq59lBDNITYe7
amVjJOVlZcAJA2Kj5HQF3CzLhZh6hbPm+FuEGXiVOOP0zML/xw0RE3iL1rDrHIxaHlVCDbETnrq9
0YBmKoFovWc8MAiBGWnX2t6VgNunRVRgl22uRK1r+4YEKJgW7qI4Q3LmBAJqtQ3aAyq+Oz35t+jP
Ui/Xaa368UOknPESNc0TYETvSyI1BZQsDw5J72Ifx2lMZ7p3nNeZKoZIjjinyr31Sr7seeBYCd0G
e9B0XSts57107B5wjBsXuUcaGW58bqaTBnJK+bQtppZzDwudPw5jnafa1spegHk2DJfrOaIscLP2
vJNRUgtRur0Zw5hKWGLfyJXAMREPE/9qbtFEbwja9LMRNv4Hzl8aq3N9tDUoby6aPojR2CloI23m
GyLlRB28n1ttf0oGV2ckhI8MWKNeG2chkdJdiRO/fl+yEpC8dbmEfIq7jaKN0BF293fCxGwsuZPp
PBcTmFHMheRZuthR+Oy8VpKSYtX3enCSYIp1DWrlIO8+wkjmJ1DDxo9J1t+8D9ad7BANb1QltGz9
7lGpDtJ2vnTCcmpwJ2n8rxDGlyoGbiqYSdh6ydiODSlqJebdnzUP+NAQ282j2oeI/cPZ20R/q0UQ
dsFzblQNUqmzGZwdbF6c2zH4LC03eJj3CRxEvx6XBuPq6jiOfi5jgkqI58WYOwRjyWGnzNvpxypU
hF+JfnXxxcVOROTKBtcN5RRcJ1jRJYzqE86/yI1y9azB+efsJyTNyKTl5lhCXAAmdFDiYmiGnY07
TbnklyA4W36nnZJrnK3k6BMjQyfLX5k6jS8yhhknLyht/KkjevQmV/RKtUjSUkEDZkMxH5NMv2fL
eDqahLrA7k2+Y+5bgkj5ROngbMoJZH3/YiYzBbkcaHLcmHycH1ZTIijOiyhVRnBvRWPKF44hkBqB
wHrRStgzdq89LbB9CoHsmHNj1TaZihNBof5pZkAGvtppRP7EMMJ/ZyXh6RwJtUz7cbsv9T2R0lNR
d/ECvmYe1W4+9XBTNy2BFD+T/zAN4D6D7LOe62hhDEm9UD4GpyM36NfVP96IG4U4eaEs8bgjCRin
x8GNoq3MpUH5Amw9S4cA7EQ3LYh6ahuXBvjdgJD2Dy2tk6VRL1UKtEk0O4OGYeLm3RZ6CmvSVn0T
r6PLabmnJT6EhZqll31klDq/bIFJlwOzeeJQ77PvD6Ydn4+GWb0Us9kZhtFGyYXu4k4yIN35CsYO
W/fPqqwAe6eka6HwZpNNGgSfJdy1RTWyd/oXUf2Eu9CtnpdjXK60G6dCam/EFk0Vulboonr1jq1g
/4idwl+ERoGwYOUobW+uyQvIBsd6RihoC0lgycDWLj4WhkgZpjNpBuvBMvLZNTgoT78slmpGcksy
TPR0TJ+mqjUtLanavOT1lFG2yVR8MaVbSfBodICnMxjoZU3V0TL0ePHnuvOhLjBDwzt1FIFvakv5
y1shHnl6fJb3qydl95vNHU1ix3gelB7S8jbV3BWR4JQ0EubAc42JNXxjhFoqSsm1xj7KivwJaMvI
z0sPjgH85t6u7cpMjK9XMWIgEYQnTOewGPooxz4zkXK3iHQulI8sRdlqgI5O4T84KxKph2WzMD/M
2sujDAKGSpW0c0IBWkZvHG9z/xz9H8U0anIuoob8PMquc9w9dsonmoGmZeNUtcDmM3CDakaBAg7d
Mlx5NM1x3KLk4a6xM81dvrNfFeg0fkgb6hugleIFJSQOAVUt9pGg6AFOqyeQszalvUtw0SG7zkFi
H0FBfnAzJU6jD6/B+HmiwicvsVqVGi6hmNSTDGTDIGAAX1F5hA5v/2uv1NoZGYGpOEeWKn6bv9Y9
DQK86xJ55koLL/zESxlOQp/fPDpqNtardKEtl5Yhks2UDGt5SVKGG/pqEe94GCjRkzS8qUiVBm/v
3A3dmjXL6b+3yOLxFdGjjVbgXU/cp9Jp5Go32JWu8DGfGS9g1hcQBbt7v/5qcJWyUtZFTvBiSWdv
U/ibf+aT85f76tcaCfkbbQHXPtEUNTCGTSr6ErPDWv93B5dzG9+6PW1DiCDt/1l3yfI0GDJatFnM
eAi82ByRlBybem//v89n4iL+Aw427vJ3aoKZ9Qyoz4tkqqOT3is67VtHBgbWFLQY5YHmBmg9RpeW
3m7ugGDYtLSLHLs+bcFf6PrFLr/jOdESpCREmfYsL3jPvtkBv0d9A3NtVfaxcWq3jr+ErfB0Hd7r
hPVhbh74vp3ogWkCm8qw4sMboDKb2Kr695d50rUaSQB0wSrVPmcJQLeWlyxbaoOotrkQERCB6LsB
iI+z7K90SHiLkrCOj+TqQTYRTzWQD4kRgxfSa/8UpE3Oei2QkkEGkzfegzTE3FhKmNN51TT6ZJ1Z
s5WnmVqErtDdPa+QGWLEOPCln3ohcLRDh10AhJ39H2aUFUcwkJfxJzHKnMOW5XYxenvFPFJDpNzd
hBx56HSrQOaPepkqm0mT33flhuMCBNEHKXrBkUsYsVcbUCJi2xKlGwY6NuZK+kVJFeQjiRmF2ygi
rStTwAndf7nLNXFk119ZgypDPoG2P8JfZxB03jBkQ5tMtQ3qPEfqaIpIl7Mw3ssJcEcHbvBL4Fv0
WqGcS/3CBQvia2l5fqvem8tHAlf6bBqBhGgqT1fcPje1akv1lmZ0LwsYg2Qh3v4xBnlQ8i26n49A
7IRP7i0uPmbsx9zytcjeoJzvLAJMS3Mv3TZgkXPlgbxJ0fSmESFZ2TWodwRuO6jYl0S3VS19nNeu
Wrujs6WgXLn9p1KqW7/k09JSVrCu9AgCdzNa+m45i+3dmzlkhA82h7FQAVHRYOcwxyhnOpS4ji1G
8+4NaLDlEnBPc++XA6VnYh5vjB4u9O866JQkLBGS6NNqkpZj/ZYtZoHZO/sc9lJqJWMYwb0JX3WS
TiHV3/sN8XgwgUNV8IBIKSoCbrQ07nkPsPsnzKuFBGVehvzQHh6RuNg5JUxKWTHFpYLuPm463/Gc
Z4fdFRB1ZRH6OxgHfqC/YyysbEFD6NdG4AOr9m+tnSQ2L7eL3MLH/B1z0Ua0d9aZ65hebeTka1pD
bn+FOY9bt/ojD7pQ36iGvMFXeaxe1xPekgzQmJPRfOQk0qQjbIJ/o+bBCoLTacDgr7FVmxQpyZ7i
Q+uuqfoW6CpoSVeoJGQgNsWxToDWAxUMnuR966EmKgFxk4MTdr8BZlzLGyyM8Zukc+NnZmtPKgq9
tJ+B7VCYQC9h0ubdfnX1GU3I6LxWteeRh8YCG3am6YVY/KLUuj1t7XXZtO5CCQyP54tQqI0Jx9Jo
c4eqNu3Nu+/FlxPNgzZj1df45sZO56RIvnzRbY5ZefqtMQ/RKaEorSeW2IP85sLAQg7qyrgjfi3V
+/LxBh9CZbJx7WIRe5KteuHjcjymd0DVOQP65m+HYIFc/Mg4DjYZYuIx1ZyBtEWe0eZZqfUP5bEY
aN6ArmrjwUjmZIT+y/7SiNCawNG7+FbZNxsMEf0uueUB4p8vRGdIhtY7EJ7cbbMMkY9nrgfG5pEe
0hf8pkLVZkl/5xyJUq8veh6K1HCZjqoiUWaATzZ8lD861ClWJhObZ919oZfrkPieWHUrz6hCtLk5
VMb9vYdaSc9a8ZZbKxdr39PAxQIR8E4febKl4Ytdq6RQ3RrMrqfdGgAyk5ls1xYcvxANRykKlMrB
1VReZWcgmKabSIY2Mp+m9trsr3SrHbFvAYMUEa9OHznoTbdsQZ4jfHU+e9kiMpoxTLa5JUVaGuFH
KYUaDk7Fp2PaqH/9riOFvDbYF1WROCmgsU2cD+wxfj0O1UTBUOIrKl1WVgELbI2l1iNhhMTV1w8+
wI3fQDglaAovlcCZTJYBNBEJL+j9UXZzG+G5vsr2CfTEX3KgPFuN4XOZim0uoWhucok+twZ5QOHc
Pir122Y7xraABYPq/20aciboLaYsj74z9ua+aC7gz6McCEYLkIldTXRQ+qrVNhpHtZ8fiaUU043o
PbYJBQnNjuLIQ2GqbDSxy9YDcPUJjXtUFptZGafMuupxB6ZSBta/hvlCSm7lpP6xWygDBBmSrJh2
9DIqkzoog/aIwlQi0PvqKNhGDJf+VvxJW80y77QMdswyZzO5xyn2olF+l6uZOUXXCHEhvollG3ca
sYa5n1XVNn5+YDN7QClauDsaMDicw+7O6tepvdyzHyba27MPcEB3Kw3LjV2/faCteVZw7aprrSTI
NG0pn+RlAlpV7qzd2b2mU/Q+e0yYEEboQIf/jmP5HFuEaP37MS9hbkHYNopcLVC2Mar4fYz3YR+L
wpURULwm7IEDn1uxe0TpHagxj3FMppNodOtqzH4NeBcPE2v7mwFympizq+UNaZlfkSLCk/XzjA8/
3B7QweNbpC4tJ6ocW0LFe5tl8dRRgQ2rIYlVBOfW5+iEyA3kkwUqD315lgpqXmLGM+utRQWLtnBu
JFlzkw0UEgEWLDD014rZzpw2WrjWrC1SYTTPCjkia00Z8Ub+8K/3Bt5Fbw+Aqy3+mTb/poKcRvbA
53dwn5tMwA3ISiBWBN4PLiUAMa7H6etzJg3VcYGrDuLhK23yWnT5y4ztFT2mXSGPD0OzBNJvabuq
RPNpkDp56748gtpwV0aHlgocoJl21pw7VXGOD3Wl0RqGM8u/bZxp4dktNAH9EaMILTVsL/rVqZvd
tf/O5nVjgOQnl0xxmG2bcN1qnHCdfgUsuvSzXlYo2sYLFW6/N4JvLtc/wG4shSaHMGG8h0Vs24So
uiiAH5fnYiYp4w+dm/ru26A+NkcSr5HzkexC9+JC4IwccPlLOfameP/7tTKiTY22RIU1MOuh6e1k
aOIEJCi1xuQ23GIGSzf1Fp9uT7j75M8iXWJ79nYro0ggE6tJwxtNO4ObfEaQApfg/P/c4mMzUq6u
LqGEThI3wIIkRis1+VnCrW2FzQp6QliAo/Z/KhgbGQepfik82rkxv8lFCCdIS21H7Z529o/mjepk
04vvfhYCgVmHN2A4CGd5SG19auBXQDqS5H7ApBVcQg+VOli+ye3iiAtOBP2eefc3bKYMPcSKKZo+
ca97j97gWuLhviZ2UjsmlI7Aj+ZnuxhgGgZ4OZbGdYjZhpmR2HwDzfTpkRNEO9kBcNAjBac6yU3p
/i9GcCwE4mmtuUidDtf4zNXUYFZ6I0xb8Jr8uKC8ZMmMFog0WtSVzAfLNAdb/L4hMz4LDLUh4+s9
7R1F4MlhScIPMfRBRvvRCrDHEpW29hcwdYrOmLNP+i7/13GUf6WFFZsmcwLCJegHYUEXBRIvd2lw
9ZMk4Y7xHWwhQS1/7936KIbm5HSUDJ/jA15qys5yrpEJlcPTIM9as0DKYu9QN3Qu1JB8PI5q+tn9
4l1zALFmzCJWOHAq3J0CuXa5IUfAKd1QAdXfRzAzoAlVHF+3bAHDIO2LoLg1zGrPlmdjLnGifMuw
CBITxlMs6KTlaoCeOByL1XepX2WSzQCRVni0A6xAiOigi/5oTnF/lGvwgD8ErIwal27maasHj6Ri
AwCPGGHcLqnXo1tVzEl/bN1OPrk3usPQ+wwKGYmiXCTguwzN7hmOCYyzWshLnxrnrXp67yyrGRnw
MMLl04JaUajqQVvXfwtOexnozd5UoAw5ZbMLCRd4OwAz4qY+GirkwkkuvMr0tA4V+lAoEFnVjphx
h4Raww3RmvgwpcvClp7kKi2luCk8P+GsGDmUEEPuOAxJPBrodgzpLlvf+QPQKb98sKH0mo+a6sz5
vHsUzs1mMD7MWgl01aS1ZfYtqJMdqt2mdBlAEwbKHDZZRg1XUtkpCQLxp022mTNxqdUrKTRbVcD1
EnyaRqqgQcyhJ+F6qdcNFMG1W+QIfYJUu7ikZh54SkcFRgjqUoBYxCVcUPDoYwUwwLrsCgAa+hkA
u/dyGOLevWHI8Y4HDXBS9/jYFdrL8WRvVbtuuffRVWmmQOA0AGJxMNX7H53IlKtRni3YOl9/q/kI
RIRkCD5h9zwb5W7FB0BCj5KcIHV5fxCiaoyD1gBC3zAdcKqJjitbHaNhLIJJ28yLzXienQAa68QW
waNGQ0X16e1bvnTGrtK/dAGNelGjg7egrB+Ph2+jqd+x4Icc3FXwEGvWTqeySbdy95jiTCllyYpz
RctACc3oyWAL3sD8L5+ZUfQ//VAS3z+QhbrSnYSqPxaOZqO4RnuBKg/SBXn6xl2mGbn98cGp5cJB
qr1gGcI+Eh6tVbTW9ZPG9V8VjKHuCctaiYK/+YYlel/2K7rpIAVGqsUOLuaUmWnp90+FSZhfOzE8
VH/+7Iu81prgl+cERqMUw5zYz21R4tLxbTTfrZbRy7tBU5ahUY1agNVVi/xR8WpgZvNWI1b4H7ds
0qZROb60Uk9c66LtHxMtGFlxP0aK3sUTNx0haJhK7lz2L+Ltm+yokjT4Eoy/xfl6jvgz0GSZI8uY
khI8YKGAW5+VKqprVCMEeMBLKg3BU5YqhfPjtKy9IX4mn+fWXSb334x/BnahMtzIvR/Hs24+mKbT
qInvzc9qqZHS6uwCwR+yZsQdottsoGgqu25GJ+pGsWqmhconrU3USVT7f4QlIUBRjBSv2z1JGc8m
GLgGlRqjR6admdwkSGa4eKtTsTI2lZ8nhQgPOj1nOryDhMiqqo6BVocvAh+KxFEznFU69RyltELW
L8Nd7xXwWlRjxOUWylil8p2yWP28YyxPAktAPvd3DtUdvdNBUjKnmU1EHB9bT2Gi5izA/6O0l56O
6Ioo2jmMJQ/bgM/5OAsjqLb9UcUILwVKTufNb1FQf5v/gPNjAGBzk7RtojP6fXBkd55pnjjWV/JW
wyailLQVYK49dPzTJK2hOU/WqtmBVohwlGKUxWFvfXFQAmerITBEINDKK7tiCIL2ujZ42jLd0ey0
beQelZKfL6RERJaBehVd051KdT+HKotbnJ7zWFWfEDaaWnRkqYhgLgxuq+lsfeBBEhklM/7SNW7f
tmU1o3eMGk1dLJ0XmjQ46mwZKN1U2E5XDfQyYjJQxJlMyGDVrJzBOj3277p6S8lnLute9K8Ufe14
DidOj3zfLbWuwVFe9K9dDB3v3kXs+LIStNJGUtUiGYrPsRZA7QcL7CHTSNVOGwXqsQp4V4S8VHaP
J7+YIqkCuuhi9qimWeUzrMnARCnYLDdcjOG0kRTMBUJdAD9H3KmpxfTesftFtLZFXwB+/1UdRYBE
8Pg8s6+Z2+YyUsSwXKtH8KZX1q9Jcw7pw0kZwGZXhN28qXSfSGCwTW37tmhBUUYmsMONQxaHQotW
yWgbqq/gsxFwfX1bukM3RbVc+SLo/ebkDpKQrAWWlPNvl5FrSrEW2Qaw40Vez5/bgOBf/sL0Q0H3
tmUOayljG7rkQsBaNB67jdswx9fpfTEsWx8/7a6MGiKbrWjyA2hE7gsV3NzEWrse4Ak53lg5UbRO
wZF2CMuPeYEGZvbDulLdTG1CF1y21VNzw7feJZtAndYodEMWdMZnCxaFSBxxi9G/u2AwT87P9GzH
RhlPgqCkHT1L63gLhlUoFF8Vo21Y9iu53qEr/mgb3pwMyXpGJMSq/ha5lhmtlivCObUcpJtyqSeq
2uENmvIJkxv+vD4QwAJbqh6uYwjLGHKGsMA/h0vKBoJhh4o6aTvV2R29CjV3Xsv+HvKDxMVB+/8j
zU928UOADuLMrYmYR+K15uw5KlFKW+40ok5c7Ts9tdU0oB3iRh3IGChuiPW684eHjoMhMlCg0enX
OqhMacjZfYtJ51Cm0cIA76uSNyIkGKhcSGwt/JTQD7Q+yMwwGHCfiAwSYIassSz7WrKUB3S8XEsk
kGnb9UIuHhYzqmxW4KRc0f52HitOSvl7Zh11wQ2vtr09jnLfE3I9bmCtFki1O0T5KM/PRwTfRD0x
sMO1j41fyzZBO+/JcX8UJwqawYQlbdBHYSAMHlRqgavmpt40f5vtOoL63TY3fzKqg8Mu2crcZkJ4
sqfxXfduDVQHXqN6g4eLnBglBnx6PZX9ASPkS0TsogtHdG2icB0QOUp55EwO/cq35QRU4d4NUJ+i
1JKtiBc9DZXqkzupfPD6TbYD4z6R6Rf3klyeWhK4gqS0HA7FKWar74zlcCbcvGIzo3FlMeKpxut8
JcxYSinIwYfy3g8+TlDYg+sXhQPdxWjufc1uh0qNgvWbsU4xc4nhGms0NgZ3DBA93WTx9XMEO/to
4+ORdAumCUPdimYEYIcbI4RiwEf+ViSGqZslKIMKX9mu3Rd0g+t22nMUjel7RB4rZb7oPS9TW69J
0QiewDlAFRcSBrWDSL9N1u7FwBK3CqWzZpZ5O2eDINdXsDtFJFWR62qoiuo1VadWDOZY0vEHDIjB
SsG6GH9Oy9l+wEAnjpNPhD56Ci8HQHBZQTQSFpU3RhrpZ0bAJ5Blnt0X8/Uxhuq0UlxZZWOdcFts
uplnjoYRawXyUU/obw7brQoroQcrgqNwnHeVFdDKYdDOkbNl7TldXnaS4vHQjv6BI7qSeVKB4X15
U9hjVYQ6lhwUGx8nV3slJLpWdNAXroGtCErqSNS2g+SxBAZfyD0gaMEkoZBEbrZqFXQauf+S/5RT
Jh30yWoIqWUEtOBknDlqmGf3HmeG7DqYIN/co8EtspsrzRc50yMqcgeapsQfbnu6dwctajuTZI49
lLCc3JUZV239nv/vhqjTSEz30UJ/hXqPDjN5ACJWT75P4UZd/nkxfuIkE/Vsv13X43qZpaV+2XZ8
eRrP/F/cN64wHsfGFXlgypDT0s6Qs+JPyHzn3y8kBXFK8ztEzIgKsxGQdeNTQDJPfX2y4XIAFMoK
7A70njGIPFVIrZ39Mpss0RbEXL9pD7uXSkKYMbKgiBS/wAURcG1/EAOfVdYWu+VfRT+bW6I6ZeFT
wQYftq3HMdSEWtxFClfohqvohSqPQtq5SMCv/Mv6jwocwRX0Xbiy+pev+A8wjFKrGGM3wNgBMiEd
STkMufy4iReUm0VJbZyBOD79ae0aabqdOXSAuISznOApMS/LPFF7Aq9Q9MlJF9T1V1lU2X6zCghS
1602Guj1zW1EyrMd3xmrWGZF0fO/fy9Wgqb5rsw7IbY3oPVNjg9M+BGjKS8XF31P47jhqUa4asT9
3kapy6W922cULfyVPzmsCypBA0UXYk34OAufbkAD8ZvE8pDkS6yGY/OFf3dDLEZI6NzoT+XGlehB
pNGUiyhyu7JiG3Gwp2YMFpGFRhBHbl4UHui0BlUq8g+eWHT6VTwnBSthO/FBDWYxqXVb8OQxkSp3
diEp9URbx82MrpvzkvEI2QbjDi8MUy7f4Z/jPr5bL7WZ86vK2iGHEmpN1LciFvKvYjJTD9/B4wNx
y+Fkfm4/z+YZCCrpALE7XEJyabZz9JoVki19gOyXQAWNyUDFq2AIijyyhuD+cSx3Kvx2oSxVbTv3
VUdclgiKa65T4Rb5mbs2W4q8q302vWbDe9VSl9pmTWdtjjWARWpZk+hhUrWK4NWewBGq4Rxra+42
Hf0GWPhWnBFpLK7kEEoTVHMypR1wVYVWVIf91zPa1Zbw/tKxsn4UewncB4tQg6JN5gghGgAgYn3c
Ce0Q9vbyn2C6kBMgWfJk7C1e08+2M5uGmy64EJFtBuKwho49gxSW8CtQxWD2NFYhyCwrfhchyppB
MFTb5IFXsI1ZANf/8emJ845cL4QY8oSplpZnUe2/+4Y2+sGaIFpyRpEaefL6igQ1IVrahtlHxOLj
FzJZlGy8jF+CNj3crc+Qwomzk4WgfbrOdhvGrUejchI9YX1Vt15boJBJykY6EXIPHoZhOhCZLcGr
DakO4+PQB/g5C7VAK0lkK6EiUTJpXfptvew40UUHRmAENNCjPwC83qxtKmOwFNUfsxmQ72W9UVkN
DJ/oMsZ/Ks4+fqa9a30Iq1nhAOwOJXS29xElVUdbyX2BSBwl3sk6LooUuCiD3vPeSmwGgnRJcVEd
P/JVuuDHF/dvRcPkNuwMN6VUjV0LQQ4SIaO7rWe6YxoMmzFAd7CtOqWhel/lfdJlHl1GNVJQKw5G
KUtJpBNQhS3lvIlqsSHX0mX5G4icWJIOBZWrE4+nR+8lzJv7W+cNzm6arv6l+PPcPhpRJ9cLDS8c
gxb5jVOF3irNINNHrzmRBdWpwGCOi4Mk1y9mTeSucFtr/Q184VApvqAneM5CD9ztI+Gn7VCIpkNm
f17muX/yHLxVXo2gZ5Ed49hIA1ycLMWaQ0IT91eu2XXraOo72/5ECHsWZOw9KyOHbCu3ryjpgZxQ
W2/4TT+vsKZTQ8otr1kIsNqawwai2GnAXXEiwnWq9szO5B+wsDVTQOqXECyLu5fLlkmwPLWWZsve
KvhaGqB9vjw1hA8uhL7D8+4HGpXK1htNxEdxdb3n4vnck33fXhVF3aK2WdM5P+Rb7B5Hm095Fmin
iXQOfwd7UqYRjcfaf1JQKWawkUyjedOzr9lZlHkRJW+REtuLuyPzmh61UUyE8kEBfAWO5HqfsmUW
AqvFolrU2dH/wRaPhCK4K921X5icJ7qKlPA6Ue79IXnLF5fjVqQ5L3YeUwWHFepO57ipF72CIomK
vvfB/Y81PdPQrOCb7I5gVK5D9cHGuEgkN6WFzKXfEDs3Mlr0079FQoxfLBxqwdoXhM3WdOTLTWFT
yOk4d5bdWkQHkjxfRrJZWskzXqsuHdg/JXOn3RFCplU7dkAZ16XiUpAFCCFoEUxUmqg/++eR8BCT
/2Itbv31n5uGiyMuWBdBjC6v7M27/aNzxrPzOidPgHihgziufTB56yYRubJbeQGn2TI5aivw4Sk0
MieKcDXPqZ4Dl3gPrReKrMUVYO/Sr7jmUIFRP+DJwLWxXhe2xMJLvEm7u9QTnN6LZWXBmQQPDpeY
jkQ3MTgM8QgxEUBhb6J4bGQWdIOzcRFkYqovWamzD2zvIYtp6qSb+sk1IdGjHMq+aQPxtZbuA1qq
YbR8lKWhWy6VWT07imzrR+ImaNHT9MJSaUjLwuYszXXWYt14vjtxGKnX2oFWjiLV+bR7lJjMBYew
3qhMPBnrSIshoLdEPigg9eKOUv2OvF//rQ1LbwYD47DqWUpts17LfYe7F5kqUwaU39I2YQ2daJ19
AYAll3dj56z/aWL1bFsm2ywRx9dmxtJ+LAwkUlbgPY40dp98GsS/qtxJ68poO2fA/57EhnlXUqO1
tRF77SoG7dDdSyhawxrI/QprN8QxOdBZqJsdZAbTuJ2lS9Ej7mEw2ZCA3hjzcUZPEzfu6K0Mf7ip
sk+jJENzo6TvDzPZI4hVZlkRRv5E+tw8wudRP+qTb7DnsQc+nQkEgAUFFQjKhhQD1GU4c9fUZfzu
jcjPKFD4coZ6h2g+RHvSzzlooD91j8Oc+Ky3Es7GCprhQ27w1xlrWtOnq7Hqes73RgcfWmvzZDgd
cCmgw3qghzqGNx1anYx55qeg2S+reV4P6YZSpw0pHAX4rIDe1cv1PUWjofm6dhHPP/YfIdM3c/pH
YXxuhBFky9Fm8cj+OqTopI3krcs2i2Q8LeSug5QTmCMLBAWRaKWhAmAV+pbBBFtWo8zyqbVwtc78
zLkHVMOGWf/liugskXpP9tzSWPJPagcm4lY7cRxTW7z65YlmzXgR+HKSKKE0ULpSULdnnhc9iis2
4QWiIGAMhL+ZQ94Bz8YoJ3t5I3Xr4p1uvSZUo1C9WkcORxR2S14YMyHT9las0bolaPFkHpcoUN93
Rezs+d9ERDzMpJXQQW7D4YY+V7h4kbbw4OVlqeeAD9zkFWdM8LS1GTVqp7ZUTquUE9gn4G155cQk
1DZgfzN7AdfvygxpqrIOkjO5GXPUdDs4JxEYqHPIlarVL+IOTZoJLNlBpnsBWNQSqRcKQknZdJYo
SOttE5DKKCD3ig/de+3n0GDwC+5kDwkCmOH3t6FagD2Fqi9ziTJjdf/3Or20OEyIws465kaubE08
9kvNfpBDhRqbolt8Sum52HHxYk7A04Xw68WOnYmE8YKgejhtN+bcO7o963syNnt600Jhf7YsMbgs
/4y2rUs5PZJMWfH+ME81PdGE+4QtrojFdckFatT6p19wpYPcUdIRrCEZqcjpufRsqbMd6Z1WFdGZ
ZeiFRCz1zWz2ktiEj/irhX0CiYE6ZHddueGMiyW/h7yasD0RGX0Nv0iVzSzEDcKgXy9cVfrEM60f
DTh3+KBXmhUugRSSrvGPzvvRghkMBv2Ql8rZig/d5DAGEre9tVEMOugycrU0VlFDekH0qHhLkTka
AdQrp0xS3B5pCBTArDKLLqnF69YqJbfERqP3oGzU+Gu9ZJEFm6v8uoEPfvkYeAQTiIZtyAqf7xOT
3qjHJRXxN8z6UFJkc3yoy8+CVBsWD8vwnZ5/c3ez6VY0vPKIww/Yu65dTdtYxPd6x2UkHUEaWYlE
P2/uGL13yrtDpq1ZgKGqgtGOuVga5Mxe/cdMg0FqzzDEuP+AwXwqV+7H9zNhIcJrlMiGLbiPDV7L
dvxhG87Imo0GCBhe0Hkhm83hAyN9NWhiZugNT3pzIwgQAGejM1qVx/YW+O5i2cYG1KPWn33f6YcY
O5EN3+q0LgmcKVDjMspp8/cjghU104n/4xekBppcUIBUzK0tp/IF8wXhuBdIUU8daN5rX/16kcug
9Abfq8vCeS5aF8SCrAuZAljOYi4Ap/9y4F7A/au6c//yRXGRCmSUvUXaezE+4Yc38LnLjQQ4mbwx
6SZLTdybdM6a2WKRXju5Nwwz/bqLNbCErgi8pjclvJoYV17+IetWeswapwmj1ozmCuORYf1DhkYZ
jTe3YMlHzdhAj9fzPVhyceu0iHSThMU/CwuQBEv7F82u0xOSUfxPgY3dpddVgmR//5Ifztx1BT0S
xNTKl9HotUEipsCI4AwELuNZPy6uhWInSQE0V+ZkSrQACZij7gLPIEK5yLgOBum027yctMQeRhaJ
8Z96JXNSgRTeJkbY9TlGgKlSjaHtjpIZo11OqqxIu+5PFQU9OpbLY4KwaoXWLPYRWGLT0zbEGkQ5
McUsGQPmUnYjVX4LTZTCEqR93XAwi4yeKBasixZJbr01MSpM6oJRBAfH+wWUxBTQ2XAkCduoU7u6
+hQnThwE6hLJM8d26Zx2aBo5DixF4KFpS214P2FzHKvxKTw1RaAZpxGOxAMg3ofG/jAILlI93ese
1gr5zVXC3VxcK+CvGeC0fK2PwBDklCeIgMr6dfhtH9eyrYgtHfD0GjDEzemIb9G6LU8NwSdh536c
am+lE0WBAC9iFFlmKauOATJH7nYtB75aTYzkV8PW0KOKyzhcfttKmdxNeoUCLd3Fxcv/CtRgWRs2
W104VQf3FY8vcn4hLkbokMuddQtIER2ymXb+E3qGL6+JNwDGmNDjFr/7qR9Mg2F7HlpbXsaAEwBl
RlIMd8gS2DWxJhzn+mFsPmlIsaG7+i1lYPopuciVnw+Jzy8PsrIUQ/RBFGFX5VVsL4qkIKqu5iKD
CTKGG04sRyFl+xUXKQPRovQnW2KweGFKjGHpPBeTnnJjCVPpFiqm6rWfGxapdD7XvZkRgb+JHysA
ysbKGA8Alo+zMoUYVpM4MuwYZUeYJHw1GxlNOVVXfUava20dgz/8aqCENE6SqUCYQsdN4Z8QZpPt
lF1MTsA0a7P/aSK90m0T3nV6RkNnTxuuZhk2LmRWZzfGqtX7cUqyNkSDH+Yzf0tdYg53aZiQLJwe
P+i5BG3Pb+Ltv4hpIb3UjckceWr+zDQ5be0d9JsTM3tCqqbadcJAteG3WBWrWvLYDXg3Hd+0hKYN
lMCRwegEq5AWGNVTIzEmGgD5qz7KZmuvfJbo+vmRH9Z+gTwy7aIiO66/IB4wTJMtjI/qnOyzaeDW
cJGTLVhRI0CGzEUdsHoGD0vfxlZKr/HFZFB7T733Pgpl1GZv4/W/z1z0B6F+GnMybHUhJbaay577
RCA31rmolijCM8oWoTGmPnqmgL+S++W6R7mlPtHdJTAUsORaDorv0+sb8vL4f8EYQyMe6JE+eF3H
Mwlmw9iw+KMrOnGsLDZRw2nqhAt0oZexw1nU/ofyAYMG0057b+/6smN4bh9otREgZWzBCOqIRxHL
C0jazrz1RK02MMPM1ktfQhMVt76IarZvscLOiCLfAmvT2ucvrc/qJS87uZpnvf4zozE8FZTRJtEz
xrq2rO10gKsLsiho1FntteAB+sYsJbGnAAuAf6cECrVQp/VYRgvEqR9Sd53zh63gEJHUGimQO2XN
HUHU3UmSHSWvK4QtigmNfFfbWRU3BukLR4kdM3GtQgvmK3o1t6g2METoyieb4m/cH0vD1MAIIX7X
DuvZgBFVolZCXyLIZzJeZ6kI2L82sIFhp7/KHv4z/X2tm/n4ogJrcZtOnp51UveTH36q0+Q+ZK/f
xt9YVE6oZXKCtOHaFMSVk/nzVlOf4jrv8Gn/bWOc7iTAH/aTIfRwgNGYb8jiGtwyGZrATJcIOltI
T1BdNyUmZsNmMZVRT+QaXsuqru3FOyd6ap9GObBLU9LpGpqq8ExDkpJTqfuyygpjd/5XmXNqKvgf
wieK39meZgQZ4T0DBrnyGz8vOeKsPveYhoHqTxVf3cdFPFOV9bvRqiW35ui1Y0EcicIRKCrRafL7
AfbmvcF0B1YdYG2fPslOl0p8/AHTSFW1u9JIxu47hoO6gbnkOk3mu4LVdUn3d0u+Z8Alqi/7gC2T
9QgxXNjmpA9NlB4CZTLNSmAtmzIe1mL2RFMb1c0MU2BpSmpdDcwFFn/RbgVwwi6cNhieAipWx+J5
bU5m2IiGbzxdSv2whBDfdj1FswQ3IbCrrj3huC0woCLndDVDsVbGnddrwx9XkRfB/oPDBOjKVzGw
MKqOChIr9SXAMHxWB6ggpZ8a6h5JPADWufA/SbafNHLbf6/x04mCPcYTHH8pITl/jz9ihHNZukon
olBK/HmUWjyzNcQUNTBzbvhR0YGk6CDTuGB6rwuiKA5VkMJdPH7pWH8P500Iw7JKjFWlAJaKdj8h
bYzA9WybMp0sEFHSNMFsvdG92FJ4z3slPpDOaepE1Mu9QHmLUiN9HYNl8lHwUXb3baUNHE6nFWWu
mUa0qNIZXezhLjglicH4rR73MqftULeuFOKntxIuXwKia1PYXsq8L1QwIlg353Mlnwn98iZs6QeR
f4rowOg+g4sWuAf2m/XaDZV56+cYATJX0m86Pt0k0pDyFrszVqtWKFdweWMOLyvBf8sTz7FJQR5H
3XUT/vAaUAQzbd06SVyvwKmuGhmR49FnwTdirB4ooPv5oCqZCAUqczP4NAivq9pODJofkw1YEdxW
lZ6KJ/gC4nXPQ3ywg11sMJJH/hjN6sBddJ9T8Fw3FXWz7d6MbmLK45W5aziVTdOgeMRHK0Y3bPI+
oF24FWLY6S4eOp2a+OFRf5rhyBYSYaY+40Phbap6Oi+qTHOdzfrRfpaO2peCTCKEfRfZBlnqiyzm
OgeErrY1kbZKFv8sX9DZphFIZzYK3xTWbTkFaHVtmmKbpXHZsqm1Ep+MZQuE0aNQYbZcaGpfyoeY
qwE1szvUR7+eybNRwsjJqdtGLzGCBcmA35EeLqMWu6fjj/aIismaOTRQ7Vb66MiNNAGcAapQjbV/
CiRMZFC3g5XkhPVcEieO8FHUhQSdsD6Dw1O2V6Sps2MAgdW8cG2vgdCNhC5Pksu18oW3F6AsCDzO
CFyorDwn/Wp9cR/J059io4n56MVk6U16z2RXjIDhhW4kPIKZhbF4KeQd8PToju30926KIaI8VZf+
AwFvRy0ofKigeU4jtJFeH2lbENmjmRQPluwlw9+yrthbPOM/kadu2xPMFpsfflPte7QgzoGOvtCi
rZbin3yszhs5Ny4R1mwolZnnW8B2msvU1Ukj8dqfDV6SZuR4/nK9MOw+RYuv1iOG8yYf60T+dILL
+y73RVUMGVQqY+bTNXG5g7rnb5ttbVVfFgynV7mYbKkSrOhE+8R1uPEBtgzkmRTclzHqTyhw33nE
aOedtKOQk7kKSxMuaTuS2MPIEOX7nQzRKzD5QDykFcoZmwianYEq80hNVe1H2XoMa0JQOefSoWH3
LIIiACOwCm9nkHlKIhWqtFF6j436Hxdtf4hNeJW/iZ2O9URSZH0i/LW4wKNvXlWuTZb3zhvpApYa
CteN+qK9dhWkQguB/FJp/e3LvGrWZE3q/Uqr20NxB1sq88TH67fRDXpozFc5qqId9wVc990Ydobg
j6UXJSTZbaERxioFOhpq7EG2Pnvcgihq+6jEwRqqun1htR7a1hywgquFCtM3YOyHnguTLte335Hd
h73PdM7OIT04ZJ1uZXJpF9yDyJsx+2yp9Ky04I7o78/U1kXnzBHS/sFV0DiTsJo75VcASUVEc0Oo
U19vW8j+HkCE2k31NLpP25ho/M9ZHiPS7beNrvhzhTZtnlD/yFpXbM5ulo8x2CI2Eh9ny38VehEV
9YSZSGAosPMGsSI1Faa1IC4dBBKnUoc9Fe0W7ZEwvjGIBANXqtDULoapY/SyT3TCZeuTdxdEpQXc
vZeI0YhYxgjWuNm7Nt9FdRW8dmBGBXi6aXEJMra31odh1pZ78hyrV5hh5U2z/+OcDW15ymBCFDrQ
3e6XJWhpPgvAPbO7Tk7K7len1cxaaE/3lPYifgqs51rF/XwCziFAnSUO8iewhiv4GibcSrDhmJtO
Yme83hfOz199h/Dfe9QTcrj1yOcbFsk5J+HMg72NwNTd2f1U8p2SgI5QR26gCkXKVEKx1q0R9zlv
fIhnkLqIRO/Z7RWnPJqEEIxuFZsSUorbUxg/1xFO85PLNyMjnoWFqgOwLMjY8U/ZMDZZt31W+NQt
r9oMkUcrPUE+polphiKTaBvojj+LquOEgqr/yM4RfdNNJmiKAq3UX1m8wrYg9n6LWkSjRrbyDcYG
LiP1lTmHsMNdWtvjyzUo2IkjgPYANzHBkxXT/mI8R5oUh1b9LUHekoGMebZlBTnNOcqwHWI0Nx5v
BEKBRwUnFqlVA4ZyuCzqsHgAfaoaQz13ImPT2JUp672vxiAanY6FmiHzaWzzt4+BgvIieIpNJ2dk
jSOwfxVV8ZfQG7o2U/eXuUisSGxRHdoEB89pPtAMcg8H6cm67XTDsMagq0prY5KWwl6xJeLlIto4
PzaRtkxK1/p1pd5gOlxATwc+foSUwNy6x/LF99D2P0S75c8WR83b2XkPAEiybonE3KuXcklOhnIH
ahzuGPPyHbGlizIoXhp+uP1xRagKNFnLgth2T+Dgg81IRThba1QjIQGRjs59PUUkSyWuS/8SfufM
A8zP9cmk5DCtrjhJL/EgMLEK0pyCt8zEe6Zu9P78QVo3dU4ZfncDRbsfG/W07pSptzftOJc4ZcQM
f3HIzvvN4Mofj8kB93GpU0dJngjvytC6E3AqA+RbtF2umSKy4x7j8vgVxWQEeXDehe7o4uPFKg60
e9fI5WzW4nqKzYCSRzfJQEzOa+GtLKqX4ZdlwDDQ6fN+Ys1HMHc2ebh4XFAvyvWZDzdrSw0WCElc
nuso3UED/lSqh1ySQC3Us75ruq06fMBfENoIDqOQ7Lz3U+136k0+MTG20ScooCPV+nMYJ4GruRj4
ds136A58tzArh8JSvTd7Mc2kORFjSukLtvgTb6GYQRdQ7WiiKAWdz/RBtEocDhkjPDIvubTgl3tm
AmABNApbTcYwgnLJYggvgBFkMmKuXUaeBdwjNT+SX2MKAjtDcCdm8sxyYONXpFGFsmecDFD+emeT
Wgc7b/UH6YF81QE9gtrUFKvJKQdt8oF+ZBQQYOPXFLuPZmlTGwUev+eyeViMPBsLdX5A4K/4zuzr
lm8zpvtdKuhqRQKlmUUlNqfcp/Yt1zd2OtWUK/mV/TC+YR4Kqq0tUZD5vdXUatvgivw0/wXSz/pl
f+ivkxjPk8oa50BWdgUrBkh2Lx3Zxca4b84XgzkuHk6PaDjiDBb8WtSckd+J8u8Pn9KayXnYAee0
1adt0j5m43TAFMeRIMD2M88FmznpU6Psqu70VkrdiXGO5l2ri/x7blWCqyo2izLLSwdALjU9K1+T
B3Ulri1Q5UyCiXZPYugwqqre/+KeWGvtXUyD/Oj3mouNIHUs7L3uGjw/VDpORIMTqnNhX+fbYhwZ
goBuq0LOcEHqJlpWVLf2SYFKB9KZIz5lZkm5GQEYt0sNTyUxqNwLAL9e3sfNhh2h/SeJB7a4YQU/
ykv6RtnF2jKha5kV+21/Sgg03pQDjaJXNaXitAh4ktjimA+DNki4uSIgAPgZrCfds26to7O5ZU/H
3aJwVweR3AL8zfdZIOQErMTM2m+RdMI45ggFzFRZOrdyEeQjgNG+93qEsq09+4X6+MzeiJyvMzN+
3CM5VXlS5ep8KMvnXGdxuF8soevGDRWFZmlkusj2Nki571rnc1yip9ao1z3cK+5B69NTIWR+soIJ
06kmoA+p+vExk17OVIQh6HfvaxeCGkf/v9fXWmD2/omA/ecEK3aPAPXARl1gcT713Dao9BvNxKqg
bqtSOd6ODSnGivLFACqs1agd0jcmgOFhZEI69L7pR5udZu9NJDYx03+8tJ1OWpcOtc2FjiFtJo+n
eFVNfyhO8fgRmH3KM5ejASTowCJdW2waOM84qQDf2HOFeH/TXzjdSP2L7C0i5INQP8PmYMLicx6v
pzHSXv9N06xVwa0LiVDGfo8WRUcz0i8d8jNHwr1sewmeF1Ou7HUzj/hi20ZgMPIwCU1ywT3pDpVA
bMDumoq2bugfP/QOtafNvTEgiJHH8QFEwS3HwJqEsDtTEtUBsSiUaJ8BOnFGn5c/o/4hC+Z3U9Xa
puGgytBi68xy4qGtJLN2yXajAzQL0IekzWXhx8YW4GjNY5oRaQHZYVhpp28YNX/cvNPJfSQ3iZ22
xPAPjY3zAx4WdrJPz045CoJFPmx9sRxwa83fXm7NRI925t4597j1oDxSKc4Gl5vC2JOrhJW6+Qdb
U+drU8M/a5HHAMrdD0nUd04AD9SaJlndXtHdapiL/jspX7m+3ZqfJLXCf1qJKtzH5IzJXSy/beUj
wZ/bh8GtYkZs5RfVk7EHWpC+gTOxJXuU3ldC1is2a82koHD0rp+ig1HKJtAVbIkn0YrVWoDEIgYK
DV3sqEjx/xVOcwFvb2R+wLiMwo9DolLLwDRRVow+J51gXQHbIXJA9tj3IutBmZb+nEc3dTiCiWtr
AC7qZd6t7LWe4EOgoaYGikCeqrIPFtmuHVXq/5W1Wq0/oog6NaYZb3+408Fo5q4YU9b/qbV2b2ZL
pavwwpuso0OpoAN7wLSroDFkjXZmI+CR2kfVw62apVMiBBpI3nM9Wwkc65vZWfKuSXTjTi3+JsYy
RuNYE/R0b4nNXMyY/Bnjk9TGofXHBX1pKPUKgmSeTSU2PDSFuYc3PRfX/sGQ5JtuAJx82AbBsijh
Iz99SNxlmc7C6S4gIvyV4TTMQekLUO+1RAoJLNOguCB4K4f6IC5GcVIl0oUNT0XOWfAOGCEDO5JA
7ZoSYR2xJI4A2bhGUVj1+SBxVDRDJFKJzinmTC1o5xDrMAj8b0HODh/EMp9dwf1UWZY1nyHHBAXo
hpeRFf8e15fRrheT+TKxtHAh3zJX5gvPURIuVMoGiEKiiOGdx14t4dxJbmvMntoFr+mmkHvhGwM2
r4qydAyvjkaIEUVSHe2rq5VIIRjFnTguR5FeFsjG5z+OeZgvoFP1tfTvh49QYJJaYQfURQpMVUbv
F/+d81iQcyXv2V8gS6zGaH0UIQH83+doorbLWKyQNx3nrKNtQT094ELINb68OXzPgzRwXG58jPJY
57dM8vS/BXFSgQ2OATfmSZwH/On3qCrq+k2N6e+BVgExqlPDnM9CCqVfgK3bstZPI57+lK3C7MTT
5q5nJXfZ6Z/S+EK6LTeI7spgelRnUPttvrCz0PoLVNeYy3Z3FMy8inh+N+qmSw90N3SpTkFwEJLy
AaewDOMzVh5UgyDxFrWQjbHP7URrv8LwlFiTBA9PsgWqP4Vgv9t0VJtDO3WojMvdRMYB72+s0UpW
l3mz1k7ElidD9Ec4De3ngml1/wJ6MSSje0NbpVfgkQANH9mc4RKUdkXt4/aG+O/MgkFSptvyANXj
m8KkdwHdkcVsO74z7y9vO5MnW4OA+fg1HkEn+PqySnFPPbfG4y8G3VQISH0AMhaLpUjaldY6o3Jg
iTG/0GfYMu7cYDyqh4mBTOiwyjQXrfj7GXzhE19zXPWgd0fZr10FJG2QZ1lFVkYRt+AKVNIVE7e2
imbG1Sv8vX/MJZLGXqlG7r8e1vuGgwdsOyQ53c/VQuOJx6xwwVHqx3Kl6dgcYUCzPhVXkDXADfBM
XwI2l+Twd+94bewXc2I0Ji4rW7QPkwu5pds9DkpF1b1EhsR8PkNHxAqwq06Kf7X/8Prso9B0DioO
8+J/EpL22W56E0NJmg1seWyr4PKa4578LXUitUrH7zsc6wgvlR3T80Yo8B/ua605S1z8FSR07bl5
o7dOdiymm+/2HToPQ4ohv7winF9EeniFUEBPUMcgLMN616R1lvgJ/ZZyCEgWv9cmz2HsIFlxOprg
LMepi/M8vnQJZKeEVDIdlUaFIGjRc24rEfuUTVklQTAVJkacHkW5CAtJxqMg/wzHuP6iW+Vpo1lt
JwwdVxMz0TQ8aeD7ebFIO0n7ru/o3SvLrzoh9FDF16JrrtagUJOIg6bm+Wvm+gLcHNs8NSz4tCmh
yExACkUXONoDQpG2dApsg+DJsjpVZHK52PpkK/kTYj9p8h5aJq+yS7M1doAtepeko1DJiAbIwxKQ
4tS+cge4hxcdN1QQj6QrNZb+Jm1haSbXNvFvsOlln8EoMuBKdTIvLqZO3tfwzop3QXLivhYgIsSr
wJivXUgi7OYzk5fTr+0+prvhwiRL3VtY1QvrKsi87NKxIyuepK8Q93sE3cdv8htYuBv6Y/p8bAsn
oNi6NI1+1kmq+e1sq/clQ3PwJk9tV8jTC4Ttumt8Dky1SLoD74APZC7aOSrUi5LkMLSuEaneI3Hw
SLZ/UCM31AEYV1BxhlsVSZxOMIsUy8tXHDWMVr6pXRIF3tuE6eMjcEhDfVdW3so7QIy8V4S6AgBI
V3tdp7APdZyHVN1oLO4PZTt5DbOnDgsak8QCFeBxVXvk91WgE2xuWgaCcg1MlFTLs1tMkaBdOQRS
fBkdoa4HCkazGYf9DAYxADj8JvVimuCz7NDZztjO2UFGMmpIp71E4kz1i7K22dN6g4lZLYLf0DKD
kdOjXwAO05aY32kzzS9mq93wH6nvenSdBlbhnGxs9iVwyMHu2v7feTYEe6Rvuah+H9fuuszMw/Jt
IRKfYQKm0hPvoQmZYD3rBNpZJ2Q/tv+GgILHTJXQl+sf7pFTWcC6KejgPk2UWTVTt8paQvoo+q+Q
c8E7isKy4d+m53LtGXTZX7nl2adlBZgSbMeUWnTZitSlAboEQ3sHhCGHmT+1EEGbVEVoGLHvRBJ+
fMIBub7KSIGG2ggNUo9yyvQ3m+IR/jOXH/QLyeFU6wKg/0FOD/fT3WizO/6a2UVT7+K+U2qECvhn
SlMWVqIwac7dF1oKxaH/XgESPMSb/Ze33L1GCRgEhUr3EXBdHu6+nziHypADDMxf96hnwjuIbW7j
O+TDx6mXx5BB1flE10yoo4t2xpfFBOkUNVD4YwOOEgIV4l8ccBEpBkzySXnfAE2aned25tvY+mJH
0hTnzZ1GqJBJz/uL4lbSKlqGzpwN1R69SQinj4gIa4UeEwJDbHpyVhlzSRYi9IpJu8owdFpmatbr
PcwqXdsQ+iuRDlJBSMCd2TqCMB5Pl7UA0DaRxrsVjuXGQ5dLrZ4cwvPk/exQ8m9UuXDzPZNVhmzS
4/pI3qjrRvJSh5/uY7cX00P+LPKlqIBLmVXM8ZmRtn1yEELh6dG4Q/gtf46VUhUE0HKFR9V8ER8L
g84s2mwv1lRkxmmUMnHJ9Q6yw4bTPW/oqCjf7A7sXY/jBLhBbqkC1wsqPrRHCx+6bYENSlAHMzbw
jSHmsOc+2ofkd7X0nWOIaWHyEP6vxuTpABZYrVbw/7Uo9KHAGpSw3DYZ8RaiEDO4IIKOjb45XJX7
6r/esHZLGIQwySTLif7kEJlIF6uIs4O12hd/EIImQtjbpdI3MtPsUCsrl4dNLmBokTnFzRVmPl2e
vX9KMyo2ItOzAPKl8GnD9lMEFIisiJIiT391SaWXrnsO15WebElIIp/EULDf/IgPat9v+dnFPOXS
6ZHAi/Pdz8IWac913UuaGf++S086okxhErJUawj6x3Vb336FqDPFBjhvumhWgxho4lAIj1BF42oI
DhHxJ+t0vEmnDTAi1J3TUosZZWX4a/7LOsJIHQHWca5bNalmgNzszNhQEXSioWDA48UkG86V4Nh3
2Sm9RGwbXuzFTDdyJW7uMkM7mLeb/GMvpU87QZkuO41zSI3auTnaHlgx6DZK131kiFgfY8kRL2+L
5LE5bUVYfSnbotFzSK+9W8pbEszWOVm9KSVUAT4XBStUfyv0uGkXRZo3bqMJPUtnTHu9v4m/I/i2
km/MQS5Q5823/Ab/lEx4Ov2+iUTkeFgh76Xz0K2/Osiwh2TMDVRpX9G+l9l664Oxqtkem5nDWaHx
RsAYqbbzmqVTcB1WZQIu/QgMPM84h0VHyj1q32KnbSKfhwEduG6Y5Wga6uuylUEGG0E/sSn4LQ2o
zueMSQOg73MJxp3Fnbpv3SLX7blYDmY3uEYFBv6G3Ff/QvDgrcLCyrJ4nkkZdcH0oYLWoz4KiKZK
UstmsJWTfLiTneVjKxCDyat1wb3pL23Bjo5OHFXSK9385/sjZ6QCBlRGKYJklHPouU28HHuMF2EK
sPeKUxachAnJIMTZV2y+Ft1bBI3NY8VZ0i5pp/PiLtBsQCeF3axmX2bF09dRTmeMmUkJCn0G8lZP
67Jn0M6HwLrR7feuIvLeU+Z5ItptdcDFc9F4qn8Xa1Fl6Yug7Mv7n9g7+Nb0oCqF6fMWZJO928sl
ycEZiWm8MntrutUqk4vYq2nxr6iZ4cOLprMcUR44XipcBxWYbHt5O+VSfTSMmWvD0dh5rdjt1SP6
n3pm7A5kcnV8pP0A5Lx2aS8r7kh2pWQv8r7ZUzdh30+qFQXuuUbSeGdGyGP1o2vf+R162sEiHtnY
BwnSYCAOebd1WgEfWBmy5kk7SMcxvZUTovq3OYgcjhcXaz8b/WEpiSCrknJJHBm9a3lQdDfKFOeB
74KrTCUUbcV2okavHX27Wixh2s8ipZCEfdz8VT5tHA5CbjhSt7/ilWeV8rP4EHL9XuOsK6MiUExT
O0BBuAdmj2x3ka/wP4ncG76xn2nvj/6iaJbm6TKmRho6EOUN5MEKD3xhWdu0I9qJkB8I1jlQsssq
EuGtgs2aXMc5NUlkeuz4v0pbGoJSxTK+rRdzljqdqhcenHLMgkMpX7eInucPGPf9jxtYg+Q1r9Cy
nFvkHNGLgUhU1ejIYXHugP/I/WzDoDAe1uApKFjkwuXKNBpHDrRNDAbUZJPYLHeB/4i63dphpWHf
QY+vexc8Gv3aw8aSmG//5ndNgHP4DrVWDvCnuTpyUrfFgU/G2FTlyhcIIgou/jNoXg4pAvinny52
uNXFx95CWKSJY2Rq6PdLxTyHQyfADw89gpnrKwim+rR7OUgb4sf99V7OxdYW4atfgViHPP3wNKpp
YOI7gOAsefuSR6gQzL3iUPEMBfLmook82hGEm6DQBf9bj5aHAnOz/6f3D0toWe/LBH/ZDDHtgHQW
HWcThMLyrTiZmswkv5vPHZgkRQvPvRI0KQXBjjBqwA==
`pragma protect end_protected


endmodule


   
