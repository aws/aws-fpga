`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
C6Y8nFE7/2WhxOEJYmZ5GSkWjsnFVbwsAHA/IEFb3EN30DTpTK9v7mBPmRNycqYkIOvBZz5EhOXw
050+Ofe819T9p0hiK2wWtm8Y0X6N2YIF0dmMIOE//tAYFh5U5jSeSaIa8hOj4OOPdduuJThTH9ab
r87inxeE1EIdTN5bBVNgIdjZ9YAoL9RNO77J1KTNDRGQrfjBpU5owBx83PUN9HQL94zLAh49cdsg
lm8wElDpG05EAnhHCeWqLCbDQZ9h3vaCdwoFTimmkAgOQN8kS3Nhsp75xo247WWJDM5RSRoqbu20
A9ATuH2GCb5E+WaRfPph73vomuCSZRNuyWH14A==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
4xlHVyt2yaccNP0PANb0bdAqhdaPiqW9MeUYbHfIofy8g5jgwyxFUUk250NdraSBhqksb9sm+Y+H
aeHw1tAD9adpEfu9WFtrGx5XrX2oFpUw9NurjqZUaXBDY3XxWvXTWlFCFPlw91Y+dw597jLfxe8V
k+FI/P59YTPbqx1/cKY=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
nGRMirBzBI31lAMp5SiKUS/iStyn8CIz/NrlVXX/KIpdM2ILE2UA+WgDfLP7A1EciQfTvMXOjEQb
eoiUmNTv2jUEy7wPNQgZSt2TofaRZr6p8BpdQFeILf2FQ5yP07xFmlNLNE591bTsGRjpSAcHl3k2
F56f3TK6w2dQh4N9u/s=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 704)
`pragma protect data_block
yeDrOcCsCbxcqJMkc4nWhzqQjivTQEjpQyaHVVj80ibtM4/9NhlKABHfdGa352l7u56HY2bj9ZDV
VOepdraV/2BSiAuADPPlNBkHupAHID1FT/galsHF2bzPU91iLkB+jTwhc3W1671DlPcaPCkYsBus
78aU6DTuWVZxY1OQcMsQFhRy7RFPsPUwhaKYAP7hRKMyawJ6X+wN6HTMmJZH6OdxFQ0ugg9pUEaE
BSZmo3bXDC8KIfoTxcqtJzGd1zR63VIPydoqaeQs6QDi1HouG73T3udXaigF+fLqWHTWdLqJ5pJu
oa8hWJPvBVUmCMFowK3XRanJMYce/vK8v7T/NVHv+JHsjklRpQX/6S0/udS5s7NRafV/VTKgnt/P
b/aIljJBpNXJb4+Bb/US+Gbt0n34CxokVDirbaioUpwZ4H4JC+/49xXfBT94EgV2ffLSnfZdr3fq
jjXO2KwOAXRjM9mdFfGQGHAMRmCKS2GELQBnT2ADHJfIy3JE+iB7svRgpmab9RWUyVfjIxT2BbLu
0+NA2ocJNqCWGnQNUxMtl6RR5pdrUM9B1AeFw7k9oxpq6AoreB9A65PZN/JH4KBA+UzY+Ogxo+W9
ANVu7JQLGSQAaY/rEE3vYt6JlF/dFmEsC66W0dBp7Se0VPhf03qwLimqIEkgInuKt5ANltilnhCm
xp/hBJ+52Pl5NVvUFF+tm+aFMm10epUKUOo/8W6kBwdWp+oJc1nSKGj+VcMSCaNUvdGG4dgr4f6W
M27vhOjYcq4WtwGhLwc+6FUSIxCPxiL24kGCernht8kf4+/WrcDTf3Xswc6+s5tf8ScbksXV5Qwx
SF2u7bszxwyNK4vF4w6A2FxxPCnnMXuvGEj2+dV2hA2LArh6Pd28DqCvfShrl+V/F5ZCTRu4Okpq
JvC5Vf2b7QMoAs/XhOsRNfP43w0=
`pragma protect end_protected
