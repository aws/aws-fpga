// SHA: f463fc25b8464dd6c1672ff28a603eec67bfcb40
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2016_05", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
QAB4rDjUzv/yD2xw3Pe8jyRAGvsJyNtu+6Y0ZOgOqIg1dzL0OjOjPPxAqpIDXwIOCDjKoSxwNgzh
fGkdI10uRJPZCzUypNRGojt5U2EYhQ28OVzdkVDTyT6hGdeTsnvdRQWBtZqfOHCjlEWFnObUh2qx
Wvd10C5Xlym0moBuh/tlUBU8mWVWzzG/lORuRoq8BfnGERGyv5282rGZZ277u5SrnyDYZruAvatG
AF4CaCMxTs2aQHBydCcIrlDat1hIIPlgBr9047osZN+HMenP5XFHrCBoqFE0kXPjDWOxGCj1P6/6
phe3qPD5tbjSN8xkKbrY5vWC8u4b1PhSyTjw8g==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
NSrB/UKdw4exbf1MsTjckvR0NOD+SKkYr7CxI+jamjTugz1he2xhkOcw3QwLQVeljg4zRkoewCwE
dK+dBhSpMWXiwmnWZ9na6ttpJUOyEAHCPMlpPL2MTFxWFD206T3NnplXs+PMU8hYwwUQtSGGjE7+
dtq2Ari7HTkWX3YSqGo=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
GmnYhx0fXrZJNQwY+ft+xzMpcHIST1sCELD2mcPAYWAh0pfxeGmZ696o9SoLhgC4YFbYb5cYK0wr
HeyXguh4j2rtNdMtyyoYznbfdbutndwzljSqt1yrTSKb64AP3T0pMP7uSrjNt5CdLGuY9r4spa5D
VCW40Zcm8zu+VIpOyDk=

`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
kUEU1iIf0554SMxbaFIpGy/Rsw8A9cclJvF4oBsUCyDo6scH50GJ0xLNAyuSoifEswpVl+NXdFOh
97fNCux2Gg==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3504)
`pragma protect data_block
FiAQ2uamKXFNLRpvuSY8QOVSz5FxQ62qJew2P+3dpXUxo1wtA0O5vHq+pVQUZ90GrMMEneQydGk+
JAKLokfver/BwbgTKDmiO5lVl3GI+cUvH+R5chja4I8TgIppJiHdNsFZr6z5ZuklE8ImC9v4zFyA
UE1uiSa8I675pDHq0mfFumgpJhNaUJDzZlWVYVAGymUoJpA5lEIAkXCk09jR/v/T1YHdcJNWRw7h
MW4DywbdGF/HrjOWkIDqMkMUO2EvCcU4Xwxm4xT/QeOH0gZ4u9B6ioixMB5+oG23jxvcDU3MZ0nS
ZU5S/WjapU7r437hwTIvDTFD3XYa8oQShiLMPGCIwDMUtnfz7isjxDCz0mEecIzojFxkss5IOWzB
nQLD+nk0D02rlejRR6gZu9Qi38KMm8fJnuBdDSwrX9mBRI0T5YR/HTELy498Gc8xh0M+e6OsSIdN
DXbp971kdpJxY0BJZDmva6/wmpFDLgANIPwGdU3kBIoUcnuHqpgmfCQfztsskWKBC4vKMuNcaTQj
tTEzGhmK4Y/KWTy2mWGjtfpMpGH/N+ccirxn9o9bn6pREGGxhEcxJRhurto5OgdXOsbCNXW7fRQI
4ImidkElluwnnp7Kxk/atkUdJFovDFOYnloST58CrLR9e7S599kHLj8AUYWtEmMPTO9G4n6iADBJ
T70GQMMmbQbTJulfstwS1E/LZXUslXVAVRuFduR9kxkGFw+qrEIT8+6KGEPxvx4yPg+lVveqtB07
/Y8b5FqclAm9/MMcYuRrD02m7llO3MHcOaVMeqoYMC5t85iKmnaPVZd0ZrSJgUPu2/7DKdEfx4N0
oQAImPhRzMGXZ+8Ft8x2MrRUA8lWafVvlDcBkAMDqqd9wA7wpObO9NNZ2pSnAhr3FpFapipAriB3
kteh8olJF6oKPLf44bnArpyorDI5czOnHfnMV1bWbJ42aTViRsK2UaReno2MV/llWzGBOqsusPB4
g5QT2xNpIS4mePFrpPiJ/oB958EPMnSV6D9pn+ImnNQ1tzGSTMYFAKxwx47z15o9CdnpI7A9TPyU
6ItB4CIDoc/323e3DpbQt5q11UzuGhDUQnefEwxrQYgBqeiScX+pfgFGm1/vZi3lhyxIlBcNCxkH
8AYccnQeCc9pi0d/mkRpW2OWbdRdg9/kl6Yw0NfdXmIz7sUSNrcPEyxDvfusMTMBu+8XNx8+MMgu
idf7nnbLuuklz4B0gwuHgUivMAqtqllRtOeSKTh/jF3uYyzJ8zHgkPCguaV0/VzTb0KwoNgPpUhO
OiD+/zHemQfl7g/nNLllwDgHE0kCIpii6PNSpHmJ+2KOc/HM1pPuSSFhXLyAVEIMnv85uJuZe31Q
gBQiPMhw6tf3FQeBj4JT77DZFLdB41KCCYspftm5K/3fypiSFX6Mb0r4MrAh/4BJlNvg3LLiq6sr
uqlMcmhMmVKTom4cNBMJXNILVB5s1w3W9pFa/qDP0cCchHmVljYov/nUVg0rPfTlwYhJy3wZADaC
zluD98lNVpUBriVgWOM5NlM6FLrkqEEY9RIF6M+DNz4Vake3LSFn9qvCVCduOqf7GBtvanvX2LFb
ckRi2/3Aam3KVrRdNs2MpybCejRSCqKX5dFIT8uoLllSEm3aQQDDkCsN7WPe3zoKu5Ta23nu17Nb
2/dJHu+HdF+RWWVpW7S0rZMmf47KwmAqC0kzW6CcHIbFqk2X4e1TE6OsWlIr2BcudT/97/qBX+S2
m5zketoTEzrseRL63oITD9SKdfKFc92vR3p7eloKbGDfKeu/rXCTNOJ/G5inXs9A/FxMJAm8chwm
68nDUZs8Ifm/2nZJkR16TIhVrVM8t+1Y86PvKTzk7qhWOlqI4gq/AmaOCT9ItCbTEuC0AjFVNoQU
Y5d8+u2aCnrGd/FDYwRfjQt1J1alZs2tfM6KrCldt5uw1aS5eKm5sOFodv/PZGdN5UPrY/Y5GnAm
gY0duoOIfDhM71n0TdehK0rxXClr2YGkWUgdQ+O/mXQNS8AFk7zQBFFhxQm6lGP/GLY1nA4UzsiD
hg8HG9IJs2Suio2KoB05Z4EJ+pw23FCxd6pmI2983PR8p/Z4+FTnV4bZ7wSvB8xdOIW7+OhpVwtO
TOxm4nFnucCMBHr4el3EPkuhH9b0bg43yxd0MmyWTFUOhUMw3iGEZwBIHtK7xqYvoBxVzzp0yIHt
4K2frPQCbGCT8cjd+J0Umv0SkQap4ysw2bmUpt2QjkL2JHIPF94/YLhmc/0ev/RUFgSqhMX5/47S
5lczNCK76eE6k4N+rKbCVg3Rehs/SJ0nmaCCZj4MCjQtpJaY391pCvSDJkACQlGSyuRhtjSDGwct
hnAXvNjtfPo7pgZj+nyvHuzFCG8fFuWg7KaQRRgPuaOP44Xtfw0LiTZrXX7esM/OBGOPTOAYdD1m
/ObZubMzjirAzfkXn3J0gN4SQ0F9CmNL/uwUVSZG9Vmbo1RdwuX4fY7XPXMaLmbltN0pqZUmqZCO
xuSiAbzkLJ6u3HScn5hj6GrwUW47Qpw+fUb8wmrQY/sBQwyKbcE7snPDLYeui8jVSShPDRG2Y3Ap
G3lPaXZ4cZsgd+NGUxqXsR+brmN5t83mAzt5cy24hBxNvQ/NS+HhN8e6v5zVQg7VRaYa5MtXH4ok
wSsAcam4VXGnDpPfCspUV4dsK8KIxDy3zgVe3g7aDiy1DacrTSWDDxhBQ9ogMMxb3Q2Lzp1gkx1s
yXXHBX2CFDgDyilTiBO9UfDE9+QHyQ8c4yc9STA0aHMgJ5etbzN0i3Ol/phSsa8yI1ElKEeUKaxt
cw05FL75YRGtgLE0N7YGTf0gkkNjl0g4NS4Xytea2/aopb2mLI1qxxLlw6IHu/emxtU2+WrhPhdX
xeYeOlYIwUiHKJPKG1+ih97WMOuKQDWccc69v2chaK+s6LA7OJKYRxOgxNbFTmxZDabumCpqBP+g
tt+M2Q2DJ4SpD1m1y9Nt7Y4RjHSdBjtAcNETlOLEDSczycNiVqilhJxlLtrU2LiRq+isiCP4+Lre
p2Zzbxu4q5XiydWfgRNrIOgvdHJh3UiR9DPto9u7u1gAltSvqTv4CLPnV841ufCpC8xe+sew1XT8
a7uhLSdSqBnYivkRjWoetb07zFkXLgAp+e/u7qC+Kbfp5uNxOby3I4I2P5EK0sSRW5rNwvBxBDiF
qxK5rSGPJZQqQkRB1m8iKvw+cknvKVsDcSeCOuApDQI9Xk/+VxBL0TuoccIjkizhsyvNosgwRviU
WvNbV/xZ+GEfwx3Y2C9MIN7mcodD+wolZUPph9sof8hniD/EkRBymJy1GtLNpPBIQNQs6uAHiCoC
oUpq9LPk/XOkZLOe87ib/EpSXQHT4XSGxT/9c0FH4xah9Z4KKsicARNKHEe7dL2n6C7DjblNSwyI
r2Mxe/bLbcMHoa4c2/gWnpNmmfybR7rkKzpTOHyRvs2SzyiuF54KH7cExXnDjroxrosLWCY7wvCp
stqjVf9hOQwTrAPKandTR4z2woSHa1kgX+53g4RN1eMnod2nLhu/uAq06/Du9xtVMhs/V9guGHyK
Y/r+Y+l62RgP2NzYti8XTQYW5B9pWLqv0JtiUXPhZi0NbMAMOi+vAev6okxBLfYgSOiY3kaScshq
dkt9bctmTHvvAZuy2mlczvWfsb8qvdT/M1bR84znXJ5FVuOR4MNHDL/WEOpD6AY+HD4AoUcSp5Xq
GctWaTEyXBqhpu4xQ2nCeHdHCnjNwxihkmL0NwOzUBa/ZfGyq3JrBYBwejzmoZ27EaZ/772200tS
TloJh3xmzs2T0wbxT6Id5UvbBP0o/GJExgtGT0jIrcNiLKJTjxgAiX04pco7FzdvLWufYLRfG9QK
mjaiFwORDFAvunjJ7iKwCbcxMveKH7YAMhQeHqG+7AF/zdTvuMSJIqSNhtwKP+wmPkGYxvSJtyeL
SJaNnBlGmy2HOI3fPqoTcVqvzKcZmWHXRwPmIUxLjjkU8KhDHIsSiGuDBHLg8A8EPeg+7FUnb8On
Rr+NHZEJIgTglRSMtno+yiOiTAix9bFjsr6zSUOEH+ITTQ9e0j+gouu+DCnuS+mxqFpK6tHcAPPc
KTZZ46VmfetW2+DMPz2B0t3KdSV7AQsLDRZ+pEsGs3LJR0INMpdwKQTpHTqHJqOSQi0H668zXsDg
gt1Idg+iAPysKA491gJodRsZoQ7zUTBpJ8Etge2tMBTCFhFbPgILGtye/g7GTnG9UgdztW+LJRUc
aOoTrfqvxfbXG8sJGQD+EyfaEpAWfk5pV+NE991hQUhSofZvD4ZvP+CwYkM5J5UXKOiapqgbeyiI
LPqVRA0h74Pvlsolo4eGD3cbTBsgJ9+8L6z2/6zQLykClfuJzkfeOeTPkijlbiND9xx2Twfyk+8S
aNQGL5jGxEpyRIEJE4jGq32ZyUhrZhqfWQu48dLLuC8g9+9Tv9T3Fc09fZYtWrpVJzp7+X0cNbKo
jX1TLRJ4e0LjbiZVOV5x17SMSShP80/wEjDVl6MYlNvg4xRZzuu2c0wLWw5h0hp8rYdGzPa8d1tX
6xhlsk8mffW7ntTbq1ZrV9agRALBxI2lfiqmka65mqebMkSS3+t8i/5/YuN16qDmnkm+bVIJdSJN
/7B1epADZvS98RZ2vzFLOmBEGRYsAK4Ag4xn
`pragma protect end_protected
