./../../../cl_dram_hbm_dma/verif/tests/test_peek_poke_len.sv