// =============================================================================
// Copyright 2016 Amazon.com, Inc. or its affiliates.
// All Rights Reserved Worldwide.
// =============================================================================

`ifndef SH_BFM_DEFINES
`define SH_BFM_DEFINES

`defines DMA_CL 0
`defines SDA_CL 1
`defines OCL_CL 2

`endif
