// SHA: 43f4f449b937011c34848123159f70bd11b98098
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
gilSA/S+RcbfQ91oJrh2hs0y9lp0uGAsaX67NFrN26ti66fuBJaM2QyzwoNz/NvpGOY2eGgSQz3Y
kk/kiL3mKauFeV/6W1IpfcmlJdAaSCbcAZFED1SNuyLFs0YcrKHI3nsHZnYftg6G1RRlO6PItPxd
gAaFOd3lQROot2VjOr4JKkPPThrdpdUDgSDfGML3naneApTaZjCh8shj0omR2X5ifLAsCfYG2NSN
B2y+8AYdPZhd+j9cLHdOBedPrBsUAN66V1hmSTci2N8cGsD9/BqDm/JdXYQ8p+UzN40PnvKwTXJ4
+3U5lclL+7+/iUPAYjDiwxf3adjVcVKswQGuTQ==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
B+ynkNXGSpMT8TANBXqhzMS+Tmj9z9HV7EJT6Bi6W1KuwCj2W12kiIW8t7QUvjexyfNgw5bKolbm
V1fwYPyH169xD//DGqseYtgdlHpzbo8Oc/gEAEaak/z3HHx+1x9T3d7An+6Qiw6XunPdIZW2aWjw
k1/Gh09gc2OLm8Qojxk=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
mBT9VDaMG0AYEciRHjxiH7d5v0MwJi1CXwk57TS05Wrjl9I99l86YvR1QpVaDOTEUcOjcnV5SFT+
/mc1bsz2EFPWtHqYJQ7Ze5WW9CelNmufFTbVaCu4nPC45R3zYybhlFiPG+pAC3/emE6wMCnZgQNF
gMAWnJVckaOaGuhP7nU=

`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
bXABHU4bqxO0lz6VxJWa2VQjvVukolCI2A/xMevhysbs7or/1IG32dyzAmrkBRrlcVwI6V1/vXXD
7YT3W9vKrQ==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3056)
`pragma protect data_block
ywefB3seeEB0/qtRprMPYTEoM4QYtCZWhrU+EGp6sgOf3rJIYMKXrx9ELGq9YDtWbr5LyHNe11VD
GtRo0Bi9o2hJxk0kpz91EZKCYX7fYPWGGWAm/A+4uNOZNfzxaVVJxXfJEs21b/zPhbzumtPb+3Co
aesPgpdbFjMcFiXFZkuRVJg4iiAPVYe9DjurdzU1lIOLD86f3Ht84HgQcPsCkr1/ADeg6I0GB2RH
t8Z9SIIXgWK25zq6M5eKYfB5VxX94SFwKv2SnSF6XbIE1IWOqvVl228FyjFkWZh1XF5UGTRsw8Ms
UxpVhacpsjotjYYZMGqU7TT05x7XocB7AyjOG2OrGySkC6ppZAvNQZihRf4Qz7F0w3nde7z5Lcqw
0FG+WtI75Ff+bfNmxevb4c/alQOhyVxDyzBwtDklf96kMi4XBFX1cX8P75iZfKo4aEiQTvXps4/P
8o32CkBg6cv5avrVrhADrFay+zq75n8ztUUByFSNWw6e9vnT/G6Qg2yrY4W09EuTgdIwrKhKrhxJ
cPze4GXKxet+Bp4UpNteZsQLENgWS5CC1Px/kost7tCrGU869aURuGY5ybBpDjL33mvjapi50Dq8
0lMcqGfS8tmpDzrTs549RS2Y28wIaJp8axm1cRJP+Ohj8CdvY+eKyHOiQfuKasAzcSMnT+oy7Muz
+o79QsvoPLhNredMLUDKTRLHghP3VfrCI0v6r2ziE6Me9CaKpb9kf8s2STg5shKlnWMUsFUG9l+/
180ss0FH9KDFxWHGw5sMW/CcFSbBsHWs0eFn4FH7pfWcNNH72F+5dT3uswMQOTI4a7tZRcRb4IvA
m5aT2U8olbGncVjdA5VcXqZc3mQ7+ATQVkw+NiHUcfSiGytLB4OAq02y2WZOTFHp1llWLu35MsN6
uUsfWtkQ3XVebmASqGqFU+zj1liIRVfmaF1sQQY4+ff088YF6lbGwQrBxCMpvV5sBA9GJK9n90gl
+CZ7zY2bFX7JplcrQCDO7EY8viqRidPPolZd5bJQBcpEx21w2tNCNWL/bR+BE0cnjj6dSuQ/KVpn
vbPwCTVyr4VpHhNZpYFXUMcK4yZsXl3ng7FhERSz9QX9ltpfTEHuQKB/7lkMHwQrZe63VuG3ItDl
g7vHHoYfcRrnbkaegQ2os0gJuGOXom2WE4IeN2crczeE69fQ8MgTsW9CYtfCRfR5dAzQq68nQ42j
4CK188Vp4GGB6p7Y9Rma8SY+GYIhBqr1e+zjaW9iwbpvcaWDYuAjSF3X8brchlKj5ApOCoemlA1f
x+Bno7UhnNC7ksQH7jRCvMbabXYEtzJFqK8ilou9WeKPMQ3R1SsfFCS0sNfRttD8ehOPHJQh4ohD
6StFh3qi+SecHCdL7aX3YPaKv1VkeHlEeiVroVIgaGZJhQgW6RvG03l2l+2UIfvMyhi1bKncilCN
X5DWX4sRzFp9sZYxq4CffXPNojCgHwCDUZDFvdDZxxp/rHAHHkLgA3r2bGoHDv9dHYfs8Ds0un0S
yzkDms5vJyHl0FrhA8joMp4c8MzB1ovRyfxU+sjX7x9KCZXZCv9Paooy1kIF8Cywe3sOSKUiwSGe
V6kPB8RVmjfkyNBujIY7usxuY+PboZGVsDVqLuhd8tI/tp2SblQvm9O0m4zJkGl1d625159Qc5Wk
PnHisWQ0F6HFOxFgL/RpDkcqILWFN7kVRy9ivcHV9ddjze6npv7TvfUKnx9DesDs0txxitrl6igC
rOsW2D8/HlRejCE5cOPxa2+HXdavmuFGe4kgRR0+g6Rlp9H/dcQAwk306rpZz4Lv+5nmVIGq3sWe
Ve0lboaqrpI5LfA93Q8+Z20Dx43zwq2sbK4jkfd+KJyLXsqIy8nYdRUJ1rF8YOgZI8l6qW8RuxWl
CAizKmhdDf0XfEKb++nukF6VCSBonkVIwgzMUXQ7RS5V2R8JBN8HCzOh75i4jry7/6qCTskcuG2Z
JPEJz5aGM8EoCvlwoi7WwoPsaCl9lijp2CgkuQcuDU+2+zL8CC4yFvuJsj8sc6vV5IhXB/hDYkuj
/6gONhzUg7fCcig2E290sAKXsjY3pZwvAwDMIKH6RWk7JU9HSaY97G/hIi8OUlTWbBodR4qTuPWx
9Ky2GTL0UNbCy3pazqPmRrisbkFkLqKOx+RfyuTg69C1TvgO2dfg7PFfPj6gk8P3tUYT/QzSjUtG
S9N18nms+D6GoGJW8B1lLFTKhwIWNsk+5Ijr0+xCuG2lIISFDHfbYHa4eFGSh/eGiaxwOqIcRKFZ
UY4+KVCMGFn2agBkUaZUMhkoj6VV1XU5Q6m81j1Z1908My2uctXL66cPS62ss5sZ0F8ahdgk7Pad
bKQv3IuUFGkZ10wmFx05zARewtxlkwpmn9fvYSPNO3BEbWKX3qIrA0TPtSUA7uLffvEBsoMQdM7L
Gj78nyNXaYVaKQe9KS1SsNYiNYYWNP9aywyPSqC34mVk2tUN/B3WEUmW6HmveYTMMx8jtuf8g48X
9q0/wfwgbEA5zjU4FFz+a2QEogdemTr3uTIZEkwSJP1uIGAdzHxBJMaSDm//zKQ7ZqtqTsN8+SaB
hNjEcYmcEtKmHhlrQDm75vYzw4TsbCXRcaSY8S+SnUKk059+LZnGEnSe2Yhoh/Vuo84dk+uigpRC
Tyw1egZiasDDqsuY0R5frGL94MEyl3e8FiQQFok4tOrYOtBMpfJyjsJuI5/wD4RsJ4mDqJ6mlSAH
/joQ320ge0po2C3CteXOqNJ4T9JUMyYzi1oOsyj30yf6lD4QV78Q9Q2f4XuW9pIJ3mDDCw3pGFdZ
vpkBsguEoNpZdEMPoABbGaBkLqW9gDjbgsAe+HR3H4HB2BG5xUseOTTIslhZTY9ZPc2RcORHrqOp
x8NxbQATGCr1ynTdzB1JCpFOSLA14V0NUYS9q4PvxMJHQsZiC3IBj5Bo4xG+FUVUqAsM8ReERPyS
zclgHFoBVXEGwbWIL80D7+BigyTOuhtWvstx8L51Thrya0nX0ykQpMNtDlFiOrKouVRilFPgyliv
PzoBX5jYk/z7OFu/ODDARK+KCtcEgNSWZ52aceBJ6SpWZvCtq9Z8aIWwkPSFSsxilJOlRq2+TCcv
CgcwCF53ugt2dIy9SyZ/DB5Z0/78fv0wTukDyrFyPOY9Y1NpXLTo6dH0JEg3uyTtctqqw6fKr6lw
9LuDAN2Bwm1hfP3m56WOkTM4UIoR/GR3CPKcmS64yGpqtscqwgVACXDl84GmdI6unD2BhP43jluQ
Jp+CvHwk7cEGBbvwhMd0SegtMPyookrJQ9UyXYNCDeUUAt2pP4+UhJLuk3tZuWmZjhdFe4Fsr7En
Z4KLS4t4V+JQ+tUMa/UW4lypqFokV8Dt7cKjbpySkbzJuaQQAFoyNCAJ4EaBkQ+JtR0hlT/d93y/
wpmK7BqKAsB105JX0OWnO88dOtdpQ9Z6rDgIJuPvLtygt/mLmDdexkKoP3E6t4EXQNahCq9rz3IP
Ee/XDi0SvhKFKxSw4WNp7/dYwBabHBMKhFO4hzrMwwsq4nryIImiHM9jVTP7jSdEz3LL/ALFvHpJ
/CFFTfotG4UUEk3T6UxgStP4lwhUTw1gWqApSrZlvcjUMVjZIDSwr3FbS57Ki59KRWv1e1Z+EwmC
0JjRcymVEDC7jMxiThIY/6MY7xxo21ve60Y5lmDk3enRcyCCSk58Tm2izY/HKRVECdwCMX5nxu7D
RmzArh75vbWu2ZjQCiDSuOpcEq5fH6cvk95E81H1Vcl5aOAx5gsUutI1O+sTved5kIqvejNzk2mj
P9JTJhwN1HfITTwwqosQBekaS9ofdAoqrqmo0uewCJTn5WFpTMERQML3D9GkwToBouK/1e9Nh30w
0CPAeAv34ZJX7b/VEUnWmTd8hgqqL0sNYOhohieUjm+h67Vs2MqMRPPhIRxqeYuE3JsRvWkJ0hAJ
spl8VlGwv32euqC3v0FQgaXVqTTsEIxLJ4L0BesEcWW7u1hHoSYnc/FBY/h2b8WVU18BTXBFO7Me
pigqcvTghl4tVWHEsTHShrl79DenfLOrERCV5rStE8P24To=
`pragma protect end_protected
