`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2024.1"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2023_11", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
mpELdXsUsqDdaTNCPKFoRJC6P86KVNo4kpQ4ezqC17QGB3ZaQt30d89t13CSStLRjNnOSCIljznO
ffnNe5QNzUwh+fqf2jQDQMEoNLP4Cyuj7axDlH+Q0IH9agshshwYT60qnyDVsoqeGdeltWd/6chF
8frZdWc8gp3R+Lg+1U/VM57CtjC2CY3iYHimqLHEBCinW3Ov9wjGlXVJ4i7rt+j5y6yA30MBNWV4
Rl2d0Mn1O4Z/TMoQIQuVs4Dz0gA9JTOuVsa3uSuR+jCiuedh48KEtb/T0vkYk186R8bfQSaTNVaQ
NVnyJAKf/Sdj8HePYO2G5qyzVA+ncvrE2c/ryQ==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
mmfUdwiB7xjXymhqZfXdlhJAcTD+Wpy8yAQ+hmTYv7OaV2xxA7eGYaVTSpzAPGyLwHT6fr/gbz07
IZyBz7i4YWqv1jOIxti62I9V/HJFP6Bokfge9VmKqpPx6bPgM2qOEMBJiJ/CG81QVAwx0TUidVEz
FLbhuPQ5wuvLtqHrB80=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
EGfoQcBM3Ah3UQjaRsmCkB9JNr9rvDRALiiMNj0AbQ6TJ+eSUY5hHdufJxh+YC7ZYcqQFZXlJjXx
/Iu8Z6JditWtxrEv91iMmxlpqNJjjULklTfL6469qgg4lm9yGVwWmKdwa5ZLXSHEAHq6pDILo5FK
YT6h0FOv9Hdliq4CuxA=

`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
QRhfzJhqQmYbzy/2BeKu7p32l4ANOz9erebhNoXedAbD7Iyej87zd9LCD2uWow2OA6mESRTWt6IV
i9Q28g/ZAQ==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 118928)
`pragma protect data_block
wIAgNAQCH7Ijwnf+ePcLhMIEQzzgG3iJcPV2vB6kSSrLcMgZjwnQ4FnNKmiNHfRj+2wiswYydKSL
sNcq4uNQLCmzUSmPPaLgBaMbXiV2wCafyZ10c2BWDRWvfsP3O3Pyy5BMRZ1cZcfAjhwtIQNlKjCH
tCpK/goJXHnJAG5O2wLqpAuU90CKjGIfX1qgBhEuZfeZ3IALLEbUtuaqNWm9VrfLj1YWOg1tbgfr
Mc6UPV4xuKmIu32Uzsu8PD4O2E5TeDJCfdxsnuUmzbOC2fze6Lbw2//suBTUZOJpK0qwvjnTdxFZ
0SRqo06Gjekc77ss3XWhjL6FWLQwb10BlPOuzUzlbXL5tJud1UGAHirelMwlcWotrBWmwBnAfcrA
pAdd/Lap+9V7SreVkH85Ia4Dey/1jakR6fFHYa257IBz9gg36hKK9jwMznMbIKchXeMaxFk6gug8
LW+Yz4SCNHPz2tX6JPoAZU28sTP19r9YqZolctkhYFnn4zTdJ3eNLhivACUW18WU5NdweYFlQkMs
i791BPmTWBWvjVwnTpfNypnih/Wv4wyzSAPoh4MbbnExwNuoUJDd6jjEBOB/S7zc6YM+uiFrDbIJ
45TvEuMhsMCT/G9H1IzKhCV7zB/VrRqWrvWIRKVUTpJsjAvA/PPZZ5HL0f6NQhn+2QUbE/GuPATj
YgO089KpNlZ8GEXyi1LfW8LSg0PaVBMk6tsi/yrNr2rvx4r9x1TAQByF3q645QQ10mDp+b2qqSKD
lLNvjWSBsGdPqnZ/PbRPNtfOG+sAJwobk5RRON+W+qYU/BqGQu+rqNZRV1NMutZ2OqJN2OjmdUHN
H46aUAOpWHhzsqNeRU+teiDhnpaohJtZzx0bplcdRLsc9QPCuZmIKmR6V3cUly7z71forGi0NMZb
hrERPUzxs2m3pRiIbsuiu3yUtUl9SeM7Mh8w+eSgeVj47qgAomW05K5dNLsDkHq+rXttrp75hg8Y
QJkpY6M9k30kx/k7yb0B7DnIogWzWKmHSX0SJaDtIzYmkDMwKTMsFOKP2RDsQKQJVO/7OWhHDnx9
wPKR0g+PqFfF/YxEqUJYZNA7r/7/Mtb5CvjaUt1p7pmdkyRno4u4uumjh1A+5bGtCHSHaAl54t5w
lUXlsRBoy3FvvNYGykPaNZYRu+EgOoEUSM5jkqDSFuUMworj3TKZwTMu7BJcuKdD+v42PbhyTsfF
H/RvCIcPo4T2tmUy2BP87O9OlcX1MuWOFXpp8GmhpnR+N5ynhcFSPisiMLzTp7daKJywMDBnhJ9t
IogRe0Qn4y+RxbBpjmkXOU8u7UGMMEoZtqV1GtgO6RP3890NuQWus0kWm2fSn7v6b7QaAfI1Gh21
GgenONES/JIkB+3WNio2ZNTq/j19kbTBNo+x8FgqF4OKO/hq6QAZzGdxqHhqB2PtFhSNWswYsWB3
uc9F7F8aeV/S4Vn1uD89QDFwC/tHPaA2vDWY/W1QsGZ+eZISTEaG5HPcmX1TXHOjz6FrKgR/Ieks
vYFyrmPEJK3KWmGPAFd+mHKt7E9XxxSPpjhKrxKTz2MyL4CqDbWOrLAz6i7vbaGA/ntXqjz3GEZe
LyNs5VbBowKG5NVnIMK7wHXOmVhuZWpCQz5u6dADHCYOW/cE21CNdIo+xSHkmy9ne8XGnDUYIQxz
f4Wcba13zuKwzowDUNhp0zIGO2F0XJeghT9JOYw/I/ZSaTApAtC7YyHVZN3wzwwlIHgB+mrowL+D
P7THQuhBIRBf5W3kpOQgg0asv+R6k7YzJiSLMoFRf4xvnn1ySFvNYymedoVkEyf+39t/aF8l8ib/
zTuprD1CqS+Crh9m5iGwkTTAk34ygm5kmVzvIaQr+qv58BZfy24hpxXnKBAfBko/xCzNxpkOvzRy
mwdzTxyOxrJmkHxrqFNbLppMCb7DV3BdcXcM7ZzlxGRlbw5qULNPReWrGr0FBsL7vKzO13cGV1Xr
SFnjzV8DEwdWEIhuYdTTR935of3I7qOenjFYvF+QioCg9oVbWgl9Ud8Gd/cREh9oVHfF2kWEk8Lp
5bH7TxnsAU5oV/Tp5XpHhCHItl76vjfN3pmNQyiaVKDSeMv5OJj8QQ51R2XKa5+FAbggtHe8NdVi
ya+xqN0TvWa2RYOYwJdEpe7zVPu/yAefg7MAbrwYRyfFohm6bYaPMuS3N5buqrQmaIHzxs5ktdhS
P7+208o3rSFkiC55DghUNxMMhj0Vj8p1b2BQGRV3rX5FJFWGoyYrbrdP68yoF1EETG9/y2ToWUVT
WhvqgY4HfRnbwRKvDlFBpQRZLbi9BaYeh42/ymOcOVj5rzxIytD5W5sUQnH8AVud7x7SSbH8W2lg
5DFJG48EtDDeuh0iHRA4F9w47T/f/eQH5o4Lly7TXWPAif9Syp6F+76Pt7833/HgGZIe4+HN8i+R
1XR/FeheE4JvIMSWGqsInupxwforHWB8OuL+XNNPr7oAaeRE45yVjYTpwERkwSLYS6n0xWPzl6SA
HuZzTjlKEIcef0sOxpcP1MVK9a7vLSo9aOJBIWacbpIYMusz2IGPQj/5Pfi+eRBIgmKK14v7QZ2+
w+cVW82Rs4vb85aJTSjuHSNToKvjsFq7SnzC7R9tAKcoGyhcH+vXa4fw1pKxt5NlDVHhIu3O3dla
WRZmZoAqPS4TMMMs6ot5LeNaZ4JO2n3AboydNftmSsZX/LPTbjSgwnogNmVW4HSiT6AdVZh/c+BE
10cuZTJBi/XM2nMnocLvBh9A+S9YPRkBYEDn3Pa+c8uq88xnOzjVWgA2q3jS9lMyn1KZ5Y8PDaiq
sKocsoPpE0twqLJoSoTkQBwchl1eiUQYEaWws/vOFqtH5wyVdkXtZSF7ju1IfsRUJBmrt1gtAH1Z
qoTLtmVJFsJXRyGsXMRmCKu0rOP+gVPlVOpWjX07sJ20XEcR7Mxnhe+W+ToX4qkV6myPXKu5ucod
aAhrNMArlRvZfxonokUtNi31MGYpuq5kNaW6R1txTgSadgxnnOBhKHnOgclN8hkrAPeE7dVZID0H
aULQ3kJNIT/KOVHRfdsporLboo/0F39YSHCk72W16uXf7L6mmVieE+r5pvkFc7zplGrGpHrnW4CR
KCpyh6H/nW4id6e9W3kYyxkOJCjaZJZEV5XBBAbguKCdjCFo7WzLv7lfvt5F+N7JbhpCJVUnSzCm
dC/4F/ZafAGNVqn4uhhyhGIoK1SAhWK/mvjIEr3BPv+HUqzR/Y7JASoLZlRIyy9OXpogmmAAuLlc
RlePyJJDxig/tWfuWgzZqlhiNSZ+5oVQnKpd2qL3GjCaCPacttMNodA0DkZcfJfj1N33dT6a5mGN
s4cnd0OUPl8cdY6aqsSxxajIjynuZdiVabJpC1pJ40zGyRz0gSgR9yLK6tMPNxgkgm82P6RvmYSR
Y1eRLhtDUHk4YSufu+PJ/0eugdircb4TRnPgG3eajedM3vC+jdIrCr8asDKT9YGk8UAWITX9knCH
lKu1Rr7ib9dM6hObT7Vbw5pkXjaX+wtO0yaYt6ofAxSgd8Mn8jH1xbMbJtxFjeUhoehGq7cB2RBV
xz7x5jfChC2OJujDD3/TNI2tMwexxSO7qDoNUoogfqCf4oWgwdx8tI3GdsgCMPeRu0T94QsNLic8
+JVwQUQRW5mWQnKa8FNCIbEB36cWsO+s9b9CPT5XEfSqfryuELlV2D/bJU9qY8cUtLKCMXaZtiiI
EZEmPUlJZiU1MEk1sJqGZgoC19je/4N7p13j9XHdhEDWbUmXhSs9vJ4ThI6xSDHwKxuv6/XHBFEw
YX4X3ygF/85rMO7gX7veLLhsNUcsdJq0GWN09PmmYtho05Q4vajCfF3YkwGq9JRuy+q/bSCD0n6b
P3Kup8rNJqzaXq7g8JOgAo8DPVPuHnHzO/n8VIwOlGZGzlqjKsMHs9pJ3f9DjALwNWYmUfQPSM3V
P7eUf56nN0qjQqx9LTtLkATugJ1ovJF3ntxRkIAgIeE3lrPOS0SM3tjeRZkIBHZhT3oiznLzC8BM
WKr2dOXGtOeT57/4cskEdMiW+Kww14pnDVA7iUuO2/sMTuQnHW2zgT83rA7TPsjrhB/1+WjkqC5i
YWwFASlgH6zBe5TxRQ2vW6zF0RMj/YoYfY+CV4Gzx9fCaOQc7EJVq1hcnDcVzcM8eZx/D4vF90Z8
ruRJolShsTTyOKAgJKTYDckwXYNl56nYETK2YcqKy5rYlMf2s0b1e/Ael4O6V6vGwLeLAp2MivMx
SxtV7Pamntd20OsLIBEz5QSUydk+4vOK468tRq9AAeZbibnvPW4OIkeTZL6VcrEKCcN5KdCWtfqQ
L3lEaoPaK+lvE2M/81yZJXEt2mqNTYzmHHVZixMsYKuFL8pMJYHTp4Vpip9veG0P6e5AfoYDqXUh
vo/6SEb7CO7sOJ5RcDizMb2mAajnVHW4tnE1zqRsPGes64Ud+ja/a9zWKRgJJhtgtHLgpg7pvg+G
bHCYX3q87jbM2Icnbh8AhUPsABlyK2TK8hxe2Oa5/OJwlaSn1nHZ9x+vf4AsCIh1ygTnkSrnPZWz
t7UWlPL/SZwudJjkQy0fdUvGBSYZUjJEzO/Z/6KbrWLpyYCGscWTikeW+AzQCLpcf0y1nqkV4zKR
a31uA9MxrlOGfkFVYi7egLp5iRgNNeBZY+tZYfaC4TLX1l5EZEztYj6W/AUpM+ml74fQu7984OUA
n9END8Vkl9mZZZP27ivjjy3/LOelV/MZSxJUMUnHdH0dr7w+rcbmdBusAC4GTVTZ8YgviEdnSIsI
NJiatCZr26mKTPnPrlpklGmDWDW4mHGb0AglQVEt3TZrFDI+zisn2trbtbG/P8A0aK9uzJzt4u4r
c6Fs2uB8EXxsFDUjXV+xF+r0r9wU4eJSWYHXo+xP61xkNdbv+mvoZHL+PueSVLnCYhwjyPwyACvY
XobuhzLecUqKGKSrKg3hHIxtDjVUrVE3L7vsTr0u5JHowceXIL33AxFZIykC+ixuGEAtry5S+Ccc
3bk1DB/J3ngmfL9sQ10GY15gh6+2QJHJzg3sH04QceQL5J0uh8eyJYd17j5RCvmjtNfMIQyvhUk1
62M7vKLTAN6y79p4OxI3uJsTRpfJUOAkzHqp1gOM+6X82Iu/9AumP/dX92NJ/NiVR3uapsVzUPgh
sLha5aCHGpVT9Vci0TnoLgzVONLWGVmxRuZ5cjwk+gNxNxNZ7CQNvp9tIvE3OJnn8c+mnZcbqutQ
z7TPfVymbDI9Sqb8rzQSuC8nrU2RoHJNwKGAHbdwed4KnXXu0kEsxfk2VCkP4VcJzgdTXNPUzkCl
77817HFzOJ9vA67xDvkK5T3fwRwYM26s1goZyhTql16xmgWw6HRSXz5U4+ba7Yijc8Cc539bkw5/
lihEmmqcfLxKDXDTpixzHyu4cnwI1mreajeeoyWZg/5pSxjyRhmEDtnYt+0MOJ+dnk+md6FMKqp8
aLcsQSgjcfcEVp8WWMLrHPV4yVrBtvDAx4QMMvRC8fbzeWIEALIBqJrTPtLZqotSPhPLjPv4Zrua
63Hj1v3UacSmGMd3mOPcaWCdbvk3vfGie2NqJQSkzwWpjnOIRWH4kuhzDHVUiW2RgxQmpfcFk+KD
KPFeiIbbfgARzK9RPDczkJ66wGU92J+zmUoegFGGVZJ0bNQNNBKtGfo2FJ6Xp1KpqmoCPFp3ArNW
hxsyE4wPLNhHQvKtczHlzUZgp5QjnaKyl0DtNyUYZfYbX3Zcyl9D8JVxuj8IsgRspMqGOL/pVZDO
I8ZiXeiHyWQZtChfMtjwX7UKXdKgzEucWOd3T2Q43aokih29RiCZHsdgiEAl7efGGwXcnxbxPQBJ
ZLyv2pt2tMmT8BFYoFv1d+niGN3fdD5p1QL2lvmJLWOZodoigjcpUlBJbRchCBf2n+Orp+z/Gd+c
7iAmozx6vgszbzIKWvNaeW05IE/+h/shfYX25NFWWQ4plV1f7QPnux28tOptkDTtpk2VscVEFo7J
GBvGJgTCz9wwLZw/6+tbCIaoOLMt6hHXnAdX69HCRY+IM/dB5jdsHo8ES6ejjsnCE9x0Rsw8m9Tf
uASnHpN1J0FC7ASl4cTUW8PWHW5OiaqCpoaQcNOYH6uDXajl4rj4n6NwYWxgy/YGBmVt4V5GUAio
QtVSSQXewnc5iUxRWql86LFHaGCxr5I1Pm7vSAgxG05igaPgzoHEx7QPy/X/PxQmEt1ZfvvPgIzq
TDU6b/KJPCZgzX7J3QgXalO1uLvLERtEleobp+npihjKhtWx52ehGWDvTx5qJiDBJA/MPFdufPlA
IQq9yQgyj08wz8cecz9mMkBXG8XXKyMtaNlN1y6zPcrOu367vm15WxWH4760zsrFt4OiaYCamMU2
FGVXMQuVEwkXtFcJviXvZKCKzI0SBqFCeNkj/UEDZAhaRqKMtD0jILqavONgcW0HpoND4iAawUZF
UTL796jHU81SLzoSpu0JTWVu7xUeJXkGF4vjChFnoS9gnKH4U6m97fJF72h6rTUp7f8bRqWZXolL
9x3BAAnTjgLiMiUrjgmJkqCjTHOf/3GhCSzPxuPsB4qBhn5UNbEmlLheO3j07a9a/ZAnse7GtYyA
M+jYpfVD4AEd5Kh5GsOgHKj3hWchTblY1qUj139WEs039Pt065v9Ula8oxRDM5JbJ1atM8Pat6eV
05gkzeq2fiajr0GEozChM4/4MR3J9I2t9wkeDt5NWE+bjV84DefCsE/111Qd2WK0ggg8m6hKxi8d
IKeGbUZ4hCwiblnFkJd3n3ABFR9Klt3ZWkXYQSEerM4OBLjtaFDWEusKPuqsiSUxAVSWnn2a2BlK
8so2zOsl49fQeHYbVd/cExbafQpirJ+ZYCCL1zdQ6ODtNycXgWDu+lfNb+5lI47cjMGaem6Rq6kN
CPy6sE1j00PnjXhh1eUMVvvTTAxLqIEDlR2pE7xRFtdctAHGNCwCF4RudUXM5m8BbEb3jLG0EsdI
fpLeoqfYyFV7sflbtx+s8qtRTj1PHtjhrvetMPh/TDwiz3DQbzDjGRamUv4gQ1YxKubmI7FBgjv9
2QlcKPWKXfTU/o5LhISwbdl7H78lqStvkCQ1mtpFxUkLpYsAku4fTuuLQcdao4yg6T1ZYT2BN87f
y3ZVnmEvvN1zGu2Vbp9+ccBCU3wK4/NhJq4sewJX0dMY/qEKJ1Jv5nuuBKVxhCo5obAH7R2Di0/u
1GGvoY+hY2wRggds1dH1EztD62vk21odnteNs+gQMDXalMGRTsiCmhpPA67ye8dkwrsZ6Rtf4PSa
2P6TH8d2Rt+v9waYcRmMypKHitTZ99GP8KGEkleySDSQAzWAb3bpu1RY+zfkkIGjni5hrVTOZOQy
e7C91L9Bhr/4wUvoe8MbuSzHoJ1TgK2vNUrsmFv8sqVwgbaDoIVx7DIsiqspr4ESptn1R77RLhas
0IKMFbkDSaj2II8n9DhUDvpooHHjwvvsxc6SiNLbRAuqYmybG+mOOAEvUPGYMbhwJmHXQY1RJV7K
tyOIk6QGPGzPpXyasrJHo6L6Gc3jz6JwSoWKRZDzS4rRx4ePCuOsFGe1Zj3MiDTbnE7Wf05H7FlT
4NtrcvaaB+gJVslSDqeWUFQRgfZSVarXUPnaHDROdVgdY2r78z2Iib3CUC6ES1O8IsX8pkEV9S6o
EAXQPYeME67kSY4mD94ofZd2/1t/wVyXkgbD4hCCVKgiZS2rR/p5hlh9DM/YfvQ+0kk+VDazMB4K
VaS8X1gGdLj4eC8gkpEasMMUaZGfoY7cbx5UTHNRKfV9WLAt7MYLC7anmovS9iXCdCj/pwJiALhg
UZ3e2x9eUP/OwJw9Q8Wq8f4t1nfwG7n/wYIpH+49/FIdNtjPN2pXTYY4A3tiRB2s4sAAJ7aD0bIp
29K3IXVXI68vVIad0xCZOEKjg1hPPx04PxuJ6EiSDB/HO6gjYix42A0IHe7zRZZvYyHzeSd8VFkc
aDGtPN6+63RWWrXKxumOeM6ZpB2ZcKl0K7Pe3IbR/guBDKYVSmuYavmG5ugbiM3CxVHJ04AxYAAe
uw0MLeh1mpvv665McUut2h37dkaCzW06km9CScS3iDWsNpTX5VW4r2VbKz+i6ZRnpOe+2YV0iOYN
mFml+Q+YdkhuhUdCPOgz/7v3zynYKV5Sg+EfIR54qHinuCxaFQr65ChxpPQ1cpKKVq2pLl2+o7BT
qNL1DfebG+sWUKoq18+VrdGrSkAaDf0GMTmjd7Y12yGktpsmgMw64hakV0Zy/wHWztK2LLQkI9za
u0wGVIouCZPAkilcCOQKNjqG+ICyxEE18IDoSbmgFvug6Dnmr+57AO9STKDz9Bdy7FpUDMJR0ABH
IUbbearmoj8kTdy5H95z8zuxY+FS48XczftHfwGqm8WD/Id0jK1Snx2GdkvVUbjTdp1KlBPv2In+
vY6LHKPo0HiYuFFQDXGq3iRtIiF2ZW8Uc1MzcIEY1MjRLPi+IeSYA+JFKiTfLTB+H9K0aXpNodlI
zI9fMqg9AtB7VrlTE1W3YEyyjPQM4kov+ZqaEI5hRVj+3JkxLJgK0v9fGwiZupQaEkH9GB4J8U9l
85XTES5DCHlEFerAUUButW5bOO05V2raabMeGqYeJsBD4MTWfEL4jcbzuV2fITAwIv1aa4/4vUi4
DVYiOOso0ea6uldKcnEE26LlDWnMn5ZlSivVE9nhbPWVom7qZljJFeQQCXCiCLx5HksfZAMm5Aom
2E699hrt7fTIiaUiUpNIqcZebjTFIeZAEkpby3LcZvvXZpHlLphconZeQZmX+6XvAm6v9lJUL+0h
KqQLWswDkyULVfK7EOOLnw6MnhU8b9ddtBy9Yx/PJqEeFWEG6UvB8sADv/RncTRzO8GGAlsTCqrN
oLj7p8Nasj+qAehWHPmphO+OuNyapOHyPdUFxiC7Ov5ND/Uu2ekMhH45fzKlca4q4s6JggIRzYl+
Gfa+Y8hyL/QTy/cZ3ImfRTYdrsCZzWyaUg/aYn5673rZEh3CJG7diqozEj6vQhe6jsLYVGxBOmql
zwIUGrZu5TvG2qconD9NMz77rpTfBQiMacF/3nDnoog5K+bNkQzhMStrkJ49187URnWHcBzB3PM4
omD72HLQDhvM1ZGvq+xy9/tV/KkbBeYqRYNzYn8qZxW8ippaNHMt3Ec1BWVxgHX1qRE2NOoOKFws
GRkzCg0Al5N9mINA0/jrWa0vyYiKaXNVQskMtzKXviITp+BvWNjYE/ZIXQuG1SgMVZWuVS019pvg
kp3fDU5leIqo9iBjHmuR5VBJnM/8HKDpKx/kBHslDqtDJS6Skf8wRrgz6YlX2JXTQ3SOi6aHcs1+
vV1h+29ssq+ri7UrxDLrUGxwGgRE5aamArKNJF3aSAbabltnAQlJXP9QwrQP07gB6LY95PEIBKIw
kZjI3c0TGUaX/TkhcVAe4c9z5Gkvi0smBlnpNsuJAPR6BFL+B2bf5thmsDAH1vMjNI+RJObYuc4p
drx8E3ex3NzmkZQUdB/v0BM/lE0ffwIhNI8XpqxK7uqDLW25VJ0Qan2y6B/6bOZJj0l9zjPtpllw
vFhwUOZKD7zIO1yMVMpexGzZU9pPs2ItgaTrMJGmucZ5+J5L0wCb3rxvKNoIfBb3utfWKpp0E20f
NUndrN/7wtiMJz4KAhnrlQ9gRd+4JcDEmZkti9mkgxoEcLEeTrgHuYXOTcq89/ySftIJ+WC4zGn2
CUWNcWJHXCC/dad+gLTQBqPH4m6DTq8IrGpghPcJ+MjkHE9OIK1C/BVZBV746CMqejo17zGOzsTZ
1MtexuOgQ0Y9kA9q3VAUYd5Qdjr7cdaq3+mUGNra6V3fl74f6Lqg8Di55A8D0FEBC9oaChlstlgx
ipEejyxdvDXkGt9Was6zDAiekm2TXE7thBwdm6Zy3is5gdm4sIIZT+zg4lbplyPa1X3j33UGM8Nr
SpWjdQd7TUzFqgjvll3UwPRnqrMne0uFXLb1ZSLlCdkqvpiwyaO0dYHWL5y3bljlaGcnLB/VrkWI
N0Fti4BpF0qyzqIoEC+FiwMvZMwcj6T+ApdAcpMKM1ElXlvPkODqInyOkoRP0+GSzh4grSuLbI6c
kvk8zWKCkuFCUyQ4pZJFfuhiDOysKq0J9k7lvDRt7H0OH9ivC+/ZC/48jJze9iZE/ZlNziRm9ucW
GTK5RiKCTDmiVZ+buz+J+E17aBra3CFgiHt6ZumHG1L/WWJwNFIfcn7dnGW/+/tuwl8Cky8V+JdF
o+o6n11EPjsMdE2ItK8kqmJv5iuexzd8h1Kge2jvPBS/Lq5qIz3rgH3XyBSVYcna7W/uCjJ3wD6b
wehgJghThtS/T8xvMLTclqsTPoMlDqAGsnbfWMYyh02zcV5228QUlZ+b8Da7+pC4ZszHVEdQRzIk
QLs48W262rrLUwTXZomUJn917Ys7Fq+tQcFQTGQUFJ+F12Lq0HDcvRPVWnniYfS/nrgg8LInrb8o
9ICpJ7gRUB6b7QXvdTyk6SnYqn27Lv5aRNQxNFGKpzswgRAZNd2gxMSn05tILU1DulgGzjchk4Z1
PaQI3Y7m6GNcN0TJ7KsIg8OsiyntnqrqnfH/JOtSBWUoCiu7rbQmt9bGYktFQ6nkbvBStsqEsROD
VwJ73iepcYxXxsoJveycpTAoa3YO7cbBrELXfjNXQjMXcizIZKCtOOA52lv1y4//xgA6qBJfv8XF
QAwYpIjZ7R6bOz/W2ZUzU44SpuRDfBfV5VMKYr1Z0PKDK4I3hZoaXNoBJP+GBiNtMKpNmz3Rmwpz
kX1RypdJmJDb2tOr0Bw+CyS9AX18mL+awsjJC572SrGounmFaH5o3wsW3EDNrD+obu5FK7M111/Q
u+LfpyM4xUxgMtIW7lKVt8mpoZ7iqdj+YB7Q16ExYKeRWmOLbD0QFF4b4AaxUociEzV6UlKb3Kpu
peqsM2ay2o1fGOGfDzKlAKJQUuWlCRfvF0sdhGPaQVx33H7v6IjVr0aexcITCZyw7QhzwzGAi7qU
J+xwlawWlZTrXl+3inyHMmw9pxfRzmWN6BlcWA1LTLJLjnz5BA7MFMk0gLZbOrYDqTkfaTWTxuTO
kb7lxJenUYMa5bSUeMe2wf91s/6lmqT81zvf0ExGzQVseABKfiL4wVSTmaSMWIygLGeQC3BuWG0N
1C1x1Znq0aKo1OjKxAF6wpZTba734vmvIlHAHQ5h3jGRfmegxVoHP7+p93OmVZVnaM8/s567XPaF
anxmt1WDckEmjnqrRRNJ+97p3P4GtMovuw66cDwbYZFen6r60MxAtk+OMX/5mbjo11cNmk/qZE/M
nrsLlCs1FONveauZDfT+kVMd9cFrAwxFR0EBLsSrcedOoaflhWMEkjOE8N7wTOTfSVVtX/N55pp1
Zvf4Bx+ayaeRxTRfJi6zStC8YryhbEDK/S7Ivt0D/ChvFDaP7Uiv/Ho/zN6C3oGfoJ6aJFD8u289
DsiJovxoKlj+jZHOGXls0/8vnvez6MmffwnksC0yWMMSk56M+db5NY0nW+8iRx1qOH7zm7Y3MCo+
UOjl2oQJCnHQSWEnmRmKpBCssxeuC4D9EPOLm+K481j2YkBmqME6L/cxva7kL3kT1M6jQemw7Qiv
47oPDhgbmQ7napcBHu9VN5R3uOpCf+ySYwwKZXprpPliQnfn5/sgaqwavLchTYnuEyths4GgpC21
WLpTdQrvsSK/Lb6g6piSj4M9AuN+fK7ZvHTkEsZAKXFU+/6ko/xHSc2uvRtmhseLn3+BGBqK8B/I
JJD8asgAj3fma1NTfkFgz+U5hD1SVATqOReLu8NQaof2xQEUiRF5z9odEcuD0yI1temlT4tApod0
LRqHcGle09UJDwyra8Mb2I5tTyr2UgfTAocWl1IKo8YvQaxlf81199O7Ws3DGXk4565KKSYJSNCc
3//RxBrCyLGllOntBIQkLF/41G2rEWOJ43BoBDgh+V9rxXbeCH0Cq1LvXL181oQgX8vRwSHgFIra
UaVAkbIfBRFYsCwozM7WfW2xcEwnrucePQH9uVSlqQJsLrnoRQUHG7QZe0FBpyA2i7Hx4CLJpq5D
jRtXj6xL/2/Oo28tconwx9JR8h8pjuGZOeUWi4DSZQlNw10s3fV1bCgjz7KMO3a7vsn4hfBKaZKu
wp6yyXVF7JCnu1NvJunDP8bhkYv4b7/OhNyEgczcTVF1dok1SYyV/D2GUC47FggPQ9X3eQevKElS
pMW4368NN4qRqQ0KBQEYWNrDg9yZyssetWAmhqyxGWOjhEO9L9CLlDP4EYtWl8H3Mm+AIr3HlJ8Z
3zsJWpeWxTES6zE+4clH6uG1miwDgn3QPIwmE24VEIfFSutbPYyDWofyT9Z5LsfXXoeW+fpW1aQW
LOoeCcvnCTXFt4dD0TJe/9xa5jTX/bVoDg6E2QyQ0wyf3+hFq5hTRjQfJCB6Q+aJfm4oVF5EqoXw
owulZ7Um1IF431mPitdz8Vz0Xz4O0hLROyMELp3FBgFjHIO6AHHouSpfwrfo7+rb861mOVPJebM7
Ze1QWH0EFV5v1dUCDl4fcuSrI2iwuG5gVWz1wvf214oZ2wOd/H0hf4oaw8+qojQ6U915EfDWP8ar
crhyIVhOvslgIMXXP99lfDulQBoo6wPrIHrLy9bAU0mj0YK1NqshyRDx98Q0nZKZ4+OBM1DTtt6U
cuITW3lq6dLo/B2Qldzdenu3YzqD1/aGKBhYJT+yWecEDM1xbSiDk2Z/29ggA5ej8IsWSZFXh0Zq
7Yu/m2ZMlHAD60ihGm5xEk7bq97wZW4GhhM3YE42jh+cIgraGGGhdddzmf7BnM4MVcUfB0MVzR93
BEwrEEY6h7psa99jIPCCidDEa4w27L9jcZNg/sVUGWb8cUtecN0cXmw+yNINrbWtTdF4JqBNNw9b
xkSg9YsbprSl4EC8+Hx2xIDKNvGrzIfNzuesBZFiQDa7HBj6rEPLJso3u+bit5olx1rN57SCpyVt
U4ji1afgonELwDoA0Qt5ONTqxAxxRM6m6MUhIOhhKiDnUKWUNdQzt6IDHeJUketTE29BCSSVNuQA
ayyaZIqtZPisMF820iQl1WQREKji5JKg0X2na7IJe3Ch2Dru0qkmbG4gasW+t+gHBFpf594BXkHe
waCbKP6gyI3+e+/99my/sVYN/K+VjcXd0Ufh9VYPj5LpgqndrymfdjKxksJehWjGHyltN17BrdxD
6Nw/+bHbG0z4SlhZF3a/YX6q4hWKMlAAyvjx8J1AjP+y3y9sdd16Xc8LYQUdqpRKbAc8Memfc+h2
+7TdFMps/RhyPPKGnJl+unReLdRb13dPosP40z/acAtfCLJv7oo3rJdaNW7xzmonJzHr4Q+JURSU
8lF3ky4Sc7Z9RHPOlxCT3XNFUU5riTDUAMYlNjpveZEzADIlUauEuLET0ISUku1Eoxvf6ZqAgH57
DYgEGi9ZN/jAiMFCBBa2NSbM8eoWgGAUu+uwyExBl92EwTIaq6ZRUut/KbLQsD6io07ykRKBY8W4
U4lLmsl3NDIHevR9w6CnoUXCqXoWieUqkKw9DrO7Y1rj83DZX/PMTs/xvP2fRrCaR9YfrXVtjo5X
7dS/8XVAKJKTUo7HfoWpT3GluS0+jpafI1xK1hRhEEkHvvgiRdSbnVXtYqMZ7mWXWOu2bUCPLpVd
ULMTxDGeg0LE+WRLnYLjTNEM2L1rUi+vcxabWEI31qmhZBQGM8FVG0kPCr/yLu0JqcG4QfjQwcB5
yfFN7P6H9v2FLOQjvG2ENB2S5S+W68V/w0rtx7NhVc1za7IdUo7PUb1mLJRiq786dkLgZG6wiApg
oLjFVOYjHIKVNtlJD0MITEA+BGD81SjPhyo0pQqN1qeSnNB5llQwDd05cjdDcK+PLZ29yzvcZDmB
7Z+DfVZS0emnTs48VeXSpCZ/ZfE1jt9fCl5bCA+CpIh4v2HpCXFtZz75Dz+sMpH0JVOhR27vye93
jFU6Ij+T99zRAjT7aMxYHvJbFVKkf2/GqLKGpVD8z1kg4k2CdaDGFK7KL/33zgh/6KSkXRZtIcZ9
Ops6PRj9H3+5IpqlzZIoSkQzmpg09HA62NKPGuiy6IXADBAErthPFG/PvyPmNIHJVgMxoHrzU9sc
2mlEktBDHDTp3YJBC3jQLsOQu9ohKwnhISWaaTIL3oK+c7TXynHle3+sSF5tjCkFmaqz8mbpH72H
PBnjb52gktFbDBUITvQDD5udTmJd3WAx5HmIr+Tinmc+a62j4ZGDivViZsLrw4izccyngeitC8DP
O+Mu/R13e38zBDmXtSXtiQLlYYr2oGv9PNNCZn0yeTn1uIGLKcfmcfoIYaJdLCEp8RgL1iSOHQE0
bGXTrZzZenNtIt98OyN1pJ1oF9QtFQraPn82dnglmtlvXoDippPq/gHysai1a17/aC34G17W8tTC
5rNaP4tyaZyThBY50qDto4lybMPJNWYjaEgdwsKibRUk/EEvQzyiO4XpjMZc3zzQ4dtbqlUFpWIj
nhP+IZ2VWHVg1v8cZNP3FspTwNhqkRwwtp0fumDFi8zSMfbFsyBNSbOtFQwTfDAgLNHSfh9ExOkW
jWQZCgW3Vi+IBT5WlmQvMQ5CWTYm07LivXzSDT17YrQ/XhmXn3285fzn+cZtmFM1qPgiJFSGrv+s
gLzay3Laz5j1tLxuwE2L3Uy0jSbxJGyp1UOAKl/lz8OZwJa0ibh4REdEflWtwQiWkVkIWQG8ZOQn
YSCh6f2FzjQOPmxR2XZvRC7oo0gN6LxNckDblEUn/tt5eDY1l+OaPL1zMybFd/+78vftNUdYWFpT
LWoaCpCeJmXf6R790D63blZQSgq0tBa5Rwi4FqfuA2GGWVjyw6BP1JZGyuvZUbjaOzqTdcfREXwB
JDTN2Co7MkC2aluAJDWIxTMsDzEuK2m4aB4Nd+Mj3GNduLkeBtWRnYjQyge9PrbMvh73gX6b8rVI
hsZfFHavaJhQHXBEH1zeh/0YQoX8k4s1JfHPbaPbUd8mOOSlo5/cmWA+moL5u7nqkEqV9IUtZHZL
KHgyyiYeM+dZVCm2fm6YvBUzCwhvwttcxyZov5W+36Jw7BgRjWSNiO7yWvPSQPaVz//oEyobMFGj
gFIeAdi5sP25AvWhUZyBRdhy4g8JCuZgblcFMF1ok8NEu24RMz4bt779jnI5876Ghda+Fg1hXYpN
4lxUhFzqwyWuAKBPsZHM2N2NAvaX+Qosh+pEO71+4QkV9JdBG2dzH4jMRXL2gv8bLYnSjeHdbRG5
wfYiAZ4gjabFPWz2SAh0yxPVCScY9hkvfCmAq4RwSNBhixHj+sn/O3ga95nUXLnFX3Y2NCasMjjx
p8CRCYPFX6KrjR336HAq4OYByngiKVEtnI26Zcf8a8+mD779wEZbGsrSlNHp99I5qqgHoRqVZJzk
uS5t6e0e2g4tMc+m0kj49B1P6f7JQPP+Skg6yyTu/J6XHga3dNPVmfq86sOJGThHg9CsDoxK0lkL
P/ylmczMZ7uGda4br6eqpdNL/52gKP5XXZThovLoGnV8gS3BpznXJfxZyKzPv8K7fgtjCSGOZ6SO
ndHJGaLR2AhD9v1UjWkNPDRwQjKPubmmwUZnGjSxKVVhDOfdnc+J1vGMXc4TvW1REv3vaCZ3goXC
25SvaqQKxaXPEN3ZQizyB9UWV8uAewp0BLe2KCr/7WGuU978Q/wqM9bYJJjjVprb17fNeud32JTF
g4w6WZa3D6il+1WA+vI9bpsAwt42Gv4KSFsZ2qfT5GUR8n1SONoqgARbyxPhvf/qmciKA2Sr2dmY
KXC+6y+F/0gS7uuz11wlM9cOauy3cXYEbsFMQusLSO4QkRuKMMDjxguHXh80GSFV8NisC467cK1N
fqVb0IrGgaLSAvjyJE6ZfrmLmI/MmUxVWRswZTuJgBH0gjNkGzvahot1u02cYsLywQxg41Q0XUCj
rh5APtG3gs4QdZNuw30itbsgCOBEm3uFdC0QTrCNkfBzGeMEOQjBHu9OtSsCOIh0beQ8NJJVGe/t
lEG0O2m7oVL4OG/TOIB9RvneuDQIAKwo7MJe2sinC+JqeV6H0Xqmp3zs3mrNC9gRbgZDEZOlExYp
5Jo9zoQ8k+sGGPrYQoVCKwFlHlv+wpyHv807P8raP+U69zkhbI7XEAEHYdr7j0Z51CZJupKh2/Iv
wMo6VeGie4k7Br/LXWc+rF2nX+9Ir5U8zzmAQytJPEhxk2xi/y92OiFoZLUqiFo7HwMKi+XfinAu
eljeH1vkEn0sq0dweOXkCGNDNFISyHOB4OAsHjaWrMWj5Uh2J5GdE2vRDkLBs0t8Dm5nkP6jlNH6
8s5jwTVpxFYEuu1mv763/akTv7yNe4ch3iMxWUHrWSctRJAhMXrlUAQdqJNLIWW2gYJnPNGKMOTI
dG19PWUH/2MuSaVbI6jceVivE0gJwZrZnsm2vvpc3VLhyTxbai2+s1XhIOEQFsTLbrfJb+Ea1xst
+CEmo4Yk3ONdH+5lXjqMMoueYWKYGiDptJVDrrL4Z2u6vGGkPF9HveuqioicwUjVDP76zvTBUQ8w
ZS9RfgBI4X03db7qpoVIaJ0GsU3Naz37U59RErsGsSD8cDbgSZ1MCTZ7ZDK5lvCO3Qlg2d2OVY3a
fWcdQChufx+RGFjDOf54VwyyaqyDK80xFFAK5Mzaz1o/EhVi0AI3QVIFwNCn/N9uZnUtsO5dRG37
DzepLk24WDtR3wizmFta0mxQgnQQI6dlrenvR83HCBfP5QbDTZIJmmbaNl9eFklFdZTuYvMLlbl7
x3cnAIfX68ZZKwv+8EPdB60+tdYKzi7VL9v8MnHZp8zu3vie5num24gnfoopi1Ovadup/RptxJzU
rVlVFCUJaPZDcz8G4h/Dw7uZ5uzJwAXmj6MrtRwXcVFvXpCc4WK0Ti+Nwb9MZ8acDU9Uytf7X2OA
dpXUCinuHU64YY3GzfWyPb3cfXZIpxkTlySdAPw2xKRvv/Hh4AOGBjWj+zIomIa3Ta+UNst7uhoU
LaYbqm7hQhhTkeK6kGZTedmBY0gjfDXQeoeo80SvoZ7GKU4N0BwT2w6iL+eH1jJdnGc/dZI6/RhD
kpH9oVhyBI46EX5x6v8khGeF/a3FN/b2nPe+ziIKdmv+cLvyfTnvc2Oj5+e04UleyQc+uiKbOmuJ
vyZWQf0mFCXZu0snP6xb3APrmTDcyOp5ySYgvGABHNRoFGvuugY2Vc2s65qMmcze7eGSJYLvky7Y
cDIZEy/E5hM4FmqtI0FS1AihrFJulHR5QL2g/kgmd3eGcMBMemq97PHcJs+mVDoQpncRcbQ7jSXx
aW0I1btP/MmQLOGHCEIHzLy1GdhaudZKLlrZWCjdeW3CNAu0WmOTF/gtxVQ0Ru0tKmGhmiSTGzZU
ZMyCAzeRB3ZAvsxhsOnXPAgvYYH5qax+SlYeZi+qe3iVE4aSK1bRCVR4XEL9NAef/ZYejmzupQyp
YQWO5lnAcHiEkQEzYrAIec9YhWUnUztDhBzxG32pdf2zlF+H/Z9nyAU1/eBd2Qn0RUVH6qrS+eKU
V1ZE6JWeqgLhX5uiO6Uqfp0A3qaPv0WXx9WHdpg4rTHjS8YhZs6PQ7NKFZyPJVGr2EbXrRL7f0Vk
iyJS77mNey53MNUqypy+q21buhDFaoGkgx/VHDCkuGwDGNL7cLiC58MZYvCi7DziEJdtbgxpjYnt
AzQW1R5h3h+62QU3hApc34rHe8bfi+183FS9c4tuWRdAEcDL1DQF7728T3bkvi7ZFNZtJTGjmoHV
aTpD3VtSxWTk9HqDqBx+pH9DATCzP4HjDznupGKp7mo/PBlloZKlae6t//GlEHQZJZA4n/CkvMGw
7voVhgIReSE0mB0mdLuQxesWdTD5qr25/2z+uMaSE7snoLy1PYMdeR0wAg7bqs497RK4cM+B/EpK
r/tg2MHeSiWpkKIUPsATXygD2vJyecBFfgfmD/KT/Byz9/FhgkXUL60RYowxDZRrS6CvFu/Ic6Cl
n9ADP7BxKz9zZIBLTy0TgdHKdHPNgYyayEOKMSZYSvsfJzh/ImMTcvHKiQYABH6PKIddwJK+PDgp
LfjZ5uNbcZagQdJOS3bdPL/sOJEqh3Y1V9zVVm5ERDs9jal6fz1adTB/r3NxYSfzGPZcDBO6lxSj
28ZjKx5xPkI2DIPenD9wrJcv4icC9cejbWfnKA+3JWrVXExmJqfOCph5x2l7yQgCaMxu9KS39GsJ
0VNilzJkSrNu1ttq97eqUyTSGNP4QjOqY0aj3Ypr5tZucvnf5Q8SfcJ8j3CpDd3CIaHA1dL4u7lO
UoQ6//lA+leQK+w5FcTr834sIab1qW7lBmqtSgI3HwqaTVRPD7avLpWrUIEgzCyHF4NNmkAimHux
BkAkaqZ4MIPfZ0oyGoe3KJftPZhsez0WiUoR0XSyyyfkzK6cZFFoKR9lf7YMY2ltntGcYnCV+L1z
ImZ6sQOTKZzs+DqvtXqdY8tdC93Xgtw12L//Mbko7V5u3+dT5UCugGcH4a000gISRXFyMm5FC6K/
siNrBAaxm4Qgm9Ct2ZoLF6ikoimq3OfuqZIaDs4wvKyGY0nZi49xhcgfP3JqHTkSQEURiZjIEx9d
O9Woe0eqq5wyYzPsuKG5KDEDIzTv/7E2c9RziE4OHOasFJTrci9PsvlogEWGiQaKhJ7YUqRLXBf1
bL/EybJ+vpj4m597EHFM9DTjm3LIuKUYEXCl25NXAXe1D1tLPfA5szwTTVaXs0BifZuqW12/vTpv
PBNqWYY5ahhiK8qY3ZdeDtS3c2An4OJUbbVwAOGueQWBvlWWpxdQtJ1KSr4FxheptixYrcxZU1XF
r0p3rJ60bzkIKuyfwc8z47OVrEVCXPN9i/KKvRcF1jkpjq5/m5jKg1Z+fIokjGVm4h3LiFpGZUq0
5Feg80K6mjxYhnEHiw1lqYaktE8gpm3sG7Q0E7XQaOb94AGtmvy+u1mtXu116SoJdMReDPiwvJgw
+PrxYymKUQCoY2Uxy6lbiRv2/hj5tLEw4kozyM3wrlo4kyCYaF/NAItO/9UY3aGILUhTKVyR8GbY
wQz9W8dXyQLfUVU4tSW7CMd/euRMbZXf1KBFo7SDJLAkfD3zpml/QW8xnl8QofOKXJB4oZ6qLl2B
5DAMcukL7QFuJk2BJaWdhqWGd5wT++3iqLpl5/u/qZRQD2ZYHOb3u4ZkoZRZTYSnLE6pcq6ZQo3c
kX7EWG5wqoe40bqnvwMstkT/6o3hfg5ikcyryKmlUEUywoX6EX8ymmsHFGQ8ZjSbzxnzJ7rEYeRz
My+priMY+77pWSguex+EKbN39UYDsIl44S2KHNHZDa9gLgA4sjpkUtURf/h93hHv2ui5epUNPyRm
LZRbRprtd2rTOln98J6fjlG4LmXaX2+wTnzLN7HpwgLTW3TeSQzAeccX9yeUgz7WfPqurYrZ5YeC
yB9OMSw7lghB18GdBXXTTbhmMOw/p+VIqTiBzQboH0FNeRVRz7VNxZWC3vYEDels7AG+vECuiGzd
LOp9iJRCb29J8yryjpFN7PldpbhcZ21CJdRbEyNAqxJk75XigH6IMT6PbXJNyjARlSjHej1A8cfQ
2K74AxTQ0biGOwhBnKzl1OF/VuVIiOK/5u1rR7eT+uTrDTRJq+rcMvtTkYED+93ehGvQSbhwunpC
IOVG/poqfrMcXWWoegOBR2II5QwuFbMYwd/X4q/JCpy3eNjdLmz/cheD1vA2VjTa0q2zLw2XjxeS
MIpR1LfTyCCxi6olAaYYUkeN36vmh2tZUNLbDcmfnKnPYWBxwkNqPP8IiRHVGl3g3wmY9Irg0OAX
JR/XGiE1Ykdm+sbt9PyHteYIWwXquFTNCD/R8L1CAYceFvKJl0F1VUi/zV2N4KuP8Br6D9DMrB0X
/a09wlYtsP3XMLMMLla4BBP/XYolc4e8gjEnYXm9RNLfSSA8bd8AzoeflEV+Kl13kVHM4XtDbZEO
0a31tDURGUB3A1f/mFcwD2PLti8/OzJ2WOd2hLthRB0pH1Ht2P/XSnyZctIZUTnOkqEKn6QJZ+zF
WINDhnLG37XAejEayg6Tgb6xJ+G9SFYCOdxU/QEjGos/6+tGcb6VG+MpezcY5nEIxJ8mh+XUCb0r
TDycoBHtw7ClLKA6ECQzXD6hBV9kmAOdPFJk3gedMRWoW49jm91hKpl0+d5H8FXiyH2iOp41biMZ
bg6EN0zc7F3caLc5xl4Q7XoSwHtIKoVC0+Pm1Z/ounxWZP/N0Y0fzzpV+0JWKeBHvL4AWePf3k8O
GDouT3K0rzADs5cY02nSxuIB3Gh98/5UcQb+B5F7392WYbspKmWi0laBsLLOwRSTkprcX5eyWhwb
mxzFFVysylxUfW6uSj1k7RvVfH8H5oy6FIg2OPduj9HUwylOUrmezqs9+5Yd1D6B1Od4LFEv4qWZ
CRP3NL7s2FRYVgcexArrmwNi+ck5wMnqUZ6NcNB7QMuV/PUt0tF8TbHIDikdrWqKJ6ki126HjZH1
lPM+kbNIkGIuYdyHMgEbUwIJXrjJecg0XGpQ42TVMHQC26kOBNJMNcJtjSYGjsbvot3AWuevYcw9
Ug34+eL3wj/NsW4Qrt/jkmDCCRjnGIeaAAk9b1jUBEDKXLfGNFs35Ux3oCvIELZqANS9ejySByED
pxFDLNJMhnA7inMn1NCpOhnSmq0A6BfZdthrb6v7bEJppx95hSIgQcTLcKbPYRAxFPdt6q5R210b
tDc2csSKz4FY3aDLCdMIX40JwG5gG74pzzib2rdLa+UopCChb5X/tPaYv2xfO/iEFxHdtsT2Xm2E
xiYUqg0wKYHYe6tm+4NOOt1lfkXgWETR2nywgvv5fPfIXDA9tcOB7Kr8EbyUjtxml65PscTGFJ5a
hMyj6fuy6gW33GxO7xWpejNr7yBTA+628cC8WpbPBO0gcmvOiWcvUhCV255U5YG7HWnrX3v/qVPY
rPtUcXdqrmPM8MXYaYjpZBftbJi+zbt/VHKkvLUQDmgc6CFbHyMrz+b5RU1tGFt6xMu7ISIoIrf2
Krqg1DjKLApg25xZ9bwN425SJ81i9iuu5eUGJkmSSz8mvVKcWuQ+wyGgkm1NnYVbqYN0NGXdGPUz
WSDYUJth6uE4GRLvX1aYMXPwngWwKo51Y+jV0ZPRv+u2Y3+mzGjl1MiLFVkjUEUPAw9edQgmAeGw
FIb2hwZjxOA7ZaGJNy9/YdYp6IlBnbqzFQmReGt6idwSUl081WJoxhGfhgM+x5OObptMCaFXgtPV
+meRTqXYUJDTxA29NRQdxL5nx097CnCPoT3x3i72bt1bHaKYGW9jZXCI8M1VwthRJ+zJRZWc0jWL
ZXRQcrBNs+vt0t4lY0bR6nmKRCimzVK+mmnyDfxZngl8WhV3ZDAGluFGnQb0wcJVm1LDNlsbhbin
ZTlJWgYXdSM4v1XPS0U18RZh1sZgTW1tZCtxm6LPFvM6kVdtvoS02vKFxX+RjPhDPmFOluLjoVUU
/RAf5EJ/ajS/ProCu4uup9S2inmxiuxqIluUqkIK/bbWYTerzbSvQBMFpfWy6BY+uPpUPjdhgW5Q
eyNEiuNjc/jQNGGsMll7Wx4SyNHcU6P8p5AtW1W9n2imX2/aoT1B+xXvKD8EA3JbXDBMbM0LGTDV
cYRtQh8JDhN1DFYwTieCt112FgskmsKvUVtulSzR6mIXigBFItPq1OQEPOzlmogqjveu003CAtpc
b0nE/2x47B+yAdqSJL5l2Sky7GakIpzTnRfwDjnYk7cOqbGPed7/Ua8B5QCdQuLCPzdG7UBenDfh
WX37Y7uJxzsrf69CaR8d2CmPXpwjNnylS46Nd7KnKDLOU0F3+Hb4Yq1tqPkYEVxyv2koDMskK+a3
mmeDA51wLILBUA7jHIJ76WsxbooQICeFUG70XpCi1DZKCUtw1OPkAy2bBAL7gTtRXAqQ0SqDJFiU
eiML8haerdpLiW+2gNoyG/c+dP+ActJn+OJm1PP3eSHQBdpKvWBkycG7SviFq2ECWjMsBcLsp9DU
/BbKP5u5ZY3Xb3wPXTKO8WFj4uy842FKVYDIpu9/6Vj19I8uSS7wWoXN2wK4qe6oecyO0ZrYk1Sr
o47Z7gij2OslvJQxokjYEC6lYSvIGBLpzszvzqlmLiHvX9lE1WYR+j6VwLHlV+uWWdcinqMeYZbF
m8ebVAZaZuMKZMY7sJni/5HRil+PXz+WiCXCF7ouJC+LBDF1MSYWwardoWduETHR0RCV3e4cxZgM
Jx8SknXjVFpNFWeOHciUY3m4kr9YTCfNoLR4uxkhJAAjPXghR6geyvoaGFzw+fh8X//SOyTgdXf+
QpDcNZXakaEP7Mxjm+4dfNpzvNYz9YU0CVbyjAaC5EfsqBbmX3ZvRMbBiKmiScFdqG4AcMy72oCR
Mp1MPyS8bc4bETi36vc10r+6PqHMRsaymgCDpyBkyeEsTfZH60Nb4AeQLQ6WuuuTWVkqKURZD+h0
Fj5o5deo9I/kWoMZJAqYbuUGvws4Rwn3ROg2+Q+Yiozx6/F/sQcyNCe4bRBwfjfdW13Dtm+twhBE
JywwLQ6NpBK+YLS86rVCoN+/yKVE7zcJYVOv4BWhHXZSbDc+Jk+Qu0c5/nJhMhL3Ad2AuftlD/kw
IXY2gkTEbE81q1rr95A57duA39dxBX5JSFJVS/ZnOHRSx7nFT2MZWDX2gk29+8L2uFpgAWcgLG0p
QovmD+9wVdcfHdj34xk9vBrHHDJLJ9zybcXdtxVkTmdFYVd9DZXnbQbmabpnp5D0xCjo5tIMiO9Y
dIDIofBKgzlQbKQw6Fpsfp8VmtQ+Y1XSuMx6Uo4HXZ90PAZSPKwjlKqG7cMgqB91cnxcjHfbC0sg
Rc9DpwxOTj/H4tdVzW1fAcCsssPzvuXqPZOw9NA6cxSBXK+RrF27EGYSm1ZllCoqhdQgd+4yoNe7
jbE2eG6EUc5ElmxFiWBYZ9b5ieRjZCXTXZUDh/SIClZ5DGdh1H0dmNKDAAgvKf6aQx8AaL6tKzNI
/t+KUZsPwBsaPliOuVq7J1NdrxBHt4Ad5VdgptIHEf8KtxS7ALbE0977Wu0R+dHmOKiAT6f1dP+A
lrwrE5dAqWMeJvA8mooo7Hh4H7szBzEQ+UdXxfnFRKgnkJPhwGhqVNiYsWrYH5QsoNISTTLcz0bf
nzH1tIt/Fq0dKR3oiWVIxOMqdT+9n9bj8Mn/whCKikxN8D6AsVrl91AtgLgS7c3e5mZAwdaB0VvK
aEjnQVxnrnLtjGrcHQ2rqhIgSVhNbTHBfS1Ez/DxAYTGCBfvB5gTlOXTc4wQtlMV1mupbX15p/7h
/Fq1LrdQj9TnofNnw/4KY5IUp3P5iw6DZrC7FHh/T1C8NvEYj7TwlOXU0QpTTRehH1/NAgQyvzGU
6480xuKttHffq7r4BEJ7kE44OOfXVKrXg+NEPeCreUjM6RvAJ+/OIGXKFBaCKBYKDIj3tm8yvKnt
e2Wq8A/URxVrCAhZdObXsqkAq8BojWuzuSKGxVZcbgsoQjrshNE15Su3cU46FMVyF1c1vOd95vwb
HZBMxR5FC2WNPBWmzdMfpZos0AlyT5brK/bkYBT2svtVKLEvllfOa5+SK9uud4nkMY70zgBAvKE8
/yFIg/6Me82SVwzpW7AW+HlLGCLdYKNC1OCPSim5IBHLExgOTYSVyfncDAEMLN7rY5WFlUXp41Uu
dqJwX6NRJHIJCKlpgcggCc3tOQ25VSvb9/LzwqA4ALAsuc5Pkn+TX7sMOpe+9oPUqRyr3tw8/mpa
IHQhMbI+o52/Bi3zNaxo3owC/KRthhhoMvhTKh6WigCU/QL2JedMO427GAuWc5W932jp/rLueJdU
Rb11xZ1XDw620bHET2K2ELAtA5v02olNgKeRv1fQnU91WPDHGS5f57M8c6549PuLjOJwooJIIrHS
odtcnUdMWqFS/vtWC1GnqWEbjcGtlzJFL636jhZ2AT882ndSWXOa8Y7xwT0aUk0xfV6Ress9/ue4
nn7gRrf2aoavQVWaZUehwv2uHNoKiir5QO2WoMgOi27CqkHjjU/lZJNNVbs9WOQY28wU7hyNJ/JN
jWo8Id3C2XVIfpZTvca8ki9Jb8Ks3YBU5IYzdJlNesXmQGZgxq5u38AHxdswD1WdiB9FILGOOLPY
4FlwL1KWLGTeq2TFTMnKDTbwzSOvrRKarC3Zv8mAVMKUtdaKNPELyTx57K28Rh5yoSTMgXnoVqyn
XNNWnQjLhzKJNoneTVeT4+ZXWsQUnBYzCDmMHLhSdz2z4Uthm4RGCPG+D9gCeyjL/rIKwuKx/AJj
L9zPeYCE69B4nMH7dCwQeeOuC8+jOwuIxRGKwCHnxJ0BAeGCCBEvjBdfGUj/VD8bfkTLsSNAKvRQ
nnxI7ILFmApwWblxoeibylzVWhjjEKWFs1eGEwCxfNeTLOlTKrfRcu1qse4jQJkM9thbJHo+dwcX
vJw2y7isFSOjIuwLnPfYgGP+UfQsk20UUDqAAnrjyDpjznvJBjZXO8gZ6msz765EHqGE9o353Rda
O2t1fCutcakUTBmnMSvzi8PkhsKRO9FddULd+yYih2IWyTE8v/OLrsPmS9Tk23UoT5bmc4Zq3ww4
9Gamg18ZxNz6drSxugqFRrpxUiOODAGn4sNBGhjpdvA0mBmrzaI9I3TNCDUvnLHIMg8tniSuk6zU
UQwbuDJqmm67RJpga3hU1ic6x6L/vhsaozGatWY5XOG4WG+CPM9JbRgePTroFt5pMY0T9dfhVQjw
ypTKYz8eeyZXnDmXIKjF7zTOGPeLuoOw4x8bEy9EZXUu/axQHozsQ/1BshFa6K9M9Rf1Z2DkUB7q
WEFO3ao5fC2A1TM7MVgQs5L2gpmEZRm91KyC0zek2F9ZM+3p6xKeczYYAeIQ8uPRwLVL+dMx4kQD
pGzEVIaTmDjlPaDSrvR7OBM8foRMzaQzgGRuy3sgHUU38dUJOsy2UQ/rzIw0yNkSQKlGHyAMRWHo
i5Mfi2iepuajL3gwQcm0s0cfECTwaK6nzsSFFXFJiiy56ZH5dB11eciAAMlPfIG/48RNyoFtQCGl
Iq082oFEekZNyF9TP6t+LWFpuIa+U01ShTR/YADS3VXHvnRirDRy6lictmZHyU67Ac6o/gEJNYUv
OZ+K2wWgQ1Q3RLbWlxo4vKsStxRjCo0pZXfm3OvEQh3pRskf7zZzXi5gUEIjVlKBnWXbzMZkIa6x
ZdEtep4nrx/WAXYNCMA3v8dWTPFDz9tFnQND1cF2uaI6QE+IC+P9MRN0Mt/WyaFLlSy/IQE5vRuT
duJLiPIE2tgOreMtfn4Z+jGzFSJ3KEenjwbL0j9Igumlhl5d0IG0TxQ9yrDooZcegWfopWemb1/Z
+8Zo7P06XCmTJbZHVAZ0phNCvBbIFPKshHdUf2nqCFwlZBercmjm+51iWMS8ypM0Drv49Y9z6+Bk
o1XySOVALhJw094fS8kIaReQJgxXQ2/kSfB9zs/FV/Kzp0DNr7QUZsIQRG3jCSHv2qnyAVL53XQY
yiGd3JrQqc1uTkH9aF3UIxPFqMidxFgqRR2adNSigRV6Y+zT6J7+swYNp6nnwFMTA9Cg/UCpQ3sE
XjXX95tt6V9ljgSK/VNrxPB1hUYmOcw9IiuEcpcRxGuQIPae8rH4HIo1i57CzurUDm9i5X0oRT3M
XZ+jBNgbxGufyoDNZWFxuxCXhc4LIvV+BCP0nj2JyEnCNDy0Bkcz24HKj90lY+3eGhqrNZ2XeaBz
ovLKewN10KRaSJ9zITvqjnTCGgPih2GjIll/hC3vxRS3p3RXgQRbAjO26MARB0mPramBbq27Nsq/
O/yl5fozxpuE1kR55WruBJAYzUxQWik1WfZzCXwZHiYbPD+ErscfYwcXje3hDxMVOI6H/CqU6bZw
aJnKNfE7wsVuAFMepcPUh5wwODyAfxsFYYPO3algDOGZgUEDw3D6QUsE8jbSAvUs+8wujUKHl438
BxabPfTWvGbhbsW8G7QibB9b+Wwh8i9v6ttY20Ov65dtG9+lwwsC4LQsBR+ssLqT2lvPM9zAQKZT
tNVobK1kmGYuZHDc/g6TFVCwrkZURObTqSALAkgn35I++M2QEOau/KAdFtZcqCYbIZq8aSVkoH/D
9dFsH+Tdat+cdWAAb4whdY30DtM90yVz/9jzx9EH0L+dGXtk9/ts2xetKGmLzkpnxxEkTp7WJ0FG
0U0NQNTB+g/wi0H9Cjv+RpnzdcoktyrDPtmsx9Tm5MIpvqDnezQUoxatm/I7U1MRiwF261XLS7lF
xhv3/BUZljLBb79vgL/FbUr2lsERqc0G5cvKSbVXWYIUYk0s/Nfp3KpnMofnS9JcNRqzCKSO2/ds
bJMWixmnFfE419BOroWVnChgy5lnN1LQcbEzNerFEymaMgeXe98DBi7Xlu8XMaeIDwuvHOeQeBVb
CKTG0ufOvDjBh0SaIzJY/bLGycAn2sajSNQaoPWasD7KZ1HJNEyJgWkP9lsqmI8L/yzWFtsN0iA/
+kWV1eTlIRSBt1oOBF46BrzXeq9ug+iAOjVqBrcDUJ/9vZv08IistxdasazeRjxjOiekgHRBBTI3
jxJr0w6XkHTJgmW5g/WGXg4/OtmXPjukGlJ3O98rkfo4BakLTRBT4UbjZQlcreQpeIVWGtGHCsts
8uk9OYCIh5wYKwp37CHLg79Zxy0YaAUngx882B0ig3nXBpLPFGiU1GEEnTF0PFsSsx6SUHSrEbDS
KZvHRCn+QmM4y6jAYtUfeeDLlfGQFNHZtCnXZ+JLAUSUplwSO4rfPq6Enm0WuIVWKoDhAZr8qXOJ
nDZxDRlevFKUWOtBgkndpyNQfx16mVOmRZfIl7n8pPcrlU/CDMxB5k8FiJwkGy5Fh3AeOOhJ8ek/
Mv3D9N3hsZeLdcQYyGhxg01nQN+26y56CoJqObHU9WBUc20iD5TQ1WGcEVHiuEa+8GHfZ7tLavTY
Q98UtyyMzOZu61k3L1BUcicYWGd1XNufO5elmM4fI8ay8YEKMT9ctdex2DRgD082dP+WSUxS3zJD
YGAN5atCxDNvc24rE+c3O0p4oqF2DncQKZyl/S2dumVQwZkT2SbLk3pLDgJVTg+da9iv/MPcRaCa
qh/Z01B1lRD1zJevjEAPRhyUeA7in89YAUZ1KR2btc5DBVEK10IU7190B1WOqsWLY4P7pfr5vAjo
iCyz6AhNgtmftU57B4YzcwOn1aZG1y7cE4g+h/hEGlDbEE1tVCLilBbFNmAqYL1fipE4M2Pm4mf7
9pSJNyEX4ZUtWSksEhGS42/YtPwutuok6Xo61Fg31SOQK5CDW2u/GJXalILsbeGAbMjfzISv6yeQ
y0IJIvY3KGKElbuQ5rCLaRW90gYOz5PyLtr7B2y5qiSa1gq07VTLtRelUzLAtSIbX1FqLhIgC7x4
a6N9wY1a4VNn1Z9Euj6k7y6bK1xxh3F044PBgmwNEyhU41JYuvBaJE76EmDSw8F9iScGWh+zqztK
WgxR6xM8RqJP4txGcMMmUZd836dwTy8ahbvdlC6sbUBTL8j3OAueNI6GC4ERlkIIQEYQlvWsjEPs
VZJjoLVokl+zN0aDRqsRQBCJR6BlLEWIia13aekblGdJMVcrDrrxvn2cH6PIZO8ed4Xw5e/iwYZS
/AbwWk0ldIF4TNwnAFXGKgju9/ja32lDJi5yW2YzAttSJ54/J+ksajHwuWoj2hkG8bE+3ogsoafH
mEn/HrzFgZGLJHZHVYZ6T+mSTcgWbbdqf7cnKfp6S/YfT0izNZVPt66wg/9PQqD6/3X77lotV6lx
fIHFHWyWCmDpmmk0FTna6ULAXX/YTqBw+OLm2yFuaZw1DQ9cnv9utwvaGuOaHStKmuF0pRdKwXcw
77EI7ES648v+SddlvJ0fHMcowl7kYSysUjogWD5q812a12HEb5UN/N7aMn3VW+42jWzHDDol98iv
AuZeNbTkS1heJ6ESqU+0SgI5rthxmmt9QWJ+iDnfmMISX+3atBlayHv8486LwRbu4MF6e1FSZ+DH
PcnTK6hgt0I0W59T1EtPq+QItPV2MvJMicWSbit5WM0bHvLniQEAHa9uK1Bz9DVcO9Unlc79L7a/
gX8k7A1vTQgKm/dsVQmM7obw7wtsaGOFLuHXESvgY2XlBGjH91k7hElW2FuUQLrjp6go7BVcwZGU
PBwrJSlBa9eiQ2fjn2ARiYnlWRgbF8JxUU7FxBSDHGlc5tesOXZogh/sOEk8tlXkI2X5huskt1Op
HKrx0WVRR5GIItbvel/JG544WfB43j6zyuUcpr7kxVJmiidv3YPy3q1hD2fPHSVwaZz4DmUtyWKD
ZKcxX5XR2guzLFEMN1FOE4qXmVp0eVAo1Qolo7SnMd6k0O56gEg8Gma983jJenTdClEbSbU3XI0K
FHlTA30kUT4xti0tZHlbn72rF53xNUFxwLuu4TMFsNA1Fpq4pUizIRygRgGE/beE+xOTEydzBGhK
DL/fmEg++82XJMHMChidpqrO9ezQzrFNyG6zTNJSTq6k+d98mpZCy7uT7ZNI8o0m44WuT3fp1VFW
ZYqXgDcGV7Qpq11CoBH6mMec8bNyZn9C8nPQtEezu23TNdOeLrLVIh/+m2BkMWK71ZrUHN1QGnq0
2FCDX6OmiKpshgPjN/8p9ApXJvrV4Q27Fo2vgFMkjRVqva4CH/+/BsSKWzkZi5QgMSbvA9gwYRaL
BRlTJBsMj6B85oWScAFzct8ArR4rI4quVLoGiZuHmeDvzmWAoADK5cprF9TH4awwFE8AP3HPo//F
JGeZNNa3HO87i1tOVB5z3PQQ7AYdI5FRI+/qDErkZfGpc178/cnW0ibHGZO88BLvXtXz8SfGLweS
ymRLvqNB17tuSVT/yZzFIlGQjs7BJ7hDCEHKRPju/RVHhG8vxUHIjCt134MssDC4ddqpCq9+/ocJ
cfyvGu/A6PIUCvvHp6mnPmKhALaT1vxpu0TIiEcNjy398PJu7NdZk6MkepGyCPm9dT6E7E1ba1XY
998ailuUOZeSFuOmdgSqj9Fu31fpNdMts+jZCp1EAWNQ4FgEouiFnMiLPWmhEzBdtjz03ZkS9O8+
0cFdNMeYr3Vb6SvbuFixpL9VXNodCpx/cd30shyvpqADBk8hbcc+4MD3nARpODZTwIbKNMVG4vGE
nw6NVNhtqwoxkUY1BO4+PprfgzEupwDIGnUP/L+eXNmHUZdCFmjgio9SaDr5/lcSGy88+hZNGSzV
728ptkKt0vc9JD23qXvkvGg9tAN+3qLSLtmO0HqB66q2tje3npm6WGWUt2zQ5lXwiVFRbKXCDHhS
GwV6IhPMg2x0/yhKRbvJ5uOJS4jPxrg2wSDtrSxncdgr2WopjgZ0z5uje1FZxKGEdHyB18xcDcBd
JyuAfWRnCL7Ck+7P3xqh5UBDXwDtmzNuFd+GVx3HHIjnhyRfIzSMteoPY7EwgSx62SLLqHv8Fj5D
SP569sldyshfnOYxxOyzYuWGNeJQ7Zl8TOAzH4YzAVerrAQYnBKAiJhpA+gEFmz3A3/2XqhWUnxg
SHfM7U9PrZE8ZFu5eBN9u9r0AArE3X4AY4F9KH+P3bQU2w/h2lwHGHHH0MCisLCZulm3GYqx4fid
cKcKqepsX4DBfo4l2Uq1JnqwDkVAyzmRvS1tO3SU74ModpYg32IfEuBMZIMPFqhDRA6Xvl/aBO/O
JkN/t172JBbGc8g2JHJlB/RS8mp3Icw9kL1eGVADHWxps/crvlHfelZMTnMGp8ee+5cVR4SOK6pd
SGHbPy5qrOao2wRB5upJCQZ5IFP/e9usfybFWgRKySxLjHXiz9sI5uaoHXS/thEMHAS6ZfS22Pdf
rsezuQgLYPEE7IrQsNfYzooieiBaPdfnsB0h1EiJlXD0/jCf/MaQ7KYNd9GGagcxqWsspDmkHGQX
JazbEKLb1OP20jOWzXtNowNKZCWaYazLDk3f7t5418lMzj+3EjYb+DwVciwiYXVKAfXQhYhlemhn
Wqcu1mz8rYDMV34+Orbo4SvqtPuobUG8b0u6ju2AJ4gdDbCh+92gqIQnzWExrol49Lk7YoUpVeF7
a2zJRhBNdC1IcT/O1w5fM4l0wqQHFROeXlHEzOem6UT+X7sGnBeXUiDDTedmojwVJkCo0x84J6rU
MHgTYwmdVgP9VHI+1VRrYgkfZTQTuhalCZKjy4Tt/2K7Yqftolh9UR/TiBLHPzivyNl7my+bhX+t
koB1PD5XAKsRTbu5+jyx4pmNOdQ0qLS5j7J3Rerv3N+8ITnKD4YMTIk3BgJlTYWGg1VIEFFhhedP
6HzhvJbHD1uP/R2RJspXZ0pp5MG5LE21BeppaeO50/dQfM3vF3R3QuNZhiXgRbMGKB7ztwtZsGJR
tZ7oT5HlbbxRXE8EDnz2Y7y5SCwI1vQ18OyRvbJZ1vra09hA9HrkDNHygF98laeEr0MAXY0zoVaF
l9aAoqGldz+SSnUnVRJ1jp9vY1YzeTLFBwr1QKt05Fn7TNPRr3iCyn6HuitQQOkDGY339dIEEyWj
RlJEgGlKB7U5MQRV3UDl5ZpQ2Q8Hz9bDUwHGu2+1fB0mHrShMgAmHL2OofyArlwHVVa3vj3jKEEZ
Kln8DIa+xPgk3enx8CF7umMupYurgpm8eEDHQVtbwNrU3bQ2rrqUgz3ACGCGLSPOzXECowl2CTy6
hIykPbhNVYGJH5ZoAOZHm/oJa18LtjBBRLG4fO5DvPfwEytI5UN627iJMmZ3C82k+IrKpi4qR4yB
V0slzyiZDryKDglhMJ1lAOzK31QJu+r1ZoxUDfAPClFF5uAtd/T3j0NZEeJlZ+vrqljQD400U/dz
cB3bzMx2uaZDHza1SROca2UQ6dAt0x+wgNMIG/toobbvabC7QoMm/niY+khE55UIfehadpeWdrrz
CHaY7GixfhafSj0uQl8K0ADHqP29fW6F7Benuzdu4l7bIm0TW0rNswYGnIXHSlMX8gzkLHcdHwiq
bagKsgLdCihVVwnJd3dBzisvDOgazNSFrNLTXbQoZNAVP0vOxMJapj4HCUqSi/7c+HrDcf4tYm4y
3/g/t5SVq1aSDHebSBP+6yOy6yDDo1xS3Kjrnj/UYKFdwuk12J6FYwrSJu+qWOoa9xBTDuaCSfxY
hE7cYXy08Nfy8Ehn62zyBfJJnu8v9ZCzNWfbDvMuJK84tSExHCa0M8Oic90ow2HwxAMkI7F2c/iH
RuctbXnNu/C30s9+E+9K2PbzOK2bbNhrwflgkhLQZ/pqnJ3JQhTjHOEOrf48QvAbubEucXth3OeW
oAML2jLTB36dZbDdG0z3KiDADyzIG39wsAX6IHe8vAp7TzQT1s0HoNkPqlQGm95fWfsnhvTAv14o
uIJ75LiYC1DIjSVS7BH7yF4x5E6j2OmTVH3cnWtlwLGpd3cKJOOFeFVmR2nJ2LH0a//i88K6zR1W
eBOVdjAoJYLkyceJbCj8i90fNn0QRLvEV9JcP7psEUS1Rce+Tx4JSoCLpjdDHvVkPn1c9Zqjt4KL
xUc7G0mi5RBGrr924SqzhL0ggWUWxScvkSZoQ3suKg5IeqCbi25o1QRb5+YURtCxh40SbkH2eAnB
5KEp23Wd7pHGiDC+FAwZLYqryeFVKNSJq1YmQeURh7P6uUrxYMUCdZ+cO3W9V20ho4PIzYY44EkS
7Qk4FBIjSAWlKlIgG1KE2iZxCD119uNvjjNRLHHJEW4S75gIQO0lmnQtR4SN9djGNN/aR03fph21
FgzkTEN4gaK5SEITvBnb5gDfplCDUNQEDV6xbA+UGQvms6rN7H/YZyhV0kt+ggYt9uRbtj3xCHNd
cxBZB7x5XhCxNPkZ9LNJzj+2RkMcFeeGqWXs/7IzkzyAkRmeIjY+QFuCA2SkuK1x76XVVevG77lK
Grw85mg/oSgBi2XTUOAPp6vqEflH/3E/2i5P4hCjImGdGnldJrtmXUbCJWuJ80rqH0TwNYtUrHHO
aReA6HcfVA7z22+VojjWxkW0NzYKV2HvphrNZhUZMThg86A4yHLWO9z2JIymvhQZkvU0jSmlhixx
vF8cdfspmrMa8j/N9UhJoj5RCPJJx5haMqLVDqtdQhIt1Xg/k4a+Mq0shCoUXd+dOIh9K97/w5Dr
gNn+oO40ietE1zRLLdU9zxh1cGzMTmGY7XpPVK2VG0clZM/TCMFNTj3szc2kQx8y0xVwYemlrptC
7Ynx/bSlwvWaO6bXCDAEVD5RGdTSgROujSL+tm+bFSiOmhl5FZ6Zuap9WTsXXk+FlxfmvGdgqc7q
5Y9g6Nhl4FH5Iz2u3cU6jx/16MA1Lu3QY2NkjwzZ4n8cuIXMQZNTWzBUL5d8UejFegFst28S/5Dp
9uFY7wOOdaEj7QZRAi+0hppZ/rkILnBzG8R4rUuTHh0zccltDxVsDhLTu+BDPkGWc3FSBJIZyhW3
4hOZ4/iKvMjcgx7wNLsKqrB0p9+cyFVnexORh43UPlfeJ78pqhbaaV+WAaDW9SPOchPVsbVHjyuR
xkrz7jxZiPOJ8G1ua4IWiNYSiEbGV9jbBlyr8RZaLNnOTKM86JjNvFHd1ZB2uzUzVGd8i7oFxi/B
pjL2V1w4dtkUj74PxFYBabQytu8Xe85qVjIBF1bFUI9Y8XaOGiQVUScg5GoQdJcgfm9qMoUu7OOE
7AOWpFXDqPwAZp1A6vWGqGBGBa8JZxqbSxNapiNOOLNN077Xf3pUDQAuuMnFIDSUz6xhtWiBZm4M
/JC2Y79Au7j+guFyIyI0TuNxHR1rJ7IZW+OpiN+kYiv78aLqHueO8oPEmvgRU3ACAzHZ6IJyat1H
X0lDRg/Si7m14eTFbSpYgbfTSkQFG/HuP2PEHXPoEWVnSGmLeSmQDCfaDGlqZo9mo1Z5lNpprTOe
nFR2CW/UFTPOsqr4iDOahaue6JuD2NkT/1aDuN28/jTZaT2gFj7Xqy3c8Mkzj90uWoy1D6zKRBI2
pM6eiXYeGvxzqKuDJV2IWpXLYFaTtH8FSkQTNAbXTgdpYmGN6WErD+FlXJg9OXntaRM114DroNZ2
vLOK9JWzdbM/vZL8vfgDPsKFkA4o/35LTvFMhRaM5/xHezMtLue3lPKI74i/07OX0blKUZngAxHB
mE9UOYWJt3Q3qKTXo7BdWwv2xaXnKYmebOtohafuLay+TZALXdy7zUpAxkn2c2bAjV3SqEtZfjGB
NmWryVBZHbeegO+stdl0+AE9pzrdwn1u2lO/0e3NwP3TPHb4aFlLRH7POBn8UUtzLEA8lpFHVwzh
cuUL7llw2VhIiBBB5TI24h+QusYISSczSfaEWR1nc0gGyqVv0KwACnZOQIz8sStIYILfqve3ICbh
rEWM2nbTjFJ+VVb/LaJjqj2cW1DK6JGOUPCf8lyQIyWLcgDTMapCn/8z6IdtxHyuc6JR7JhgHKf6
F3hMGjOvbQn3GLOxDGu2BavdnhAAIMeXEuu0Qn37ZwoBmuOCTZbvboWppvCD8el8amLB/uNW+eSH
tohJG5edp9/NdrkH5aQMjQlL0VMRzAWPtmr1goZA4mIlYcJHsHBVGD2rxj0BEs2WsQrktJndTm/o
Ox62AMOlfianhLaTQOqAtYDKJdoB7bs+YrD5t3pYjBbIB/xmSSz5wgJOwdqA9hCcMWJDdNWwGbId
A9PVhgcX/SZzaOv35xVwc+QCKfiImKr0Vnl1IZoQI7vMa3c+eLjxlRb8lexsFr7QPQ38oFB0nklo
ry0akGPL0/4G5H+Zc7fdQprnJBf4VB2LdDWALu38tjtSGgxH0WBvEjkK3qEU4dKarlgkLinX7VdC
MAcnRMisiwugOsgfMzn4cdwzmXm/AM8FF3fIRikQPqSR6gSDMwRImJDqIw392mveQTxVSmJ0xiwB
7AJRwjLzzI127A+Ca9LjOQEs0sdht26KnuhnEAHdRXo+SUlOLyjRGdieIouOqtPdcn/r4hvXzvVv
zZ5yEq3J5Apj1LCYOk9d7y70nO94hNcDkq3+Vg5E5k1s42XeehRkt0EfCyl+1XNgTzAyBSd82cks
5CqSZhK0NL3Tld5U0QKwHnnkHgbV+0F+KxdiA+dYr2vjQOSHpRZuSw24ZCfHho6QRMFFljK/k9qx
zQQlKaaAfGG0D7SAECWoLvrIHWYvHPNgvTCZF8asySpENCFT7+2t8HKP+YPHXl9vuPDvFJeimQXF
EkHZnchFXKlut6ZsbJuN7UhCjoGRsDkkdrmfy2Yl71tzG7yt3QbY8uJ3njynIw/isifdr5cCrDP5
TIgYyF/DYnGmRnsitwTmdNMhFRGfUuGtgx8d3dze8FFVoV5foj6zstlo3wISLki3RGbMEkzRYit8
byQtVqhRU55mYYutCwqKkzbG/n+6u3z2db9uFlAJW+68kZoqYyojWWFcVk/20wtsQtfoh3witrj3
kkjTRg99va210LJi2VU55lhGss9+zOTQvtemJi+Fw3a6lTeNzpo6HKm/ONKkKdW3k0pSoNUFuFkc
NtRXVeegPLfDSx2II0r9NIf7oEdDfoDU+4AEzFSoTmwxhjBBhCKC+/eOMMCjbF9LvtzYSn8ta9mJ
OBuX2rxSXONybFwRBwsAT8mQtwAwK6tRVCKeqxYRE2+fzAff7+tHLXZO7TLPsZ/Pl2+5eEDrVMS9
qzc/AyC7YYbhk3bjJEWFxhmOx+X2gNZ80l9AZWohUXyDcxkX7zG4O6b8ZYKGUXHN6rrt2n43NJjP
ZjuQrgSrFABOVIpFGxyJS2Vuc/1Jmq5iFoad7TR5Qvf+AnbsAMc+baiYJXXiawq7yEdaQHL8xEr1
0dUCQ6QF3xoGp9y0OjQ8wiH/shI1LJipORj/wM0g8ZYYaTADzeDPZNyquAVuvhfGWJ1LNKr6+x2j
YxjFii/wV+gh6UDrgOOk8qS946xc0N314aqlRBZZbtToweypDCFTLPHLRNw8uo+y28wTxblerbru
hxwxY9liFc4AtKiU9Z85CkseKl1aF82WG6CCu03GXWyPGyZz1IL4f2/IF3SjEb7v5R3B5w4dB/TF
NBqP/sbfNXOY5sb8LGLhsn1r7Q4eySMbLdawXy1e/yS2Eq5NE6hQzMEFteWozUvmLFVWMqZcuXsG
84u/vDFJMVgTsy4eW9aXj5m0swhnnBgMK8fM7GBJ8c8DwEggx/6wziSlHMoPIsUd/XRJ5PWxUs2+
RGophEJxOZXIyyEupD8bTjEZzc2O7lBjlHlaLS6RB7BRKZ8rHr39pcLl9r56HzuacH2x2AvZumPP
trYnKUJihLxRBriLfICIN1+J6fOK6qgfzaqYd/Aik0egabDZP/2pxjWjB3XCiNh/DKBour1kV5hL
A0TSoNqEZM+ZMPQnfipFKftPvyqqM/mTwH9S9zQbKEx0t1UoqeZn5RGNB+Zg+kxjSJfrxEMcRc3v
pLocksxUjgH4QNdhQMSc50Tdhbogg1D6aaLjdWdGoHNMEyiHZ6+eMpmSzcxNN2Pz/o9sQFJb9Dpn
clRnAd2wwTdlAF4sXB0m9G5bBmbFnuYTtO+ogszFFKFFJ022aZEasch6WkVoONywJ29AX1Ges/F5
MtyT5idlQ2TOO4qdClQU7H6C1Goxxo1jq3+jHMib1oqa53HbpLq3cCmNxZXkHEjv54KL1eVRcvgk
nXMcNkfKgt7UAma6K2GGSe57GrW6yJq3BxkSqAGF/4O3+TZ+8IzyFqbwEXM39lKmBRS7DvQkrnFG
OTAVESzxcONJL2hq9AjxUGtFfHe5S80NjkXynTOT24P+HfafF8U3nlUmJKE2Sey3z9VPecaZIhZ/
NVpvzMYuf90XqSWXm6WVFeuQ9cq9ZjCNCPNVj+YnJYqO4/Dk5H1KE0H8bKjmiWFWDk/cv3EkYuur
4BGeXef1ohIB/VJHWUoclPqRByyFM8sUwuZPEmdKUkCgZRZ2ZoH3i9UdjHO3kWUZEMSmovhazRk3
NP5KRhSIxbabrCu64sneTVtgonp+bJIsFGZt/P60o6YimkoQ6vZ08tM1FMFjAqfDIfUGpfMbOqcU
iB0H3OmQGHwOOtFxklfEoOMkfJ9lQzNJYh6ixcvSjDrRUiMRNqjmkW/Sy18Zsymd06hZwFumtu0r
7i5TvRepbpAdvkgpdbTV6xKvvkhUGcQfr3WJn8ZlVB0trMmxbZkHuc3xr4dTDEQBN3b7He1N+dE5
1W74tRzYYLGQ1LdpXqYEpDC8/uXxwMGIDEykm5SqKwAFTLGMQ/gTXPBNUW8dcZLb1xYv626Qv65i
IAfJ3rODd4+eTrcfLxTsbD9tm0WIsCiIq//jk4PFeHN0vXqEiwdF2S/3AbbC65hghl8rLpBmz2/m
uLNJd7cczqUfE9y6ud77NniXn2F3UtmLApJKrARbTxv0SKlXz5/a45WMyF87eHzyIHLkPJHK6oM0
+oaF5o0CqXhLOmkC60ucNSPduzfsEVqw0HhmHLfll/CN7/HESWujezHGaeG+NN1X/1hEl1JFS0lm
+I4ABryMSz2OunddafLZ/CEIvDYDYxzR3tFl69NmYxVEMrpL6ekpEdzpnMUUsAkA6ubSFszznt+m
ATr9fgS8NaOr+fMtidwWQOPYpk5xe3R3OcboxR8/uHqoaL+X8Dl0qC3Qdp67ZubZLzmQM6WCg3jS
k6KZ3yj5/JbHC72mtrOHaJ0Z7SNApTKD7zLTFIIY00cr2PrGe2o6rNWXzjXcrnyNxC8HPLTM4Qnl
oj/NIkBpN4xmKNgEcH3rNyjLjyj5XpNPa0HlN+AmJhDMf7rafzLvrv+65XeNm4GCgH3pXyVe/C8j
QGlzoOKvUatFGegjJqYf0/+/isQMbgYCgE+RuK5hEx3rbN6tRD4t1h0WXMiKeKgxu8cacrNTGpe0
gT3Yp5mfTWErRj1WtSPuDLbqTnu53TJcasv0V7wRrnhXL+kKvGJPblIrcMxUm13Y7a+BgDsVUiSe
5CocgFl7jtPas8QYIIC/HtAzLCSfERheo4ubO8ig0rxLhTLH25ehy7Gc8nG2/jt6qHUx6eHWNhjF
JXyEUHfsUb8qkUtf4I/A1VQ8X7ITtjMaQhoT0CGIg4eujD0UwSFbvWglzsWR+/PKRIJV4McpJhHP
aP2j1+Cf81SlamX5dEOdKT5piQKx973DZCqTM3mCywC4tWzhrZdFDbNw5EKw+wn1+2a9egjliqFq
AoxijmKPS+q39nwWJk6pVSPMn0VOtJ5B2cdAmH0dnCUr7YN/zKFJn7Tx9ptxpwYFcnMAuzBlKtRT
zK+wEIrwIzduLEk8XsW5FJ535BVaLFZ1VGS+UtwCOd7rqI16X7Lc8hX5TtgNLLzsbB9+32f/thFR
RPJVyYA2AWYduS+jHqdTdLKAN2yZVYZ9QgXuJ9qtrbEeqO87zDkHVEyNcLOYJ7iXO7SHCUDOPFy3
RZPFe+ZkUN79smroPYdnLMVQZ31b7QiB2P7DwxiTbkArqnXymZsIddLgj2jQMVLTS/oEY5wS5XJ+
fqFO/5F1DTT/FMkVsuFJSxeFe+FoTi+0b6hDWJ+gqiwYqKcjG3BMJjmILyE9oxFeGpaoTuclLdAe
1LTJqdfw6iRvCy3fStOKzyiVOkNNVbIeWPdPFTzNDGrZQRvlwzK9+DHCFWIF2r5Lp6yY5tMX43DV
AOA85+S75hdZREnTcB7pB8DC65yuiC/FtLEhEKRUsCEppJxnqYoci7Wy6Xnw9D5tdm70WXUmRs8p
Te0EfYuPWhLhSawq3eP408bNFeo1ojzB2CCyM4C9GG9ow0BsePbuc074/oKKO9OXkeLh3eVDXNtf
G8DN6dPqO/zo/c5u+4Q2kQ9BrRY2Q7SG7SpELd+lUoEJ/tcYk/alSNwTVVVCq5nZlJfRumweU1+g
jocGp67y0x9Loa/Nr2KayFkweEZoVVD/R5KZXgXrGPr9DW2zqUsARPOES0NnN9gudfpMf83XkvSw
/MBN5B2GoioygNm+eioWy3i8bs2TNQwE5kR9UEjhDFwN2Ddd8ZainEJ9sLxBOwBBxDf5sT14C/2b
uSFLe739a3RDTKiZ+0hA+8czhKPQj+8W8pYRYXN2fUmaTXeyZ2ZTcQGdp7m8kF9KsoNi8BTCtvRG
+v+i3h3NrBPHaWI7Mbt+26hbyI6Mxs4lOjysD/rtwBnGOf30Rjp79wK0G/dU0iUNP7C+lzWfRgFe
d1BIOblVaZKddZ6vL6WvGlvutt0BSiyyuhkWICySzznd/UtR0fEfDVjcKePtMkKIHgs6OY5htPfw
Me57MRffrrjCTrnVzcECTp5m/p8m2do6C7yF464cFVGUyEz0SptuJs7G3v5vpQC3MneQjtkNUJ0N
ApZZLu2Hraud2Sy8+e14/I7P2H3oQuLuUwxTJfBrwbQn9sb39YjWzadBsxoS2XIoqm3oO6pAaX7g
UkYiIqNpG48kmhgpzLye0NJr/wvfbLDEDiAKWk8s1faAjz6DxpSNzmGmd3fcfLTBY/w/lAOCUzAj
rM642JxJVEPkTgF2BFevgT0ZCwkvxMRKHqRfzkfkqoWzraWjb1p03G85OHDvC+0KVxESUy61fRfM
8/r4mHYgId2dIODYStBbfRwlHX7hKMP673U4QJY/sDyQY6RkI61LDDlWCyqoIHnky9pPZgmaSAPB
KVI8PrHFzxiEQ7u1c7YoGHihCeAKS5fjjx7YJ/wWVxwPcFC9NDl2xCJbvz4/J6mc5gcKQudGkD+t
OVM76zPesszNwSXC389SjTNtwJqu3hDZj/zsvxQd8i1LD81ZA+GTWVOQnIPSALZwJNPPGXbCtJ4V
RKeA8wKMZtXv0tdc87UfAgoIDJ/8KyXAefDGH/GgUegjpfTug4j3TD4LHq7SLl/I5gqjP3GhQlCb
oJ1KhwvJ7bIOjQquP/DXGW9wJu9aba7ieUiQKWDrLbwAZN0zoLyjJebfIY+JE7PbjkhjFScmPTgd
CIaGPMqi8i0GA6RtBoLYKl0EFuUO/ePARwj5mStNBR+T7WK8QsipGTXMBLgOgi20kCAiYw/Btt9C
Vq67C/BF9AGRpFANFoDqP23QA6fGA+t8WmSi3ozxHNnjrbzu9wDDtn0KMX9U3IYEeu5fsVcoRpOC
NvIJiNGmEYm3o4uDB3H5rAbRGPQrAUjFiSDZDbg+lrjtAwhHxaBpFHcnSdCCc3W72zcO9J9PRk/6
rF88STEyfPIAxqk1P/VlFNfpHo5zSsO8qy8hb/1KOQvU+sYy5CaXOm0j9Uq+FiGbtY/lOIg0fJiK
khBsLINxNtBx5t2vjUVt5pY3aJTHE5MlzFW9NCyht7vvuG13qoYwk7nDmRmgeTOPH+wI0DVm1zBm
zv92xoKGk4vWZZAbKugmGPUN4631wn66FBNopI+8VtDS+iHqSqGdfrkX2qpQ596Bcehd4SOTnFku
c+qAObJQwlIYgKApxTOkItf9YSZnF91+shMVeScNe0850wLvE/N/K1YbUQyAWsj7AggXVI4QRdt7
UtD4uafcOzNQ0qoqc3WmZGyAqniKCfhZMl4uJ0ZpHeLNZDVv8VNuA2jrBQAAbn8zEMWMh9L4ejGQ
E/cbimT25DLQ2LEqxsQvErzw2NPYuV0rTresivotx7WwP+L0/Eny4aVzRaTUrVetRIbJkrPJsbuT
Hu/XH0qv6d9P4MkH/0B1WoxPVgycZbANPS7wRfpZPui62yMNYPoYUOlKUN5xQt1iWcWxAx95RTbc
oEjOeyIgpaiZP1ztdG6fhtocemUBwZSazSHI3ARDTNEI97uHmMeBVF+oY3tdzPuWhns3tYd1+ZQZ
EC4MZCztM3P8UmvNvphcLiMEia5PXmrPsGJm+32rxEpxNvfaxIS3pxgCmUfqeo2lwpE/mBmrLYCO
I+0qjyDFgIXrvVEUPe7FV2E3J1txYWefkz5yCp0T9QW/79xDImcvDKFVyjBOI9BunKENvlDj12B1
MA3lRiY67zgetU765lSBceAgvmbHy+V6NmSBw5eBKk+QtoFf1Bpmk88Jsyz5kYjDmXO9DB/8Za1u
5CP666ZEAdMKyF4wCpSRHIVNM0eMWRt1OeROd52fJdhRiIj58WG7CYefYNA70ttcxxfTybsBiQDL
Y1xbZCe7mqY2oPNAuF2BmhAxiw2EV2WUHXCzGkaG9dpH0tKkeKBSylSkE7zhOe00kdfNWblMtSl5
f0m9UZ1aja1BDo1L2fWs0nt2yl6qWCYSmLpU4mDwVcd/mYc5XYWS41pVJAorYvwpXwE1LMsre/EI
zuTUiu+ub2VgQOAArcUTkGR0eq+J8abbmIfdRdAffNrJCYSxX45ANLEJzIFEbsdwJ9ttW8RrWE35
KF56S/f/xwq1+OnRAYmIXm9j450FLt78A8o6i5dLvlgRGDxAaN3URhnfgoXqIEPzlp1a611lx+on
/LktkW36Kpi68x0rs5ARg4riNDMS5GHIcrRkNS89h0HcfCoE6BFebHKGrVI0mbH3Od0Ie2VnZsF7
d/0zr+L0hQxGEckzhoKTZXIWofg9lXN47SgRk8DlGusfamxQpKmNPZB6iUW7hWDbRiawYjkM5QIb
8yME23HtQqBdHYa0fVVOrZrTVbti2t/jaovMHBX1j0HmhjhpTSJu/D/4B/+2CkReWRqjw2zqiDnT
VYXt5oJKEWTwE+RFbW9hQZ8Af9HwAj+aT2d2EeHHfxtpK42boV5bq09WGHm27/P0cXhrHGYz9jMg
D0OF4ot11KqK+06DeQzqL09MmBqn07HGHwc06E8qqXKirkgfkUMUg6X/8nY9MDJe/1Mou8qSWFei
cDlpxkaRnu+lnSwv88/wIoZHx24mm2PULiF5syxEVk9uEPpzF0eX2eII+/P5Id028M/7Tuvm5AWx
XS/JjYjNPZRY+OTbZgo114qlwfVDv8+7K4tk+SB/9CIAfMSLX1rj06tmYhsLECgjqmPcQuq7UA2F
xq8D6kd3fwAwbdBFxdeGDAKH+jhq8jxmwmbCA4Z9bkAHpWP/ldzJHE+UA9bvjo7fnTKNyOo6mArS
lahLrJvYynpSiE/vfIHLkjlgm542W+H6b2vD1qJ4u3XpLMER8XXS2fW/Qv2rSe9T5wCxdLp6Hm1h
ArLo7LUb4ivUVyAoqVpf0yQtcTi6IyVfLu9nLID5jVYAjBTovXCsvbHczZP6lWuAogys5+rP/fs7
k7IkJX1soB3HjAnbWLghQcNYGE3bhrsDN8Dvk0l0VGLqHIaBt1NcuhABGmpe48DQsJ+hEXwCPYtK
3itT/G2Rq90PLVNSdG2nvM2wK9OrB0d3Ml2qUa59ZHuNpR4u/um7dwf72+YRcLPJj6G+kUJpExR0
PMIE/iBv4NC+hG/IQ7AI83iJZQj4r8odSNGBkuFvbNXYGjb9tadZxrPAzcrwZGLPadcwUf6ql9Td
Xos3UxbJiBS0qGVh6nilycSfEkxghPWj0FF38McOIUswET0U3SJsHCnaRYHXc5e9m52/VEFprjmU
TU9VuTZcmhRmn4G6sbqjyLMcHKl6LBGMeS+srTwNaRIAcSs4Sxfha4iRuckoWJ9HbmxNZMX8EZAx
aVqK4KS6F/+R/Nt/EisL/Bn8emlgF7WLyzZHXhImxBS+O2hyUiEJMlu0DdkAoIz70GnVTAw1h6fz
W9Kpbn7Syd2ztICv2BUCrcJJWzlGIlr0o5R0rMFAG3eHHSrwrHeDJjR/GzXVVQOqp8KTa0y0dRBx
zFXey/5x7la63gJ+LaTEYFTK7BHNCWVPzas0ECdpnox/SK81ODPysa0UABplNiY2FZKudioUUXUu
nT2M2sTVFdIV9M1ClTUYMONHx4uWoLiSAcQ2cgLxtwZFGOBzgHw640PBdXz2+ZcH6C4roHOTXt6x
ggfYiSM1RKCqcTSLCMxtLT5dW8DabtpiHgpnb3GH9EMKIo7RNp5Ub7m2p8U2+mEjbBgXS1RxdZjW
bZhnTkw/jzZXgznAhjxW9QeUpU2a/iZB3vHQ5jsZ84CAQNmt0KDsPGazQE95oMOmehDiOCZy8JIu
rgArkbWwdmCadr+rVZ6F2RuaxtXFavjDAnWygMv5A06eLpX3JTh3L7VaSu1K7UgX67tEbH+A+DD9
aWgvrSCOd6GVktQjiC/oRAPWNIHrpxVpiWJYAc2ihevqqe31fmCqAh622PxYC73Fpma2TmDpHUXH
fghgBRN4MN9cq39j6MLcOuFecbtLHVBuWhpryfw28pQr5ljEqm+CRaSfvZylaC+ocNJi3Z5lz9tZ
fO0Lxff6I7GX2lMbzoBJtJtdV+CKxnkY5LP3CofRMoWAA0r8BifDJbioW9tEr3POndcTQrgnYalj
gJ0Rqg0k/wHNOAcGcSCqV8IDU40G3G+ZRcmLfhelaFdeJSb+L1Ys5r9T0QKCWXs2ebclHLyiqk5g
oNoMQ56GWCoWYSLgHjvr29tSZ6duPBG38ag0UelqXLeUvB0vrhDJ5ZML9WXxseKUDsbjc7VEam5N
5UQ+tmVLcSJv6HRPXSymODLE3trMB09oz4Z7hpd2Pe/zXBA0fxIYrKeV3vHDFWX8bhZsSwzjA0eU
7e2XSgWMJdpX2YC1d9S1/LlPNkHGzRYjo/x9Z703zUFNAjQ1rH3WOMFqmkZFVvn0+wPsnt+amo6z
nsy4dpdHkDxXiSYG5gegcM4b7kKjrqKBnJIUaZU0++Xxsw9XNWgLj+eAEWc42E1MnrENd1/oPNW1
9Okj5tC61X4ace0F7F5J+IOhEyiA10pvTFB5QkmTBqQIm0x2E0tqBlkOPOJoUmTpdwaC6wB6s/og
ViJXte/RG649a+0MJ3QXMUwyC4gAFQoQLnhSwgRuOJ4QO9XCtxh/b7DLT6GBqMdjhy4RLq2e7q2i
hk1z+R91tIwqMXMGWqWx7uUpKUKmJmuSY/EmupFagbatW5jFLX5vGRsdw1G5T/9pkFO75UO7H+rR
3qeIiboenKNJcjUXYcQHGMxXc/t2/uMXqyLlKBiFYHxN8Cnn2p8bPFeWN8kAWFgZPIKxyqSC0V+E
MRSO8CrXQkrJKtfY6NTgVtwWorvy2paol095vpJLOZEFo+EM3jT88K4Naqvmw4SmjutVKo1ynRdt
Z9hiCPRSnLpyEPuvYDAFShw1+zpIhgjGAs1GgiLUOi7eoMOyvyDw6NJCBACynK5lWKklefuMRYls
HJa0RQh2r+Qu5U5AS6QS95Ns5UvlYxaohAeejbPEh8Rm2gOrmRZa+clDYE2eH33u7zRkmuDj72xI
jwAgg7IC/p8qc7zTH7YePYDuMsL4frlOk2KONH2fW5P/W4cKCrfm57bcj4n49iqcTa8zuHAMQhxz
jDUlFZTEQhk6T+Kwnt15r0aSLc8v4NJxtbhPUhkAtlUka/yuSlnHO49L5Tu+vtxhH2Bjeay6aTLv
XF26MIfD7p3uQdvwO/Xf647P/NBMncjJp7aUamrPn1UHSCYHu88euDeAilRaVAJix9mpNnQMCTpo
ajshF8RNSLisNRGQf9hHsmAJqFWEZGHIlWIynOkzoSKeaVfHkYK3qbbwKlsTi+ImlRta8mjbGY51
xpU9mAAuCyGYmZbbXsFtBBlCGAiX21DzOAvAQ1SOrSjx/l5QZdLD74LhdbfRvX/+iepgrdc2GlhT
+zCjU1+5ri6sQ6Nas3Lr3Rxkm3Ihieb8WaSDIYudIPr4W0PBkvY6d5jMldtu9OOpLWRwqAXFeR5x
P/kKxa6xXmiMJ1udV1nLJCO7CF8Oy75QkaACxLl9BrUFk1Z+K1B3qIfJMaUROgIa4fxcW/GNu/yn
IL9g+z5mFPtGakPD3z5EyjaZMeV5iFid8KbIzSEZ4etheMHIkukhhzMg16BRoyLl7gETuaLtuUBe
y22itihEXx2LHOJlixDdh17Twc5sZpzyBBHV51cEg6Vb4zJ9p0Ld3KOo9EquMjteSIobKIXQXMXQ
mh47IrwpDgcSv4PU4W/y3Ci5ix8fHCR9kyZ5dA6ZPZ3yq6qUv9+eWs4zoqAccVU1gDSicCg1Q/ni
UqrVJs0J1Ge3ejY7G2DncIgCL43gB3GYAAWHmmh+xtkFyqax3JlyeT51IqGYcUMRcpg7ojRnfq9L
x5lhCqfM5W1fLZ42AtZtGDMMTi+oi/Xl/q/XqLD0VIdwLyFMao8Nwy/oILffEMm3tGpDZFb/SOdB
qkjzxFsEoZs0XmfOqVQ0fFACZgOUJ+sxPK5PfgmAeRus/DQXQQvOsq0WVTmgz+A6sVj5Zy57yzS9
mkyCFNNrBZhFtPQYkVvSHguNu+Y/AfYTJ/J9rmcFqFcbfmeK2jkQOCegoyVMVPLSEIvGJKuIInv3
xYgG1c6IoYUvBxH1GuNPBM7LtoyfGtLcRv9a5zenIkVCwg+C40Riyu5kRNtaoGEhsjNywfjd9GFV
S4L9RxK35nxkHF4VEglVePaoi3ubF6PVfEA8t4pjVULbKRKW61Z5KPdziiu1kNLYALTyVlrSx11y
oEl8gsNdThhTWhuW7Fs26dwHKMaZw1WWfi/jHU075brXbesKsDJyrTp/MN7e/CHCaDEjz+gDrcSO
0YrRR1c7NCC+OidjxD40dLg2gl/QPYtIiVZOEzBQvN0ikd8jfO6olMfzWIYdZGZx9PqGZrlZEG+T
0uZn+YnZ0/t8bdcekxix3x0azaX0WQGJqYUEXFkhA0OqiX57c2Ny2QUuxLLdJ8KTIOrvloomtcin
chdrVXtvB28pjtRAnlnMMNJdI+k8ICtXINaofkyRgv4sKdqLr5d0jEdrSbFuIwKKCxawv3G+e2Nw
6sXZYloyfgxbqpWlqmvSuyESc0EBd5aWICre8EOuaJvdvxOg+ZCLoynao0aO4+g+AQvqxvd/bOwI
FPQLu2vxW8Qw19ssgERNg85A85tzaKb/HuqFPAp+tMcQ6ypKKfrQHWf4SQNwTLYuTcDtpLdrv67I
5zAx1gVk0+68RdqwkDLiDE/s2hMu9ekxKx/M8gzpT7zJRe06R5rcIQsP553VQzST7GdnY+eZDeuK
DrueoumnSaGinW1UMBr9QS+rMuFw0Uz/6YFgkYQJUbT1/ncw69LosbQS1zoWo/0A+yV47AD1iOo3
Bauh56kdN/y1jskn9TSdNNQKn1goHzzPsALPuKljbAs5wVGFR7cdH6IJ8ofNcdQkYNQxkqcQ5fKb
g1GrA0iiYXPF1liS64Tr8IIBdskakl9j7UMFytrgc28yYxEtkDhqaewyb/szB6RAiWm1WJaexUpl
XSn57+P2TDm+3bfClDfA5DEfEIS85GA2CXSiitUzS0YB4TT30F7QN+Kdm8w7dhnwqGsqGoAYkc7z
UoloZJES5whncAAuA0EXVyoEkgl1ZbiS078TtQYFL9M1S0zuJxQgAn76X+KsvoB592pxaBdXvFrN
l8U5wboQq8HP8LZ/TmOESYF08L0giYHj/Q3W8VDNvqD42y0miU95SWcqEH7//lN4zHVRFJ/AG8Wj
l0zcDl0WAUWw/mM3ZWffhHlKVY4Il71tLBzsvoT3cZ8zyBIMxWmlUTrJgLLJqIbqVMb6srgvbI3q
LG550mBoCIlC2YLnq1su6nncEuhpttDHSsBLB7KUrNhy+D5SQQZIGzD1mXA6BO7h3vS81oxB8AAB
N6KGjqm0QMp96RH/H2v2M+UGcND9PtwGcdNxQiTFHrVyAskvDLPp11uDFQD2yF9XtYuOkxwW2Z2u
QcqLKO3j6Ma/AOoWyse8NnBRjuhoxeps0c5EMjloqWk++iVADfTLRYGPoWvv86IL6X8Py3AztxGL
j9WW+qenPYn/dmQClDUpHCMTMWX7I3x72rMmKkxrEicX/DTzwdK+jfSFCsRiyt+ui5tik27QC5Vo
LGVRuZ4lj5dL3re3r16HQwIuiEUJlpnb33uP4HjBYgIBtZwXsP/3VmQ5kHxPIfIQRtKfZV0/XBxD
PSe7JgktlPeJzkCo0hETo5gqp5v8GoUxbqcWMQUYoKNSi9UH73ZVDljpenm1BVb1CVUg1nNF7V6A
6wBYzz9wR3tqicFB5czs3fljVZdCmuDPKw3q9cYLoF5O5NbqffZNbTfmphYgO00FxuS9B4O6GL6E
H6NptLw6cK19q+MgPT+xqTg8b9urEbbNF7KMCSQosXuWqmUrI10hNv26azfZGAHQze9U9GBAZ3bN
yM7jAtWoQ5m5LYj0DkyedcDCv4Ok3WLbiJnSzM/BZ9z9JoMxNdBlFW+RjR3U0g60gQ3/ISa0fM24
OJ5UzUvCfxwtCDfS+BOmAelA5MPF2eHAWsEwgqiFxfGKq+OmWdYMZbcXgSpagBveyvG+mN+GG0n6
hu2+UWuS/no23KssMzlSbgMgVJkT8HKdchZfeC9wksV4z+G15EaVvcZiGrCbrp1P3RAGSOWiS2Uu
8BUamQ4s8pb7+J64xJ0g03oyvvbfUT20sWiJOgHE4Mo1VPuPkTMu4ff2bxZMW4kDR/bEAa+dcyeo
OjO1u4OJDSQ/+h5NXLsw99Mg/LI2vEP42LbGeWTPU5OfFndiXmG3weYE+rvq1a4pP4F2+Am0obrv
5dkb5k5C05aD3z8PCWQXZcH+QbTqWd+/VwiZ+lNcBR43Lo4FN8JeQR703c98BbSLl/DWcJmGdgSA
0MAcrUGy/9u11rt7v4W18O0PIM7eelPOJD1RDpHotcs3yu8mHT2gRoVF+jmsbYqc+yW4KRMGuMGY
upxtu3PDAQwXj27Oi/hVnwoUQPRXcojfUyNJFIklDoR6TdbCCy+x7aWhl26X83qout0qq/dbZ75b
D/MkH4cVPSKs1TJKKs2V1gJZnkWiVCLgFPfoAxSIIK1lqLE61ufiESzGWCqdtuURhDvXsgt1WJYo
FaE+B9xc5XVJBzDOalSBRcwFCO+hZN1U6Z+ZK4NEHHe2oiaCKhbEucd4EOtxghV9GZPEH21LfXcN
eIpwUG3vqR3AJYRph79Vx2wzhJLU/0LYCsIpukXZoSOvRk7ThUTQY42grPxpspf0gzrZ2yPCH2hZ
GxuZ22oTRoS53oxHdmoQ6bAo+drqFOrazOpjOfNI9SBSLVvFA0Vih/oFaqpUq521zrJMri2jzsmT
ETkGdyGgkROyDSY2/5EywuV+Y3jwDT4/YXcTMgQA1WtTlAFVni3ylF9HSQzRd/bFXKXC8bexwQdU
tnnA+cGVI2+OU6xPO9pAroWA6eZ9BiWgR4AZzfmfUjFA93WTxewnml7KrElSCwQzrRv0sK78EMX1
QHimU9fc/LfH2uqe+Y/PcZPCt0uDoEXE++fjHtHdpTX0hEGKqEgvkNSOV84xQPmCMtVNIylsxtPJ
j+BcYSY+ojPpKn6veECJHteoy3scBlJ4I10HeplkFXAChIG/63EJEbaNlSX9QJK1ILXqlzgrGjhJ
bvo8J1Q8+f7OwyGohMZetDBJ4d+4pni4uE7LFSHtyf2X8rBznckwmagnVOYFOxFAyWh1RYMML89m
W39nrEz7lvyNpxg8jZAQPzi8c1Db7dQy7UTiI2rJVmUHzLoZZqw0ZfDK4lQMXuPeFqvk5ClJIQAv
KUNlR+MHkIizbyk0vZWKmFMJUbwkiqeebdWknrpKBCERFG9oDVH/MtRFe7EwVb8qEESgqUlkQbb0
xp3fZtbd4rf+kYI0GlEskKEdbL2XWMcSxnefjE4tP7rB831cuOHU0WiUv/FVvYJvA0paxmAlm8UD
wahRw3rlyBi8V6Di3FkLqWKyI4AmbYScqo4uzXkKDWAXJxt0gz0okRDZC6f0lP4MWuSmxwjzI6yi
OfcNpkxT/R9OI7eubI178FRzfMo+iFaTPVEp6vgyhSEXsLBdTtTdvPXfcseVHLdz6K+GFtRKiGeK
e72BULISWURXfJYjr6YZQkEVof5X/D3kQENRbDW4n3fhriddJIeYFlCpPE4GeZVtLx2aoQWPGZ7U
He4fUMB7hMHWR6JB88QELDGf7EQLRamQWaGq0PUL9YR8WweogjtBsDo6knEBSjwNlCZsEILwz8xO
At/ZfMWljWBNWpP6fqqmyX+lx8P0DrfGI6FHAzW6Wv3SLZ/3IC1/WB467coL01BBHRTpIaXW7Xfn
Uyl0ylaxLicelcKDmrznjRaC73vsoTVuGypbpMCPrL5IDk9y3jqUextQTemYobEvog2YrxT9KjqU
pS2uy3KbcSDDTjxn7TgenYo3nAm8TnIEQF524i5T65eDV+lva+GLFWbOTsbHDxjjIfoY7o6HXhmr
3WvLVPJ7NambFts/dX/wFXMXzkHn/g84qSUWEJ1WeGP7sWD+bIRMafk8IikmYztt6ZsXdTMOCi2/
z8r8iOq2iyaOaoeCZDS2nlKorE1xK4UD2RTcovVQV6aCnEDkzkGhxsz5ZptAmF43DnmKWoWi4gsz
A88KfimLciz25klaDlvoUtkwuJt4Zc6UCDY/uv8icSw5UMLkWo7ct9F31sYvG+Of5IVZX7K73eE6
4TqqzH+atVmhuqquzTf295ir668B6sL693nvCoCy0EJq39VLDqn3mFvUX1XVG4IKY+tEsIdNzS7l
2M7xOD3YYMf4WrpkybSK9HADiu9/ASEchaV/IMBwcN47FmLf3y0kSdXy0ecSkpg8JYeBXKvOt+/J
UzbcpbtvcEd9KkqPAKQjFtdS1rXFPy+uo8Y9Mlu/hzkGy5qxHiPHORMc+RxtPhUqHIGJlnzS3JAB
UlXDlBRAUfKkL3VVRCB4WF7l6KEG6CaoWiNlvLpiv6QHLVBEYQiaZWLO7HaPcynnaPPRVtD2AQgH
DQYtS3Hb0shJ3wZNw4Tt4evCLRHJbX/uj36tp3QGV5Ru8cXtT/KhYbM1T7hSAn5vSNrBZ3sDy64Z
X4PVScOItQyCeqOJEweKsEZqk2T4EO+7vhQ850QYhOcU8MO6jHWJD2bkBldLAEQ9wehgRu4pzFT4
UNmRBKnNZQtzXgyNmCzhcEn5KQwcbPDuUQ65eLa0Arz/XUE49J84eBPOOOlUon0XC1F1ukFkuDGY
mmWPgFhL62+tr5avReNtIl12dpdvrCo65yRFVqK+hCj9RG02g0rVOpt1DEzBdS4ZT2FMtTQuJ/1V
++RaGvtsMnAcvtVXLDICP53tErYsUHPDcEJIzIXkZqzWvqnI00wvuTqe5HRVd0VTkFq6OVYmsSmX
Gjm+9HVjOw+pCWJLD8EXxFQo2KuB3JWOfwxZGhdC1qrTIUxeLhz2om2B3fTZiQTTswazhZTNP1vT
jN/gRHHbwlpDd6rPq8Sj/lynV0r6GOLRq6lVQ1kObBlzsOyZol+gAJwFGQ3Dk0ScmJ6KCMUq1TPj
1HTGyWHFUlU/SbAcZDonM5vsHAK1UL8kKgUoLz08d+67cHlHfv3fdsTbOqZg5CF1nmspuQ2hp1/G
S1tY7guTH/pPVq7+Q/gQ8Wqc4sY0B4whXKp3TlhqY9W1NawZ2ymMvLpTXTPb7hMNaduLYhtYn+Hq
KJR5l9vRVR3qmZwtVcbh9rUYwgRgTEuP1whx7DVsPAN4zRBtzwByx17xhB94MduXjWEPyJ40nJod
T7VDxwVjkp3zxewvOZZ5u/sAm5+985MNilmxoKc0wEMqDjILRPJ1Gp7aLi06nkshRUTWJXwsSOev
Of+3IWblkm5MoZFKNI04sCFkHTF4b+VDGajteuaI7txvDmwoSI028+ee8xzOnxT9Av9F73uKN2Cc
iEasHkE8iiqj7xCZnLccm0mFV+aWURdVs5VjKe64ZE+jo99IrO7iSr5QB+b7w4sRouRnTtO+ITAq
mhmk6Xrs8BoDRDGSU0rJsCwcrxsAal7FE9BeHYVouTM/V/lljrFJ2TyLr1ZnuT9q/5VM4IsLps2N
e3wGhI7u6yLfvPKvYj66OPmBus3do2tIlAgwKusLIoDZvx6LYl0r0NNQ8Wrdhrs4xLiR0MGExsGA
XXA/zR4Y7E3KY8dRJviiNdfrpva+ZCbR7m7rA3lLInKGp/DFWlZXTeEDZ0oPpXZIEHcvmeklxR4p
U+Xmq0XXgbPQ0gxBguZnzOBq0xwY4CL/3vIJoE9ZSDaEyO3Ot34O52yeqX5O9bi24v0Aw+bhnW7A
DFWupQjHUvpnbeGGeWuDk0J2hcLyPf0UEw5mtq5Q+xMtJn+kV64Ib6cYEaqEw+QkF2GGw520YKft
8z+m6mburQnrG6v25P0E+O3UVi259bxQ7/jdhcrEgmcAekuvX0bHdOzagObv+3HWeJPiBLRMVUso
3eJrx2P3Rr/hpacq8RNmnIGUh8Hv8jvWQ1sWZnoGQZVs9i3LTT5XW6tFRgwuV68HZIvUs94ooNxu
ccilA9SCpmPysqBMB8oSmdDs9DdiNJvYQXsNkKrhvKWiRA8w5WL5E9RdUw5Q6L2j0PVXSbDaudjC
FUSh9zC449js3k8myCcpyzzJC4f9gI/8vV9dbd7E1N9V5ULntqWX4Psctfobs9ewMOqeEo3Mjsjj
7sZ3QOVPBfPlE9MuQQJGnI74z52Kt5ou2Lk3dZ3U5he0CwfNRcDfxseyFArR1fIAdTFZK6blrKkL
rwhEg+e6hQdC5kyzQgOcq9X0iTQNxA2bW4brjDQpc/XkyNFl3BEXFuJf8JBys3O5dDYmhjGUzO9i
lqAdlTnAwdDDDMZIiXTT6ubL49SUnq0n2YaHzM5OBeAwi4bqYaG6pKRszwQu7iiUN4/k2fLMOBic
TXNyo2edCMXJTq0gcQZ9Ow5p/Nw6T2si0ZFLPuuwbcs7nBrB0bb+bCoQsde0XfxWAQSxpcSIwE+y
W8rhkE4uRMnfldIbPdPM6ixPsJp0vs0OylWmiXIcc/AH6xifOk+REbHNA19paor/MT9onc7Z4gXC
OWtiPTIyVGe4dxisB1FR0OEC6yKpWh075If8hLSNuFkvGq7mEeN/UDDAalMrQrd2P+DeN4zVLzez
4UIKw71ex1UzfuNsmI6XT2N/qJS6XGUkMkj+v23nIrqIXSEnadI66vbYlgwkt/9Gm0sAm9/aAVfE
zSknKoOeJboUXeh2AzGN1yFACgGbquYcVt1I8H/BShZCGAnM+CGLaOAtMFgBouG1VFyPys0BuAC4
WIDhIA7FducC6DhLJO7MPll6SdNRgFt8k3wzj0j1FByBGnpJ+U6WNOsYE1niayXvKnm+Y0n1TT17
tvQeh1RT07JdpzZolZ3jpB+293B/HEowyZN0uGyh7/6aofhs8A43ebgdXHzXWmQQB/vFvsMxwUfI
07YS2lT+dNTS/bmpgJtKnLMrQFYsDfXOUjKyhV/+jjmSzyY2UJQrsYnFhE2/iakzGZANiochBePg
d8TXT5JhucBnp9OFiFf+k3NaollVth8U0ptBjY7nAkoKEPJenaen8mOn2y5FyOCd9bjnQjGYcho9
niFxHnV5S8OBuVjP4MgJfTacUDNc9Uq8u+Gf8pAW0RCyP1ygaDU30eb1gOAfoi0c/nuFZfOz9TWk
KHAuNHRokzJBaMn8MvmFMbbZBmnP26lBZQ5k0hhZ1QZS7PqboPnkWggAOfVW+3SCR2E/bNeqfBDO
cVTHMn5X3csOt5MXxjUCEX7hxHGKbv+Kx50Iz+10hdw6MqZaR4kThyY6XBDOeOU+rnxc5a1WOt2v
s8tu5l1mUihsefnc4nAGhqMNBf3NfR3xsRa6NGyl0a/A7k0BV5/IwXGS5vECtaJevQu3Qc5hw1ns
Eo79oEnnjZShZYQxDAxUZn0sQAB0nz94fn5SYPlPDJeYuSG3bf7AuT9ANYKT478Uv/UvyqUdCWlF
tW/gBQzEiNLVcIR8pB2Q6F6dk89TyiHRHHUgFOvEc1zsD1mv0s43tmzvtuNiwx+L1DO0+RxO9UY8
h8yHi2bc2TitStpTO2yMysPDzprm+mYq44pj9MyGOTp8On9MAuo3WjnnBuAd5+io/hgE9uGIO65F
CnOYnoGceSF9nCY6r46pBEiiDVMsaZ+UBPRbnup6xtrFqaCO3clNRrreDu/pA2GreXfyBjR4QZIS
dk086uq9Palz2iu5aRQk3Us8hfY6iDD42b9zVz2W03dS6hXrgh+GabwemoICSZQqKHHnL5irbotW
jy7k9MKVkDN0MItH7ikYPhl8k3PP5C2npj4NodsXowbtTdmrtH3Aq+HXd+nIk5TrwKEav+kllfaj
kjRcy9G/F/nXHLbuo9QDJTvwLNn4v0bOgwBPzJTM9Bx3Yt3SVu+DOQ/w9DS0xImYiEEUZggzQrXZ
7m/+qH/PTTTRYNfrB5ACwtzCBipD/PkF9k/Rlki6fwQoInRSxMkFmrPmVYdgnmU9B6ACFrBJJwH+
+Zx/7CGidmITgWRFJKgG8b1PnAbK4zdK0jqugAbbNi5NERISR4sX5EXdB2XE3cA9zFZBP6/P7Emh
teklP0TEnWuG8txi7JO1vpoiVVKs24OTlNvYMeJZ9Uf7UVlOcyRqFNDSibTH2vB151xCTSAiNJuL
U5fIB30FlZW7VWXQnR3ijz7V7uOG2q8MOd0IW8gSROh9ppSjLSsqT+xxOM+TfoVAJX9WZBKhfnl5
wqVcDK1ccLnVE2K7/3VesZpA2jg6RYiDj3qkVIPSc5lILtTXeML3/4rWIJHoDxAj0MG5kqXte+pq
XhGXrb4Hu+fnE/gtkj4QD0KobPcPepsrMX7CWeCVvtaFGYyczhlbK7D1Cc27kGZlTykMdAbrnQ89
sf64JLI1syVZVQo+u1zHo028Nu5yusVH3NxjW6KvLgJ1kP4iY9sOakaheqdpawBsixJpzA5fblFM
0FLzGCY6CEvKVNGYPbU1aLejbucEivKiFRNNaKPhMnJDBYfKz7a3A3f9PunD3KsD0hcAK3Mh1ypD
b5jLx73BT7qyZD2Qu303jBqVpeThbyCzDwRVPZCpsGWAIynIZo5ppLODMGzj/3v7EU2DxO/9k45f
Qqu9TywHNLkPF5XC65cAk/wcxq7NJ0vqEgk8gD4S23TnklVWR2NKqlpiEHwAQJ5DSOi/nrFw2MUx
GaUFNPjV3OQ+VRAdQENT6SmatmwKCqOWYn4+z/n++/nRcMFgu/Mo2jHuwiRhZfvk3XdEtQJX91RN
KyChUgzvmoj79LbGgHIFuRiP+t6lSkQiiaGZyWASympPEzClDK+O8RUg52mBlJNHgW0kSiE20Lps
siDzo4e0bwUtCgLQ10cPEFIyq3+7d/JtC18DyJSTxG2brb1cvVIZMZbNfOcoABv1/ghYQILTBuyn
SEIIXepnbZM2/tUYIoBtzzCcuBo7WZclKLtwnVinsaRMl0ir0Vohj5FyQHVbtiAJL7K2ZlkHSCjz
pVGoGw+x4M0f/aXIdfhGTmAJQQV9fCh0ov5WYeRBktGJTBGmzYgF+S7my2GBkvB0J91fGkfNVpw+
ZwssxX1ShYWUM3noF/IRhrWt/7ZAR2EhwRIMEpSAXX93hM1QSFgdum0cNIAqT+KpOeor5JC4iXgv
OLezX/xPijIiVYBwDWrEedsX01AkOc9xv7tm+ikTeSdrIsTY6kZTshaqAgJfryesnK9mjucDvPAp
lHINhPAzQnMRMy12CumOD0eC/MYWo4TVFtVLB6k42FPOMI+CIdGCYeeyTrPyqX6NUK1ctkxlxDgb
9CBL8RQT8tIy1/pNvgOAxR7nTHU3ICBJXB03zRe5s6IJHz4y+guX1IKvb8q6T8I10fKnRxRUxJTn
XYDkUAgTxCUJQYQOqYkb3B9O/caLqeFm/nxaUMLVYDt+9iuZQ62dUo+gli4yyg0LtKIdv4+5sIPm
x5HHyIxXiC0BtncW0GQYfVg3l/aAXOSeH/RTApvC7PIGQiS3GMwI0QiQH1MY4D+G82dCvmkQqItz
F9vNS8X5U6iHPryAJAfo9oHh4KVR0wYM1vsR77xlUDCS+Xsf8Jmn6URjyR9qX8NBWegk3PJy1HsI
On1ZaJdscDW9gbwt7WylszildASXNz4+UQWWfu7QUEMuhUuuMlyJh7PL3d1Hgl0+I2V6bLAFQQb4
XfhDU5fdR8FYtn4432blvhhDr1r9DAyyjvXxG85VJYPCqML6735411iF51nSms8hAYf5D/7xFowB
DxsuD2DSxfCHRGCiV34uLH6amcwjMCF6+Va+X4KlTfo9JPF4izr1juGzsdgW5hjB3V8QgG3Hb9qp
cGaPecSpx43eAcEgiITso07LJQkEQOoAKfUUkd4u6pibGDxyn5PoDbxLoJH767hnVeK2Xooc/hWY
K/Al/BeBdGyzBbR9Y8AjQp9d+BEQR9igwlMcJ/mhuv2CPYjBM4ReNugI3oKLpMhe72v8vhfbLtYW
xTI4nI9mZGLVExFtyWCkAcjJjZVXTe/JZALfeoGkiun4QSPI0TTGe1HvfO0unNmy2zH6MyBnOTqZ
gHCKkkDrSq0Cjf2PCM9gzu1QrmG8TTOsXJaza3YJPoMIsZ+C3P/EQ+1dh5m3bPq/o+RHsQueceWC
UYQHebUPpGShxNA5xd2oQSq1Q7ipv97T1vvI2oFe0x+64bxbuv22sQQTNiaI6Au/QCeXyafxY1NF
XdYuG14kKP8edEYF69+Cfl6aG2fEk0HTZEfPGEK+uwdjdsG9LMGvJFZsvYV+3VUFNTlwMjfakqOE
4VDVHkuqNUiVeNHfHWxFn78DCsaxw888HsqGvhph5mXK2/Jtgb0SkhcsUhcXKPEvxVtK8o3zNhpI
fvjMk/mgsY0DvrJROZax8ujdao7azIqullFDmj/XfA8s8+GGM1TFzFcAqkGF7BOOAhkYCJt5KTgK
zQs/3ZClf4o8XNezJrhJyf0G26U++uOV6yWjPCCtSm+UeUnpsV46/aSX9WTPiVHWRmgVylsfSBc4
RZ2HQ/yUzavNpaNDpVQnI4mkKa1/wNNImoqzWva7Oc8dthRe11JuEVO7LoIkf0s4OVd5aqwgdjRx
HtAvvuYRCwoDUxdlXpeEp5HeFE8fIdKQM7hrt9gvuU2Br9NwbzfltU/X75ydTIHKiwnFfq7+P098
qI5mb7pg4aJoaFQZXmimAlw/nP9S6nkDyXpZygTJUTMnYa/cTqEPsS/bP6PobdzI6KnfP3Fy380V
sGE8/SUcM1FKYxtaWb+kU0NJuk7dZmgqvgkhM/x6AXzdr3bFnNzuoKjl8ad54e3qLDNqtm2fgSoM
Z8Rtf8icBb0qN50dVH7720dW4DBD2sea6p/aWt3+i1n9nwwKsA6+oP7U6COsa4BUCoCnaLQar5yf
bW8HC3M5CiMEIqAz87GVh21hZoARx08hgnem1xqDqhRX1AcjnWCkcCL1VT0I3oHuQ3qmDu7dTe7m
oAFJHoczmwRNNfEyWalObxjVCGyvr3AQ+Q1YhsuK7dcbSxPSXX+bh/ruXwYVQ7ghc63xN7v+FTcL
luhG9y/oIrDmvu/aP/ftkvQMTJHD2bzmrfwitPwHLR3MT6pIOFcTTpB4ZjtdcH3VM5AOhORP8zB+
AagFRRenGv4b27KE0f3UaZ6oMGJVtozloXghJSkgPmrUX+Kdzt14+vSkQQ2cLEzL4dHbJjT6OpqG
/Vy6FjpphInjjyQxXCaD6g6LLYGnREGucJs26CGKkicJOoYXywQDjxEERH65ktdHBykvbrmRZS+y
3x7GotM4CcvKaJS4t4adQHpVtO1+/Dj/6OEMpIt3Yzhj57S0bOjzx/KYv5l0zaDZOsCIECnOj4YG
SR16sd6tUM0LSGzn73jh7EFmupYvDMdV9o/k/lpEN1iB2q7XiTFDxg029KsnQaVFM5tOC3r5ClAY
RlzeeM2mfnjlfHVkXRFaYkxEz/+M2GxzBB3Vo51ltoNBqNsJqpOb3o6HWJTjqVFA2124GS2YneYn
DQufXy2DTTe9WnUF3NQ0tE7Lg9iVYpyxpgL1+l10a/Q7mKerZjf74UJ9LaQW+tmGdEaiROJJdqwx
mPF5m3jlxObB/j0fp0R7UKocofnYUPvMhEC9sFC7T65RsAZbFoSCHNstK7klbGtcelPNC1fIES15
k0n4z++Zk2VYBJzDnWXxQ81/PHwYKStSHI8Bvt+BJisemruVvU6bgJ7LJhO9k9zk5bNQTHJU50/6
jwUdhkPmBZLpXqq607CjDLUsQ4zEs0RCt3T4XduSDqy2VxWhYBsaPVNIpg10J/F48SDD3C7BtB1W
mMh3wDvkKLZVUdApnZL6B8jIkmds+/NydqIKtRhmfKsa5QHmIu7WbIMW5qsSKjdl0pz623oxWm7w
f5V+/AxcZFEzkCWMG/HL5+lLl4fZVK55HIrLVl7VnK1aHXxG2ThzXD9ifpNKlCw85mhYVYXJfUgY
3GeCWkt18Znaz5jKD+hSeDhDy1kEpzECFkM6btXouQr3dPwy2HQ9agzf+TVW7WXgB9Z4+WvsTvNt
MotYhfnHeco/PJLbngWXEXs0xMKcofPFNBQUb4Id6jjW8yr/w4ExHzE3ppc2qTxpCSnXL55JpW08
a7D9m8x/AxTkwFe+dQEE4VBeJjGNEmuVmzE8jwAMLefAWv8OINh2IwmPbKp/An1tki1zDdy8IIXj
0qhXMnjwM94CohlfJWBYdEQHTWdNIYAmMg5VAzuhv8A44thAwfWXrtq2o0oZH0RsVBWEJPiAjj9P
wdMdIL8qASLk4RU7Lkmf/DYxk2oik/HA3H7gxUQd0tll0GPrkU9a6YMbPbOkHyUR+LGxV9D0mS/E
Hh/PI+lsvAert3TXGmzlg78n4noFWavX0Y9uLe9Fhjl6h48EF/LFATuWfnpqEMHkMi8GY+x8fYxU
E+3XfxPnBN/86A0kATFKF+jT68XWDNv7eo8veZ3MJU2y4hkfFVmAZDuJTDCbeJBb53oaoED885yS
D+LaO1u6Ymuu02lIhvv0TffldlhwVlq9OGDq2zNLrU0J3gRfzWSbPKMJsnzXE0xX8hB2pXaa39HV
dFzjaWzd8DhulXKNEH0XWnPyIxGlRTHvuThOPm0f2cBeahDOyp4J24/bOstD6zQNMLpD4TIpzsO1
l8dR+yBTafPHCqwBqvE8nRRWFxDwnRgE/zpIE5ZMHoXXmrdY2A7FqL9dABtFI0Zex1/9taoTdfEU
qcZrAHdn8Se6lVoIEeDwTNZ0opm5A5YPvhPW81P8fuc2rkg+9LHgUKP/sdwFpfGAWRkrwXyuZGkc
PJ+PqceNIdCTL6IEVn2bbqO1DG3jItPWAwGlR+gy0f8bw7NwkQg5ZP+7tXA1HbVHIK1g+yM9vl/i
s0gNKRJtOJUuXkZwxAbVzNhYtErRH7WRv+VNJWTRSlONXSxNrXtFFstCCzbfmBi1Ajh2MSSyLPwT
8jl57hVeCw9iIhF4CXu18P9oxz1A+bYnAbvZDZGK0+qHuyP7gmgKZu8VHmPfqeWcvrhk9XUhNch0
DxPEGGTb5wRRm7znwr0ylL6th+ptMUIIQ7BMVuExv5Cd/uAfwwkuDohpnhULrf2k03CX5eDcbwV+
9wDfI+P9yhvwVjWOWC6IiCXtoX7YpsFX1VcrJUhv4K9L8jbJ9Gmt55bfe9VHr7Vpw5ux2rbsxeRf
YBgNjBcQrBEcxC6573x25jAI+p5E6fTAungKFXcuZWXoNMKCsUfWq+2O8Ey4hbNdDy457oi98pG8
cIo+fPpLcowl7a6inCRdmhVQwRW3Ou/T0bpVAfNv8ev9Uoy3TDWupx03Rnw9q/tV/c69f5sllX+x
CkmvQh0obpNDZn1X7h6U08raLY06mxxC6m56nZVHCcmrLY5ClHCTwTpd7dyVBldQ06USrE1LRbCT
T+vZVBiXlTCEEOVTNcBFpA0hh8jqLll6LV0SX7H+pMkXhmNLCYaj+5iXmPWNTcbNqHUEN9TsP7Oc
154/wuYQMB+rTfPyNdvAmgZ8ISJXtbfp6Q9Sj+T4StMWcq9Dj79Ba+yfmmI8QIrvjMK62x9QMxVk
L6z/TnD0lljk0BMnBd6/79rvqu0KawqUQCbM9d81kt43gay8qbqkf9KYIVt2lBBG5Oe1nebzXeb7
tPV3PDNAFMyn/1TjGZvF3yRqf9Nyw4rMi2o24hQBnFfwrQlwsuzssiU/iqJYb0daZ5umNZpp4us3
eS1ngH3iymWxgWdKuiL3WUdscL8liVlPRus7eUtSoeJrzHPFpSspMQOdx/Yq8r5bzo99lPtRaf84
xMWsUbbZAwdtKvb5znHR0u1JGbFvzDTZRcxVZyUoEd2+7XDMiDpIrTX084rBtCDxHX6YAwD5rNHV
XwP0bCANz9+Irc4eSrezwIe02B8kaL8UKa/uNxGx96Z/CdHJXVk3uurGz9h+XsZKkSxP9NioCXfp
dZI4YbvZroneIMHw1w77pVJL36tdXRZMWR//Vszb1Ar0D8QLQZ7lfzldXcmO+VTTkoSSM+qzNQIE
hPtBcC4ic6veHT1NQB3DikYM0F5AFFK8B1wEr9pCyJLcHXLmdjUpJs7hPZPMsyYSoXgOc7Z4p7sh
QeidBecu1MQLg34KAtAzkjjaz6Ay0NmdYYSciIkLezes/NtZiw8ktDjRyp5jWc7hnDyEOQX/B7Sr
PIsck4Mu/BXpvzxhDXssI3h6TfxXRgWJ/Px8UcOg8Lxhus76HgB7Dg5Y4BnDzzCzyiAPzW7J0k5m
ppKjvo5QeKdwOy1UIQosaHn1faN0r3OL9pzSpg3iPXtD29Pmd31YX6W80H+Id1Ajj/DZR5+y2PMY
8x198GSYqmodJ3FSC6gY3x0LyxvZEF+MMvMmvjGzTbJe7Q55Jt3r7+5T4YS9nJYDDpS4jaZJ8nZC
CxzdCt1E+enGenExL+u6uvpaVmpeK/aAhiY+DMSIlyo9XkFsx2VtArF26e4uvSroVVilQxOIiH5g
H2ghKzJaXYMTcZ2ovE98Ywx8viC7mhXz2s4osp8DoILw/nKFBGnFHit0quTK4bBrYmwXlsAry5sx
p+gOXvjiLo1EKtddZpczZF9BskNfn8N53nD3AerWgE13EqgA5UzcbVPwQHfpNOop/3/7UPPsZdW1
8IwaWCAqYTx/zDcgJa095fSHS899xKGoMkFMj0RWG8PwgE6gIZZbxUdS02aceOlJthLk6RD8oBQd
YRhkk94Kx3kzVz8RCol8Ss1JLtivwOt+HE3njKaUzDfZh17NVoA4Uy3qh1zOArTWXnByPxFRLPrx
FXB65T0s5Tg3GO94cEuVSwfZTD6yTubGF3AA53f+RjrVW0ruCR8+iHVf/lRDH56yWVC+XmU7Cop7
+lO1/S5g1Ord2AX20LREZSaECyhlDW3karrcXPI44f8hTfrth/r1KBpGn8c0VIGUh5Q5l+Yd/+Ti
vngOpZzBNS//hP1PTySlAwmHMVPK78CuI75XqdGG+5ga+SW0X6DCoUEp6/1TMvp/SRxm1H5H78fy
UZrIBTELK+7lR5iY3s3bPEindJV+BTCdSu4YVAsN3FeJ/x4tQYCB2fiUEJGlfstGRLAti8MCd8Zl
E/bm2vstLt7dpp9Uwh3jK8cxQ6phbgHYUznOURbfOP8VgpAMLylemn7HagPMb95SqQHYbkP1+Lmf
bDXEekdiqfaJUgCBIB8yiPH7mCb53eMZiNYpxXbc7hbzWxNhpNhd8Wws/BCYZXiRf/Tqg7di/z8d
DCkP+w7gH5YGZiI/3TYCChDj92EEfN6Fj1VVkqnRWxecT+GW2OXSAGpZt+egxY7Qoxb27UooHp06
A+IX576r1hNSXxPRC2BfZZuu8/756/ITkj9lN5dPUcv2XLoJVGymK9bm5SeouIVLIlzVO2NrT+dy
DivZk1NQP9HSun+6czl5ZLZaE2AAfIDqs6+7oWJKRLbo2/ZIqoXPFGSEKUrXKdm5SFy3H29jIFUu
VaZcPEwLV+K83/qRSZzFNrmm9Zwo8zhAqzhNvRQnvhQu9k6tGozbDqD0TaS7RAnYlCY4iPrtmQbJ
gbSlhIeLj+xOZwT3nFQ86Q63k+gmRj9/DZbiukhnTAXLEr6Hkaeq0xyK67ZnjVulD0ybUg304Fku
UCfloXT4pufa+YQT16/thsoR/sQsPn8CM6PU+FgkV+eJjvaWhej2pvSepuzmHecEWe8AhUqdktco
V8ZnxSJfkIR7h6WSogfUDhunrzQGt6pRw57FqbQv+MlvgNsT8Hq6212ndIg9Jy+hqvaSvKWZXlSK
QWjZhb7zfm9uCRzNTNDtWd8rRhA1gFICP6vS678g53aJlT83K3p4f3qYb/fvg+0cZt2WatWC6I1q
axHrI4Ed9VR+y24fX/3qCa74ZD/TYq1Z8lAOTkCFiJhK0vGq9q+lupO028Y83DLVYVPEHFcMUa/b
xDASO5vYE+JixOhjd6280FRtvo3ZmVG7PjslZZ4PEDOSNzGiYgCZjO7a65CYCAe7fq0dOdR06qbb
lGqdXcHa0s0k8MgowLpUqiX/YO79QkXz6Xj5cTvnCU9kUfLVKWhuVerFD9hyRWUr3LWclLcoeFrw
9LouiI3zMCBlEW2fpJ+antbFJ3oIEFhNj/uMxcAL/iW7TWbMqCxMiDdh6MWvOwRgZ2KHDtJzc6sU
ryZsLyPYOF28Kwn+lgIcDfbtg6dnPNLjtFI51v5leXdhF7Bvu0ntfIXHJSMFALTylPUZZd4YRcYu
M34RCD8vpDCWlz7xPOc8O7h0CigDtgpNn8xQj00nuWN4neIm/c4BFW9wiR99FylyVtg4JAarg8Rw
iv4GEnJC9AKUBNh7WlRccktffyDxVclHR/h43xS/2llgP3jSnAGp4xEmsznrlQLTx+XFAuuBJ6gL
VomIRxGRsw4KBlSgHhdJ93od9dH5+aZNJPGjvOnBtctlpKmP/VI1gdlFXuFbRVNgWFin74BAM+XC
Cit6P8pWp8jxYTRcAJbEGGU84+n26GDWd6Cx18XnBkzVpf3QTIssMVgCfzoHDZdZBU/o1/Ho6RjI
qt/2g/FwVfudOUY/FbwWReu7IBT66OQBoT51+c+1dUiaUn9zz8PIpfd9qkHa44Zyb4JMsPnpo7gz
Aa69Em002zSthShwpQX9nMyZwlUpjtQ/P/RVuwu4sZ49JalZHzaW2kjDwNOP+RvFLRbH1iPWyvAK
UUCBALqdGH8kRKP2i+Aqo4bcwGdpLexZxIgxd7x49lKQ6YGFxCRPzBC9EKb8Xr8P2neagCHRiapS
HiHfvUrFUFKX/sJvD7Yil3T8XWOfaBK4WH1oLOVg/r6940ZJ+sZ4nazMOir8nqUxlJe0F7cB2ld9
GgrngJraYzMBorQ/ZYl0HgynGQV2uuhCeUyoUIWAepZIY0ReSOiYdgq93pSAgOa87Lld4DIw6iii
8OzNBWtS9fLZgmn4RF5ZFsKSuIXUqdMD7Z4TVoSQkH71BjVqa8O0pmt95Ev+RNOdYzBuyrEp94Yx
nw/a87Vr1lXjKow3MLE5sWp7lbhe8yK1SmDoBhSMc5TlI+F9FSNrOKz+dcTZs7vwzyU+wXNOs8AA
FGIg3tjTZmXNYoWoN8I/ceVn8GILmdog1PUV5bTD6hVR0vbw9q5D2/ltsOV9hbjVggiIUyOTPqG6
j68vCfyu/p1B+iHQ2Dh48j19pi0HJVEs7WuRjb1AQFARySOrGSXjzWADLjo+mdibfjV5o4mOUclk
azsSCM2Oi42UStSvcGLesJxQJYPS7oWxmWjpK7jWyQMs5VZsOJW0LOaQkUkFMarAQiBVaCsqmwnm
acNcx6HZ4DNyj6cvvJi1PIPd805EsruN4PFwvCv7TqZUYGUb87ZzUGc8ZXkFMFif21IoCaEsTCtR
FUaw3v93rX7anur2eGHdVsYKU0VAEhGyKxoh0CLB8Bbk6vqjt2yqF5y/usLLbAw7ct4B/SsIX9QF
kGuzpXe3FCOiHr+l1ZzFi+STZnODHovpiFbR1mGhXF0wjeTwY/31Krt47fpHdPv9MjsASjdGOCYW
UWl7CRag9ZGU80nrRbwhA2K9pKf6f66RKR1Mi9l3luAMdiQ90gJUfxe+WEoCtOn29zRTv+zodhQc
bA6SiwSqA78z/V1vjipcZFTaGrfUehHzuYBlo/wx47hTEFnJfmYrA3MPDXf9AL5bJKhNtlE2AgxL
jAA72H/I+u2eXN5/UDUQwdNrDTvWSQ5m8vtYRQBawj7Z19yqPY8FGULP4nFWekMVkwc008Okr2yG
mBiBvw77I6mR8N0TpHfl1BHGr5D3FhXrtsRDon5xia0Cvee4tRjvoYxXAh8g7zacXjoDjTQM4lj3
oiG8OTS2FaGfeYClcSeuH5ukyMxOybUDA+ZkRCaDzrIwxmRCZAq2gUY92hfLFjOFO1JjfmXQcIrh
kYpF9LSVE6UD71WH6q5dFDO6XrkyD/FZjVXr/A5fexBDVpvfbfbHT0YZDMaeUC79XAW++txrdVel
doIMSBpQV6csbhQUt4I9ZO3n7uSnG+QGqx43NB5H+sMRJ5egg0eanyBVzNYw48lRDDrzmkQXMyen
ylB1JQVTs+nDTfoT1zdpdz3526E55xb1+5zvHW6o+UqTdVtzJoqrFskdvJHiZzh1P1HSeIyTl3ub
PwqC6/6Jj7l/kI7TfrTszQDse5iY+M092Br5cSpoqqkGByMBHfIsYdfKu+6d2HeW07Fuv8QrfqFf
igRZ2pKhY+M8I189LFxFB0inP2jjdH/aoA7qJl9T56R3C6PZCRhwFrS2upwGBGaLWgVcOFhCHisX
+4xEEgwF3oHCNYYwKjMu4Xc5ga9MqarC8IHffwNo9POZh5W8AGsIQPPFokJyQKEJV35LaZWr7lYk
4zfhfQFvhYAAWVSSk5gDuGnXAyAJtxP6t9A8eBgniRfBHSTb8yA6occjlidWQcP4NvHKGpcSUsIA
P8dTSoA1xfxDxN7woESfOpkucujyEkJ/4EizPPpnW6WzuDvF/mKDyV2E6Tgr5Y31j6Hb7/yLZTBm
eDikMsyy31vHdanMShc+EcuA+d8jK+CviG2f1PDOLkc677lV+xLND3Gt4E8DtJSD56fTSFvQk4mw
Zyhjl+bWVXuY6WqZ70kVrS3eF28kwRUYysB6FfpSdP9I9vF11XJfVi2WhirtKFQLTt/riGdMzGic
R+tr69qhVEk9SXjNOE6Fcnf/XGr3DDBwhoHU0nCshB5kyz6PhAE55IHGY7lMjDPAOSE0ujsgxUVe
OD9tDy+REV4S8blcxwZF9mWm39TWxjSz2YV3uWhLjY0E4PY1SgW8g5DhhW4D1Z0WtVSbc5vwVQUX
UwR8aZ6tiYrhOd58XCSoeklLV6RnaTiXna7AAT+GTRv1HXKV6m9nGSwriCquK2Xw9r6j+CMmGZQg
js2YqQdcDavqaISqA45kO6PvP9MRhj5UtGJ+ov6fg0xqFxRxODZQjCl0sflRHsZgiEJ1zw3GP/L7
SLBoBmVwC5bTR6IIub6F96Sqpl/ZiSBq9RpwW1VqoGAUfmNJPhBDEw37ypW1yM+Wv5LEWvWUXPPh
/InDqWl404tXkbbgWm3ycy0iM6mXF4KLCk5dfbLAyiugH7AE/ulXedW430oCr/WEjucW8QwRHJ/a
2NyDr98c5cxXd2WVwbwDOD34H5TnvGou5+csBsWvwhpT6iRdbMXLgREHw/GdkC8jmcqCPbF+y9YW
uIet/D7lGpB7OAoxy/2bKwKs7ThEr2ZUhufg3Pw9/2WksOlhmd8tMl7PH0tJv/kFYM1VTd1Sy30I
iwjM1Rgo/hq70M3/Fm46d7A6RrQ9r8PKSaSNIJX30DztnyMnkMG7zZENWj8IyJTTdkdVOwzVWfQB
K9FRa0RD/gNeM/UlOXzdrlJyjiezfaHWiD9Iwm4PH1YufTydbIJOmSP9aRJ6iJdEo3XIDEEsWMoU
ytAUZgB1bZoaxbbZ6QCkWUJ40ohRL2VlrbTO9ppUs1iOZour0mTeV1DjUKR9QpxlQdn9p/09LQYC
LfGbOoXtw459+vxw770onLkQrMH6K8u+buVmUExapwxRhJWgiY1Isn1w0HlsP+5BFMMLsYrHRoge
QAUCPspie893ET66k0UK/anZYGWu7XoYAz8Q0AaEt/+rZlV477dBP4vHpd8dyuHZKbqHEAbaJHIg
c0Oh5DLjk22+FS1PK8w40vnM+dujeuc4q+dHDLxHfIwSQ0xY9wUD7M9hGobYNgFBhsX7uZEZPQXZ
CBy13v8mqzZ9yeQFXWiGZLEQKPuHQB86O5ohstgy6YI46FTF+gqdzfYrtn7pZNqGkLWyAdSrz6Yx
Xm9UGODmecih9Dx6ZekG6tidrr+txQTgOnp6HXKtavwt2LITiJYHvjX4/s9gt/a7DigIRJzrcMVj
fN+QsyJGMaFCCY/WyBzDQLWIfZ97Zy8Pv9v69D0Hh5EL3KQ251V0WOy5ztrpPdv1YVBxinTzlCuE
WWqZh6jgHCYzoI0a51KO65murXR+qGOMGtbqeK/8jabxZelO5Y2ZdK/GS8lyly6nesVf7yHlsOcL
bmTqmJDYzQw2/HvQLibNrF2E0CjEeP9uAyDx5Rq2SC3LY6mVBR8V+ig14gLeM9JudpwwDjm/qhjl
76BU8xDcEluyADehfU6YXrJPTq2XKLAXDx5eGdf3fEGzQ6t+OB1cOgY1owC82XPm2Sg0DwN5dm/f
2/8j0jPcctFkeORV2YFFX7mQBax1kBBMIvnFqvdAx27Ryoz/mNvHroYf8VdGi0AaTIhikVih5J2s
VGXsrSb/CshH+HG4lAcGqyd7qEKrGcRCDY9QXNk0K6PIg6wFD3h5/b4gioOlS6tU4BRVAbpC5B+I
iW6BErBjs9fHNUU9adGjJs2DjPsgXtuNLXibPfJFvyj+NLQp7IopwN9ztLWGfQW0FUyRUvy9QV5S
AsJ6vRavhE3jkKFyj7r7A24clrfRIr/tn8h07sjy7B52gQcAuxcQdu8+c0w8sBAt9wG60uRPWSp5
ov9gfIxX6yogsfU+ay0XF8BcIWZlc3pFusMs6e7ekhQP8NZzr3kwB7RoJcXIH2htcFftB52au4C7
XG71sq264Vn9sCyjZL17cQqPZ5NZkD8wpveR7rTSRn1qruu/3v/sZPAGtbSBvR+CXaGyLLWEuj2S
QRB52wUvlLscNWJztjsYj4JADVQITHAtgtq8saH9tfNIuW2oZ6nWR8M/AqnDE0NOemTAvNR2Zh2A
GfrdDu2cczAzRTYs5MOtthgIbKh1AT9No+xlbJT60p9QTCbAVT+fQHFrdu2jIw5X5Ky3q4NDrFSY
zBirRu4iLZce564iDwX9DKvw5fAWEsT+hhpPdPw+feh7W+3O1nrtGqj+NRq5SmvKCGUjWiJ2Izfy
HFowexlFxUMjoVotUQ41YKmgglRIODM6heLP2l6D18t319aFzS6oT3mWiZGfMqoLoIaRFgccH4ID
Doh3yYkfc03Iwa3hrhmUW3uZPPuklWsSxS4GZ+lmZ2D+77SO8CvO1wbbwBeN1f1WpF0JcNQg/Pk7
Eta1pxR9Fr1LSWMUFipnfpi65wNQPpKGu+p7le4/mrQC2PyU4ETp1rV0LVGhs3ujzrm31quqb+7d
ZhzpMxSRGUyFW94jzG2aCcypVp6R6mNZKoV803rmRv0Fuu5EhEBVMmNFSDxEbfDizu5Qr0MatRzo
LoqO5wM+0WkO33Y43FjBXfvXkHvJUCD53cWib2tANqQXYDIf9y5HfSQuWtzwC/aiT8srlWyHPYwB
dkTFGwKE+X6fhIZTHV91QBQusIFjKh4k5+XQOKaMI37CfQrguPmGbxeKuWeX1rMnzSIO/DLYWdyB
fDGVkc/bY7kCzh07kIQ62VzSSZE3uSBg6+LVIV+QZX6/z/HB+bSQ6uEJpcnQsQzNqLbhdAukLScz
q27VnRj6Bdjm8dSRnFEoKXttms2wGv4GGXRILTMAiwUFlSNWpWTx4xS7nWuvqNwdXPUKico2BWuF
rzjq0V99M6XPQDBmXBp0l1xDcCxGqUCv4RU3D0Aa/4URS6GoNrhOFDLdtVdAaIY1QjoU/gIWZwNe
zXpey8dHfnTu2Ea+zSdJtSnPy/IAG3/QmTg2Hp4MoQyUUj3ATk2UxcbHizEc+3zeojXTSqOr5pkC
LIfKzLG73N0POM5iWpm72synZ+hfUDAgortfQgtog7G/HTLICFMOloA/PADHUfvtUvGpHG9ngbpv
iZpZKpfpw1Ze1l8fa4c3M9W2+QC71Abg9yj27mxHME/T2zpz70jpsr+A5dSgvYE7oSgqlkMcI2b+
OO41lY9dJCcotAwFicYVNtMtPCzatoJ2NkozsYNqkurUfz5lRi/gE/uOwPWLwg7vEO6pyarNeo7c
d4bwmMBjxb6Y8eDvEZv/0CuyW3GujDVkU/1ZHhsEAsH0+uCAPzXZ4XzV1OAMkB3PCObVmOp32poi
ANSS3Di5ESNC6U3gK5Q4FqNQF/JqxYcrcFFQoLGHaEkbftWH7eBSWSu0NCNIZF9BVQ+MS7IB4TVW
NwRbp/5v/SbvFPD9ens8NEFXE8sPvQTG9yVlCsN1dZBbAxlvJ5t0VD1apKssYpR3qnOMPUlyMWnx
Bu8cOB/lLvFZGG0Bc4UAc3BM0K46fHzI3r7qjQYrzFQsJnvj/zEJaY7BAnJJFN84fUnBXKO1F9d1
HDVVRGp+MgIv2UKQAYEM0BQiKO9xgb5mN0yzXoTvsT1Kap1hn/s7b73JdCfT96f5jan2CnQdl5b/
rukyEU5z9VXpW/jedbxlfyf2R3BIQEMWAUJDmoAzRkWpMs+qZgOCZNpr9RFInx5V6NBKlszhEYX0
/h02+oar7u/35Jfza8P442tsh2clOBvay42Byj2GAr6EUGvBCkvi+ptEr/df+UGJCsL5nr75Ggt/
oO7rXFDeZNH1icY760x83LVoNS+qEX14mBIjbLacu5VsupPCPTjLHEU/jxRwNe/NgPaByrzH1Gub
Qs5fjHXKQ97C8uOQAcTpWbEu1Gih+8+7JGvq6yDPPqeO7/LdEXsUOoZjpZawB3k6t2ydWh5UFp7Q
kPpRWsOMt2pNc5MZGfwzhep05pWbWnRKbwLVXm1uuVz9MnVQlYGwxqkoJEOcsnWFnGw0B1iQH4O1
cEWbCOdurmQxZLS1uDyu2v66mLvJHhWzomkdaG/stE7XtXQpNoHyeEWIA3ELi7rMMlQJf8SUC111
leEH2BlBlut9gHMSWQGkacwHF9g3FlE4KgM5XkiFoOTb38TrIlv6G7JJLCVfpF5Ztf3zPAIU2sTN
3HjbgFlJlnqB3o+e3+dVcanTNQinEnC/Iw03mHbaNLxW7DYi6cLsR1i6fPFc2HX5QIJNZM0FI0FK
KS9kXL8O6AiKaZ0+e032c4emu2zaN3ZW5tvM+EJs7q6FXkoXEcdWkUnfeKOasqwP40UmAwIAIEC+
i/xiSGLbzQNslLlnsyQlCd8bJhnPHXB59cKXpT+6ywrKxMLywWkWbbST1YspdaDqa7n+tIL8ip3f
jEBNTfbb/6ESX2ZbaZ7KfZdpCtDwShPCIIs/wUtvoNeAKpw3rmjpNCBDnrqgKNwp4d+MnlhWqZc5
ucS87ZzO47u0rH4Rj/HR7g8pIacflE5YtIf0Ow2dVfnzgr9bhJzyTWNIPHRuxYoTpLsyKXNrzJaC
I6z2kI4Dh6ig9Dp/eL6M/60RPK6sZ5ftQwHEzFZWYt75IIt/uILxxpC/HxtqJZhuMLD6zMfej7et
3PsCpckhHsdfVZi/60UWslgEHqtPIYQAl9Lt1Z6fpEe0FMS28lGQ+09IqOnr+4FRS7DSrE2l+Hd9
KurTXPIZ872yRITvC0qKNIA6P1uAwVAA7H52gGeY+X8ULVPnPWsqucdbAhkvJgTkOb16GJrX1Fb7
0R4k6L1/FvXrKOUINRvAP+e32TMEeGhKneuEzghBPMsl66UnI0NSqXyg/EHGgL2hs90fu5FZNyyt
7acjOi2GUGur0C3xUYKitQ9rDz7N26nNQTwIeW8BTfIXbg+fKZH2OykJzro05EYYBDEqIg/1bNrK
oL/YtlB7EcahsWGO179bX3YhPmIUDv3VOT/Q/hcO6N2/nJOrC5u0I7I2L2fToCzwlsV5yOxL3+zn
esvKqAMJdG8xxI3CqP9EX2Mqmhk2qL8u86l6jUqm4pPYEyvqDB1iXq3VqYorHEigvylcZ8wudOK2
TlbefbI5fIWo49yANBWDHOe78u2y4EES/wqmJOwIdFAwwau7U3nBKpditcnJoGNpM7AtOvPR9HUx
1g7lavtEgg5qP+8b3jkfXzYZ3EijvvEZ0WlI5Lg4KVWOK8xGNEEuldV4qA+3NUSKK4AgZKDmpkjc
XA6suOnyhoETlUUZzg4lv9kRDiZCFcqsvd4qwlcGzPxLs6cUyRi7sbBnB8AddNlnnZZvsCsomkLd
HkYnB9WCiioCPMKXuI1tLnq/HSNUPMoZOu+iM66vq+jWP23Lx/SofvHFsL8nSjqoX4hv+PMSsbnm
B5P856wd8Oqza9DhxxfZURPyYtd2U4afRkLHOKT2qRlk16VVVtaGAWzvDqbNiocKjzXczARmnTyS
4KJ0RgnEyzDyT37Fp0M4HDpT77UeYLYkzRMuFDt1fCEQUdSiwyJhn3IRda6yKM4PeNfzwLMGdpMR
lj/3eJmF7+6Z11HYnC+hmnKNE3S752L5Lxm2RcUQP+d4l8UBmItOBv8oHrRf1IdqJSWJo+/7bDoz
6AcqZVxf7WqTuyq3ZrAiBVei5TZUXN8TnwHk+YpEzlWuOCgKfBCjd/kMqii2wUQVWmfLDjqQs0m1
EZdjh1j+MbzDYzbcLFFcCRdWO45Wn4iJalazyxihjdeDwIVeCrG27fcSKMc0op4Vroc34kEHfjK7
8MgM4qY/QW7YHbRreGMWKl2Iurd2f92QE+A4h5HW/1bqG9MbNdfiJxNtl4Ewrz98MUHjNfguCGXh
wNKLvumKD5GPXl6v5MvKQmZLnSGU5M1AIKoGEsQM9P1rvpo398Obtz0TAKVO9VhAXGMCcakMG02B
qcqrkHSl1P30rjZyPyrmDYZTeeLiUxUOH/bXVCHlSIwhgQ5hi2h0aYHG+l9mk9yoXeJ01ieTZz3x
EEv1BmJL6IRfZ7IHAqs9h6tbF2D9S2RF3yw7FcIO/4v99nN6BzSef5ibB7Ed4Ip0LVDesrPUiS+X
fiv1fhzHO/XIibK0Wh+KDinUhQcb5cfFAfoAmH7cpoWWyc8dqHLbT/CvMYEfqkNg1aRZZ6itVdDT
2bnQgBCF0MGm1QqpjUhE97Sm59Bz2EgT4pYJdJe1uF0iYJxz+XFnRUHfVL9F3wQuLlrGKTdOSTJ1
lEfDi1Swh7wxu71Pzggmf5kJky0JY7LQSUIPAe2Tsq5e1AamFIfNUMls2WMEzV+91+9UNyQajjri
KonyRT0ZhUlejUvQJuM2kdAYSmrGh3VBjrNqcIA+ssxivP2LnweS9o6BvINtcKLtkedzb4xplfTw
O7Mo+053ER3iQRCDuuQ4SdpSKIG4Qe/b61fuGYy2lORjxqeMfkHCjulqxpGWW6HD6FQi+unI7QQF
AZKne3hkHj1yUdREtdZVbvHq5j2j0vHJfgEhP2MkEQKLxFDzjBrjnH8Qj0nUEPEbxu0rnDr1Y5Ck
oIHS2Pmp0W+wyxbhPyq4ozJwlVonnlPYQpPGj24vUe0az4R54yfJHsoDUbvEWF/UUQeetEUvj+l6
0oo2T3xWmga+Kt2o4TZ1Z65qUnDSlI38vMnXdFmyHKwkUlTPx8A9r/Ujnqj92Li1bUAS1370fBO5
ehCHhU3uQUwmi/8Cc4350NE4FARlLeiBqtLrvFkss5IE276R12TB8WLLv4xAn1vVDwQst0gOtwxs
QrhI1buLOdn5Kk+EKKm7K0/PjJLOsKAsuao7jIp5/DyDRKW1keitgioMrz9QXWq3aq/8U37EifSE
jU5ZorCfzAFxH1RhvTe5Ls0j4tELoxIxEkAKY4vp2FllBK/g/A5B0g9n5s40hQnVBi5wa0/mLpbV
0PIcCGZar3gckWXja4DzTgRT7OzDkPadzzTxGevyBuokOl6FiKpAPqZye036M8g/eXbigViFcN1S
HFMBZj7uhwMLn/N3fl2auhG0ROcf6qF54KQi+WAJ6r06MZ3gIFMtckQC2VyDNyGB9skeq3l3s/h5
hn3OZHAo+zE1lXrjdEKE2zV8hhttzhRkL45ld67Ji1ZbmjJI7X2a3BvhIVTfsL68AdZY7weOo5q7
tJ60H3MQamp1PjPLohJqixWWU3TX1pT3UDZ/yQisrbsfdi3O8kbfrw2e7jJUvzu+a5zcDamqjg6b
OR3vZ/YatmSXtuFYTpeY8BTivwyJ+DN2Fpsp2hA9mZQsQu8FJJlJSCveoBToc55pJrB5mzZtksv+
WhcoU/a2aYLi/qlPVGiGSp1e9rXWm5wXXoUZ0s61uCE5/kfe54c7Or6bAQ/+kf546aD/etJKy9Kd
A0ePIwqZaJQk0xVwd2BiAzAeIxux5BTy7Om12UL20UepW9Cy8Y+NW086dld7k2DNX61AznDL/Byq
a/lJgDh2HevpkuODq9yEKMPdVOJDtG6Os0ILNttq13jW8+iButBoShbUeAq8a4+nPv+o60GynWu2
WUBqK5tL8OjcPysXftqYHCq1o3Cr4mkA19EZZ+WDnsXkhRxlbwtD/FgMMJOZQqWoXrVpDvS26I95
jAbDsJolgSsTPixiZFlVuCAObHYXuD0gTJ4iNwvBhIv4ZfUj8uog1MCrCuEWfMhE+R0bhRaYj7rH
cjWg7UvTQsvkNdE0ElfWwL7ol6O75Rm6qi48pczGHDHaG7IDS9S2JIl5zIecd0xtYEuLBA0GEqYU
RWNYOfI9inScxNguPcvnHyzNkyjmN2tWcZDPIMDeM8lp6yq0FPWPOxW91lmzLtSUvhpbh7Ks79Sv
LZ9QF2+rKbhOeNC17dpXwbagEBZLK5imnVHZgih3AgCMXDlYEcfhObw54wsy74b4crsgQi3IZ1+9
zyNsclKZ2wFKxcCn7MxrYFQvgppVdaZt5zSq5bb3LITuG4+wjawBunSijfbBeZt6QqThDPci1jq7
cvDfDcVQNhOYVSIIYcOF1IEwuR7npPHdWfz0tBhU8eFZrIu9jYAX8F1eNJWQVOZv948SRilEDfnH
CFHJcj1vTRoADUtaMB5eyNBth4dA8nKH1hau1C5tFqHATXqQjLyxPIZNy9fOsVqQldAffu/pF/NT
7ljPuYTyNEXnCnyvL8Jon8aVYPdIXDglkvn9kaiZ1KKKQIDia5SgsI2nLb/ir2nFiieMdONFLJ9B
x9qkoUcHHc8E1/oxSl1LYsxeQBirbgQMAnv43vGvclozTK9Etrf1FI/gslTaAGgVes8I0IiCyrvq
hA1qQpbTPDQHYeAKwmEFYVebdOnKBpJkVPgG7xxAMmdMFL+V/4GJr8kiek8c9um8uESE0Hq4f8h+
aQV70LgE0KNpEgSu7XgvC54MG+c8HgKBZEO9ZJvAZD8O7FrUV6tIDr4Z3H1tC8HoQqkF/u8qk8S5
oqL0dKmC5Ne7gyhoh8rfXElURnL+X6NsPcerx+F5ciXVqUMYNX+yZV57KnbiE0H5CtI7WdsZ+YDZ
Fm9QEk4ezf1NhpwREMt6Tp3aSzW4L7y2SeqDRjlIEj2OOYXmXv14BkeOaT9sAtvy2V85qL1pBbcI
MZj2r8haev6bt3IMCuySKDvDnMieAc8p2Rpvpibsk8W3DhPK0SKNj/vXJHsTgfMWS20dIDM1gnB+
pSSK0OaZAEpOFnU6tGP/Q1Oe/rz1GIZsCv2cr73Mrn/+WxgsESJlWJxph9uAefMLuUAvDrdSHLcE
htff916pCUj0wZjm+7cwnx5hgvdqN2FZ9syZ68FwxzaIniVHwdZz5Xglf2nDto8JU7yWYoTwCpDR
EBBmvwD1g9ygMweRRPMFd1yaH51MsdHWRp/jBc2vviHd2ZgMsWifMeQvWnJUoaE2cmHnPq1C2IMS
4Ympk3+e6XnzcyYMDyujpKjwuVskcaDuDtxluSc99kaboQmTsh3J6gFsQQFPuzw6jO3EvUgPZDyT
rk/FBBvHMTIcb+dwztQp6Y+Aykz094OGG7KbmILmA4LO4Zyksb4UhSGxWPVvsuIv0AwV0/xgKHu6
HKpG62FM++U33kere0Ka4Zjmroy4Yg4zi6YEPmv62Exkd1LDaPsjsnMdbY+zpdIKZEe34WlK8UVT
mv8SRqcSeDYd4rldlyksCE8CTwbhIYC+bpcgDvcfBv60NKkTApL4gi2GuTshfJl0TAe54edrKgT2
KTxE3r+cJ/p96zPr7uV46o1kVDylnyRGA2tPdTGER2wDecI3MWEIZc49CsOE3CYF/WNC1z73xWld
UgUWxc/WOxhF1HfviYVSfWh9ZuOqViXQh/ecCkbz5paWEuWH5Dc6qLqZ/V7RNlqkEuKB0+Ggprr5
a4dCIMdBzbdOys5TgB8Jnp8hcGHEA5Lt8nBMZMHzJLipikkSLy3o6yHRqOw08xW5kFqrtX0/Bo2h
fO2LyUvqACoUabHgAw6xs9MTkK+sECHKprij+wHAhjOkODXK3o9P0mCkwTYEOVXLcKsuQAZ0dk5k
8zDBCPFPYsm94m9QOYDKqF1EURFU//6JB1CJczjrx49losx5+MqrlRrW4O8w5fIXeYBPGv3vhoK7
RkfRpU5dSYg0AWcaEIrLhcRw3FQe6AmkT6kfUeu5+5JOf2vXGJFtB/qZyDXBgwAjlwVd1/pKqzsf
EV5AvVJshNZYQV9c/x3OCwvjcTZPgRMwmvzfOr4oH/Fe2FjlaZqL3sBX4xe1my6gJOBQnJ7uvhd9
MPBvJzH4uJc4dycAjEvFHahCDHg1gTSeIJFhc4GPK+9iN3hfVx8V31/Bg/NBopO/EaZ5K3F9JN95
o7eIhYKtgSJdApOvHazIrSy/0S8sdST7kZbpr9B7CCA40CDmw9JsohoYI3KTKxMNfu2IvzEZWRbB
uQAcc2SLG5aPn/AeAw1y/dw/4Jui1e/nQiawfD2kbXyj826SA08fT5R7ZbQw+OzLCk9NMt0F/xlx
GsOGHDqkxXPmv0rMZ2yv/mXWzbCinAOituMEBumchvL3PL1jQfgUAbKJDlsX01Mummu3IDdCIZ36
NI0YGy1OdV4arNs5GWxMaBJYD+xsaXx+G79vseErpoOu7v9mBAJXIX2cpZ8l0M4c274w61zV4bGv
c8NdV/KUGlrdz4/GEtHONdWYMp67NVHblCE1Boa+Q/RbC9q78cWTZVeaVr5g2Me/QypmODetL2RC
vNjHyN6Cvuy9h7Jf6syCmNEsDNTJbiR3R1E3u4NXHpSsUOHtk87Urk24zeKvmYpZwtGBoi+NMv6J
PjJOz2w3DdkyWSxL8uwUAWBZShp04c9NQrSDvI4QDmXbYtXXZfKVv2GhSmAF8Tnsb2nk/IoCFYwB
R7vxZaut8BA8u25P0qdaDfAhHcjRWF1lyQVx1GiIAIAqDTX1FzHQZg8NKmK9Gbg9q5LTHFPwtEdA
SzyLLVi22tK/yxU+wUNN79Z+9s2waZOAq3r2HEEwgKfttct+lnJYGONj6HSlvBoFRNqmPQ97pNa7
1TtWbE2ilqgMgNmcRUuJ2YdiVvzOT1iNXCVgeM0+93fHOpSq4CSjBhj4YZcPhJSv2Y2FxCR2J+Go
W6cJdMPIRrD4NHiJ1y+sUBw6pRMERjLXuz03wh6qQAhagQ5EG/2eM4pfYNd0T9VQCgvT1JGgejxy
rdmWepNRZ0knoazLO8doPkPbULi6KVZZfSO7S7DvA0PfaH2rV65ajXejREEY/RnDqz/pbukURp0Z
yqvtBbCxWhYJWA9776AxbaIcqhhMQCbz1hbIgz1D6BOcYKQOX2upKTuA3Fwh11CU9Ru3biRgCaNg
fAh+KBG2Ci0sbkeh2ktzwltjclDko0fFlqFh6HVloSLM3+5R1HIkVNA2iFfNAoSkn2UBE2moriSW
Bx4SZBiOFAipK+DYCjbc3N9Mu+dsWGw39Jr67xBObiw7Fh0121g61fnkk0+cwZeUHTl8zTxJdUgl
A41uelN2XtEBeaFJGURuJ8X54ChGhIr9tI1hH9Mtxw/1M0MNSjl4BXavXNtnBZwUZbv58i/j2wh6
4x/Rfl05PlDnO9m4fbpsDZVBDCBJ5Oycuo3RCRaE1kIKUd3tPMg3XVqEfGkEcmlolbIfrqKqP5Hj
2daDLXiDQPRXy2PeoqkLjePEIZtIiqchLIfn7eHUPHx2f03LD7Usi19717qPs2N4BpOx01jFeYXE
8YCJz4lnIXK5dZqW0CK+Gcli6UoYDu4YZ7YAxHIa/aLIaOJyUV2p0ro5Ih/4Eu5wVYe6rPd0jLS4
W8mivvjl7eYsO52HjYnzNBPTk9nAiSNTKv020RS1+efgMXmJUPcVFdYml/3Rij3SKgvdjKPDfWos
KmKVvS4coHqthsRK+LCXKCjpGBxOI+DdvhDkVVvuQ9LaChNdQZKjhMLkVFMq74uEAUQEG/8Hn5az
/PxU05sAHQ/G2Qjv+ECIyJfAGA350jsBi1l7+R2aGs25XJyP+vq0sz8TxkEB+HFZLez6L38dYjLW
2rTTzitwJYcnfbS6kLbvDrMUWngE76/jgjnSJs+MKn4ur/bHDylIo1ekVSkOOX37GlMQIn3SFl8G
PV1akjUKTJiuMQW3Fx0mZqI1fWUjJD1l4gcDjFhzKTxTDNuAh4za723vyfakege/juKjpRLUz9h3
qS61Wkb2/V/h1zZap7xm+fRQnOimsI897vIuijNIt3CQfqxHPJDTuZRJ8DxtYwWlJ6nmqSegBHGL
1V1Na9wq8SWMU29WRLK6aZ81m3Fr5BhSqMxq0/uRp/vzrFsQc9Hcm5G46rqe8MkMZcSm2wAELTJ9
q0qM1H3BL9pw5O0Je1buL0HBshhnz3PZgGM6qScMxXAEUepbF2k7v2Ya/ebC4KFuuvsHdQe7DF2Q
nnHLo+imgGdFCEmQ9wepg66KYkOEMPWVI8KVsENhq0bvhiN1LzbrUSO7mbWUd+a8aeVCwotINXk8
Wqe4+hkhg03mSQstc9A6eId1JSNm5mCstg4dd6YK8weiqgup72pVOTEzF6/ms5KLv8STqZPvHb9/
85gQ3NaGBAq2iQDEmHkuvJhR7rdsruYnQClDSr6JvMHGh7OxihZloSMwGSp9uwJCPKPYM48fgNWd
I72owzy9jvwnssIFdTa+xjULz1ZZnNgNque716DnyBppnr7tx1UgoQ+4E6wdpFxKG6xIoO2V+1b4
O/kfLIhEHb/oOSCC2DNHsvtdQw3XsTqfDDvvQOhNfVxLN8QZMtFQq/CbZZRM0AyrbHzPYDw0McA3
hEWjcZoPd83F/W27ohz6xkMdqiK8wGaIE8h8UomUQcKfJp4MziF35QzuBn+z1bDNTKMJHtDo+j6B
xSDlsBo6td0GLKKxZFW8weFOo/xHmSfPxJJj8Ttr4WOBEsCL9XtNvXESI9fM7XKqItfam/XkTvBe
Hu2bMzM1RnnF5HPaegiCuVgkbXOt+wJ0BpLmY0YLceeLW8eOttbfB4uBWRRepExU/6UkH+2COmn4
8R3LJeb5o57f4+T6PV0Lcv0hudyYvPb5jeEHaXQX32/PQIt0nt8KuQb9y553vmiszxRV0Znlm+Bi
yW4eJN7FPGrl4rLLBap723Nj/yNZ6J/MANmc3h8VjpW9fEBzg//mVIpL8tD4QTc5tyate4cx4+/o
gXeAnvXxXjNPgqgTWA/qAfCaTlteEDxHBVLKnG2X7pQAGdZPgxz00WLAsCXkdw7QmPufL+7EnKwj
lal0EENSwU3VyKcn6BlLn41/yNdZioowWKrS0/IiX91MDmEFkudwB/rA7wSHR0HuLQVSfFEZ0PCp
qYkNlBnCz8yz3jx/IbNBBstgPyZadif0nJxotXqplh8JWUl45F8g80fPMScMRne1l/eKHU23dw3t
t23VLe7yzzil75dR68jw4UJ6HqGnMAtiPF8CcS/H+F3cx3I9NhxwMTavEKMcNQ0RLRnkhER5t2CH
7MKsN/XsoO75PxT/zc6Q1wjpMgHJ27b5BWCrt0kYTxwsxhO7ve/4vPj09Ua3dK8W/g26XmzUi/LO
lKk7WtS6ykf6MtEcQzk4GGjMeJ0N89V74X1Q8TX4jP2PAUn2MTXg02DMuhAkzVrqnhIdKvaND+v8
ZedtVdpCnysj7cnMc8Gu+4eKhyXXff2hcmOvwjBjuZZ40AyzfsbRbLfGoQ7VszI5SNUyvjTcV4BH
hT/m9nsbF6689vOHwZ+zZC5ivKkBnQOOsM+30bdOtBYA2FWO2OJiBWrJi9TqZsjWmmIri45c8swi
q/twF4Bez1suIQQnKLadWl81BByPM/YmBNaLTUyNxI6ytv+gNcNvQiYl+VdZDx+kkuR7oCnMJQ//
IPGBsEsYtGn29h0kyJ/8V7ZdPhehBtPtYSL/T8wFWDz1fR2T0EMSs6acBYve1yZeUZQR+xGY7C2z
dKE4wBwPd45TdkQMBnzDV12K0onnTbGu5oE1SM+xiMyH+tJJG8Vn084upkDjYqjkaWX2FoVzQaJ2
pOLpzP9pyZS+8zVw3ntzURQi+YM+VHL0ya8dHxxteKF1xmUCElgnNIC6GFZxkMskcjQ7JU6gsI36
54K0uKpegP1lRsMdy6b2gsZGPyvZRA3W84cV0TAkzV0Gn6FJhdsGE0TjnoX75bLjdfoD2X00uyF9
LCNDSdHEf7E4ANrNQ92GypylvJgwlVpi8IQzHjomQKqAPCFSI3yABQTBP/ETWPkvCIYL9zD14ySV
td3RakEd9zBqtM9mLbDlLeTb8zQgwwQC2iRl4St/FbQRCbT+HmZDCl1qUgFBE7YMcgkRnUF8AmVs
nNBwsUFSVG5y/4Ardpm6I9qOXDxXjOUthat+4O4mUsTiPsU9ckcMP7sW+zxY9G/2yeF//1Wjavb1
QDf1GxLSes8T+Lx0/41BCHzSGBhvIg+wL7smJGhP1YWrXstmcb9urjIhRWL9Tj/Se5D5NEg+NSpR
ZylmNqME2GBisImp9SBpEz+n6HMPe6YyjPRwtss6dGVBNiiU5JHS2GD4NmJKlZkFnIR7yGpdTRGv
i9urtlHnSZPLtx9nW0awu6tYnbQvoEXLQvBa2ronIN/HLzJcWpKIZUdR4P3lJSZTs8ivBofa2mBu
jRj1gHC1jHm+LXCpTYRH2JU6jk3oAKzsgJFgLoFGc8N6Eo3hG62seD6BKzOtvbt6M+ZpoC8JTH5T
nZT/2S3nOEpcAjrKDym9vxaitiR4FG1/B6UOREITKT5NedZ2vjDHmISaOdhiqgB3TMyUYiJFUqkk
BU0dWGZzCmpFu26QoGiWn3r7gvyzeeXj0CO8m/GMZFiQR7aeNVIN+0emLTMF6O3Q1qTH2m2RP53f
866I3UaQ+cvVo9wcfrjtIpKRHDqdgukK/g/e/gMYxSSmDo5oSMdsnksGd05JVX1PU9Ciirp4YHon
OPt6+d0ETf4BftZ7W7tKwNUJg/kWILKLbb7S49pAd9nsk68qq42fUZ+BB6heIhH75oRRtVZA9oHd
McxuklippXIX7ZzEM6v2mikJDkyzAyjP4Q8un8ZMEY5pVKidHEpUSjNOIwpNOT1/t72kL4exfzSj
pZ47zcDXiZLjq4dzzGUKVdPN+7eKXOc67PQ0+qQD/s+ritIxjKloRKbLBPkEjdooHa/hPHDKjG6e
f839G9sxIDji4EKos2g5sK1GLJHrn1dOyH8Q4+Kkm5Mqdm6DEchUzuiCpmQxqOx9MlN5ApGky73A
jXWSovwQBYWAqxlj4Rs3IZh7++WAScW+xBaSIS5CEMYE5YF9so2E03Nxeboa7zxMzBQSrK1EPaIj
NtbgTU27Pehn+iDqskn3nT1brKM0z81bjw64E34psmKN91veHVnnGHus1Vzy+OCAm2EwDojxJdbl
OofBtyLotQS/eLfPkNKDPCLb9Vg/hxrdlnNNdJJpcVNDR87Ze2aN3OT721icuignCJlfWiJLocm9
rdMA+i/497jSGAi63CQTbHcWa8wmKPszuqFNrXG7aaZ9cbqyaMPLXCLHHToKtmb6yK+vxKGjL9x2
RDvlsuE4xjhz8x/DGchAtM9a/n6KmGaMg+yC/gvrVFOaZTU32UaXRTwJ4QClihAILbCmu01Fh7ll
uOiGBU6gxIIH6NxVnwi80l6HpRfs17QLSSczJZ3SlUhhTrkGG+urixznaR5RC0CnnCk5kU+vRt3M
+L+MSBvnzA5xs+5pbFGwFtghPGT91+aLPxmHr1u0+gluE0U6F5odLUozcZdxZY2L4v4FUaLs/kS5
s6dl9J5QuWTxyHSvrS5UejChzrEXGGA8lYZXeW8njIkHvzAPhbuA61xIogk3/hgf/FQjArIA9MNk
QiEVrauTujofi7xi3iOgRwGmv/18HyBDgWzha/dheJM5/8Yr9ItRv0Np9poem7te/sVsYS8J4707
0VWYxHfeULDnYqfMgEhtnHqxdn6p1lVOOj2fk/8EG0oiMawLziYYM43HsTR8bgQuRR4Ffvmr+98b
A+yxROcGsqaWrnhurl2/JRu+DSvekcTm3oNtkQ4EWwhUpv63lFv++aOpm5ta4g2/TvAQXaAXxDcz
1sn8cEGRuc2UZ6ujhZ+1nkszXiQ8J3AQ3AK5/kndUvI2CaESFFWkIaweaZH1IJXO1t29PQpgLSDt
A8NHRSKEjv9JL5kOPv38tFiaJtJH/CbzofifvBV2wr3u0OuVUixbAULr1wHOIAhuJ5NzaXPowuDK
SoGE6BvVyJZD4ACP516l3mye/vcEVmAcF/0G4qYoxRYSFZJL9jRKAQTsNgGrwHtX9LURpNxTFcJP
6vaOHeUjZnR9vOqdI4sZjEUlt2yCTvFgwex23LahJcyTR6VfppSMXLzEENGrFPHbFPhX9ux1BNcs
pi7hbUoOlDfqZADYi4HrALFEt4yligf0ynAhT2i8Gw0b2xXbXVcg4WtyiodtDUCRdDv+JZ/ml/TD
LXCISpuv3HyBTi2sIEmBqT8AQ9KQi3013NHGO+PaPP/BEC1L6Pmk5S7u43X11GPBzjtJx6RLq6ts
QzcLGqn4s7BV3jCns1FwvE0wvKs40Oo2eJQRHKaUsUmU1qDV5je4lh12SXW+0Mn9dWI7ufUdJ15W
m9NvWzha0x14yYX1G98qLynV8jYYKT+KIQo/xowJnRwTs3GIHWXyeNLUsCocZw4+ZUWAk+VQeSdI
Yq4UtxHQbU7+KrnYg8PVOGOaxYJBxh/Gsum7I0m4uTrsr1fxrMJ5jQ2EgoulV5MOyeKAFtWiD6+f
gjIXprW5X9d/38Sbbky8XltAxub0FY7i8V7EeydqM3uTebkJIs73TlXRvb3iboz69qjoqeNRE0E+
Fsjdf7KWYYrLOy2qmgDh0+A/cnQvFpoLpWt1IQ6vScK2GhcTbV3c5xxwPqgvXkxCMcPnglxiaOl4
I9GpqUd/XAtJYtFUKuIfJZdtATD4aqJG0hQthm+omcE/eZuZN8di6crUK5nT3p23z8Ldo42vLH08
64sKMFMOrvjtf/GrQuvlAWnVoUrZShbLBZKr58GWEbrJHeMiA/oXxtmxfgwR3/1d/7BIpz2CcPoP
pvtFPe1Ge+9XoIYlvwsH774jiS+X31FqnfArWoNsildzc5aHVhTuWOc0BlEYJBea8uuaNvxTOQlu
whrajgseQW3bHvo85ptrJ2J/PgSD8l/CWoL0FFlfOvC4GwbIeOSWqQHuqhgVYuE5+LEcsmpT/3Nm
a/IwHQ68rWA80GLwDU7pv/BFEV2sSWicYpZ1tQX5cv2nlS3sR8KsO8/EijLPNViril5wI9T2XX7e
J3fSTkzDe8Yn9UhA6LbJmcA+Y9OEnFOCgSCuJnqZk0NupGg3yhbRcfwya5Zdenl4IeLF+Kr57DmJ
1BrmM4YQtC3rceVnLlIWYBCteqj1Gno5+ib8XjRBs0TtbHwIXjrg98Yppu1zjE6EamKkxfTQV9fE
GVbh5cDWWCPLvo5ZKitCzBuBx5VDBuWYzMfxNSqJuKV0wtMDk1rtA6QoCqC+0he7ByA5wF1fwich
2ctXcaaHgP3/uOg2X2mi+RKUVxl199sjJwJEB4h2VWUt7erYhH5OLBWZqhi0tC0RaYDnnrjxj4T+
L07Vbxv08/ALz5u+zThZhR+jwvLWVqY0ZLXERzF/rotvcYV4FTjUSUPJPyKnMsdd8ESf/hge3HKL
V1+aVVRBKIGid4LVYvoIkmZl+5gKm+R0bwrVMQ7XOj6nMC6gUXcr2vWaBhj6dTiQrcCwzybeaiP9
U27hKntquAHX3k6skRbUY9YSxJwUD048jRBW5CGtC2U4ipUzhwxe0FizOLXvpOO5t7zoSfHdWrHy
mgYs78kK1I0f+SSQNS8WDXG1aLP1DMD4kafemva7Xcb3euatzxoqVq4jbk3MA08pd/3vNXoMAuL1
zzI6dYgj94GxnVEy3z8TqsTk8atF+9dsFUcrrhcsSXX0zBDupY/mNaZK72qVlrxTbtWRY5kpBZiG
M7f9a3q7lZA5cVLGQeOv/HEWzJu9/qgpskk07Po629a+JdjNzbTVU+m+ghX5UIgx0LSUsrcby5cI
W7QUrMc3tXiUyaP/+38KEAjMVFaiSvva+aV31O2dZUaF7drHKbiN9wfRV7n1wgxZGbiurklFvT3G
z4IBpJK2xF+j4HXnLUwISAwXUalIMWdkx5lJ7QS5sIqu6It5L6ejB/iROj5RpXDI9+JDkwpocMQI
SAOFqHggmkoaFxpVbvQc4orTixsZZ5N47gWI4BBS+F7hw0CGHWkIMZG3xVofJmkASZrC0HtnE83S
xVqIm4POW6SfF2bHiounQ4i2Vtg3pzb5lGDFeqlDvZ4QKZHGWMJom3PaG1bqGNig9qU8rvncEk39
f4VlZ9pwMWEIV0m0QNsY2745hWUBw927bZ0D21HGMSUsprFYHt3244PQue0QPW8ZKG9thdd0TGih
LAd0+K5kC95IEWMRjzM4m52s+e+NTEj7/ZDckGMkd3pJ1iSV5ACXqx4N79hm5ARajzkJQtisGY4y
0PbVs9bBWBMpzEtcPkxvil7q0/heB19gRfGqLAM1D9tDrb1FLLMb7hKx8L1egeTotKETXcEtTmVQ
SxALyN1Mc4pSOP8KetTez5eyUTLhc7RaaHjiCOGRs/g+maF+WW97Ehd8SQ59I6gLyRZRsxc9JkDd
ifdJ9iY1Eawp2lDOBPBhSNupkONrtdeJmb0KTSNNDjTevk04+5wHNiPCoDltZ1yHoJN4Fua6G3tr
UL4fLnjYtahIYGEID0uvBof3Lj1GoEtkgqqo/kb/o6F29VlFbcs3iVXjrQ1tUdSUQzJygKJGh1yj
P9BSWxC2SSZGUlUVDTHN99zEjiTy8Iw7wdnlMs83MP1uJ8WPEA2buO1coJGqgvsY83twCaTKAdAj
BHpkynqJMGjqTlmzlFtLPCMxDWt0nH0a5hZAfZmP3Kj1uSyRwctwCcgMMaNHr4cvDffZbqF8mz/h
VmQKPerobr1qiZ9Vypa6LZ0nqtv56KWFdIJmyAl1zPiZAeShs7ty2befO9Qbct6tM4E416yQlPsZ
MkpS5Vrw20J5JHEUNG3vhhVDzeScxxhjgvNXdmYivqTlGkNWZFXRVpmoBQRuKGihycb7XxDXhthX
iz7j6xcl3ZQJkSD66W3f2Y9PczuDSk7lHv/keQL3LHXTMltM8A+lakRHVzHLrfamZcjWfpZgqPns
cvAvhLSDFpVC3iOpGH4x6Go0NV28fIKIRBTQkVh+YzISG2EK8BzDZcIfSSevajda6l4TatFd/Ftc
9WOpXrlMLEPYECIyf7zdvKcaRCQ9gHFCr4tSJiTH/fukEjaf/gZ8VoDNoIQYJ7F056adMVBbh3el
uM1rLgUOoYy+T3bcVRDGOj8YVHeLni3c2fOAyQbz3Ja5k6BOUVWARjAUGqq7wET/KsHnTVE6M7d3
1oebOdPaSk3SSwTQs014/32wB5xOT2Um9sOJBzQqYSLBnrTTjYUtgMDJ/kSHr+P4Qq5NoL5exWQZ
cIXhS47aEyTfGU9jELJYm/8q/0cTk8feQ8aaBBHfq4ed2JIgrSZxxd0SBaymZPZiP8drUbf4DAo6
qdyVQP2rc7LgL3ol2tTYrl8Avkgcf8wROFO7XHTXKOBgrKiSV6hZNCLoQeQkJML5gI04yAAlF7ol
g7ncnwdNJAQGsxieF0qIqC6+s66dU7hPCkcy/ScpLT8pJVlcGXZTZ3f7BEwRu0rzW0wVecxYNnU6
CjHoBAKOqxz2Hain1haqM8T+t3p2N89jN/dR2LB57TIGW+x3SYWwxdpQTKopJLGoQrP2SkTJ69oc
ojxtK1wTfGvy4haphzPm/O12xEfWZVvOU7+aKFyo+Lf1u3EAxJdS5RGzOHrekX7V3R26HS2iIALV
XXrlZ4l8+RlDYfghTsCo3UrP5Q7e1/OYPwd7O9nrCpuGMgC6mtAD3mw0KnrzO0+0MnEyl3k08z3t
eY4lpNw7XFHPbTVNx6rg/K4mJSawLk5Uu70Hfho4k7dy8LUgwNFXpVoR5rg73qbAnvXIxddY3Ha+
ONzIZTEX5PLbSVOcY30rvJpTaIRYUYJI8SSKLfnWmhCmrzvafVhLrZ6fcBrpVWPcy8KyMOTB5h48
ConhAZHexxkErpZT6bx/C+XP+pKI8KBt6uVjkgH/06grYsRi6LVc4zSb/wlbPYbmzj2h/eQKbC3V
7cltOZ95fcSyCgN/hFm2UlckCMtT2qKYN4q4rc4sAUKfWnxMQWAsoBV1+rCZrVrbQg87g/yU9dgt
DLbGezpPtYxXFRbN0INfNgBfI45tnIcUenHOuHnCqxVWQaoQRH/+57BBRnqJS6DPOFwFwgY2B34K
jQ+qMG+ai2UFBZAsP/n0VEPCe6RLPxTH6gEiysJ85i1yOEJFY6beqH7a0QZ6Tr8mhnNP1dyMy2Ii
wRMVVxIFyG4VVuZ42e4cVfe0btZ+jzqzEBmUm0RN0H2BFPbp7nSRYGuz5LbkzDe2CLWgBjQoM+E9
I3uJKRie4Dz3Tn2HLVgH/3pfXL59A2MdDtXnGYLjLQVYngLS2RQ/Sk1xsGZaS/s/vIlVDJxUlan8
L055iRmFIGuN5ljoNLDvbe6yHrTJkTpkQV40J4O4tDkyf0Y5vrK3USc8M1bLA/i9kLlVb6riX2A8
fPyEHjLOdmx/UfId15G5jO2Dw0DR9saAbpXvgaLRpKuMJgt3dhFWWF5fSgzVlZos6Fuqu527tSnD
+KGxJl6QlmtLhuAqmSyZrQ9c565PlfBowyHW+ZNrzSmX5Epq4ZLJi/BRRI4Eh0avdZdJOVzU3ofd
dWjt6zqMjpLpe2xWO9NvvaDUR4H0DvyUkgPUCOsi02+244mLeXyXVQk7HduODwbPMi9s3CJwCRoA
AYPAvRrTuRoFJh1WJv9hc3Wl30Yk3uwnNw7dwWZ0Bb6XHzra7m5dwF4mxLyCUoVS/nkrIjE3hyIF
w4eGFDUMpmTVZj+nsT2WF5CEEr5pf1wm7rlUw9V8fKiS+ekKpafbS1wopz9TwbHRCitx6Ssd+ZWM
Zrs8REFOZbmPwU5XE6nPtKjJsPxPE3Sh20muKC0W7VkycBkrXPJN+Wt9zeHMTKNMkAjficyN+r7k
y5s7bcr5p4FqUrc4NfsPI3oy+jkymOa2cLGafGSLi3tQ2WyVyTZNImK2bojYdfPX3KKk0QRrXIdO
tEVYRRR0uKxoVQNyLZMOfsQyFSK0kQMofLB7uai7i8TvwZZbT0U7GzuAiD3/zZfumOHVdFaRdoAA
U0/YsWZZTY7KMDvvnsIm9zppx2nclbbs96SFR413gfju6awgUuIU0ZrqRyR2GlUeZJ2yBUtITf5a
dVLSnk5Sxn01o/34zTs6XtswqEDmCVjh9rkwfVgwMY2TWjtT0WWFx1HJ7DB8kDArHIZM+BUuGosz
P+30B1hGJ7klcy+nVnnS0EDPFiaQNNrn2TIRsrog3C7syxLRxElIFtC5bAPrYGncpdNZGqtZlZ+7
1CSQaxYX76hNDbeykaCumvkr+QX3wflhMxDbiWXZVaQSTLbjfLZR0O5fnhwkCWu+//lNhmjahj5K
05LJUGb9y2wkbNjTPk47227P5SB1B6KkWc58eKpArSlT1YKHDKwySlTC2dfyURx80Y2zlzCeUFtE
8carYg5XbwWhJ9QmmV3n3cV9KnbWu/ZUfuIF8fI7MyOHxarTbGVQioLZv7y1KgoajIBixHMGf8uN
apJEGr9GXd8+P7VkI/MTkDtVsbv1IeG9DB+WWvS+z0n77zPqeWwAIuW0Sw8eMFqMX3fJj6CobYmc
Sa46GfmJb1splmznFCbzi36D9CisZWvOLQvSCS2RChK28ByqkzqzctOKzI12ZliMcIefptGsn1pe
f+ntGoHJlxu1WwopozJpa9DAX6Hi4162HAlU81F+eVV2edIPETRNBfIX4k9CM4ADp7O5eYwkw/It
mVPR8G19usXFdAQH36nPt71jAXXK/iwwvUFrrSXT0LEoGewr3tlh8sXQWaSQTjLHwQNopDdtPnKZ
5xXV2odx58FWP3I+Z4dd9aEXhj7efii8WE/l+Ls/tgcGvAYncIihspQ0ErdPZVONIS505Nh5E4VG
OYVhZlDu0zzweaYyUtRTHjHqR7Fd8vssJSSpKF3HWr37jsPoxnfH0dAI+Vm33TTKZcbYprvP5XB6
G2NrS3tmz3pxWLxUvNppZ9A0OLgyqng+PjuMnmL6qn1rWzQJP3ZBlmNf4UkZVbVYb1+2+JxwloNC
W0s6/iFcvqkYCrN269IoDywYMQaCWepZYFNS2s1SU2V0+D2omgbclL6YZk08RkJ9qtP3Pex5FMbG
/4QB43u3ephoCVAbjc63LciGDbjLplEQeTCoHeg1ZrliEcJN0YAE1Yche/PQVkdHU5FSA67vhrhW
eRaxYVc1sbUcdeMOZ/fIFq1IVPa0i+DsfEmdVdEFf5QA1LKDvHGyZCjkRgQBvTxok/+1uiiIeijI
1kEhE0n2ppdUPrdaL3XOaAlJ1Cri9LDisJkSodP0hPom9Rtef4tq5OZNHRL2P3bQNZGJhm6oH55M
IRQZKRN6Lf+HcTuIMth5fZxaeoW82tCgk5RKzphIUq/nNrKAbwEW3hVuJ/RMSsEjYLOMzl+iowFd
fcbSaQbLR7yq056TmhXckXBP51jLi4BQ/lJXw1j6xcPUULldAHVChmp/KE7EL3/dnK2I2pgsJEDT
yoTb1ms7ujJ2+pwQa0oC3Z5VGPFnIxMCdboGYElcc39NP8qDuIOyVvMxXTwxez1H/LgNvlzv/sqf
dGAe4oU1+Uo4QTNWu7jCbW50VdO6Cz1AxQEnVZgOfD4NsYLHq8kUNcl6nzIV34mfnTc/gFth3550
GosYjPkEhkz6F0M6aUT3vk1+3CfOBcH8O8PSM+2EPVEz/kTn6Or2wMwETU+Evug7iqi6XioTdPeY
GOlIXZLPs5K2dbDxZ15s8dlR3/SYVR7Bb3Ee8P72ZSI1f1C92PdB4NXMBIhy3KH86N+NG+JiIFD/
GqLugNgMvePqvR4KagQ/6OSc/6uR8+viO+HuCUonzyvwMQ94Ihc+qZ5g5432yWvtwh+hoHZWq4n2
S7Px3KfBc9PXjy3PVDVXwsbvzIxeODsNa1GoHb1cJd54aN0CoIBlL9+mzeS5LdtysiAI5397aBPa
/ROTiOjYS31CWxu3Tmk53shkkFji43hSrYHmdTb1TQur2zEyzeRm9uioLFyM+KxDpN8PeRU50tpv
l7MTRVKtyYMVYKpHtB+1H9WO1PM9VOF/dQL7czK/o1fMcVMS8IFFwoBonmPNSBbSKmo+OMxCyh3T
asOeXcejxRFoIDd09uzoCz/giR4Ar9v7e4H6Cf3J6e+1YnA+MzK8vul1L3YHhYgAf89+YC/MSnhM
3iJ9OukVotTHqoY0ATMwPn7UKFptBVy3m1T5KTuA80xgXhfNy/v990cNFtEePzogzPDb5nwKaxpS
b5DaropFQn6a2i5XP6B5fBhgVJxh0qvM9iXQH5vIt4OWB/sB1stul2GIsDK4fuWTKdl+mwTuCQnb
/AUQ4drW667aNH4mJfyDrSM4wBVVyRD1MFmEbyQ4DfPWvdgVuyMOBtlY03sD6f9wkAj+wW8Fvrjk
P9HdME9etTKsPNH/wbTOvjhpbVG7tQQ2nzDKZiiQmoIF9CNJ8/h5vSrnl5nmgdQ1OBrT9ZEG1+Qx
VQBnuRm01hp4VmFhdu6W150XtU4b+k1WCwS12SRTFoXjXnDDP+RqF/DnsMtE3rurI4ayZF2nAs5/
0Z8aEd9Z7pdrPCHkjzIJudrcM0U3TdhkZt9OFPJhuFs6aHCKY8ZOmbT6fzHlvqVxSlQCoYaPTTeR
Kktr/NHBkQWMse+qpJ5JS7A9YFqGNo8G1OFEzowdt3fnlT5P4qYbnfy3ZlEnmx2bXU5hcFChr+fJ
CI+kSViUdVCTKK/FYZM6tBAK/nXC6KixcanbXw3duLbhn2IjvhjjUXE5Id/JDt5n5Frm0ztwUlmA
v2codLD08ZVjHwkCetbUtocPqiyGA69EQ+pu9WfN+/f4Rt1btoyRbryaTllJG8R8IHlrXuN5nrFg
sifAt7Ref6iBdGnQJNl7GGmynNr6/R09m0O5BidSshu/S0YNKEB1wR1WniQ+k5sP2i7zfrdR/rpl
xKdXYHADc8nUAgd290R4qyNjYPicxaiYZ4wMugcn3dgdWsJFFB8B4wFnow7JndACJYW7cPf+cWm7
vTdGpO+imZ0oA9hWzbX1BDsRbiVWt9Nd8aS7578GjP9WH4w5HJfb+m35pM0yYvcPcOWUMN0UtfwE
Iw+4kvwJ0DFKG832Atj4XdgRjYgbrZQeJOvkMDsqVsncsN2hFkem7jbsmKa27dhLK56o2GDeQ4rb
4hutxKGUUuLAmwAUumCj3okWByVvMtoY9bkvDnu3ej2gDR2aCFOTesx4eJ3X0lkV2Q7Vjmqn6CLn
9PL7hj3DUHu3YRQLgIrYOu6g0bbTNnhjtuYhAfdaJWv9kPB677K3K2eYv87n8uQr6n3Chrh1fUTX
Ggr0irC8y2j6aNNRoMw304BE/24E5FQ4JBFrSc/ri7ZD4/tL5pd8+RRij64gZcYUdycf3lIvxL03
T8ye+loo5At+mKNlUQbMenwwemF3KxSalxkT7A0AJU0x59KRYB+suA0VeAb6Lluz7dzXiFSWeVy+
p86Os2HeKRyMKb/UGFidMGEHEykQDqbpB3rXl9kWpyRdBJ23b1Ivq9NEUvu5e5PC/KwkkvUPQtXG
Cj8DILsUTfLimQyI2Md0KDDuT7T+1iByD9mIK5wFXGLmoBkw4mN9+Z+Ovdzjoho95v18osoS2H/7
miylO7ckc1svEG3YQZ/J4DhWBBNB4wn8yfFJXx5aPADXTlNF3xmBXPpfdZiDZbFdlNG3g1sxfSGr
4qXOyCb2ia6p032phQAzbxa2W+QMJ7FRtK1dMNLvqlG/gnQYI0wiX2Zq7hnChhOPcwTWUMjznbnS
NrS4MnJYZyY9Ba+xPo8Yayv5794Z5tXVdn/qzvIZc4P4K5c2bqzih3mxF3+7DLaC1QeDtqx7GNlw
GBRP1zzyPSffCJlXfFAtxObsUhgLYjzddqah/tupQ6c3GoC91saQT8HLQWDzepdhJ5n/oCrVCx0H
TXhUhg0pUaJuQF6Zk1VnPw1XbV4kDviG3EpiKqRRp8CHixud/GO0EoBz8uASGqvahCKeIF1oUvs3
taooJDr8Icgq3mq8l8zaLy31SHm7r/lntk1bpGosj8XQHaaHu/4oAQ5O3TGjJbuhNLzvIt2dQKCQ
6RhPUQ93F8UDLJtJ04dZEn6Jpq3wN2Y/ZGMFNbxfrnTj+amUbAg4ng+X3t0frbooxYME72OQT562
edNJGh3dIkxO/sWcfnJa1Xew4FjOhNVjCKU0sRzwo1NRCxwwqYJM7pKrReIBa2orWaAwuoZvT6w6
ImmMkCxNn56zJZvdCVPqAttYZ8Kd+S3+3PrrDhu8zTlH+Cne3I2inadDRjmo5HrthDcHmtrR2NLs
fFv4T+Aq7Si3C5Ck5OEbVfGtfid/MtVTLj3OLBHlKFAO1L0flWuwb3kRx3YAGuybJifqSBOwRRct
NbHPc3KYupZ8jxVvX1NiOC1BGO/XcjqUMfVYcu07qlTijiDJn1Pexrr30yKD4J51WIrc1Ke84wYl
BJMorkGfqwgYZSudB675sFQMLuUAVS56Wo49ApAD4nOxMREKiDWMbbbFMuqzwgP1zvSwOZYWGBfJ
/oiSGK6gEGKrvLv5MYdppZBjPzfr0cAaM5anOqauCtE99ZjcN1dx/aX2Tae2EixzdhGJ9yEK0ClF
O1X/fn/WjzJkAoXFjuyZ6U8DDtacgFWraxfZh2pTEaoHPwge9i4rfJ6CQZMQl4J3z5lNzJpu6SHQ
REyad2Aucjk1fFsbIXf0abf6Tu4jvud6fi/aVmaJG4g7bS6ZSha6rSe+JurxYGEAxmRyn5pTDGay
OiAKAyRVqcwTGzrDdu1YUXNpeqqJiW7LbmPFIwu8dxmQdLRlYnj1/bIXiN5/XvnSMmvGOKGABWnA
vmt2fWQHP0Ctv4oe7O1fQpTKRjS7hqCEVmv6gdPkh+MJ+yQVQJVaBI0sNIs2VfqyPExGqzIqRk05
oa4BgCfXSRypMVOUCsnAn5/lWlHfC5xQVVCM24RkcIYAhFJ7aEHsIy6fTTJ0bUOHyaVKtawPJ+xZ
0CUjMj+RvVEQPF5OsmpWtVXkJBV17Xav4fDOgqHTr7ksI9hhURZlrjjxMn7wqbt1tQPk6y9arM/u
FfmYreTqfkxeKd0AEN7lkxtEkMWofGHL5CMHsVExg3zus+NjgM0zwExjhWgVmcjtTmufLv7G2IVD
J/ZQdnEcVsNB25r/UIJOQvBPKlf5ezkuili5i1El4a1GTjOO7iXuqYevhfc+psOho4+/C86RD0Jr
dVrdfzSw6RIzyK1HCWDeuqEO1PofAF15hfFCs0fqQD97nAajhNDhBleP3AhMw8kywBNDDb7zaIT0
IJQHXKME7d58oBoMMIfmg+0p5Q7Rfb6sx2RyW+v4hQX+B8OQxOT6WchqclcXZO8m0xKK2Z4G3zfM
wbp62ZTlMaZ87qZm8CbPwhusv2x7tGZo4m4mv2ngOwmIoh2Qe8niH//YqJKaeU0y1NDCUWqVy4F9
e3V1FP/9ODShPRR/j4J5iGbJLOUZCM0wKmZILSTDMrZkPtgjpuDuenRyU8BtD4+IEz3RDCgJ8Tz7
wu+/8XiXjkeVzcYNFv0BRJLR7iKOrrdpOHUlhmVyCtOu/uk4bmMkezDsuvrUBPRNOQ7DMF/254Fb
lwgkSC1xNA6U9zEvus6+rZtmRknXs7dJORRvZfL2eEYAZgeYjUTI+uLqa63d9sin+t2kDso/TY/n
1Yj6A6Ti66Q14Ktw7vZDQiOLkzb+nzbQNUBkowvSUb0NZtciHOZyD6/4gTOhfluvxX5I+zz7lY4m
eoLVCp72U3CpceLIyO1XC2sbP2++zcxDcYaP2LNbwTqD+v2MyZyzZ9nHbBItR2KdvEjExa5txExj
44ryzjqTobmBEut+wBf5FmlDPnrTGRc7psn0Kd7hBqq5y0fikmWMB7vW/3esvK7kvcfT1lmgyGuG
eIrqTL6VzgWbzqDf2tk+lOjD45GQ8kCZJ46NxToMGeZEmw2budewUMn1pqs0pMQ00LbnAvKu2rpm
Cfwuto2eVmLAaX8KqW5w6N21gMTMiBAYyODUEnl+4btf0eTBfJwfcNVXOa1dKuquYOK19letxNKh
9o0w/OyhCC+ibSSvwKS5H7v86RHXIGpWgePaUaCJ031YsV884U5L9FSA20IWqD/yVX0ots6GOnRM
JAisxnhvb3DLg+vKj0hUI1wiO8vRqfhaqmzt+1q/kPf5/y85d5qglsJ5pM4qTqOetbAIy4bKnWn8
6gPcvoiuQjiu/Lg+FqLrPsyyq7z8FXQAZK4R4f/RrVpJBjXpuxGf89BMHyrJU6P1KRJoAKFXNa6X
jvoaOfZd9kLjsN3r+gFKDQzP5ROrQj7QK9PrXHoQBIsfreHQw0CKcn0Ati/8hZPwVc4MsEdQjKr6
jlv9+G8MbGiVo3KAXK1/kLFzqf4B0VzHiwRdUNfYNtg2oksp1szbJ3kgCikwqpYBypOvUOibKAVQ
Px4sLub5IUoIrAAgBoJ/o78obhRv5C5kgWwrRhI+rckuJ5IZCWQneEypG27MeWXT7xlFdlzSJW1M
06fJnodcM/XiqHgKAH+odQ9B8evB35PVCoCCvm872nLuONxzHIpK+FtuL5iDryvioAvAEPLBG3/+
Yi2/+8ANSr0hjK0altEZnrqeD/rrOfSojoaRf5hlTj/TB6+TffJaa5FEk6Ka2tE8Ggy4nXlVax9S
NiWDCJDWwv92xJH9meTcWS0URcQSQCchE6ibvLTkiqCGeWllWIpRly7DadI3i0RPnaxbXzycZ6Uw
nuXDgRL1SE0ME8LOo1DJlzSnfPDz2qTZQNl9s8qZxWM2KVBf3P5mVnNje8RSZhshk9q3wpJScejA
3slZSyNWIZ8y2OYS91seGmhGFx232q35guu2lu/p+rSKOq1kGn0THg9Dm2zX7MiFjwOrvOuAvBh7
IFuoIPULka7ksJP2+Okzke4gJp6b7aYpMkRHZ2iathWBMnvezawvDk0TcAwR0ZmNubeBfuMmKZbf
wqORgahfKN1U3djY7nkjBakIsktimoqAmnckaBddINLiK4O8CtF6IMI7PYoNcN2+kISzS/xLK0t/
t8sHe6frSdCXuPeSXlJ+eJmQxead/X8r/EHdy5b9jjjOfCk7bkfGuqeZN/QO7/mo4hc6p9hTwvz0
pgpLb2hnOJ0O7qOp3+iISKYAMObUSyz73s8T3D3xSYrmmpqvF46rOvAehybWV65hbFcylHkhILCp
oi0i/oKAKH/MxNU1PCiWQq2Fih+UH2hbvg9K47wR2mER5D7Ok/ht2YiU193Z8v67I2/+fJZhFF6F
RgTymk89ZV4cvpVO7UEfUndMAfmu+L2aU9Jo/7r3UmmX8SHlwJPkrL3pSFOr1/htkAjbKFFPaTif
Sh5v7c+0CbDMYymc18shVR+n9VGcynQ2Rq8WV1kOtQnSLly+cnkOnSMLC/4HPHKA6F1qzkr3mNzS
1EnyCP6qjjGjlzNt2HGYW0Ewt09JagJIFcajSURBuiUMwyPLvVwRMvmg9roSdVuc40Q0Ac2aFOpz
w81I8yR61jHN43BylYgT2YDYXJ2WoovXVXygAaNMfsdPRyoubXR2FMOYEay2T6FV6ihU1e2lxZb7
qJIGTCf2oXNeeopodsBIr6yEagQ5dGxNk3SVEgK/ELB7hBTe5f3CuEyba+1bUqm2w4Sf/Rno+6SR
Gav1aio3v+1ZlXEhfyETPKtOXL/NU6bLyKGN9b0CE2YnwmMGUVqdYJVZzRbFFJtEql8CbUKxB/43
bzVCp9spHInoNLJrzDdVIdk2a0eqFMPrVRTxeo7EqxWlrRKSQkKE5mYYj6vO+sqHJpOE2hGgcbTh
UTK2MKy+9EEffSStaPddTelR1FiD48umzSb6zoV3mnLXt6bKuDNlGmMVRSkHB+7pZDNPbslOqKms
0ffO4HQGaWg9oHecVxmeqEHJAuOHukdEXWq0bzN8NCI3kit+fQawqulfsu72xblGxQLqFFNhRTmF
GJSdNudYISQoWnvKR77GhVNNuMtbSxfO//ZZuZ8dqx9w5pt0PDcJUImJCj1/YIuwoWDROEzswjEa
0RfXHyMRYcBRP1hYLwiv5niUJAuAmJTXM3hxp9Nn0PJBkmQoQfh26fjAnY+X2yUlGD9hLsv4Q3NY
c7eysNAMJwQ0SMJBGIWGL43nWnGmCyGfS2xhjsXZPVPKwP4JlEYsE4N4j2wO4De831W1w4bAvbTp
KAgit5Wn0XrFCUrtsX5P1Mvr6GrR7E4xNB35OXuBnLDOgVPzI84ER/V7B8VB8HMn0QY1cDGBpTKd
Lcn+R2x+V5seXNiRQSjYZEOlq7KnXw9Pw8JrpeINDJFnfEB2EQN38yDJBT/DY9xkj9unM/+92gqY
6KTGN/IIFAie2WmQm19ibAgtGHzD07JvHhEcf6etL5InUJrDVSIcZv9gkWWO18FLScSdgJLnHyxg
Bq2y8yIWigyj9Iq1T5+28yhUbiHLKqGFplrATmOELoSfts3m5Uroj2HPRHhKkmPk+KHP2etclXWi
XT6ONpKUbvDLtRlVNspIBtNIG/xCySkfEcOuhEs5aeahbcXNjQ9FuN0A47EMkTfEZ2sSmbF/f/gX
NxHlW8q1g1mj339f7TXFSUvl/za6oSx2+OvdAuQ/hppENJ60zSIFWEHlM1M53q/9xkxc0lVfqktc
RvFqhBfGsEEeDVfOo2rF+j5ihEjwT8VIz8Fk+pvQ7NyDCEIXYWZGEtRRLTwKfvsG6x9LvuPYeD5A
7B4/lZkVciBUU0IWrPDCxcJ4bPu7q86fA1Ko/hY4Gmyf6Pu/LfDxb2hibax5qVD+XMU/j2BAGTRv
nCLyvR2wPu3qFl1QJCT7okOjSGZe9gBU8g+aUhzNu+ntvd0uwJ8w6kk6zRuMPfTqYXGudfcQ+y4t
jllXrlptaOybalBxtjAT1B5xC6uHyA43Vw/fNePOEbxwmO+wK+douY91kthE/SmhaRPpDuc1awfw
rhT4b7jafn/a6vg8GJUm0per2Gk0kyOEBHcFpWXtJRoJ9nWr6aQ2TTOmQnyLMzgIWkx14V5Xm4k5
qp7o7sm9cleri6gxnRlH+VrxIBFZ69OeiFQy+7/jAFxlC8g57qjVTSfyLCcLSseX4hgXXlDb6/vX
fvI8qQdWvzX0QTyqXJ6mu+e8ktKiplDO8n76FDNqqLD0r76oUSA5wWzgENjQKZIbHGqEpVRjAZ8n
5mlMst7PYhlNOWlaJoO7pU5Mu3Axl8f8jDlIFwyhWPglFcuVKLzgA0Wo9EagwZ5X1y9E+Xear1rv
xVwJ0Zv2CLu4VQ8DPAqT/hWiXvijDc8sgunVJCELd4qGGtAvg1t2meaQMVsHmefoT6DpsBFU/hPY
WnXDIKQNC+SGpn95F08lLMiHhSne9b0/fmvn/FA+aLzewXdds5yJE2MfdMg2//G/9af6K1QLWG/o
psblFXo7KkDE70lBtzEYSyDpIxZqWu8mJCACAA09lRuiL17eCmJPcyKbSEp3YlQ8G/O5x/c9Xofm
nPw0iwyt93pYJPN0CRP6j/PPe1cnDl6D6yjw/5f0ZGegxKrYCucZPrquRiRPoFGGEC2GxOtRDpdA
GUP7LhPssR3Lq+RYwWjhM9Wt1kVeoo5xGKCNChjJCkKlan2D8Q0N3qIyObLL5z72wRRvpPqti1kF
OGyKh/f2cEDtBOarWmFX/Y/e5PvOsI0H5OQ6urWRrhF9X7gnx6ajvXxHOMod9dgJYLOPH2zY73LO
Erwa3HkSblGOB9QMbUxMNtYPjwytGMCPWzJU5aYHd3uh+dPJzj+LLRo0hr2ncq4qZW1q1z/Ghz46
tgpV6G4+AlZoolYMYs4yvs87yki8eUIzCohZca3dXaeYE7N4E1sN9Ftg2bZ/OM4l5nko0kFAr6zM
A7FGG3DJvYA4LInzcVjsN1Uu33z+sVLcR7DNtyFUqe9ZCb3CzNhouabsns+DyDJFMDZud93AgOZj
J3VK4mp7W06iP0Ild7dOYfrAqdDGtSmyoGurgo3I4NYg+HaNzJeMXWKsaiz5wcPJi4LyQaH99q0m
9ngBeja3Qp0jiI1GdIndvQgaomy2fwyRxioQcIQAwbFk6L5A6/sztd4PRrwHuGbXLPQc9SexxHBM
BKfJoBHD/EFVphhslsG25tu8Htor/291Ee1bypsbe5Ti0iQTqmAU8q/FWPMNd9JwpAp0iqXLwR/C
xgS/pBU4VmXJvLDV/ZRYP3GG9RR1a/+o8D1zmOqCaAk2J7L+kpVeX/nxFNjnr5NqT75bGIeIct8y
GvAf+C06OVUIonbKwisCIaD8cEtKtxUJNc7PUbRkTdZko3fEKcD+n1OQKFOUdcwBMe8eR1X3ELwO
bngeXNM3AE1RKevJLxPll5EwKIbHiuVNf3DUfylcspFfInwxh1AT1skJF6lMU2md5GM2akA/y1Lm
RAU3fG5V+N0HDAJz8580sBkFmpblCaWjpqgJ9Vv11Ui2UwnTG21MQhTMs+fImyOdvpYKYzkJzydp
uyfyT9n6yQ3nH4siy4Zb+fy+7nUu4n+RswLhyJceUXvEI4EV1E8MrjuUoDkMSpFk1hkJNP1KtzrZ
ZDiTI+a9zzPYznd2IqqScyzt1En3BBSm8Jnuf/Boief9YIQ3yoNIKTmAJaAAfTJEYDOVZtrp/wJz
K7ep+x0u9qqyZIQVBKN5pM0/6ktemXVZmev+xjIzdLnc6vVzOjWQn0EP/YbpEsd64YilW1H/EEpv
fkhEusMdYVFFFmih4GIUuLi7MhcxTvO3k5DWs+bjW6HoLLaQMHw/2LAjJvwkTwAHJFV552cbmH/b
oMMTbXKF3R5KuC2BKKQA++3RBlHW0QnJc6/+q9BL0/t+3u2SHTMlq4vBJXPBbOFnJ7JsJkrifL+b
YaIXcNjGAlHS2l+O2TC+VmW04PCgx04/d3CmixoszV19/m5F1NcUniFmFCBLx09YTCVZ9/31ewft
TZzUgVEVQXGzmQaylAmvxRD+dWG6w+FfQ8Y3ce9T8oBPOrp/j/kcOFX5LKaB1p/U+jt8arTUls5d
jhR+Is2a6FGR7L1nw/JhOb4qFro+UTsKc3JhWqdLvhTeFPCUJSt+ZjDCBwF0cO+veuEVgXAOKKk+
kjMp4wu6fotYJ2+f15+mNmI7DCAUyQmEfI7TCaVITYsPdgUI8DtG0esSzOF4QpDTDGZT6pLLIIcu
Q1uwGacKVKKL45ypAbNTQXVqjnAxHu+QDHeA1FTCqBQTyRxW7qsJoFAuSOMO+itjGaN6y+If85F/
iOTUegBsZj9LHT42QKOKY29LE9fwtp3WdX8D9gGWGwC09GrJLhlbQOZRAv3uTF5UHHh15PKS7qdA
RmivMUFlUg6De/+j3IzJF+yhX/qmjGuVkATbJztzs/4GXg1VUZHHPk+W8ojHN3w5ZclRp0MScGIi
KKeBFwX8req9V13wtfHf9wfcTshn6B8/iZoTMwMcWV3TwbaMrjJKFeB92r3E36wqZACwRUMHPsTF
w5vbLfruLGin3WuHmgLXr6mV+LH02TMvF6Pqa62oiDfPshf7FMQqZJ3ivYFM8BAWS153cD5K+yip
gXRfcwqLG2oAfWASAbENdrSHxRbxW4dAwFkRgarbaheBt5CgDm8dJJaelerPlbi+DZBJb+pLNqWp
QGgiRL8L1hModdT0tuNk8c/MFP4jeTT3Z6lRvUsQJJgmP8Ym7y84ARuQM6abjJ6w1UBVmLGBECgj
V+6GtJsBNeuxvnj81sYjg3fsUGR7VJlGANsnwKgCmhOG1g/Ei1b0gDCE5R/nl4qEL8Lonzq87e1q
NgTFnRXLpMjmBSZRauc5HrwCK731QQVu0u3u33g1b/i2kgwgLF9dX2XbN/ujfZLL8kbYiN2W/VjL
2gmEl5VfWbxo6mCJiMTSTn2vc3g88SEuErbvaj8661vXo5qPOixBUFI5Pr3QVT+F9Kv97vhypyCH
9uXAu44+XegMuV5dFh4ijBNhEYAp0LeMXyiw6iurBWmkAUJZj4V5H8R039A6quuShRiObQkihfe9
a9LtgrUKHJ4yPykw+9vcAqOjnMaSpxC2CMcA/7KBwmB+4axo7ocRz0UkyCHcXYoT0b4SiNTc8+oL
MOEkPZvTNoS4TSgCEKPvQR3BTqv5IapMvPKHZDZeBXAIVehnG4IKYZ2M3ieqKpq0bZV+e9y037Ed
HRGPzJdE5604lSRQJlKeN4a5aHez9yM2V493hFK5Je8HOJJz60tGTvbrHhNEzpEUAMREKrWLyRmn
QEqYcQAESKyVPjvEOEmDq9dYaoiYqrCHQuxl5icUZ2ys/fEsCxsz8f8YbMrZd+vNbyol6+5jz8Fu
O/hBapiiwmYEk9UOSYUfj5/En1TsYPvikjRafS/Fov1nynYuMnCrsgH4+Z1Aagm2YVkxGFpk2q05
HWwS7UbkgzxBqFNHtMDxu7KIUpCxvxPcXf+mDmck6KuJA6cg8TSiz1+R/yai9mX1vvS2xEWvQavL
ocSnuRNUn8OCBisksDBFFaj6++6rfyRNZktlITAbeGPBxm4LqbJSvQQ+ey/bzJy4Z//MAtJ7tNIw
Tu3fh4ZcwuCCDmfZSox9aX+1HuvvufSD61ozEupE6mwZpQeAYMDydibVyZcAADhczOx1lSeQKiO2
Ahydy7+M3MBMOAr0Z/Wzh0gIBUsXlJgls0Ss4P6/awUqQADKbtXGzLGrwsSUainNqX699jNCKvZ+
Rpb0PT7D9k08YqtZUWTb10H9nXaNcVg6IOkJpQS2iu+RLQw2pyjEHlmtBkBAJeHlwiLWCR4FuNOb
3XYTwR5JGgqhqeCu9pgTEQiplPtyfh94yWaxIlCU0cYRHTasYpxVKAkn7cr/Hj3FHz9m4eMPgk3q
W/pEpPye7bTXMkXze7WYXQxM3wq3eeojD+jDJ/SXVODndKD6NunOuPh4Yi+ptPGgUfd8JOx9zdEk
spYHAosAMGza/NhIPZYLFyplRVpnkSxdndrr86xXg4oO0VvzG/x+LcsH+yVX/NBUV1CCFo7qJ2gn
Y5AJrosDkEaTqElaSUxKbLvBpoS6Y2PgtV6774khbb96qjZHsz5beoAnUGpvhLE2eqNtah/O4jfC
sm1Oxwv1p3jjfZx71FCEJ3nllIcYdzcwdRZPQ9+wBSG5zz2GS7TdlX5FnOG0V0dAjyjzQUpt1rk4
6XypIN/9fWs0Zr8CWUzXgqesHrqLB074DBJy4V2O++NuBpe5QKsgRu7pMmM+Axg5OhSvb9sa9qvz
GVXC0y9hKujhS6rfNkE5nzhSoPAYuzydUlC31DiXD4g2XwKrUF2JJroZBmnUZIhg5KeyQQQIih5C
jz6Fy4I47LmL4TeEdtjHHhs8KTs4g0vC2FLqQLiYcF0Do1WTxKIVHqceil42ppffQQxKnU0JkMtB
84DgMj8ZAqyQtTTklJeOfB3XtVKAt/kEWdPkAt+BT7R3xFq8ZwIFoY4KKcbsm2U0LBhS9rKysUVx
VVKc2q9GEmwyr9a+88F6098NrmqdI2YiqRUR0Q0UHOln/zOO/bzTIodQCzy5cE/9crTfVi60fN1u
/vBBVpdCtSLCtjAYgYcHzy+U7U2d18pjzpbhOZLKx/4is0rT7qc/vravgI5UsNckF77ASt4fGcVZ
4/nPLCxm9+kld7TrlDw2mMgrPhvmsWaVHRg3BLIhl9XNxXfbfxp+N0nLd4m4MWurG2cQ5UMnCHKx
cL9yIKetY12TyMNbtFOXWUY5MfQZ652D27nqU1KC4Ia/nNR7QNZdYK7pRWWriBmKwx3PGj8f6T6q
zdEkzeYZ/lmk/Nd4rj57QyIqgRIjydx+C8VjyWubiZFFORkLpWoE6tGrxxY1X0m7zZclWUWA9M7G
sFFIwELY1nAyanD5NxQjvxjnCeZYVSDrbykVo4UTeHkdz9HkAVUW0gm/b1tkueIP+RkqrEoaRdw8
Vzkeck6xYVqvEEg5a13TneQjJO+4vtsrJ5cGG7NA7siSiG7y3xxcCJ3Xn2xU0iGhMOQXeETfHSEd
KAd7iPEyPy5lIAX62gQyLC4WvwT0+dm6dEFoixxFVA9NzLy6sHXBXiqMwxgX/ZVQ8540sr+nTmqE
AgkwlmIbUf/N9nayDpmHBdDCnDdUZgMNddNSnD7AuNgBJtBcpRdI7cZC0o838nBmvhuzPF4+3Qn+
4thn9mALQZ67pU8uwiFNmGNxwIm8pHc//0w59vrb+5fPwsyTYPkIO/9Z8rHRzbhpq7oITBKc4AzZ
gFWlLWmUYlnnisOto4Uiw5ILMAT3p0dupz8xpm4JFKXpm8scasZtbRLaT8D1V9izcwkE08P24jfn
FQg/ndyWDullDkAaGIyWsBvM8+29a5meDm3yLpCpxfnzloInnFhUeyyb72lt4qvA8e4b0qborQTd
VtlnoyS52IvfgN1dPzq24Bs6O488ZSPQBPzImtboLfIMz4FaNmyHxS4rzWjJ0uAilr4GsoFmLQcY
RkoRx9AR14U7qU77j2MVna44EjCZ8Rdw93E5EmOPy5YLxHsWO9ElnF9pQqL9WS3frY5GgDbRCUV8
PJFcazVVOYXuaQTBWrJ9JvVeli5lKPG1S47fSLGHsPfKPowu183Nsln/EQ2J3rvYN63+dZtcwIFA
sO9dTdfH0njvkinEQ+IJUXVWPXY+lmWYTk3o7pzJTMEytjpls/34oGeuv9dQOpfGGSIrgPvgGr4C
x9QmTpe0IBiYWm6Z439E8jKOD0fhg4/Zpt+71QGUvqAEC7p6hX9KRDMEb6mX35jR6jmVsY7efEac
KzuNF17Yxx6LS7mNRJwZDpkYilqCecDZZW1QQoaMeGX/T04Fqb0r81EIy3UHqNrUJ1gLAd9N4ole
Q6ALzA7xO5kqZW/ysLZhGnQMxvLic4wOsXqv79XovGy0N0DyZtDx4YBlDlV70qPlujJ83R4+PBC5
cZcdxEmZg8c8BhUDmAzv9vHkGY7xD5Mjji2mgW3jn4boR3giakEY2nt905xVJW701ath3JPlvDEP
mTwFJLafy92ooMtGHdW0JEUDYy9iSDQE8v1RyW8K/OITGwdipGefBEv3d4yIOONTBehtQAojnuGD
z5uAeI9rR4lfLKNQ1V4NGtfk91D/Xm/ynCe1mA9N0YMjDNTJALl3f9KtH2S4p18bm/Jd3PsoI9LI
4lO1mUR7KOa3y6L0pH72lopesZg/b9LAdt157cvhyFjMGW1vzdjeQZhpuIFQ70MC/nSllTzG2/9g
Fcvq5Yq6ON+QU9/vr5vNRcQRqjCbXC7i4Cl64LcZ1CkDG0kGiGWCioT0if92Sqxp0RCYFMrFeth0
AhjPZAApu939ASCjN3ULRr2kUty/wLzGox9lac3xXHkqYuQwGICfIuoBkGwEJI3xWK2g8dqJEE/X
OACuc/enlMi8pi7fI9dngP7GBcXghAmpIjwc3C66T08JdkdCSkum1233Z4oyUIPLOFzc31+1Jwgf
Gm1jPoPvME2EcBGFn8InPc95k4RdUbVONRndS88yv/+v3tA4PPq/X4LprUCbQLQqBsaGJGPyskez
nS/NP8u/F+FUW0/3ytYCwIg1cfhoB+vZh4pAivmLYjtOqQsZlH5+VPaDD2G7qtxf0VD1lneVfoTO
br2rL+eGGRXghP7oFk6a4Xpe9wLNkubyZNsKo+H0jLle9Z6NUE4kJKeQHl/pW4SArNP1t128mhLJ
egL05niKekvvmz3Y9qrEnsCcq3rXo06IAtDDvwSaWqrUDmlQlrN+tj1MApOSy+4lE/IpKqnn0uG5
ixYMgZwFNdTw8BD5qPHOW8+kU/6bZHs77pR99VzPZjT3Ncv2BKVbgPczwcSiWdJh7p/CloMfrdqg
p8dj4WvibJbXJzpTCvyotc9OkdrtJmlsHgfD9iBlr7VOEdgy2PkiGrTcNMVJBnIcvB4qQulHPYkQ
fV6cDWc6L59AWj3XkTr2Rdymr0gd7qeXfwUrdmQY6uhQjoyt8taQaHG5gazr2Vx/qnJpCnDVOvDt
sjcKppY8wlIylrv/HostHS3MU1Csdbl3bJZYWyrKW13aP1SOjSKsUcLYTGnWKvUF3k8ZkTvQQ/QE
b2tns9Wgjjc3QKrcwXuLGkTY+7lLj/zGD/Ku/jgEcmIjj0FJexOa0BIe2SVRUkwEgMMXHyZswXDH
34PA4Mpi9CDbNJlNXwxspsNchG89Qi5LiHdBqBXLAFsmTTDIZyIaSI6ezrwScYWxbAcYyPU6Juz1
80uW0vVDyeEimXW9k23XF1e+X1++RcXgpyOTXJ93kglZho5mA3RwciaAQzZFMddFRZD5Lf9r9yLP
ZI5MULA929GN0UITqmJdt3D+kP0f86Ol1d0MOfHQ8XmoTVUvhfiQAZsGfE0hyF+eQ9IVSDJ03O/J
CAA6ZfmCqshYQ3HNnmTu5Fx85J4eAFyDbDeX00DIier+lkfFhGjf5bSumRhQ+iAfQs9Y7BjlI6pW
4TWViZk/quZvjsOLANasw6BfKgOsg9yUeXH+iWnpSaZXcw/T3uU147ybZdWoHLSTGvPetOSQkUS8
+b6AFMosdAcboESUxwnGLMxJNsg/hrW79+ypWZrVEMIufgM0d262Nb/tO8VmBFD4597BpMdcOdgI
kOE4yhcVdZBR62oWiRGxHeLEnwyT5c3lv6LbaRCmpsWK/Yb3mO0Rx2VlFCDcbV/x2EWhfwJm63sr
OWe57a/RKv58a7x+yJ4MODmilAJYO4N2HQ+eli9Kx5i9ig2epny53jJC3gduaPj6oYcA2cjYXWzc
lmCECDgsivBpzDs4B2KlFys7JnI0sIeBDdSLdj0dELgQ1xwyzAe+bkXxFaJFWjPie+UpXPhI6e1V
b/iWxTV7+3ZkhNJxe8/mAuIWc3XvGFet56tPz1WjC5YNPhgNlAHD1ICfp4YliTAZMmHNNepe8Vrv
AbnZmGnO3WuexuEKvQYYEksHs6EI133MlbthiYx3pxEEicsFPr8DS/+qN51fjAE71rcje6ccn4/K
kXBnp6NcD4z554L6DvAt39VP5pbOIKeXSA7IMCEZEto2zGdBOXHOH3i08NkEAEprDVHdX60kVtyx
m9lHepmAGTjHuOtXw0oPXpP/powP/BQ699QYU+nL8bYxqgAveKDbhG7/ACOfv6PYUqjB2gOMdWvV
gp9PNYioHLqNGo5yvddlY0La7qbuBSsr/W1jF0T1mTKi8gI7oo/uyfs94W0qgjjEm9ndxMe8ct1Y
JSkXxw/AUVgV0RLN4ipPQ7+0Jr7Pb/FylolQh1Zw/DROnUnmQ8WKdNUYNlY1WyIG/d/FPGR7XO2g
8UKodFhxs+ZPXk/rAkPTzYYOLL3fKvG7/0b2CiUQOLxKoP0AmBQupdt5tuGvHwGUrBJlzeGAFu3v
SPKU5L/pvz4FbaBJQHgXFbToTORxRrRMW7jMo5xB+Vs4RvIz291XL7PnfgXPrOGK95Hxa7wOsFfe
jCoWHWl5rzMA3Tp48cL9Qx8OdYN/7cTysBw4o6FmZ8ZLioMU3ZoSHjeurnuPncI/1jA6wfQl0Qpg
W1GBH1qdPgL5UNsMGAlA63/5oJpyNTBnGcGhf3cgSsQqdQbXD7HVN4be07c9FR+Nes58e6W2getJ
BPJndtssz1l3Tb/u74GZccRUGorlaMg/HjwAfZgCD9t7okXxU1dJ9IDhL2d7Ij0xJp2nAWJpsi5E
kR/611UW0pLFBC24hlVTlvf5VFQesva70nj04f+qboVs5DaMdhW1NGuMwLZqSxsDkrsFnhZbZJ/N
Nr4jNZcpAX+MtmV82ZtHaol2Mi51+VtysRGDhbIFK/ZQuUMqVX/jDDqW0mdW5qvnh+j9Uvengdhj
NBktmizujFuulXRKXXNLlwzgo/8vLLCQJwyLCQM/zwl1pgd/SVaJ95zbPAYJEmAm7rcnGLmaLKR5
ZmecxQcv8gfPdfnQArV1PtdyFzV60G7lw5MdGJHnR8tyw2PeKcxEoDSSBWYlbB2EnyYbjh3kbd+l
sUeAjdqHsztmCYbf2QHx7WR1A+LimfEIJI5I16bv93HzClJ6fevpYEvktOLkPv2OPVAeq/iN4fzg
JQORmkqJ29sDBLHywDYez6RQxgL31PLi7nI+Ux0WyCtDiH8brqFAsuAuG155avijXiv3Hq+nB0wo
6T5/Ur5qXBXbjEQedMVKISTEXGRO9XXMm+exgJJdpjWlZXzr3iy1OcMYxGnmTrWvp/lxtbqacG2H
+w7iD7aLp/2jwi15matiftUc60fz8JkR7p2zpNy/oifjwDG2FMZdhAsJzD8DvPPOCRWndYBWby1+
Klpm7V96TaT9iNUSd2C764ZWZKRtOEKwwnqMgoJVd5FO91k25anFrKf/sot0iRWy0je1VVQnUzas
f0VOLDmVMNyuicaVosB3gCwDuJufv3/BpYmLysV7/IL8HcVH0R+Hbl5Rt4THz8KJW4/Qd3zWy/Ni
z25UjQrpyzZTGnhfCpi0kFcrH9we62UVy9VULx760bTTSHVe8AQa5CwWn/mKd9b9s7TnZwF9gQCi
sfg6eG0oXm1BMxioexALzZq3wMwtExLVe3giGt5VRdFqJv8S/JqsY2/yuW9LaUIQe4F8iLKwjlvj
piQLKEuBHy217dBQuCpdIEGBHPXaIgd/cAoniLXJnkgKMPTwsVynk6fKQijAqKGeZWayui2tEZda
0tb2v9pQJZ3BBaNVSkVb07LsKBvClFqQ0pALRsSByVBxe7IdmmB9dcNRw0glnbcgDE6TQz9gdlRR
M6JuLcFdgIUhf6eMid6CbGm/kDkx4wO7g+Y9aNBtYm24Rw6Se450wI0Ck5L8FBJhtm5kEGevxinI
h7K2YGfSn8GmLixz6nfSK+q+sFWNo07fKTy74+bpSfSKCnBTmRVc1Mh5ON0StoqjwSt2zlFooWQK
rI61auxvNVlJHu72xWZvY8rdpuP1+cVw9ok2LOSPNj1Ceyaz6yLohTuyshHP/Q+ztxrjZOwBK5M1
8Vn5+Utm5Uj5T+2Z2+VKrk7uZE9le+/+iRd7qp4ttwTeKpXzwPh6gvMaqQiGIox8zMAcUZYUvR/C
bBsNDXu6VYZIH3fnnlbbXREGZXG2j4ZUfx/0dnEVdB1jvW14ch3OOIYpoguCHAlwTVdOY8IzB74J
/RNKqStqo8hFzL91heQSo3LUvm5777AUcgMS7rV5mjVAdMIZ8JaC59Lm2uU8UykrbWRnV4UsO7RY
A8a6S730G3KVzxEthS0BYTGSi3eCnDlvP9dKUbCSvbLDkd5wK7fJxh6LPPT/lUz43G2pZfnZhXai
r/kSG/aEb/I1K3FSY12uTEISmCI643yJP7sfmZIEhaJd58UZDm8bDKb7yfvv+hKMzt9iqo4fCgwr
eJfHges7v1lTbyg1EncGK4SDZXDCjoyDwYJTJRGQOp/Adbjssks/I86BwmXvbdOLCwYZyTNvVtHK
cZ+XCKfLzKIuXeFU8bRIPV7JF/KdqKvQTKtOV3J8e+xm5XQpRlfR4DGlS3x/M9nvfKwM8b8qFVEP
fq7NaS5dIjvY9FFejesuA815aYMwZX6Q0ylwqFsOfvcVA1v5zYUZYFWNg5tQiN+aQ3tolsRF6JPN
DRMeTjkb2MOxgY/LDZkW35OU9BHoUo9TItPOYppBHxTtkcycMpA9PoYliN1H/oeqVHEsuU4pxuDj
JIxHiNF4d6jNLaZf3Itb0rB63flDWMb2x8TAw7nRy6YuDZqAY+mnlliIPoQPNwZDJLXFqt+4Z9ko
Ig1dDnuv8yd1gCab3S/lgAZg4N0YCCx7mtmN1iS+lOyVUr2mUMUMkI1jRM7daZ+GJNYpSVmt5s/z
B1hoP31tcgBTDrKX1oA1TcpPTS8uR55ikG0E5k90oPO9zsgHEwnWyv+3QE4ebpPesq8RX5QkegLC
13v6fuPXyL8EotTQDsKwMD00sqaVqTDEEoRO1MobxWTElMbzSTFfBfzZR+LozC061fE24TipPhFv
Actc0HRtyCqZ1irond3nPYKZK8BI4c3zkba5FJDC075wvgzjaz9kip6W/SBvMGIMuXYOv7R4XhPj
hgf13gDRdg6DVmxIBvgtpTCMyGHRhWu9PDp2o224j8GfaSHY66xhP5OVqbJJ151YdhbNTPzJSpcz
661AnNyLx9tx15zRXqQQxHamnghy+7hCD+v415o11xcKfY/uJGI1Oq+GhQ56Oxn7PjWkGwSrqTSJ
7UUXY0NCW4h2XYidhMBROizjF+FE7gwN8AHGp+GTLBRy+F2nznXEVPDN+9fA0kLKbjPoTYikjopZ
OtUD7iFGZ2nQDOK0BE/OSQX4uFDeePH/VPxvXzIJhLNOO8UFGwo21rGSyIwRaOte/oiZQmk7h/CI
DdJmMCE644DGpwLFrh3OPgfqi8ttswygDUKqowlI3Dt85XMZdvlMFGqUffnd9nBd0wDfOdNWkqJp
e4y4pjPtbG6Yk9knlnrlDZKNXIZR7oEf9Unns+eddplFtR+sYB7lRbOIoWhwhYxDbk5TcisJwTiV
BKYTCb/Gi0axeGDyF/73xooZ3gDFQVvLgyC+nM7LGOeNStpkG+o05dV/ZCpAezChLd5DmooAvznx
CgkWtfBHq3Y1Ze+2coyk28mOYrZqsEBVzOciz82z/4KzJvK1J5FX6+J/JqpNyLaqSpgDyVWmNGFA
haCYOHXb4tjLXHJLWNRGL2WXZ2eTsPlhw8ahAAFRP8rN6kcoB/ka+uEudfr7pVXFTePAhkNsPZxU
1fVjrnHbOpJ9TvjJPSpG90usU+GalF4bwcehFyPt1+oj+ElIR36yHDy+B8GxupbwY/7RLGzIuk4X
m3yccKV3Thf493GzCntZx67ziraYTl0/oVainPU2Ne+vSaqzm9k04X7zLAqagNwu7iXcZgfMUuXK
jDUMfA9E8LO8hDyJR+Zv84+EF93OLMaZzCUExDmXWE+Ib/V4JB8qfBo7B6Nzbwscaoe6w0XUkpzq
wSvI+IqCz0nJtSA70AD/UpJo30xDHC/bQipa7rxxr/OCQiJ36RzG+WX7srPBMg6wRO8ugLHzbTa3
nN2x57QD0KePBLDBd7rWgAVjEqu+dII4LWXhDPYhZu7bPQxQKvw/7NpjATAfs9PxYj1ZvfSDUB0u
ZVkjOnpc42crJWfQXA5Y3WwlALrSIuV73Pby0hdc+sgBGH8g47fOzY4ZcO9yZjwa9iWqER/YasRl
xZrxAEKNX+kBhZ1CIiiFT4766QjaoAvAB9CsqxeIsuvsw55DNJT0eyMP3NFMh5B8ipWhigwmr3dh
fEUqvJUvnV6EwgfUf0hFKkm5p3dfbDzv9V+leBhMmj0CllC742/i+kQGL/XiRa2sCuv8/DvZBahF
7AMlmNC2pCKY6NYLwLja3pCfVUFClUA+DKpdxkExug7cB9U/XEGAgenbR33uWQ3fnDqoXNEI0qRX
kNVtpG9sOVf3NgZRhIZRY+5QDs53YEotIhr9jZipG5S/SitpjuebL9nu/j1sUNH+pzkRyZgw9gHu
UqgdcLFHQcNzc65luG62wWYG22QhjSLyAz7dFYu0l6FHCskNBh4EG69Kj9eTtCaOfrW1n/Kstihi
1Hz95yEjmA3s8tYBub9o+whwG/uhVC7drIyhfoioSlYqSojcz31INHudq7yfG+rOPsRalD3eCHAI
LxqPFn864qbSXB8JqRihNbaVXLoBUOqcjtxc3EhA1zZI6VnkGStQEDDLAmTnUtNplm/y4FquDN48
9HClN8fEt3uHhmsEok8yqVjJFQKHqVSAXglnL0anU0iNAjEsSNeE4WFcQj2t7uEdMnxINrLZI3Vd
SeMe+wD9on4/jF3/XDXxx3y3xV51kWzq6wSHrD0VbDwqeSghrM+N9r7iMIRSLe4T8EShztm7dPBh
Jpfna6qYeV+zN7JYFZKZhdFF4KTZfzW5i3RuIJuMP2JyfSZq/BiEzgiRGTcJKnujpSe8watDrAdc
bR3FkmCoypzGrVJhZeWAE37OBYxFX9E++hm5kGgA69aD+HWMBANyk7tQM/dB6Q7oReHAUHDZNfuw
ZAlfk2eiV7N7XtIppOZHfKUFaaaYLNtgE4F76tTjHKeyEwDcS5ZUfROLvfATCgqUfiCYMwJYpK+P
b2L+63DY33wb0t3xjt2VGg7+moY593j9CNn6hRNcS/Vfeb2E5xGt5Kk1pBvh/kUoYg7UqUi92efz
BBFk+zfXhNuMXzjBtqltymiSeTzzpAFN7dtsvuVL4s4x+reNBkxlYd5/wtAah6q0Y2tihUnXmL/P
YK40hEM2N66nufOQ/RRVnR0U3dnrRl9wMzoa2ZyQyAgSgyIZmTcnH+CV0uOTb6KiZxqw3oCtiv2Z
rBU6AnF5h1uX8kEPOOnYviNJvzegj37zvZSX8KbHocGcFriwMAMbYBDVygs2YpjEshMAnbNRt+Su
v/MpNdie9rJnoob59NKQ34MzL2wTUM2X8f1TTv1mNFGHs9Z0Q3dxUR8V0a+H9lDSWdxs9ene0XI9
Dp/EeMCui+n+n6lYTjlLDEf84jOvnW3Yr1d6E7lOdSH6PA5dtfQg+OdjebM1qcSRsOcxRN21EPG1
yaHuW2k3mSyURLtXpHz1uXd5idkMYhffEPq2VBR1xTE4uHm7gPwXodSbWNjRjczpNucG1UCvz2JU
gbzEe20eCE38fW9xdDxNE0YA0N9/8Zw9lBBqeVx3I9kcCVuV0n627P4n7VWwLaLMmLvu3YBdS3LT
tK67Pi9fN1rcX1nftXx9rdOcykUQjyKgQLFcddIoQO1AuXQ2qkGHDaHct+LxuzKmfYl15gHSnxrQ
Q3uX2quA9BMv8JA/rudp92mSlXtgVyYq1Zy9XtehMJF/kID9aglaCcaEiOcgPXHZQ0iFsDEGra8m
ReADpLqh862PcP3E4Ftlxi/plFZKr1HQEiujwKdAMNNSw16zYkFZ1gdpY8/qNatCvMD6/YxnB0GS
ZAbOaxVrZcAaaOwDXaATq8Uq1lkZCkVPqcEiJqzuxbKxc9G7OqNz7fF+0iHrc62NpxEfadOTSUUl
z1HQ7wkad7bblzRX55/KmGY65RwgEnEgfB2oOV5HksIbySdmQUEKksRMUA29+eRe+9lInWLBkitN
FmSZA0QiRwgnM0Y6CNoOjLxKcsp3g5uMfyvYtuLJ09SMlggHD1WAFnBn+LeoINRd/vTezcpoKrDN
X1Bx4ArzGTVZ/8y/+P1KwyoxUsDcbBeDmczvIlCODKebwhZS2FuPxuu0h4aTDH4hyap+k2xd0qng
B/xvb3iyUO0A9O85OCLrm49AlDnbg75rvv4CSdPLCnMv1lOW1d0JX+rW2FymF96MbPFKxoQ/V5lZ
cuCJ2EfxWMS+I4jlwch1EdKxiwcdsZQnIqOLREhZxAFP3TiVCf6nRbaLkNphcZ6vl7SvMsVf4zqh
Ie71d9ij6lgOoULK1o/kgyLxN9P3AWIdVXoY4aPCz8LWF3lXjdDn4vsOmygpq9OK/VqnuzD6isQj
jEfnosgJK72MZVVvzdVd8P6J9LHioWFzuaLzpF94bmCq0BbFAQxBc4y1Gnnh7S0Rs+I/uCnpoXsA
KHJK0NfPGJajMTPODi/xI4NduotFtakkWoDnFglDycVLpQvgFNc/dj/QCDVKGNBTfDSlY2JLp9uq
G871V68xhRqiuBSAYIBCa+FV1+qFvqgzPK+VvLVtqA9+fV17FFbtGbHIeDHzAUXk4jVmp0rmj9ez
2kDmLjt+PlubRHqesSXFitXl/tQ9QNzmGrMh+TJZ6WY4p6I8X+tdhNlcQCGecowIdaZoh3t9Dkws
7GgffJNMuXKqOu/JnN0275sMaf717O+dqxDUsMIJthu/9rmCaBXAqazdRiJy5Reh55/Tx4kbgzmT
r2u/gAip8XHLbeXs+dOcChYp3kA6GRv3Na2GMzYZHAZd0FOScDMJJ+g7PzuRcq/F07F+XcNEZ5vp
LWroqxrtypJbD39gDfoOyTSVy2sd471HcdfQp6f2LpqKh6xKzjqJvtgvxw1XQT3RMWZekBH4F9Zj
h6O3i7UD8xi+37iK5sX4mxf8coNmAqMDnImA10VNVJgJjIr1QUyi2GQqLbexljGasiEWwJk7RTlw
B3SDXCxStdgDaUH8p7wsqJ3ZEdRSUttRQ4YRxb4oc0Q6WR45qRURpYMfGwSY0CHuDQdLMn7V06H2
dNoib648Vsm+4oK+QjZKTN5jGtUotCgTj46y0BXzD88coPEFySNaawYeeem7BxLLqB+UfVXWAme6
WPP2F84MjNvK/QjLBdnTEKnbUPBfGfuPFmwlRUZB/lR36nwwZV12D95YKyS/FKwotpj8M720cDUY
MC5HIG+wvf/fN3N4a9ec88NwAfJGAOYP0viIxX8eeIXC7hq38sxWtRQr2EqRUw9ogBAXcN+tA/xx
gcOUd0+HIfqXEdZeFb1yhEQqUuUtOxyRAjmpL/br5OXeraDA4011a32FlBcgLoDqC+fx5e9E9dj6
6+X+vROLI9ajNpmv01E6Pt4HTnfKBqQn7t+3TdLsyppv7Pt/nh72tFu4pzlKAwbPqkRgvEK9oAh+
y6iexCJIlrYrPb1y3zLvA7YJ9zNUloZex4Sn3qf4xk+PSmXSyWxHMMHB/8OQkSbP+hCv/Gm46PDt
I5z7JKFGrEotD+6/4mnkBhsPtl4R1iRaF9vkhheMbCxAeiDwPPbZQnpuoDJoRScMCqYvHM1wQ7WJ
+7cd8C0E6dL2KYxwM2Z3G52muVOjHFfmmdlW6jYD6rZYLBn5YRA8sCjMgxsMR6C5Hj0t4DPkXrY3
Pg3e5/E3yquJlAMh7Pl3gTvkxK097yTc6Z5O4+LBTKxKOYaEBScZmB97h1p94fZckjvTSHbWOfgR
vfh+3m+7q79BHi5RzVfo2mEjUoUwxboMQSnhGhn0AgwwYHd/3C5s9oeJqQkYGMpPtlgAruPJKUD8
qUQk6iVOCxewPHvGi4PFnipIWX8W3iu9Wef/cdgHqjZjhgPUHjm8b1xqTSehe0v+dV9wGuZVDRkP
it8p2xXxGFpfFLap6VADZ9qrcGO8Q8+X72vAgq2M3LcHqEnPi2N7H1O1na4Ueri3pPzVCl2+1IY6
r1FBZhENjjrGvySdXqNMAszPDpGD6dry8CJM9bHavwFOyqBtIbiN6F3EZFOUV9b6GNjuYvu5qYUl
NNoU6IGs84blq7tM7+Pq+Wik/8ODdVDlXuxxsLxOtitwThrA9ruAvuhCY7uZquO93IHivSPPvkRC
Wry60vut3qSQDipK5vmph7nJdpkTe707AqnFeXNRuighd8BUif3B2whLTBwSVWZvK1MzMqhta38E
ZiPbHEdgjB1jBOf6bd9C4pFdmWjjnZXQni3NX8L4l50tWwS2wLT7AmDauO5sCsG87Tig19Tg9F97
27BUU5cz6ZeCTDRhIPiKPDg9kBtW41b9Q7eVYLeFizxsZZnmgxsE9AT/0LVXDt+XZJUXUP0D2RAg
gmC85j9GA6lsBmbh3i6wLdkhuosicTJKhn2PP3lGi9qYkX8diErMAoYoy0UKKX4Meb2hwuwJTfSr
oieHB9aUZcWcDJl63+OSkvoKKO9tfH1FV7HVX23BdKk71KnQg1BJHZ5EPIXYUUCphzpUlnUrsuzd
FuFi+H26Bato9fR/N/iXplLC8D3toYjQombJlnoirRdtGkDvwn0ITTqpCLmtUqhfYpeW9+9BmLzj
TBSrEN4fGKzbpZoWzVa9Lng7Y3NFtY4HxEBV3MEIlMjpe35QiRh0WwaGH7yxl4xOtSUBt5APrJyO
UF7KuKl1csdz0Gu32qAyVT+BH6pNd3onLlYGwjOQe97w3cNavkJhLGQrvl0j402nUGFA9f15pvXQ
mayo2wg9ofjGKWp+bK+eq9QtNhdNCc1hW63uS1v4kagWtpHyxMj60MQo4IHDHGrHYQFg/hQAsjew
90OV4pTOiZHwnhNKnwRdQw2yiQInc222/9X2sys2cE0aA8YPy4TAS3JjzUbQjasHy10fMgbUVAhd
LnEZQczvF453BjZw+uLoJ6ZetT8HZiG5M41l2gzl8H6WXv4grXCUmcYuUUz4kraRZeDo2z7tKmbp
JvzzJKbji1ZN2gp/9gSLiU/SGBMoFd2UrzoGn2aH5GToA7khTtmz1oc/GkqIYawRw9k/GIOCnO2+
gvC/J7Svash3nl2p7a7naCkiXNzqTjHf1+5M0FAz41py6zIOxQgVCac/nrwedTz9f99R+NnlS0yF
tUM1wC2HVF1iESYBHzh5ACh+OTJB9S4IwZ+ny68eDHddlmWcTSsyXcpJn8ArfhpBUV5qmPkVRevB
ry23qFs9+8YH5gbdg0wvgclJbKi5LiaSHn5gsDv3Zu2auSN8CRgk8YMy3hN9XydsYlWIzE9nfE2X
AR0JYgnSW9RXAr+bzF1rluFLAx3ayWVbcjVqyKpMB9C9NAhIYK4o4JcK7IrBnDDZDDy7yedjkdIf
Q1FJO+CuWmaIh27cASL4dMsDVI/iPkvWa/VBtFPHYqFqPf7VWZ5bKGe8BH7tjWQQw12L7qwaimJV
GYviHGw7h7yXbiqnw2Muyr8gs6F2C1UxFUmNuzns8jrP80DMI0Nc7yOuA/TMKH0YclK44NYT2Uu/
UWHTFXQq7OKEmTEPOiW7r/T8NTasLYp61y51FI+ZUOA/kanxVjWHmaXlB1TpexqZRNOWGacMGvfE
JVSC6z5NMRPu4wTOaz1QvAIkdVVo+qn7KQgRxdgE1v4GeWmsdgaW+qH1F+1JZ+gulj73aMwq12Y1
uOGQGAAyl2YRPE0E0XpA+HfWRGL+D94W0DUBbiFW4G+IdcXh1glp68pVAryVW98TikoCegcxIlUw
qrxLCDVqSg6H7yIvyLptgfIHNIrpClDEpUd+bfFByihySUt/2KOlYx5lIcvYfzSHEUX6WzPbt/Or
rVnSMjFKzznFl2uPU4nrEfcnmsxKpx0+ouDSnqnzHbJDJ5+zNBBJVKMYg9Vn9z1BrSVqVuRbnlPj
1O7t9MMb/MqqzgNk3eoPJ1tIiWrwGZdADyERTl4EiE3QIpRmvh9vz0ckhrMcrA0K8fg5nIQl9/4F
PyNYkq611QpQX8Ffh+7Eepgzh6auRrGtItfo4fjqTjKcpd1MbZb3Vka9olZTTN89QdQaButWfFO6
d1DOrtitd19bBOuAkQAbg/QsnkWGiuiGKSNygpuhQ9TfqBs+W71gY4LmUvtB+l3IHIAN4EktQk1H
FJa+547e06Khtqy3czZwuWP+IPNP7xDTIHBNb2ReXbs90QUZ/eXkDcnCQyH2CCh4E46KLx9rqsXb
r0+mLxzEm8oJUWIMB2ceTvkPqLFNKTS9RBUtrtTi3B8Wj4sAGsSjBwFFZhDZmnoQ+Z9yHpNqe3/6
uBEcxiy5UhQeOE1TjQfPCuDjDY2B64dEA6ixE+L+OJgTdoXgVAQfKap2e0aQk9frKepmKMsKSF56
FRaonimN1SYX+BSYPMf182d/SYbF6nUhICBgc1JuM7EXpdGeYrKQmb4kLaW/ekPDOoDtkz/rKZEq
zkwoCewT1X9W29Blj9Wm0bZlakC0J74UBPCdt1/nEOVn1NQmc+UKBVe8cPBoJm97U28Hba51CKOF
7rqB23qZ+nxbav5f5cc0+3ZhzcK2YoN6FgFzaD/jHFKCB1Kri+B9VPSQo9L+aw2tLHH3K2U8+S/k
KQRP5AN7ICG+afMXX0Vix1sZFQ89sZXjvjBT3nhM4oEAHUwqGIk+4MhbucOZd1ck5Hc945+c9+QX
nOCOupLcD7/NNedU1gPjHkbRc3V/x8o+7AdVZQGNn4v710/mFp0Flo+KjqS1L++sxIt8v/ntOYko
QywHkM/j79X1feo1rPR19rDHh6rdqgEsXqpSXTn3H3WRynC2p9WcJL5vhZq3ksNuqoU5ZS6gQSQ6
zzeQuEAW1h0skszBpKmDrb6i4g/y6OSV50bfcHVY0SW+Sr5erkz19Gr0cZwe1q+njbZCdfJct4IP
+CN7zfEaC0EETLuPxxATiJnK5O21Nx+2k0OMpXtx+jNWFEBj3HQicD0fd3D5MQNRPhYjfKpsO29j
DMIZjQ5Bz9+ydBOg5a2q2TL072pWcBUMbsHn59hgbdZizRzbqR2qT8dOHs90z3O3pJcJ/4coojZ9
0aZ4l8C5qz4dRvc/CQAPfIPZkxiOdQVBcpvn7/Hi8ol/9MXqPoRE5z9Xw+TzuNNpe/d6FmnFgFr2
6HUlVhL2aei7P8ZC/zOEchjJYW9lxjfhQpTqpjPoloMBY2l96jeS5GiB0PkTIuaA3dc2T86LX516
F96cmBXO4XJ62Sz4XwM8NGLwi3E/najnzRtG0VjGPIMZx0p6S9AuKN4cKRwDVWI8PcpXmJJRS23/
dfDqR8Cms3xtwfCN5MVIPHN2ULAWtJSI+gHvkfWhqllPlvPs20FkgGSs97HIl/vR0/nhYpf4dz4w
yhErWW557DFrOK3rYoROAz+jafSTCBk8l1Q/aV0Sv2IH9JdA+0Do1Z9tsgzQn4Jv15IZp/PebSbk
YV4SOcrURedPp4lT+DM22ibmClsfcN6rMGIlaXzHe1rE7O/QJf1bqE9exgedwjeLpGrHAYSwvYI8
fVGpmArzPGa8fXk+xspoPo2/LUYouO9RAXC5pDCGvNmx064JRQElx2NVPwi7yMhoruUeqQOk5mma
pgcPf8uM1F8Qv6inf2586SlfhxgoXlPEKL4dl64jKxvO12OndpOZDA8suKOSr83xhahXWqdjMAXm
85i+h98tTp/qxqHBf5jQUJLD3JQO9Nqri83QljoNAIT4hGOfnsnTPGPygxZMC3Q4PDDA0EIYNvHW
hcEMPHZ2qLeHeTerOyRTRc7KiuwV1azrl14KBxcs5PZPDLtYIb8UmLRpCugIrN18PwkC5dmYCAPE
xHxBgzskMY0HQbVz3++5HsclAt+9qI7JfkBlfL4Dazb0alL1iV/zOQ0jLkRbRpqdnf8cLUJYKxVI
jZM0N4/iVmkffQFUrUMTPHeiWV6/tZxiyKXwLKOsGDa7D3FZ5m3hzf0TKN+HNT+kXXQkP6z4bcD4
fk3fgnpCgRFudwPQX+uCPH28ALFwuoTojdrnFuPqhKMgXM9hT2KIcSO9Kjm6gG4qtwUZ7drDXUoT
9sE1j+v8efBLdH991EFn7pM4yLWpr3j8DX0CbKKzGD7OmSAc64iJT0FeegtGCd1l2bJ80eX2hMBf
XbWxNg1ARIdcDr9zqwVKElqJdrvyPcqT1k0e0mT9vXSSVSn5dk5PO2f8g0n/j2+8HATHlVCEgNyg
BitODD0DwiInmg2PNoa6CRA0svywFQVWBBwYWIwy69VSC8t9EuR6TuXxZkb0gfdeCGB/Zr7aVTtk
Zil45c2LeE7TgBLsedwQK6aYqL/GSCr2+99XK8jgAtlhUXSoK2EkDgjKeamE/+2kOjxczzRpxmdn
7d8YTaLwkbfA8rtwy7O3M4o2L1tI6TzgR7ONZ7j0YMJ5/EYtkJvqpGY5U5ZUsLrCJcmGJ9JSJBOy
lBzAufvX3ppLqVSKh1eKRRC7Zjw6Ar3BIclJSxY/jyz3qkOkKdzU3RolCj9lOEQ5SZyb8lOpwM50
pYgL4ebj5hEJ/wNO8v0GLUmmNc8PBaeDmxVMjCzh7CiHo5xX61WzGtTBhiCnU/k6Yo9rlnaECljT
a/SKhpum0T4Sly3nGoFxndBaC1STbTVLLlMuqK+dJtYWddtkSPqKTCjLEeaVCIYq4dBnYbIPlACR
R+embbxEEnjhSJAREiI3SMohF2VZzsqD7/gKiGw7RlucbHqTdqbnihdLCkKamFNQxNREW+JaGKsv
BZz1vTePzu15eKCdkim5lBZHhr4Ou4/x+XQifTm1bMUQxsfv0V/IfBGGgJAO56ss0ISSwj0NZF/+
eUPl+GkpsnQumMkNNTcmyd1xcYCV6ysHq3cP6RqIMa32oicJ16wXm/e4nRBDW/ofoFgLltXUrzdP
9XNjLM5d6U7qENar+C3+igaxXghLjL6yZNwI0dWQFGArdABYStGzSup+DT3op6dZuHxwTlMo5z9e
+Wc+GCYLbaBFxZvBUt2PGrmPW7Zw62f8DVasIDb54a9nASvDwS8bj8CmZiU+dkGYszpurHHePpQD
ozpA/LqhMlG7Li1DRBIgWd7jug9G2lO+UkD/CzLrzs1VUy2QQHS5cFs9naqyVz26kq4HyB95dTCL
Zkq2lQJn/kyizjhB74W0lZa017uidnbit8s8oifgNs24Kb3Gzmh6XItVoJu/XmNvah0B3/1VyEFS
+jhftXVlxPX6EIeQT7zB83OPQENA5TbFUZzGn+Do2q58tS6t1gsvwHr6ZwgFvxAa0NvqEdSlQJiM
+P+Nr6G80sFnz1v3Z9L/0XtzDOmV7wAz0zx9xVgGugKMu1V6l3bhBqEPfoet0c7SJhsr7dNrwgHi
0b59XLI0zrrFyrcfOp70q7ozKVrBSdlxd2MjcuW89IV9RNGPycvq76kUBjH/Kfxst/VlgwxdqlUp
4gBEQ2fcTEdAt76+6WGrJKXRme1QXqhcnlQe+zpdJnpQJcArRaqAtqnS8lI1MFp9IKSoajMxrwLJ
8R6lXvHcJ9jlXliVzx0MfLfox79PJsPjVyRNeoDj2McUjinQy4tdzjwBh+9DpoMqDWkw31aPx8C3
Y2biNlNykdTuyJ4xiq5gMBSTAcQJoSnm5lDPDgUIXhNxPgdUjovSqRxS0+OzPm7hDNte8T8lZjI5
3/59sBmxlB0zR7X4wesc5S0oejFgIdyJgfHGcZi+2/5D9/WL/lGgmzAT8hH4uWHQRaU77fsJoCXn
3TcUKH8iSadbtS9R+Xi6rYPH08UaYQ0mJwDg+RBnYzdP8k8kwV7kH2Y/Mj653KFY+sEqn94cdChA
HKtiPH1JPwgSdYo2tAHz9DO1OikouWMRHmqgfVO15WXglK7sdwRiK94KQm3s2R+sBnxwv6my+1JE
EzTA1IoEEAy4yIo6yA5ohD887bknkRn94LkBbDXYW6WdZXkVuEbX0fYE2XTzW3H8SiLmwP1NpJp2
t7MZikDx4c3HwH5eFQs+bHtvkg6d86vOYgUPorcQdD6bsnt6CkUOyZoCg5+oZhet4qDT4PVJ4yd0
2ANeyDrsPK+JIcSb+V6dWdeTsWcMxToaQTU1N4Ody3/kftixvCNiSLN3cEKu/JFDs/N4Re9k7uM6
roynKECOxPy3LEN8rTiEQI06JIM/ohbcX+9OEDxw+VgZtAwSCtUkTVPBFNeL1ToJ1TueBZc6Lmke
9AJBndgGLzLDVQSpzeK/B862NExUYf1UXve3OHLeipxQt4HjeTyznBY9hz1w2S6LeTygDQJFS5cf
i6yTkdBVMLec7Mo7lq+MZuI9M8UccTYRq1xRLceYSfgh1tu4+vHrkf3erYmrQ51rT/ZuYwrtFYkL
N+BcXiLlkzOxf3u5D/J8RrBKFcavlJpZF4HAJexGsFSiPXrIhvVP6GuGS8RVVxTFJJGOcEoM2v45
NdDXk+WxRWsV/R0oN9TjgzjJorq7LGntGF/7+uiozbvlqa7u5UeIX0KC+RJDcgfU0t+sOLmTrFYM
b2lAd++Z2SmVKkm0jGbymTclWgE0yu6pqPqFMueuAzI54o5sWMGtWX5mmJmm29RZm/bzVFsMrwT4
IfIqbZonMdfmF+zsdCs0IYlT7kxkmRw7snD3FvWcAtY5xDwpwtQTnxwvuQyVoGRGkWIzPYpDr+HL
fGgeuY6R31dAD6EzDHmZfyxgT2yrRQPIYTyH3EGqHNGiqWeS2CiXTa+3dO/uSJyo01/VPVYJ3BSf
lcSIsIg4VvatM5O8fZ9LySFb3dHoIQvINPZSeh47xD0dOhQwBabSUv/ymbuACDPDAE873LWsE8P7
q1+b9bE2q+Pt9U327xFtartIAYCCplw1mE7kTvQVLZxzterfqm+FFF0ojG4Xg6QZEEhqHPK8nKlW
IwHMaedVL65Aw9e2zd22Whu97HVTI8IRoNkz7MDHNQ6a4x0NxiYB7TaUtiMkQfUpNL6W5N0gm+GK
b2gYerycdimGliKG6WIc74lGWsPRf0LZJUQCzXGaLgZgXjMZKVE8bH/xRG8gRYtx0mIlo6d+vw6V
H4/P5h7oZNEX3Y7fGf0Ci3nyYEu2bo/90NVlinnfoULNvno693Gfx9RBQDQx9jGKDZ85o6u2VthM
g4L4Y5rhgQ52fuWPwx8SssHQA1FUeL3EieA+MkQkrp/NppaS/PgVRXgFtV903jANlKPOtr1eY0GX
cU0ANtO6pjl8StNEKwb8rKmmueSY+kViiWFC2mi1WpYrMi+MdpzGNzj+pdz5sD0nBkLdI1kcHVj+
x+OzzwFAlGZFaxJ0UyueEWJdFKkSEIuepdoxn+9AJHaXS+mISkI7biiRBs6lZ43MCb5CXvhxDJUh
8EPEZwR4+ZZi83bEGlWdxA2m/hActClaKnXS2pljNl/uctbBSEmE5WsoNwL5VT3SnrpAfrVQSEVM
dHgzJJg+4+MQlLcOadLcey2oMx5xfhLwG/MD5RHFLTXUPY+fi+VW001pe0D/5FtUWfsptTNuaJbl
FcgacY902n/dN1CinXXgMP5vnM6aVS76P5sdKowEMDo8qyfvzyd+ynEPNtCfD3YYUm3zlNZL/6qP
JWa/R3xH84H9Yzb+984ydvxlgVoRC1iYFuKQpKfU1umfeJRhm0PrRR7CngrXfrqq2fL381ZrlE2r
CNiRqy4c2hy7PKm8Pr1QWCiyXtRlt6P/gqxhaC4qAOOt3z/H+MmbwvePM/BptIpYP2XUYsWbDrJK
8pXHgR641+QjmgPIvZdzd/PLZZkzTKM15/G/B7KIeA+AHmOY5W+w2OibpSSljEnl9kBHEil6IWt6
ZEeb1THrLhWKq6dCfmH3ptZYfRsu2wwN+neMQ1DdzGO/cJmH2TD9gQmB5r5PRgCUbBBaTPBVr5cE
P1fbIIasp5bbBKg49uuREMx7q+BHXTR0Pxxu1rVt2opzF9mpZzxlGcnwJe++TJWNq6yZXR96aSez
SMfTAZTz/dF2pK+X0rK+6PjwrWU5IKAWWmVWIUkyEdqLrEjoChYRROneGb3XiX1OVsUUVHsOe0ET
s0JP3Yy6PqPml+Gj5s3qfvtN/4Tt+h9nJbSC3S2SZsaNinMde0FdC+ns7hgq5k9bC/qCHon3+O0L
YPDJ4PS9XCu/dkt5OkFZ+FgIWrncat2mq3J7SAUXYGls9MVjGMrGaPaFeM7KpcGfXgchT+XDDJ5s
jDUV/8d/tSeSAfLXt+G06RLSYpKGEPTOyy3A5Njt58ivo8ui/0FUrj7Wh2RHl/AcZIW6dWcT4WzU
9ysUkNgCVfIgnQjoCusda4/kNWZC7OSxYAMUOMUSpjg5DVsSCr340yLvz8EkCoyXYxMlOy/FnaBY
xy7LgF+kOAAQUnLFNUOg16n5aILmVLRgBgbbZa1d+4l0AHIfeTq6FoNVZEA+U5oGnw0pzVBgAdaj
AYmGqgVw5O5YBkKeV6Mv7HulsJlwcov765TmdiFcrJqWEaXLprxpI83U3XIlmwpxejOnm+d5kNmi
IzEjEehgWCxz6MwyX97/68PhxR2WA34d1x8ACGqUy1p20FCodBSwxZSfTZyIuX+b5ioiOSJ5XNs9
Dc4NPxthaGovLK6msOPzHlQbSENPYu5L5RPRHN6bihs6lsfdplh28oFc1LpbYeU0HovWxpivpCt2
gwvdw1lJauWOkdqRVtkAA4pHEuC8GC4sEMszcgkkoNIg2oXj8imz6CtLG2E6sHCoj75mq7ThpRgC
1yLY5RDzxykvXxH6AuROAWJwu62gy+CaSwTnu5Z92UOywBQTZ+mqDLnLpIQEHXALW8FtT2cWo43W
AlwgoYMLf/u5f6A84b2rEaRUr2WYl4GWh9yMK5mP8bnwJBrGYW6rQVlaVi9IdOFSkw/8sVrNweNR
nOF6HYPQx7pej+PIcHYjDN8aLjz2xR+qeiXuGPAOi2JL0O4SGR/372RLR1NLTThCPpmErQ0GfvdX
oQN0cI3/WebETfVtvnZ3ZdpKA7SfK1lZXKBdfGmRJG3+MXAKBc3lL3BEk49qgPXemVulWrMRZRzx
kRFSp0LYpmqWsHSx2ZaKOt9CBZpfd65rA1a/ikXOnVFuIHMCT/PCFtgRcOvdilvHKLnGYcTk8Hxb
dqyB0fvxo+PmitRPyA8bW485ibtapM+ymEJvIJPulf1FGBQu3X7C4hSHa5wnb2j+nelp7SlyTG6u
7rtZ9jdiFJNVLrC0BMS7jEfZZ2+V+S9c2PFjKP4QxVazjG3rK2lljx8vh7RIVk42cSVv/dv9+VkP
JLCDpBWbotlNtYdqNyO5KAvy5nH1bosgRlz91Xvl20xLzffHeVJFZkcGEb24wlV2ZApuBZDl6e8B
cRcBpNKToIL82jp8ZNW+JJXTiJo4MIWBLjCF9huQZPoeahLkXs+8n8CqL4kzJK9eJVN821f8zeQI
6a7eDiXNoh602cMcy1o9UOSDwsYYdLpMgcDHZ7+6BobdYkiU87DNAX5jq8Dz+iyWLu/ei95tP2Ps
ISfN2M3Ef33/lg/hnWmmmnBzR4Z6t8JA2x6C9v30leLSwnaRI/Vxzq6hxddOCY8ocrnLp0adVcDz
vg93VaaY4kV2X15y4cmVI6yAlFad0poj0P92UMeEVvMGqpPcz/E0ILD6nwx0OgF23fB+meolkQKE
kcgic6/FLVtFAIC6iJ4trvmkQG6VyhvDkqo/z6/G2sEX1umMlFJaba/uJBquO1v0ylgscrm3Sjt0
knK3KF9u/Yqu47qhb1vqiaZPa2rpaj2VoZKsjDcutnTLpDveXG5UkJG3y1Hbp50KzRImjlAax0Tp
sMzScyhTWmwZ9n1mlq2/oPDOPt3G7M4w3991ODRgLxGaJo2Lta+kkfoAuCXQdP7R01ySSqKVinEk
3t5LnCRTMZ01udqgCAzwbfOLnKtkl53apF67zaNRk3TXej2FGophi1cbJD0KdNaxTORFvuBJel1R
O1mrB0CoFsSIex7NEZaMomr7mGC4WgBSbChz/wjIkpTnyZZwcncNF85Bw/7Rtc6MrTt2doaNrSDJ
LUWfvjTybHIsSrYweBTes+HJESajl/M32ZAYghw7+/KI5sEaSUFmJgxvybX3YzwLC3cxqwkNr4n0
tZZm71Tbc7bkzSL+MVIaXDILaTshRIlc14PlWcNOgVd0IHbYbpMxp2RqlUnCye2lhRpJ29KfdUxq
XndIXCcrOLrEfuEyfgzfXobKJcu+5guoGCwZw/bqduZ2hBJYYpPdYZWj6rO5PsQVqTV3IxE+Ud+w
Fl6m9xdlamsVrBQ6/y61JUFlBu6rQlccz5TLcYmGUyiN59CgaloYSrXCp11r6vVx8SQOJE0VWGim
rLU85B6OgzXPKh/NwDked5pc0K0+jglY1qmuS0tdIQct0qI+iQ1jl1VY4fxOFD7y+/4tfx5PAJrr
wgoVThcyg+D1V7827Ue63yelSrQyCA1l5179WfAsIzTAMvlZhnljpjTFrljH0DxSzwMIHVRHNWv4
NM2N+1AkyMgXj7kdq6X6EEfkQ8pnkSK3KJH9Jiexaan3xH1+j6r+DEUUIX3+aOzRP5u+x4E5ZBdS
qVUkli+cPTj2gDzb4BAUjgBgd5s4hWMSY/ch3hLds9dLDRBk+8uc5l58wbSC1xgIt7KvJYUypP0L
vcWwxx3alDMEp/oQMsVtZqllzVrgT1hpvIiE89wLwhZ6EIFOSER5JzDHfz9qCFRapVPhd3Rm5SJl
bJn1JkUs+GkAD9UeR0xWlgfc3Rd0sMCey7Ag+tw4E0Y9tUzsu0m8SZNi4K0fJLIV8KNLPtM5YLYK
DRsxcPrHDiPNuyocZ2hkUtXiXUNZwtzfLHEv7USexnzZNnHVmNDZ+/mOCV39EneAC6CuKmsBc6/k
HR2sUo0x5AYXmhFURxy/g3sBfOr21MMVo8YRaQelWfg+tpwO0TLZbB8gw7Ayn4kk2iCfMiObC4zW
JVy02lx5+ujtyaNBCOPxoOMTkwwZEMzlY8fIO8rfVhMmJYsSqtzd+WTo+xca7atxzayuw+RQUUuz
JU7+W/EqpbjyqJadvTp599lqV4XY/8BlqJhp44A2AHj9dzcyyhpH32+M/hVyqTPLKDotbFXiTizx
wwZZVnTbmIfpuvMk5YkH8PEiv66WJQvs0iD6PZYSyaDM5XFs+99qXvj7CKwl8QMX5LlwgBNl05sL
ox3bYadFma0soJW4oD+u356Qn3qeArUDR46bYmBxLyyWkmey4yeZSnVA+ca1EUbGCALhsnuRtDuZ
jmjMVwEgZ0XzIwmNXA3Ju+shOyNW9uuk5SvqXLoKCQH2kPi7kG7FH7a1swSQT6cg9DSsr62B3QXY
1RC9cP0/gwINly5vS65z6/vzTHFJ8CjnI12fZ9Ehp35ZkppBP9gNWNXHjpuSqKb8Wi4GR8oKXl5b
w34KK3ncA/Bnves0zw+KdGP/YR11OeQZSLPgufIvguajeH2zOtEvqzESOYcSeJRDbtAlSRKnyhcu
LBg5AC1lZDBk87oDlQ8sziDwoa6WdcTCzbPyWNtiLaSI7zUoAZHPG3duI0DCu8AgWVLvW2aXDe0b
xoR/StQgPI7bgZKuPpOKft9AuE7RcFJvPoFIGHB+0s5L9WV23q2yA9PkvGkS/Pm2qWfWFk5S8sKP
hZDK+cA/4Os+M98E9mvNI6HF8qAy2NoeiC6wM0GeTnfaPD2vSQ3GKaWhiEJzlzMfJqPvsMTQwU1r
YiDSjnNfVN1ql6ATeFY5aO3J1zQaly8tpF769umusuI0rahT1P7HsDtnaqpsZm/XrxxVjLJm4ekt
4sBBrQ1bgbEiRkdeLYLGHryqGh7DnyYANJ5/Ohqkz8u/zT6XJFOLeKX90pTESh+zgqB4g0tEzt/z
3aCK9xqiKem2WwH/+dJaGa9HnIQi0OvATHCR2VR6NgT3xCKAtWYrydZor+9JsTma3ac9p0sseMhQ
lZp5plgN6xLFpjw0ba1QGHKmPldc8zTLMEC/8Eag8xeGMVIVbGdBQJdU+x/gLdqHk7WOYBNTkDmd
QC0m4rVy5b9Lnd1a4tuS9g/QFwNYOyXu87hqxU8dYKH2pockFlyj6CzlomsDFXalBFHhKpGnPpRa
MvcUDbCDMOqhOWVRzS+zZU1/64/W8J9qnodswXo7sJebVtNgQz7YZ0HUL2gPZRHhu30ByXgvoleN
WtL0HxFbKjLAYc7BsPGQIlqJYe4cKa4QI8EkXSTBv/KjHYI94j9ewiE6E2t0RlYlEhM3WhtcM/y1
FqKr5LvbVG5oTvJhuOlw0748bw7qTjZ21y5OKlDJQ2mvOZ/N6k7N7tzbCc7R93FJOuKmNpzTq0/6
TUs6BWSC/eSoxah+/0QmaD5YlLgvsboM83MENYI7f/G2FyJJ6xPC4/U9hrXR4d3zcDwVyMj1grXf
YzUF5XWJqqrsGbYv3V6zoyQRVLeofOqq/bUx0a2N9LLX6jN+siKTGFWGvGWSlFFfjIWFsE/7upVB
vDgJi7hMjOvaMtykhOSevrWCYoK4ej078/f5q96Su6JL2+Huu3u+L8jO1RAguzb4d3nmpKaWmCn2
eyZn68RM17DCZJA2cy6DhGXELRIjmyhLKV2YnYadITb5uYGKBAoZIsOJ1U8Re1Bp8n9/ngw9Uex/
a/G8HJsOLcTO9DiYyxaVUuitiHZHdG+QIi6FMQ7uKUSGWS/66NmPSsx0CipA+C9q7xwJvpN2khwp
qiKWhDoQhjRc8IE1nCHv7tbZHenIwflyZkrsYzCi6JPlQwQWqZR/qx6cl5/8sks04XhyScokRYCU
OQrepo7yMmhCSdbF6eGw3jv5IouNAdhITjdj12ncV2WvUc6Te3nDFFRev/a1j0f4XSkrk013a+5C
W0E8Zwez6Mu7WZ1RbGGcHyq7N28n4S0wO0lH3w4FjeQq4TrMZRN2ne9tkWBxOXQyPtSJhZb3eg3l
B3xUp0Xi/ixUjq5wypfsLIVRgLL5DQ2ZWDgAXkwtZaHr6sorYAG/yA+L7vZ4qnz4ar2nzUohgojo
EIrMJ7H7Skcsvv9sFS3rIyWEAN6ALuXq9ZkG0zFTgfwqgh4JykjE1W+Z9Qmr+QCoZ4DlPkRqM1rh
0RdX4M160qQ9rPhb3EhjL5hV1joCPJrpj3Sv3NpVX7/emyKHCBzuXkXUgCWPxUWui+jjrgkOYtNj
oxols8OzTz3cOJXxHfRjSpwyYIEijnHCWUQXdJTjKKQs6klhmxRS4uBPyFp61SnMEbx6fZSgWzXj
ekvOMe+wYPX5Dw/MHXel2H2iRtKXgfwzOxBcvZ4cCVwhzf3oNGkz7W0/Icz6/jRZdi8YppyW6GRn
Q3G4YmD4B6a5usH5on/1jHQ4Pfds06ImcG/OV+OQM8p6ZIUWLIcdxtgzQ9gphngORbNv2Oot66oT
P6uqEeT1CGL5MhpgsfaZBSQgsmv6M1tRPB8Vbk9VdfnhzWmesO5x/jGUBDn1CXkxcpNpl6Iv02fN
2wnKEKCo6bGeWi3sgAAPeCIcXNIsKA8obKPfa6qh/XbixKVnZeOUeB128Pedbbrld9GCYdTvfU9Y
m8uqO7vdamTUTXfCQhxfAVhuselSfbE6UfUxOxfPTJ0qnUrrLwlr2g4r3b0ZxYcGFTxfUIfrIzrk
3bPwBlclEI5s30nEsqxQ1HVlC6qO4JRBlPAoHkduJQTMp5hPyurmCcoErENAmkBZS2EVWoCwEK/S
cfAl0PW8oQW/ek4fnLg4drrcdqCYPbIYJZPtS/I6tHXsahaJG0Jmd678du8ioZOaDBzE3o4KYFz8
DOKUmCFstjOrY0GEkm4/oyM5fUmcTUTkGwcwl4uYenlo4sMI+/LVtSAu1C2faSboWVhyV2kXSOu+
Bw/Bv04dZzq5w3kKgVGztOWwCFJWzU5RjzDT4ZboHtEYO+qvTY5Yv5jTnjEqUX8r8Yl6Qghy9lJS
Fzn9zXzCsZasg1Eu8kiIsmXaHJ+F9Q5It3lfXolzmSGRGfaTDC0UlX8bbs2ZDJ6hESgwT7vzi79e
SW/cbOb/AQzUSIu/8H+AJ1hJki+YJwgoDOXeT5eGBtEOV4cEmCZWiPz3r3MB9tfFjysAtcQV1Kor
f+OHMr0S0HYF1zh8ajzBsk/82yPYD9nTlkfeBT4ovG69acqqkcyrXpmBIUcV5MTR1Bwh1pfTmQqv
zThf1KKwouooYPmE4MeFqIjB2OASLmgOU2J8HVXqi8qL/rTTG0LEpCOhIkJsMAsSfo+Vg3/5OV8B
YsvtzkOtWXhRubhqdFC75TZbUnf0hAkKBi0QuWB7Yclo6Nk1Py1XjPUaex6EtTeQS8FDIppnsDqm
nEtP2rgnxKbVfg1HeP+tdWlq3pcDKBSH9smRohKNiLWb2eakD1j8izQKep+jLeQPn1QiXT6wSXws
9uFj6qweVp/A+wSYs4yrSajP90VL7nv4dZsZdjM8S8RwavMogwroC5CS8fCNmo+IYhkk2Qyum7oC
v2U1sgT9lLaltGOqopDZhjXCWPTodatM+ZgcX8/bmoiCwVEXkxV3I4AyxZ15vhAJLHHhLYas9Kcg
d5UkBHW1665y28z5cGuTC8SwKb+InFD34JvOxKczWqX8PPxn6ZrU1QLKt6QyBb6tggV6z0EsY6us
G/5Vf4KctsqqNjziC6Ow3TZy3vwyzsbmSzOe2vQDFnVLmp2OH1jFgHZekc0KbNyRtUM5cVXQrC41
lJiWdQI0nFhSrcsvjemFHBVA7QZY/4moAa67fbAbTaAH81vZj8BnZgyGAdGnEJR1SueS008zsOt4
ByN5M1oJTLydv6scL5udT3FXktg1K92znH8isqyf1erEKkYyGmAaYu1y4M7O1QjiZ927H97FL94X
OJypJC8Eb8pWmtxeGr63UlvnguxnGvtpBiqFIN/6oPuhgVBBnMs8W1FPtYIzZWe0a+U4YEubodgf
Npi1pJ6Zoq+VGAFgh9mJsYzXwQN9MZk1dq+dARmVU4BB0ZPnjiLPhyGQUvFLFNQhtfRTl/sbCnwW
MKQ2irvN0cKQrfgIvSG0Q/RAoit4B3Ztv+rnObWzb7td+Ck33fTUWgN3B9we3Z0wMs0XC2g2W3op
Y1nEQyY1f9nVhWNjHqBp2pLEUKPXp0s1C7cbivp1HrSWeeeMzXLlzlTAEaqqSxcsUkZMZGjHYXy0
bONEuSXzJDpbppiS+vsQLIbToZzIshJ1lJkvxLDgUHbfCZ7Tf0G6HRWlDUDsQHKxUtsUg4/jjdZX
SqsVfpZulgkMEiXGubAJpeHhxn9oRwHUhi0TsZM3HhkillVGVXFFjT+7WvxVAjIBQFJoKAfl4n3Y
K0bwE53dwH70wXb6n4Mj1WG70VSekP50amdJCdrkOcmXXzE06cvLqyjIAB+VEOGjaZedwEpIAaxu
irE16RZ8H5A0/MgwyEQN+bIvJxYqdO3/Fh1jdKZOGz9W1u3/bSFJ+Pig9KZBK2AA1eKS9IlNBHXL
vJ3ymcgFDi8qh5Qcvu81C4LXstK7MY0cZp7WumfqKfZbZLhMExJ0HXVFuMeEQKn1tP9hYqqr2SP3
59ksCF3nOctgZEki7JfSPoNcVprK7AdL06u3mQHvfR3RoCrhUNOoSEddxQ8HLVnryhMAaQTQL5Ug
hFGYDhI+ukxQI6tbjkVnL/irXYrYekt7X1OOu4/jHIZWTX+uJo4iYSOR6IzXGJt5kFLPQSDkD3KA
mX+tjNAJR1aszFBfwjeJXj22wwLpVE7mSvBmqGTD4BxN8l2EO4DKJRO2ZRFBPzzIc9B3ocuCDhH9
sOowoiFjzSg7kdiaOEpS8jomiKY7wwgEM8yS6ohc1XFReKPLR7Bv1O4gYmi/VLcVUok29jfaKz+6
ENAOoA5IIrjG39ai7fGPFuvSRioi5gRp39HOAbWSX/NEMbP08RTF32m2M6ygkQ0UbWR2Dpalu6Tm
JshDKtdgONUzq/inEbbqZgtz8tkY+GyF6BCO8Ejx6TE4sWwuKTnA+gDsEYtXw/jX1MpA6UczE0sx
yLoCR1galiqIpN4sxXwdUs3WZf4ctFFfSWyAkwErjVv53y9KJMXUW4491RsPKMC/2Hm+5uoYxiab
D7gsyJS0XLLSEOXy4bAZMa7JBmXSOexKmzXgRiMFcmuccin7M5CYbvDt/AGTQy1M1HbtIsnTPggX
akeLo+jbXxOU7iekrgdgIR86jcsRmqYql8MkC7rOJoxGEKsbfk1DBmsy2PLKPAr+Dzt3umSZWDCd
KjxZz3ZLPiEyHVBmtc/mTrAUUC8QqZw7F+J+KKJgRExTePm3OtlDhYEaTcPDfKuZRM8eSAhEeSq0
yb/g59ZHHP/qVNoeG/+YHBEHrKhBSBNuJjmS9JW+mpu1QzWmo1NDx/DJ5uxKe2VhCaLVGuIsDH3f
M0EX2JAdOAIqP+qOEjbE/7Gwv8UGLf/Capz5Mgfh0fO+ioprCeogjTBw4TiDpQ09GnEX/PKxObss
JCtY46jM11sAMjxj5hAqRQnud+VDzr9LYkkJG9+2Csh1jPVdotUwRJJKb68k6nE/PZPfGQh6Abu7
89J2vVD7rsJnVQnM5hqa4ef0dbmXwWMznKDaHwTVuAsblE7gYZPK6sfG1T6JRUMjhhAZcudR6uad
hqCH3jdIrpFuwLTqAN/PPEDEMjzsQl57FboJZ4W/7J94YrfKnd08JY+030+jghSyyiPKYTQ3cnZz
Wufd9abZDbYpBqGPVgiPgkTP2/ZP0jolrxOzre5+WkBfl1Zy9sMaB+LcF7y90f0CUEbs7aormZD8
DSv5+XTxhPQH6u15PoB7EsqV+FooscHzKQD5ziGBbyoN3Ctg2Jqjnz3C4vMEYJk8k9nuNLqUnhrM
M66cRfxvhftBtHrXM8GB49t9gCQpbxEQrGF9m7hvBPydnKqiJwg4Y+cpBYFH60viPKKkCkIa8TPf
w5vXwUxSws0E5DaY3jxZW2talrcm9+Ku+SwF4P+wkCwFN2Bys7j9qCs4cdEFxIaETHUuaF1mxJLV
hxHXOhwFxoTPBxIfSY5+wy50Oa65qbKhRqoYXK0BgYPvBGDJWFEyZ/qDriLOpDZ5uuZv6SxVtsKW
JtPmym15K7K3NF8Ebt1qqx0aH7TTaCDvPpP6kdtXtdDcnQqQvQ22q7yDFEVrIsVRcTBxzLlU0TXQ
ehzLP0P3WUTcWuZKUZsZNLSvYLeXVdrMFRdcnBq9EQlT8Mha/WwmkGvV3ooQbSvevrmq3MigdVOZ
s/uEw8VBWp7vLnop5gyLlKu/+C/CgwbSZhDC6OcYKc2B1vYt88BYmLrA86/PuOzb9mV7jXefp+Sr
vR+PsC6sBQtyGocD7kDwAhDxkJX8rqc7iFLR54Px69BKgijaGKWhyw5+gSwuSkkwAwu7JoKWKXVj
thVPUJMzBBXg5oWTn4dVJnUQ8U4sUkSocVhhgjvLn28HpTD2FNIGWzsTVE2bssf6M71H/FPeUaSh
/SBCfSJFg3wyOO7qkDWA06VkbJiEXeSPvoS2BGeIbIHV+BeVVjS1Hq4jPQdkidquVEsazHclfNim
vpB0maSn5DtcvhJGcGq5wSZ26Pdh4VILA5dSreE8gI+7LMuiUYwY5wt7wp537x+6wc5pUNCtraEg
ZZze/GjbNf64L1hnWc2cFqhC33tkklXDIuJirb7f8IeceTzXN0xeSJASg++TEwUuTjI1zOXzOnus
ocnrzMgHOUldzwQORve6U3o/h8ItHehIWttnHqMDpwQIcMJEPcLfj9oiuU3x+v8JUV+Qf0wFKAwe
OoTdE/SWdBSF779xvkH2XQpKUjUAMlaBYppbUDQn1tb/F89wTWKJ1ZgJxrj9c4S1dg6m4oiA2Q4U
L2nOWZUZOR9nIEU8HuDen4+534KQSsWcoSn2ohsZzzKAAj9l/CpxMiCY7barDMAN7AnDUWPfXcX8
MrCL+F+fr9rkf/cPk1h0MC6+63MQnEn9AELVm+vVgcq0XnN3Ahxjq+9vK+UQxJFGk4tABgggcAlq
aXLjUBZwJbkJmIvfqw/mw5euaZQcTZuL6LJmXxio1+dI30wsfC+dBURpMWRp/4IMhe2sTJ2ZGEwe
aYmy/K6stRm91PaUokA7fKqw4fbPI6iS96c3MYk9iKMTITXvwr7exwsO3yLJ3bUV3393AzjX22ZL
bFui/3f8N7rWzNepcXHLJ9EQfYamKPRCjlEDOiVvK/GlQkO94DF089scbzU9aImX6/Pc9w6paIwR
Gd1phAv9voJtrPhBai4mFCyul0dyWhhSiRhwdGtV8GezRyloKYVxbPEjc/HG0CcPQbKH941iDMKq
GZtxTqg6V0z2Vcu+dU6tF8lfo/hPa+XvM0xIyKd2HibALmNCc0T9YcC+b8gMUSAA37R26HFYmNq8
XnJuURGh73vgI8yv524jObQEGvCq8nkDhg1oQqqByO9+/huRRaQbgMxKYQDJ89jr/dh9VhBDptJb
alBtz/7CX3LFcMLUTec3QIOa11vMmBKhbWsmCyZLqTY/65IZnp3jY8Imdr4MW5YMxLM2v1iYBkUi
JgaZydUlkgH3yKrRBoAOZGw62bMLN85KRPkiTujHKHunjECWnjp/u+/Io/3rbAO4bsDqwp1PffhW
SFp+Pv2se0bzEtSj4mLC/cPFhAERumyJJjJGKVP7z8UI/ft3vdCj4cXPjs5waEK0c9xPkDL0lNdf
GaPjJ16nhXqP0J3ZqMRfl+XYXW4XGU+oV9PKVn2s9Ewyru1PMEi/8BtKoNPD2ZY7L1v0f3g7RsCY
cCUfeiahOyVEx/CKLYLp8U0fXctsRKb9PGFQkJ1eX2GgGT0rh4A0tUPGVfZQi0nWiq+zg5d1VOYo
9k0HaS32YkNSvJSQeRD5Se+48UKBAhST2yXBIN6R7O3IyXB8+7UhnTtDD6m05fkwn269PkCtJo5o
N9RFSA4awCkQi3/urOqeyCGLcipiP/0Kb9LHggIwizN3/0S2I2Z14ROmfFsbVYrwpTbzTkVNExh7
5zA40xDXS53nKRQj6CHv/nmGB0KTDdB7xMzEqbAcdSdi4fGyl6W4H1AMs18Hs8tVaXVZpW5pmLtb
CvrW4kUdVWjJS3fA3o4xGxSN+Z2sWDAU2En42TgKUUWSVCeuirRYnGij3hkYzZKFMgU3/gP8sk6O
9LSiTqzfMVZvNCGaRD5T8fv0vGxcikeNh/Sz1kK1cjElnaho6kP+Vw+c2miCWbh+9X9AsBeTULOB
of7ep+SX8cLRt9sfP/O1nBvri5PtHjoBn5ABH9m3V5N7B44/4YAWASiF7Xe4x66uq/uWaMbgjR2Y
OwRPbXnle/qs1SvYRMsIIQllz9VPddaH0Kazitc/i5t+1oLHvQw4ICTcK1kr1XAYqPNHzhjO94ns
H3tHI0aGlZYOBaGZboqUR2lKTRjdzKbcj7hbAAlsmfnWxUOcd6LqJwGcenaZcT0EPcQ6JqKJXVlh
UlIYw2nuzJwpCDpvP2XJ0WAV71CA+OIAmJoIuc7jkubZ6kN8CEUrGEplLMHdoPiSAko4kZvlcs9+
lEmwYBtqs17lua3kvbsdMVHCuiIhT+t66UQyJzYrMNkd7bHB0Ao1l0fVKp+22s0ZRBWM5S5mlcev
laNFPsS799yEUqi1RxU63JCjOSnWEPtkehJWc3hXTsr5vQRyDJllNvwXFP8K2QraXvtbDtSeyy0Z
Rrc1xTa/W7AEOpK/LTVlzkEPpPN6gC3bqvab8EMOu3vTszIc4EXESd7gX83hpbDTpjjyCh8r/n5D
GZ7VpSCD+dNKvvNtg8PK3w35K6J/iJfb9zUV9qbPVcTVdhi7dLb4LDMOLDjYZ5xbknq+O7Pgx8FK
pb6s3U/ESdeXn/SL+TN073hBsVbiDUGV7oJuXPpyoKArzYUz9RmzvTULfpIEmg8/JlHoVmIDl+19
LPKX1fX8fP4A1MQ+UmiN76YhC+qRAfLlbIcviqwj3krxUB8bIKpiqUwG5fLVTjKZdV6VD37pDpf4
A4nALNQpUiIb4IkXDtaYDZlI7Zj2ntWnRggAn0hXKk2BiMZRrM21puRflDhRgKxXllmMwUlq7nqd
0+BbbmqAgWHbmyfajV16UVRmFsdaxNC3OxIiNEsWXrK5/adSFamCdGcbzv96qEC2q7ecNavyg8qo
x1c0kVCPaFaaol5PpEFrS6XBFTN/6YXxDQJmqHzwR3+aecNBeA8vtapzIFt7juIOWxWE6pVfBmZy
19o9Tj5Y15Qn7a/d2+PU/F0o6O9Gwk735kAio9BKTb8dC5K5c4AEbbuwaBdUyBOY03P6b5OKVmgY
5DCTXMc2Q8UO4wRMSMC1EBuOsMuK3IooF5d/Np5hCCksaLPiQfD+eov/Hz5/W7948LX0JZJMixjl
HHhDe18KsKI6QkVeMz7tOPNNXPk5bB+8Q9zb6wwGSs79hCjzry4ES/TXcNTax8X1KIx5LrpD40OK
dfu9Y7ZRBz6rLKsVbBq9qXJtgrdU3hO1n6KwLyotMNgoOpQzTBN1VWzCAz5pSN62BoeIkLTx6Hdj
9k9U2a/osanF/a/EdjTfnlexshiAOXqbNT5U93rp8lJimIbIEdKeosRtScFuzDAPYPN4RlhGdFpN
Bxi/RFRkWYu3Xv12zoCnjG2JRw8mADxjKqBeShTlODd2ICNOll+u/9Eh6A4rVlPKs4hREimulPde
blBKarnUnUwrej0xrMQAQhVxb8s7Kx3fFztf6DTyeMadIliukw6s2gBmOFYxuXBtr+3kK7sVg+Rb
VRtrRcAA+A/pZudhbi7hbAOBePwU50iHcLdytcc/lnNBmnqNSg96JjcMwihX9SDxros6bGFnuIRB
K0kfa6p7NTKyL0JflDo810mKkwOPkwbA3lwiWkPalWIJWF13vqIlhebwkvnmYbecXTb4Ld7loFQg
fgv2s9S+9Z7JCRzTCNUYgZFuJaVA3pdhfRrHGs2tUjuHLpNBiYq1uUuxqPysS6NjHIRzya0i0ija
GlKWVOmuJNi74LRSa4y3ia5s1bcRrttwZ4QhaFNFjoVlnb2LL1bLx61cVUgqYWbVZeXH9UEEdpqB
ZJ7G1Sm78Qe/FYLG6FYMy/zBz+4LWOBWgK68th9+iQTluaMh5bD9two9IYGev9ADxBT1PsDIZ80J
fP/+lbSuhgEoW9VybwuZ3IkHUyFLiwiK1b2Fn1WEqKnuUKG5jvUPMDxekajJj9fV+puoKnxLDTkX
vS419fR9szZ2QySGeglWf3BqYESdJa3UjM2UvTcS83mPgSXpthWXxUT1jbGoMscK4KdhthQuCIaE
vJlkLosRQjMZYG40JYmEscpBT5yokaVFegQdB9wvzEnuoWH0hCJfVYGNi5F6g5aOQxotUdW2fXb7
59Umal/cF/hbZL1EM8b4SlroS3RNEv1yJtAo5Qs9suK3YaN5kq2krEBn9Zsmskr+zdssrhP2QXg/
++694tke143CtUuIhPiXjD8GTU0lRgqAZbUPWxfuk1k6qfGbEIMNrM5IktwFW5oJN35kTOmxzrrj
DI8IlO8TuCnbl38uYXwxE/ECardKEgb+rxaB/D4PUL6/yu/N5vRlz+9snUOnUzNHaTWN+Pp2TvRu
bgXMnY0j7i9CvzOCAO/xXul9yWNSvRrIqE5EhIMHxflHdsrNmE6j4q2AnXfGMuKAtz4+cqt/wUoE
Fn7Zy6xbYWEOY6GCt6LX5DoY4hNhVF5dt099TceeKbLHTSXiOdT1dEQcwSt/OW+1R2Wksh965zD8
VnBYxyNvIvjBmPOhzpYZwKrcutsq8PiOv8nGc7KpAkKEzV6DXnTtFeudBGLNHRZbzEi7aSp/aQFe
eCqxt6r35ghB968bMHUohmUAAKQCIefzQWLi0R7cYAwdu8jl2W51SW+Xb+qB0LH+sVFbvDVfrFhl
y+Qpigfip++lmjLDU4AV7nTYlJa4eNhXecldHViPqmTfo/hXDlFQXKVp0+UD+Z60nBED6HZuZKQf
cASWrLvITcSMdxC2OHpKc905nO6Fx7gI2BY1Sor34YNI8AIM064Q7B2/9AYqrYeq+ZllCrfd5sSj
fDQe19D9pMVMgLBo5v1xG3YciCI2o9Ab/IB/tjx/bRnYAB3IZWP7w3vvxhVv6Vd6WxhiB2qfhC4h
GgaVplqQAvPSNopL6d2YMv1aOql0yCrml6x+eXfnNKmGvPtGBTd/Enf0Oy2FPz9y+BVXQhbnDWwz
6+mf37C9sDxqXiGrkwHu1TxteOxaEiOerC4uPhQ7robUrpiJyeA2AqV+qE4dBymd3aETE97NvD2b
+f5CbrCcMGPgX/P0Twy0xcy8fn1faoIpfz6xvKbTQYoUe0FCfxzD+XFw4jFTjy5uDyZWGIhhV5DK
x0GM7p6eC1cpZNrpJqssJ/Yqmmsw+OF9blAvZR8MHrnbRnev4eue3QXUCia79t9pku0v/Ga9NVMg
NfmxvW2jJSMjAnmozRh4OdaDITkQ/xEG+QJAP5NjCU7+bn3G6jaKnN7jSRjP2pIBvICfW0jquCoS
0a/4xCi4ZgtvD9PGP+YOf3aReKuKrriJXRdOm5Ij4xy0NJfDFhAO4YgkkWldqXAFBSAMBiU29aGX
8q3F2Q3NXBpJzppk83Jfr89GopB671KO60pKeYo8Seqq9PRN9P+U47Q5kYmDsYn1WNat2SmQltsv
HK+HBvlCyVpCnBMkX59MXZ7spI5HVgJEKg3x2LyzmcDhn1+VJY9DAkt7URLuAIMC027j0IsnBTOm
TmSUNuHaXenX3SrHIFhslRMeBfV5Bgok0AVB1wC+c4+jevuvmyiZvyB4Ue58Q1k8QMrMfr5EW+Ho
U9+2+CfOSz1pAz/pBUQeXxHilANgWhRPUruvyClVwkXV0lvZYrgewfxOeuhctWXcS2T1hYtqM5MG
JaJnFZnJLV75DHex8BF0bac8/uIxU0OMS9YknGKYfv7Ii8xZbub5S4wyo6LuB9TLmjI4Rf5UQZa+
dIfUCJLG/LkrBQR+SagEBuW5zKONLPo5XqowskQt0SYxhI8/BK1616c/lHZKaGYhuYTX5J/c9oyD
FMTSE4HOKjnCVKj0hPUmQSfU+25UDoGagyo1eZBRQ7RblDYhLLiUgIUlj3weGNhyz22ZxGK35w+x
CdUBiOwB1Ofthmti4tgrEiYOiw0m8kMBaO7fld0FAnnUpzX5XnPwtjBxuRFU6RDCc0cstbC4RaHF
A09Dhjj3JcR85mA4a2B0ufV+p+aXSVTK+j2rvxpfR6em6gS7tcTZ5pBwQoluu06xzUObdX8aLNfg
V03LFFbi+gB1ltB5D6XRBiVUkzp/dmi359+Ss+aEJxT0hXJjwMQrSPW/NyfX+MAojwO/2bDtKwjr
N1uOsvD2KhiLlJ4ToHKkyaqKV8unzZK10DmZYo7HAGEZZqdN977bHMrkIDleZ+U5JHfPyWQvezKF
D9xuNibu7tOhexeU0KJIcIyBFR/G2LuXvjkLBW4fyISJnFi7qVEsvz1SqAIriH26eQ8IZbxaGx0/
D9ngBR0g+3uaYtVJaMGb/zFQLnYLUhzeHWgVeRpfZWo6qIWjrEmU78WuDlIWN435J4hVVa8Pdiya
57sKGuxcbczP679B2YSs3ev5GtiEZEy/qNDxRxMyK3m5Wh0551ZxZFB0TxDzD4Mxho2HLs2lcKvs
zNv8Cprl8jJCPcd4AERDgixQ41srq2/LrA8CnI2DlJSph+fSOz/+8YuBPd5NgcY/7HMiQ41E0NGG
xs9531B6658KB5GS/vryquP6EpWhe/xDbNDnv6jbIG3Vh//tDNZJEaHORIvXJeBrcCGOmq7q7XbU
kxMsfEIL0+y0i1Psz/HXQYVNizWUV1RUK9LZUK1L4588hz2fLMVKTaTJbWR0nwsYlK0FHTQCCoAn
uvbyR+o4/8AXDb1C/dkcowEdc3dXXIXxMFovYmnkwQd+de95Ep5pUOODw4gUvC72nt6TXj6QZzSz
SobHb1Et8peeWGZqkU/pU5T/ro1jbS8SH68ssTQt8+RHlk6VjTwUHULO0Ng04GWIaqOB6tDyBzde
5GlLN6UufQqBjiyMtQWlQZMQEQLMu17sHf8GihraYt27O4S708Uc6Ax7XumSpFRvrKHU4KU46a4d
8+dbUqkYr/bTSYeYGwDMU0nCij3B1t80WqGp7c29A9Ia8rInd321O7+BGguGIZHMv5j6gJpfV6Qh
lKudqHjhZ8/HcyOZP04J0Ou/lrbkQgFDule6uHvnGPPZjaHynwU95kUHZWfBQiep+sSgKZU9ZdsY
7IJcuaSzXGPJKh4JRftgYEKHgqgO+SumXIudlEnQYob11TJoFPKRb1bQdwvt6LFgWaF3KgeWySIV
/J16JyCvrN9YkzO+UFk9KfVF0duz8dql+ttgcZdI/VvJk97aU//0jcu1ELqUo2c9RUlKuaNhS8O7
AAZx6H0Vrh9w7ZlmcIkgEnAyIJ75rrBn1uIyq6vNjayCO3TFB8N0UkpLTPt64lPBYjiCJo9VBbVC
boylhBd6Br1mO8YtCSQawJNCH3vhNJthq81rg3L1v2nLH443NFPWHtNNKxTCTEXyNty8TDEh1tE+
eZ8I8sDM+UsABQ2BGxQUsCtdQD+Liac3zf3yd9N32+isRk5JnROo7JP4fe0fKcl6AvcpV8ziWDXV
oIPuuMCwv5UfiKsX95MLzNdVqd7Pg9rPzVlEQKdCOl+C8MdnksguNbRseRUM7HzzkqcgxMGajg8n
c9x4SHiZ2b/zfP7yaef2dtBHjTjSfN9xncDWcnCUWvGEIFnKO7TsfW9BUyZJpAyl37ALHRapRo6j
gx/fDIMwDAYrQkrKNaa0Z/2SF+o+BNbsHB+hLiuner62Wtnb9hP3itBPwW6xGuZucbdIynK73rSd
t8kMAXKO58vMx99GVJ5JNi4BEvHWFJg8g+WqEouFBmLHn3mjI13IgzAlCufO/dfF9OVAqAXNyD9C
SC5FYe8kSxWbBiMm1UPNYlRCaDbhYGRuY83L2DedHelK3mf4RBvNpjHysPT0krVKoJHKZuNGJQJs
y871HmXGM6cIdqr+9nTn59xGvIS0PrriWhoFIBiAqkWWfAzG9CLwvA1zf03miePO9q2IwqQz5s6k
Ecc0y4OxEyE1NOquPZ4HSCydmDYk5EOKEfm65dbHSb2ViufN3ZHZrY8gHdOm+XcJIezyhY1Sj8u0
eyoV1j2xQKliSeAk/qAqfLi2BWSAfM8wvVSquhb6oaZ5q316zf+PSRz1lF1DxEGdT6SPObwEKR/j
6FRYLgQt3qdATWoJ4JhsskIs41lPUShHWab3kI+YXegGwXaaYEdBxraA9MmTQg2VgQzJCHE7u0o/
27+Pcg8537ojRoQ5e04uAPtCzHMBfImila01E9FEn5cIQ7Z6m5lE9RQ0izYf+U6TdOcH1rrs4Ln/
YOzQKV7aY7Yvlv13V9+uvdw68H77PK/qMQY3Mg6twkmhIyua6Wnhbj/Umz56abdCVTKO3ylYAfnm
+278WmhobuCeB4XPUXZRudU3tpStPwrrtY+DUZkAUvGHoX8MPZKz2EGc1itWR8s2bdMY4UVymS57
L4H9EjyAbDQttHVQIS2XLTYSMJ4IwZtGlam3yDWTKsIgZE+OpFLEIfqOH0T9SQednLv7CF40njox
6EVWvI2FXChQbrovXjhW/kBxDYMCwZRV6Psn72w53g5rBHwvoYauWGF1l9lntB48fycm0fAJKkqV
qI0RMuo+UQ/QP+Wkcae2mmmA9xrVfYt/PmGRPhp8ty5ZU5n0+6YxSHQRFzGajp/NqNNy9dv/0zrC
KDQ1oJPobyeKW4CtZixDZyFCjU1teiW4QnyXlX1aQ+rZOIVfB7YzLJxtjQPqurkjmdxxovCAHra9
egHSxzEO6hJBwl9XvKrC4+kwtXSur1+R/eO1r7Svxs6kxcYW5U+lAjYvhSPujAPJDE1bUXaMClAA
fa/EoGd/3komXEzI5SWGbrHW7Bg2XSThhw0cPDTVKmsace3f7ZGEp9qKKJBJM5kEYyaEuuRenR2q
I5ADotzJqFPHjm/yJp3psqLfUj2ixwIIuIVZaN+NwMrRVcd12g8rbn5OghhAqxd1Hlbmg3NbHvkL
TQnLzSz8FPcVabP/FDXlVRBPa1+QDVIQfYhsypTZVHMIZZBzoJBHoTJn3M2Pt3iJP4HnNrwbFcW7
qHBYO9Wc4KWhDIRNwrjWqHV59fVbTH43O2aHZuBuYZxSY2wwwcaKOKy4InEVSMr2BvTnVwZIBKta
Gq/g1cabdi2CZkn1wz7eb3ILhUgljbOnvLVU/saifRy2yma/Oo9SBxdDEMV2cC0wyDCierjRuSPY
dRGVtIOiPSMRc637c8fy9QnExPxo72R+YGH+iBwVWOLildIa5fWYRwlbmqW+OTbB3C90rqW9/ALT
bxmOvUTdZDWz1Qt2YFuVGkUMP1m+7LizdaPO4bxR5TQfxzV6g0Pm666tyohfzj6NjwYcfqd9lYtP
pORU0OH7EOXjjS8x9ZdYkYZT5lYBpY2lm3UyYa9V1Enkab0dbS71H5WnlcMcRNaYuSg/ueb9sEKU
1c2dPnfo2Ca+xUlG2wAECxxQxZkFBHYNXHk8L3TEqz8hm598mzdxG882luMPinwofH2HhRUyAy05
r7aCCe1cTBKzYa6byxpnlJRZd4DUBdn9GU+o5TvlbJ+NGjFA9F7dIyQM8n9pVxW3zCeuGP46O/KY
Zd340nser51r13X4Uc7qTx4f1eBwF7tZhMlWkZ+tJH6a52AxZKw/hBRzQGcCaOQerRE2zBL4VaST
c7NdLVg40BNi2LPRvCi97IznWDHriY7P3rYj23EN3qwLggUZW1xImxi2g2qiMiU5AmCgK02qP5Uz
hlpKsr59UA07U31EW7t0XaOg7X6KtBkq5w6n/udVxSE2IOfkraHi90jank6mgCDPxdXIR7w2QhaG
jet8KvrWW74rRGA6io18tWi4wjxJqKh9WC5WPmzzF1lr8S+MoyLjWkHsUYePwrMRTVzulUa3SP4z
csmUqBNkLy8SKG8LZSvIZxdOdpU/qUXjk/aTAj/xIfugz3ZOCDPswAlJSwK0aRq+mq0PLH2uhQKz
Sq77ZSa/1fN4jbuA2qn64GBRshpE6TEJPCXeDbfIyWymPcvZPELBmid7UJ3Wpw3EtbkM2EsoP2A9
PKwlF8Z+Ldwl9q7ZqikEVQNX5GAutJidEOaw9sc260Cuu016REmhyM3SBnhXE8mo/9btpUXvMT0+
O0OzDx6t+ZGiDeA1UWCuRnqLkaeKhdUMFzzS9o0g2eQ0QS6cvt91H+5GAVT43pw+9PB0gws50K2b
ZoRKhCmssNbv4PdU1P4x+LOkVmqndBS7WDrtEqQeE2JwsuOfTW0eFpA+9ip0qOlFW2N463sFT8pd
u8L2Zdd7vX83p3xQvD8Ydg0gZZ9Hj+ccohX8fxjFzFMsz6GDh/LPp4UdYZbRbUWZurW/7mOXBDXn
RnqyAHpt7F+t58GNQcIwGLuzl1xh+FVi5efljj8hYs+krLAHliTkoG7/gB82lCRAKswlAZa8s7Yf
rCd3sx3BrKTW0gJP200UxA5DCihdTawqvFIPkUWdegbcfp5ZqEHfexvPVNRgf/dIOwJC7KP39mLd
X3Bwz9sE2i2fnJK40oZMUMGov/CYto6Hf6VemSFyfwesDMo+jOM0rFTicfOyx9OCDcyAkHZXcv6f
UQ03caPlv6aKZMGtRX9qs7CrjKsMMPQRJ1aXJCEGkq90G6vXFxo39seWaFZremE2AyU1gA+6e6Dz
9E76RALbkzroVhkYbwW6VJ44G6QDBYIm8mb07uE1+qbK7XIeRtp9uRvFIHZ04XIMsZ/zUHoLdQuF
tFyTZpm+SNj0g+EsmTYtzEn/rWxtGTmE9VpfP/Q6oFpGHaMWuEafjhQ2iQlX9Py8KMus7j77QnbG
1FWIMmptPxDJiyQfNXjE4g1gOB7fYt62W3ggHkb6PhLpGvgp4H9fkEi/NbFmOQ1OX418+GE0/uIG
nvaOPcbqAmiO6n9ue6WfgbSV0vt1Fj8FQfS/IWxwDYWN9KEZYwgregWn/PS0XlwpwD4O2TXFuUkb
UfdieMTazGBn+x2KZUP7cINcwM4BVx/hXrd7ajz5/bONZcQ3NzEbgmf4y7fMXoGjeOBK0hzNeDRf
XI6WGkJWDMK63MQKSuiRdKrlQp2vRdIHDst1Wt4d7+qC2yoM6Cf7PijfowybMAtZ2Th1I8Pi1FER
qc45RwvmRnAknCuH1mIkv3ZUPmo5XWsG/8GjvF25c6M+Owf0JjPOHjLeSatHd94vt22VypzI43rw
elspdh0Jq4a4iihhIt/vBLpzfxchwqH43aQXG4lO2o/y0yXIB82/mclbS3mLFi9sn0sw40A8Al4m
nzplqzFWDs/qOT8b66VGb00ISTPX/lwZ8mRFgBn0CVW7miavFZdt23aP9VYpytRny32rCRzmI8nZ
GEvYbYQl/F8M3qW1YHAb1JWr5wDsBflrUstqSIJjs6SYrgELZ5PGNVlQUdKK4bxtg6D6yprhizfi
RSFAi64btobPmiJ6BeTCOAOM225E3GXC4xInTzUBJR9JsRW8yTu2wvWt66mh4Wzb7SwVpccJzLo/
9emMfBhpB0v/ihXAP/m5Im4icxCW4bwJe3Qf+8Hqztv+9RhBqgq+ffjXwTwpLn7jMqFF50u/xmSD
VR5agh/Qvg0PCAV98VOWp3dVRT0lkDy8dTHVzCV5dIDDlAvXmbN7JqBHX8c0QwTIKRjLxoF0I8r8
/t5//AFJQLQD2tw1GsjmB5nyaV1KoyHyrt6dM54a9qJ+sDaUAum1DWGAf5sLMHM/pypFmx1l+tX0
aor9gC5iWRbP3I06EHYjig/z01w4uV+kJdXQV2lMGGVENuxm+mXrMLeEfLv2bJ4wx65iob7dZnNI
FGgu+V4Akw9y69oxkO71yc9BmAMo0X987L8aPiDUNMfE1EtchXaJMlb/80A0AYiJ7YgJTklIK2W4
QqN+T/u34xAncapg/U/xOaLGbE5/h3Gzlj7NZwwR/+86mMfXZSLNoQhHBPeA93mh3F4uegEKR21v
6Yz9KWGXhpUVg5YbCdTV3V7biSReTp0Z1YukIWPwxsSbXiVPa45Ed901T6Y/6iBaq32qEd3j6Zw2
VkdQajmof4HrZx8J8CgSy1Fo/rh6FIMMHNSJfacVZvbvbVg7SUCUQ0NdVs3e8KFcP4RVFkeRBm7h
0O6PXNczrIOROj2bjnLwhs+s/B1KLbP/kWXV5tRASf+bePmyBzub+Kk19GFG6nuc/bXeVsDiVNiU
qkSXQZ5A90vXqf0O5tORjjkYkE17ql5ceE1EscKv7mVeSHqYp8775Lh94h9T2rHK3RZkLE2qdcEn
+OO3VBV/jT7Mce0bszHsrHwpG34DvKw2L24+j41bM2xgeXeWigTeeFItGf6ai0ILCrIxiY/mCyM0
Y5ZnSvikyqQbdna5K0Dvb1XqatgY/bqvfpA3XO1Gq4nSocepR/EpEyF/kiWhy1VchpyhwfVZpU8E
V3BliCU99/AQqqPd+JWrQ9S7NfP+d8BnzpPvsUuE5kRbAvRvOPvUStp08HVGdPFDURNdWnQcVEml
GnlvjeuP1Q3f74pq1j/8p6Z4Ejip1IKyJmq9Ns8wxCRv1uX3Fzee/0LgxsoxIUGdbBKI51pd9jkm
UOIb4x4lDnPSMCjRdm7kZS9Fg3QnMwAQe+BbOTDDbVP0jsxXT5zodluCAT6ysAkE1p8VxN+C+3ZW
zpwmLar4nojqR5u8wAX9o2LooNvTUjW9EZE7xaoMkpZQH30aZ3zadYXjqYZxWMdxy89whlrwI0Mj
08dTDYVz/t3zuKn9MRbF01vzsYITKgxLhGRkYcVewvNudn0L/Wt7TO9x1XQKV0i26f+oWWKttrcA
YLK3vuY9jB3urwiLf5xXrG1YUmz0N4F/PePbga2+gDsP86TNgI8xDDSRfTfVw1eiQCUeAwyQapLo
tAGe5YQJSWBHweN0qtyiunvdPmbNe7OYnU7bGhvXuAgBL0NlQ0a/cDCf8/JkPu3CFiXK76JVenvy
64o0lcA4zWENhOgkxQK7Rixp1RcpABWTYFh9KvyLQ4aYgl7rO7zqeXr3dELwUIBxtZKzATKX1im4
oWYD/jLKJfseJqgJpUVROULipFLYZJm4Q/3NA14TyJURLqR/JwNsHkbbbW2C/VQ9oTR2m5zb1Ntw
Wky6KMu151qV1oyiNjC1oJhruVMMO9QrHyonpW+4iELkFYNbGl51OsPNQS8/MrzFwjHv/UzQW50R
SFNRASwaGBC0YoL6lUQMJrES102JlO5EwS+3GPmE6LquNK3MhSEZVjx8EhzNpO4ZytX3xm79g+OY
9GxxV104knK1X/4vx7iMYVu4BrZ0jMYDMeZgNFiWJNdg3LPS/S1V44GSwt1gIm8HHCEgBGUuoXV3
eeZfjb0awTQqooT/ewf7Kc6pg/nZQFr4PlzWXaCT9psckml0nxVPdtk52NaXkfVCmANmo0Hm46+Z
Te5WAcu1FoolvTYX0P+NrMX2ou6HtAYUg9t4xSWYUPyz+GS7HFnQLFY+2PKMvg3cK1PGRreC0X5c
MZ7BTGtIhLFqcUrGzosaF0ekaOoZ9t+covSQAPZiibY3+tl9KsoH8INmI4tf6SbfP/phPxQQ1ipC
B3jOLYHcjBcsN+/3mZknQCl8rkQV3SweoNwQ/tvqSqds+7bDImSD3ZzwCrcTfRjTBnTfa/2ycCxL
+JhKgEqOzUO0yS72uRQSiH2acFh6D/l//VlmSvWSnNLSNzbIHguGZE21/hpXwt0rLvdM5iaY66Ve
6sTK/g5Ae1uunqmD5n4Hjq5mL6LRW5YLAkh26RW4yzeWgW+a6tRs4UxoQpjV9OsOYw7QQt7ABZI3
TMQlN/jTvV/jI0p7ttLvw8qF+PBMkOAajgFP6Jn26BnhB64/RT7JpcV2SRokSlTv4hOCmprf1xLg
0pvUiQa0Jb2TvLV7lgt/OVKeNokhOJqXJdXj8cZ9cJ7gnTEDMWvIZcTdqJIQoiYErNaxW6c0IQW8
xe7OzouMsDQ9ZIYiAEnuloFBR/jkaMrP0C1Njv5z06CL+xnxtQLV5cMkLsXr2fMQ3PENPOG1BdWB
/ujm92TacpE+7MtspWlkL6Y41U4nWh7817CKu74YMfuX889mxTS1xfIfnPAgqWZjabwHf1nG02/e
8s3ch0MfUjTWuwR49K84fILyujRAD6gyPjvBko7nO6aYTZKqbwfMBWUa/AfgF7BVTZrWdXK8wieM
DqetpI8HFQtFtu6vcTUs8wF6ZSBVV8GUa26jKom7UAuRopRc++O8Hyk9AaWdYXDzAe+S8Do71P1R
fuhuLQOwi+FPDiPb4/wm9VUiCC/qYwkM+gJMgtrDsgZp5U+5OZ0tO5m1ty28TDvMhlqNl5GlhXvt
utq7NPQZ0SEimLhaJIccJdpANNuKWF6fyeM7XUmGOmPPntYtRcOkKoE6f+VLVq+LpVlU1pnCPJOV
fxBzlCO/maRRQunrCNwLi6mtHX9F01+6ptiooCrdiK774+oD8cmk4vKyinYnaeBczzKp6w0/bVBt
C29po0bPUid8XCdHr1IR8uy9et0nVzfJwobI0IS2DzmSX5IyAu+75G5yH59/bUpzLdTA9MR5AhI6
FJEUW/jpacAaynT4DnQsgz33x2AFCPBHZDAZjidnX7TVjLvkiY+vi3LzXYUcCVO9VASz22YdosfL
pqmiSPnHOdPQN3GEDF41w6+6fXQEYmezx1CovHcc6zZgG26uS9G1mWEAz1A8BH8Op4QaqGHMIxmJ
vqRyMDEJhe2M1BzUa131QTnwQwDuPHrBNCEy2UQ6h6IdAX+r8teLTn3VJTUYzKC7nxYpuauYd6JK
TIrx+lf7hklb9xI0eH6yM6ZiRGyQud8fXakn1EHEP0W/drt++5Zw8sYWtpKplE9tqbNReDWamZ3k
sR0Fgfdgb1J4H6p+64q0z8AoEjvijO7eup5FKYYwUPSKE1g994WxLxFigVlOlk9HChfQiOmuao/a
q6Yr4z/fPaYo72Q4BfSp4mmFUunRiTP2p4CKX6RzaDwsIkMOXu984Y81feaeXGpczzAl6vs+Jwpo
f8pZAwIwcjsGcfvQbLa8GR8c4TxFpoykx3eAlGg4w2mfSUnGClLY65jAqgiE53NWHboYvtqjAPsB
PCpNcUiXokGH5HJi7JVSzZWqdj27HYBjECk/JhgDwTMZaNe60HFiVbCn5LIZHzrX4XSH6RMEFkyT
huuzApeip1JdQLAPq5+vToJ2cs5qlyESv80fclhygTQeXud6yTLoCkdiubp9PiTi6P20WPq3iMEl
3AM8wacOZFr8PperM7eOd1CS5BNP/nG/pLRqIO2XIWWq6PNjoMcDthfbd/CEtvANA4b6iuNeqNFR
D5pGk18J/rmoNxNY+ezTNUyGAMIJy35gkYjr1YGmUwrlrMnEuOtKCvhILsO6uXEZtAdv2i2FkZJc
2QKSftevw7YtCdGIUkG0KusOfz2WG8ObQVYEfrr6Ze4Wm/B0Dh+eubHm6+1mcegYFjKixCWyVfPs
Ntn4RlXbpxOe/mmxExqn+jQqZgVySWh0t4D5yYJ4jWOPUgP2smtg3YH5zr11FzJgNnTmKE+buE+D
DV0VE4/jVvBoyD55SsRmYGo2ThRaUHqRaHivmOuHtX8vtHLb3v1aIHTlMacvBFLjVQV+lr3vvn1z
A6+UQurj/W8+eFm39/ooECzbyTuJCKCrmtW7tbhkF86rsTkjjoT60QAM1LjA3dKgfQPWF/3eDFC1
otnudhH8k++LXqXb/Xa1ipDCakRHtR8PaLb1NAik8ATomVshwPb9TDAW3SJwG96egmVBUmO0WJmJ
pFB/YMIc0cHp+S+zmXXCCVbpWH807Ww13MuwKEh1GDZF6DiU27bg1AddutfZLsDBcbvRBGiIKiWV
d/tf4NCGHMX6WVpLTW+CP5uGccOTWzU8Bg5uOEWZqXiypxYWLesqfw6JmkUdgCaRosDeR3CZ1ccO
A7LOUrIWGyNtLTeQ9L2CFScs2rN/V9/bM4LyNqv5PE8f/LtUpvHGDr/olaMuk0u7nDbmRPba1cp3
TBWdOkgbPJyuXcdQEMli+6VP/H2tERwonveH6V0OnRaeKuNmTSAgeH2JhunMeySagoQmfbz94nX5
0zw7hs4XUUuldZONt2XuPkjuNca3V5bnezG90rFDTehl/5TfPXx/SlnO1G2Ag5hhs90EqLLO5ImC
uhTExO5sQszumvHCcAcB0kUni1Gr9cnFBkFEP+hGmsjv4Zaz0CU7FqiaEUzG/WgT9UNN/0jF2XUM
rWJBI7QM9I1Bml2kqT2e4wY3+YaARAotZcP+2rVERPqvfAiI4bke89nOLao448AHhzBt9kyGBoHk
9ecpRUyw/bEEf6hd7rK87bWWnKDXnquS2ppnJY+Hvr1L9ZRwKR0rTeAfoaN9B18LyQ8nlxvBos7W
oOvrsXDvL2+jb4Wlo0YM2Tbx1uoKFrBJ7+CdqVaAXgSQOb/OVTekgn/fSMa0YS9SLjOFox6g/SCx
pNy7LaellpJoZMI2wr3/yw3RgxeB7RFLNVjJQ8M8TYaHCkDdJQ9rwT6/WCbNQFXObGTF46Dp0vhC
k5Xn2idxpvpjcrvBlkITGLsIxTWcFmVKetOZSkZUwS5I4YlCvq5AKFxk95/DTDtPGlbAOGGLJi2c
R91rku9I7KBzBWQjYMnWFgA7AcjN0yZyzotIZvVY4+CkjlGQSTrQisI8CW0Tly7qF14k1vrL26rO
pYviZYBfnhQkCaHlNpVWdFmx+Bm63uvhze8ZTD59MXWSXUUIEvE9w0Qf5QlgjXdaDVB0nHGKiSxn
0lYT02MkzbMMyIwyqh0E8JoV5myemNorxRH/47d+VWV8if9mePUIHM1+zBM5K2LYBZYU/iysoCwR
BFhR6m5WMExpEuZ2ya1xgmq9986txLZ8U4tzgJfiL4lliJQkLikGwdeSzC5/Plb92WERloR/BYhI
8Xb3fuQcwb4pR83KEFqYqPwIvYzFSjyPsUyYtBpQNo2uDaI0+ItFAXdqzVVKB6hgCwlKrW/ajRPl
izK83IV5yOU4TyxJeUnAa2L2a+HJiQAFb9jZaI2S47qcT7WU+fNpnG2jFBXrT5Ianhyznf8besIH
AP7YKrtU6OBKw1lU+jwM8HeF4DLeRR9Sci3vHEWUnwz1OBn4Hk81rmtmew56sjdVyowAUvfLWfX3
XO0OF0NdSuRCDQEWqu/iHtKOUbB6gD/LY2J7cqkzx/xRVe8Y5FGx09PCig5y/kIGlolwq5k+QAIo
lQmW1sF9iRCMLUc0gzWObFQSWNqbeQ/+BFFIDwqIX08wyFZA2jYwbGLR/aWX76UexHU4cP+bxyCM
o26wIfAjqiOWH723nUEVAtkB6gnm2Y+JKHp0RtNC+x6Nzn3/7dcLr7OiNqx2HJ+E7gxsEv2JXxQa
eC7gpTsH7C2zyVRAdctYts3LBQNY2r3p8oq/0sERdRCOZdtRg1NVXkKia9B9T2rtK/PvIlv8GN2H
yBak6Ftq3+mHrO0Uw4TduDNey7kVjAZiKp+Cgksj6/0r8Gp3EV+jCG503M5OaR0qn5joGXBTfRnI
/W7KUU40H4GkvTgmw25WerQeaNvExTtXxSmmJEzYvpCXGyu6oW6OigAWEbu8TggNH6FOA9Vsl+9p
Zk1Rk66DktS0I3XDa83y5BGK3Vp/RSP334ZEIAegsXbHHGVqnYkP5qhBIZcjDjLBzaOk6sDnn1bQ
OuGHjNSsofjkwcecu4oXmGXB/Wm4y9E0RP7EGv5Y0sRqQ3aqHoBzUgg3W7WKGay3o6nsQ2dg0mzb
wqk6yk7vae2dcaTbVDJNb3EZw3kM92UH62Lj63CjSlKEQ3i3jwI4m9cxErd5aL7VmcLdd+iUT2K4
20GWnhl88g+gzSK47Zr/uwJ3HIa94r6+t39fyA/Udw01zmG+o12qOBhwAHykNjBinXxtBx1bXz0w
Xrfdg6QGifuK797ivqV5Vlp+rnkLciNZZm/Ozqz1v5upqeRjveQmCj5NY8T16xDAsNv9xBmB11TX
nCTHPzJ27wDPMh+8+q4zKIq+B5WuySlSq/ojcyoOxaTFjf/+LwKs+sC5adapwlvc3kqlnz3PX41R
f2/e2pK5RO99zdO98n7fR8T4Zt5d3+mcnqar5b88//MCfWvK8hjuGlFrYUsj8JbdNy+DYHuYFblm
HWWLgpb0GUis8l1cr8ciRna8R/iZJQVnS5W3PjszMJg4hxpowF8c+DFv7VF4DIERR41mE8CLqYay
SwkGWPiQNF+A/caTg2IXX6PFJ2CiqXFqjIZo1SbmJGkg7RAyooiWndZHYtoSC4IKoXka4Sv9UTXg
DlNxyWEd2zkk9MLYp8R3jGcRPhi4hOV6047gMqebx2yUEdOcqU4hmRZgLmJTo63zkepH6MhrHQ1b
hFhFzOx9T3RD+0XSvVW7t+0xHF99hSYX4Je33p6sohI32JPrzjWemV9TYsVITj+12gHyz7Or6/Db
UQUnFZPMXSgio4c8nnmTgZXDqLiWZ4UdssM4Wrtvq0qepAfMT2WTMShokhAQ2MusLM6GpKUj/tIQ
ONB8YQTRCQL0nwbQzDNnA7ZDD93CFffqdCUYLhczvv9k1YjTRopBhsl7LkCMcHsHE3qCcBhBb3Ge
adWVbFCrj5FOhNCvOsSNfW7YTw6UXzlFDzN+a36hOb3TdSZJF4tTcTcPWbyjldDgdX+4HEZoRtdL
SxUsRy1Qm134IijokMTDixxm5i6Ly1BqgXJgAvAP0aOlcnv1LPMhKw6STnttkL/vOkGIsTnV2ZFb
zkNL15AH8MVvN6SHLr1MRP6k4dKr5i1BzMjXBMuZGQy4bXSjbhazvqW7s6kTDnofTYiV/881WUAU
pzGwI5g8mKg2iFLsmzeLKY4Tf0uiEYR4k3K8uqMj+6+0fioZR7slMOi1kw5dKkWIBrvJm/NYyZUD
oiBUmWfv6ZqUNV8AL3V858KyTylskexMt2Ksr2OHOBwvcEnedhNW62cVZBim4SS+RkovviLU0Cta
nVPOfzgHaopcSxf+tUzCW0Gr9+6/GnV4qvjD5B8+uk+lMMHR0ZwVNkBErwzqOaYQMRGdGcDYQIKq
jR27rn+Bj+nopFbAcR6SsZH/b9wgRfWBBYkLtg88vi52F3QihvXHKjCe1f1MG6ma/29+g/FxwsFZ
eAthMTpJIcPExbSpZsMljpYE94IDVHEvR3HRjl5k9rftMuJdWMnhaptjWsFjBYFiWTspmydW1Twv
WRNWgv2AdercFYb+4F/7JJo1OQYRSfmtxk4Ymr0ewgcEzkOnSisUIC8Vnx5Hy0yUSqQS15MKpkRC
MAs8dXlc6tVlyNsej5wC3ki5uhnX6OdIcjgYAgRAVnhr98nFRP/wu9C5ghPpFBXSrHkFxjW51Mcm
wUqxzIVjlbXeb4dLlkZiRo7T5PzO9rWQY2g3hFY+hYiE5mU+Y6GngfByIaXF6adjcT7oCp2SOTWY
RkLZKd3hlTeCo/INS98Oh5MMvjTTyPCWdsgNzQDEoJvXM5jtgAHZWw+Rzn6EGI2i3H5JUwDJfvyX
AqZ5pUlSRIdGsuO/J538JjCBKvcWGzGUiAVUTAqENP/mUCleY0xzJwb5eqa4zoqBoiST4053059s
bNoEdvKS6p60fCps2A7twZ3bbYjUNFPcG213g1qotRGg4hwa8TIz/lpOkihzWMEzEshpxq3J1Mvm
7SMIXhoUOrrTB5hHpC8VxnXdss5v+9CwuDari2hV1C7nyn3IHT3enBg6Svo+OGYfN+sTvdHnk5IV
PXCOrzratbYFd+Wi/dMdOP7exkSGhaptJhrRimMJ0EToC1d0IVReCGV8jgva4xBIYCZmp/hxFRpn
Va0kDEl1RNMCQYqR00B2mzGkQ3jQLVyr/WsuP/wHKOhn3iURFOGoV4Tw66oTeYAi9fJvnzHgVf9n
VfzuAlgUz378ppST4W8d59DBpBpSS+OCkaz4WjsI/XpImjpyMAgaJo7qxkxmuDssG3JrDnzTk0L9
VwwfPgQCqmSghK2b51u1hXJG8GfhrAk0MZPWHF3ZsDws7d3Ddoocv2Qu33gO1BJ+wc16P+Dfj5ql
63A+SMm8qgkSQKyCyqG6G3yXGKI5K3APWepKBfBRgtRCxbupN/5UaFvVpCfMInjYa4l7tX2iTULo
JA4cIAx5AnYeTdfoDkXmOTHJSqsT+o8Nkx9sPAdvzH1YNY//+gDFqhS0cZh2ClHmtfHns+sWlpoT
MFxRj+3ZMQNcNSKxMQMtyow+zT3yKW7a5RUBLX2vYjDWc6Z8F9mwB4e5CI9dvvWDIwLvs0iMyzmy
31ZRbOXQXvgd34ovMw74zzx8Zv6a7KiYcaQFT2mNRfRY78O/5pd6mLpI0fJa1bzjGgKK1o+lW2Eo
j3f+oXcSKVL16rOqbBXecaBctL67VrR1Bwvh8KVleCRbdlELfH5OAcaH8tloAS4P78n642XYwpBz
q+Z26eDMTRyt1wxcgb7hd+FdXG6RS9C2j8w9CXiKi//kGziDTaxy1vKg99Y4WUP6t+/Q36NRS4N4
OOZ/a1fUKVD0BKMmX6dfm+QBbNFiYSWsZuNtu07HSSXEj1IFQQGs6Swm4s6EriMa8burBAdbad9f
0bzzaKKREHJviBq96GGjeRdkT26KG7KtX5RuJIUgEx5l5pKWnKlEVHKiONN3DggoLElRlwpqVhQo
dfbhyrSJq8GxxGDyFoAifG7NAkLsqaEhR8R+++w+aR0+gtIcWyUtIIeW+oI4Xu6eOcY5i/f539nk
K4Pfgo+4tHnY1P29952VypREMmOK/9/Y8iupkEy9yra/z9qL0JRMZkyh5x2Lbn8oF14aosWXaNn5
myZyeQFrNKx49+Zo+raElgpAR70TWkC0qxeUuTDwLzilFOYNCAbEgqyd0dHQbYvCLCYjvpkWS3JQ
ZZdLEQRDW271WWE62ndWAZ2p88Nw2M7svsoW38LYS01kogOnpKX3pRP34PoNY7oZ2ibPomL4tcUP
GtFqEAwQblVoJBiKHQzGdxxTWTyuza5rDG6eSNUEJjpZObCrx6dqssUyeu8XYxjXOfJ5uiY+68iv
6+m1mntx+0r6ghPWkkL+CcQPIgRk3mX+6g3Zl06gZXYAo6DHWTxdeF2zF9JGSE9UHC4M4Kr8vm7n
Vuxj7QbIwSibeIAjNoS4GCPQ+ozUiP5tmV5445XV8skoqLnq3J6fkT3riHB1ZgZJYlokiyB/z+KM
ltug+2GJo5vRSV4bTN1gRBaN8TzpVNDwbht925kettB/rWMJNy0HSOU6KMnOG8c0R7UphL6KlIHu
0pz0QUytwZma4ejyDxSBrjxS+xltPSpR5wtB/wVBlTykpRvd4njYy3Qf5J/ivo2c1ifUIn23ll7r
EDQJP/Rio7qaUechfwBGKpqLUtkjpSf6clEsjsjDKQA/dnVcpTIzwuz/YKTzN3vD5ZhLzt1KyI0j
I8lSFFZxsP0CTbl+0I7Bo6ZwSCxyqYd10/6tLgtfJ57k7x5E7h5gzQEMdyF9KBxbruSZL+U+2djf
MYlqg6+tJn5JvAV0F+HYL0h9id95hlVBRC/BWUyMrH5jJX5MEbR584++RpVxat+9FJFCPv06eOFh
e8uZ/EqkroKP6wOfdvnm3qrtFaAA4wdOjSqYEgfYUgm8AqnlAKJUfDCKROJUnQD5gSDmm6yMUpuk
Oha4A0dLaAP5h2AUmdfD6V4T54xjhM95WSAksXy8z/qIIAUBpmqappk9ZxNM5WTUEmDreGaAn3gK
JO9G0l0hE6801pu68cOqQNczTsA+MW9ThDkO+KPo+NTA1hvhCmLTQLN/fuYSRY3jV+haLAMEBO1x
HSGNnaXSOysRuYk7K8xrkVUPc/c5NCuSHHeN6H12u83ubNjzRaxTSrqPaoO9esUoD0rhB3DzsbKi
gV0qWIVJuFI5tePADhcz1cHq2W4er58Rr0QT9mZABxyQVPlHUE2boFL0WVu5udGqePla2GSkoF/R
4mFL3v9ZC9nr4ldZo4e0cN69iTBxCocvtzuQiKst0vy8iVXju9JGU/xg3oGmi50iKo091isjQ+Mi
i5vkurjp1T20zuyIpSm+Pt5D3azyw8C6PjMH0BshR9NSFQPXQEq+dtBMzwkAcUQt21yRQKe7waOE
rnXxuxSQWWAhRpU0rrEfdn/qvsoa35RA/8ZB863859tfuBiMXvOBtSpryjZ4gn0O97rbHz+ot9S2
WaUTs/9inOuPrA7WPFPWLTUSR+g4rG0OGIVVP6P4AHgtCzCWwfOm9XAm6FW4QBA2Aq13f3RItgi3
fRWWOhabA+gvWy8s++fkUZE/jXiCSL+8KBFqPb0lczG4iDaEHi7i3/vF0+1Pbhua5dAxjXLQigv2
7Wj5uYOI0R/OZj5XbKqgpC3/gr6yqYrXKYhOHn498ekm3p9R1wdD6kK1igH43sMeDlexGPXYPajl
ojiLVyCfXdQOIhwYyYIUEjbK3sLYFMAFeSgHs8uRxMYA0trkUiHmg3j4SZ7WeV6b5pS+QRUo1Meh
gCDkJWsknsWoGxFFpQutDVh5iCCDbt6lN8nS8wbcntmEq86hazOHgdlaoU4OfEQYWY7d/3mZzeVB
HWiuX/8DIrcKZWQbok54C8ZIbYjR9wtnxABlGVaGTBPdVowhjRMi3+IRSxLTgBydiBVKxc/79APr
HAt+1Jb4CEvTTxfRBy0ARJC4B6iblgR1e0nhq7mvomt6Oq3PogXwAdYVboOODpLfzZUWUxlSdQMh
+lbtPn+I+Ed8J1GUOSgbXhW+GG8k3fmRg/JCDX3F57YzVcr63uTXvvAPCFIKWtyevCEnMABT7pyX
rCdZXH53dG5NBvWXpDJDpn4GMtqgRRDELNa6SLXEdv4iz5HD2a48YJhGfYXf7/4ccPZEuwxvaFXO
PU+dg/3vcn9LTnJ/h4zN64y2FkzSBB/3wQqL5h+XmUGULRmY4EzGXCIFm2C/all6kO7gNR2nbARg
kY/BCbzQtP6/Ex6Fx4TH1v1vEl6IKCFDlfoEtYOTwKqdzDpHOwx5XTebmDUy8Bp1FKnKuPEABRBZ
JXD75YscX3M5+iUuY5q6RaNd9R9Lr3R87Dny9dU63I61JD+kOW0tJGC3Hi+2qjBPdn4g9lqz7YQA
8ZtarHP2fDZiR3TcTJ4JTGIeMYSTIRRm7lXgJbUzC3MqoUEHKD1KQRPgKoem5qK45BaJmx//aV4R
ruWnF2UlN3HxvacwC3/58hv99ttpyuD5x1iDfyM1w9sBuHLQq7gfz2sQeyh+w7/LGw+RpjNSX3JR
bzOuFBazNPOgbo0MIGrg8nZMCMxPdNbVRLWwMj7NiHOnEMkl0bPaZX/CPtih2IyMxkWWzHKi+ssM
XDra63gU0uItz79rpYKCFw6hgtpH+T/14MKH+tiyxhLoro7bTgdUguzivRcBvOr16XklgETa5qqq
/Ox/J5E51Ea+Dr5PLJVAOG7/y53I3cj9Je/wOE47hTIri+3f1mbICwOh/rCiON+TTQ65nzaU0nmf
w6ErKH9UBYNia6vCwgdS1IJT8qTz6y8y6S93QeHl+POFUeLOA8U6+mtgaohoCOpUP+WvMIJI3vFJ
uuDvZgkpurJ39Z2dXqVUyW7dsQONuYCjq1l5q2iu8RArRj+18VuhCj/YKk2awxW3tPp3KsydbxF/
NgOXkHk1Dy83Abk/1zz7ddI918iD858u1qfWuwrY145Oi/LiFAglpYu8zstALSuBM+SX1/ebwYNz
k48Dbr8UvPaSZc/cUaWWUq75pwqmgmjo8GSk6b16E6EMavEZEq1aueBZuXUBcR6zP55Xb+ETvt5k
z42mdyMsGIogB1H2ki6QSuqlWsabGZBvn+/zDl+7wA+FqxTU19SzY0rsiSKftA1foyXzYp+yoj5y
DS2CWYJy35Lq/irhHdBEB61HRDn/gJx3iFbz0pS8vY5k/IyS9/q+ivPMb/PdPCB1DpfGHINWh1X+
Y1+I2XsNIMyay7k8z7KLuXlXVvu4B+Tz4P9UUQPnwsiucN5Hs03BzdSt/OJ5YBZWYy50p8ay0UVB
r9QlR7dCMNCbODWExmss7cGM1lFO/DkRS8/Hxy/xotS+GwdCXPI6Oe0DLm2XWdxQybsST/5yS51r
s1zjtQiLdc2GbBek3SfjB5r02teKDDVQifNdLsDTgeGBdInshRbxDnPy7+qr87aMsDioBDHPkIss
n9AFUbIUmJgID0i53c3qTKKFyPj+BQPNxoEBnjflpKV6/ASj6VfIdFwZE+0i9mRTpEiOqf1cMNxI
ZpPTogUbRJeCbOae+6Z/bQ28aCB5i81LqfDXHLNXozzn+zqRqdKuTBYG91I1ZphMw6hAgE1b5L8J
jDiGnje3BKAut4/O/7HgRsEredDo6UUNiqlqUSm7icmZlNzzqY/KqYLWb9Swa2QksG/u0jljeJG5
Yfq/QsizjI2JESTCYHAAmdesUN6KlKPoP0L7COUhKE4CDSli7RXvMG1Bdz7mcj/CYZT4o9xzi4d0
u8vk/1S3QlNZXeupoFWUrSmlSEOlMSrVs4L8cDXJsrbmJuaPkE/ZuIh58TYADVfc/a8dJzE8YCZE
mLE5TxtB20oFsUaWOSHyIllVUHmA6ykK2dheMvUrBeuCTXw/xaqPCg3a2G8g2/NrFJ7c/i+/pBS9
vKNpMCFcpiMMcQZbwIhA67IWQnqN/SmaA/3hg3oUlenWc4jeQiSWAYTpe5n/OvbUYOYzvHMO3Yz+
M93ERzvZEvIxU4E138+d7limr8mFXI9Q7o3mw2AFvLSCJYEER3e88AuGaTCtUFb0tbWaMXugCJSV
PZnOccp1HB6ZgSTBLKSEFe8Ezg3pOWBIxkm97L2H7byEQ2x4qwChdqDSeAr4Mf70cH5aBrTaXTzd
w1K+IBgtq8TVu+/ErzqcmPruiOowLBCVABDxtudgC+QmTUMNNtiaPBQjPOyS3z5g2ufvMP6XUIR5
SCof4kdqDhwnmHnWKL9x0du9KnupBLm9JIzMJK/XQ91XWvcB/hVRMS1QYBl/H8kaJhyDw3RqnZ6O
lE67QI94t7cVHO9GaIujrBJgoCtcsep44X4LoHG6n19wdEWwfFGxmnM1FJeWsH0wQ3PkZwd7Rrgv
NGmE4AdtP7MYiWueWbF0A6PWa/BZWkH3aFO9oo5u9nDiuibG+Tq7wm0X8oE/kG8xVFhovdtV/cHj
uDBNCka9BaujxSWrzkHmopPoW8qsP2XXqSE6yZza9LEv7VEZ2pGfoSxgVHxkPjw4TVBuSbcnXHa3
1OPBba+3ZFCoNBKUTLtR0EZnTWUAkNzDL8bgWigFmnX0fSZsZ2MLXEBcx4c6dWXwBhkUUj/N3FdR
V/3qC915MvzvEhY4BF0XJKfpZGgjl3EXubDwmUXULmAdC1tNcC+PRYKfhHsgJVmMzTFuM0+7epu8
siHEyyLdo+jNImwEYx0LIgzGM007SEBs7o2BL+rShdAHOCPoOJchnsAgjKh+NQejKQDclJjrh6Ft
360isJw4mazHLv5mVPQBjE6xWPbVkVTlUN0TjaHspbf5C5okN2fF4KgrNpRHwxci6E8DiGd0cSG1
9tZR+VM69uf3pFFBM9vOF/wftg0qe8UUGMXxG1mOrlFRbJiCwe023R9/d/LlPt/rN1Ozbd0p/e5n
dupHFS2HIcCTbQwz0+1s2BxvAo5s+ozwSOh4m/HNsYFypZoMpDPnRezvnwc8NTSfjnuRb15Hl7ns
RnOLrOBw9BhpB1ljqIR2mx6Idt9xisA4mXsX0Lp7EqGbJlc3rON1QeBlAkREx6y8xYjJG9lmSGap
pR5yZg2H3tH62h5FP01EzcsPyagqjWOs8boCV+ux0Oati2n458kf2ONTMoZA3v1neCMI7mEmKT34
lZLNRpobqRtvQclRlR9wRxKrWCPxFCBzDLhKkqBDDoYW/hk8yLHqJiBNkm1zqa9afsOZE50vWXUu
tl3RlJ2RYK9JftWO1sJgVMMGyXMNJVJKdj5aIHflq10v/xsD7onBkHr5udNvw7gRWTaQX1bffVwo
zis9hmfKQU0yFk3B5umjzzDVlVTiQQSxGtu4xTTUyqTe39Hpk/La8KFq23G77127Qaalj1Q7F1bk
8E5EUFDhNXaDI1RaQ23dIGyGlYFRT6XhJyappE9g4Xzxo7x4opOLaVWtdTY6dWFTe/7Vsp4Qy335
H3QkULWKAWzRDI/gDME02x1uJ9MdcHS/7d3DEZ7SxWqUpmJQF2QcWUayZa9XRZTM7Oi5PB20pJnM
4K/jNR515jgtGuxtmPJvKLHWab/GFvfy9JqN7OXxyKXpdXh810JelVYz0An8sWTapNAU8JMhC2lI
gKuuyQX+01ncaFcljnVnqL+LCdL/ZvhSpxAXKGRNCky6wjw3PPV+s83U1QxohnGVo0hutkhH5J3u
sulAUSmqNo2ztSR8d17VJmWJELl/3XKipWnyc5FsEnr++r16XyPH/YEaxvyOyv0Wp0n6L1UPJprJ
agpGiF4QqnIQWZsib+YHkMDkjfL93QO9BHs/v4n0Zu53gs/KBP/eQ+hqoz9mGJ772upinmR+JeIT
P2wD1oVrXPiMo9t7uGCqp0yRLvoLY7g1zBHC7yaPSf/aCaYgyq4a6FkxytbxJ9EqGxgedLcnIJdg
C3JAPbP2sCp54hQmqJiIJQLrDmhwRyeHQTcAdAfX6fMp0o6Cr/JEXHprKk9f9D0itJuVurjaFEB8
jgU20t25+fqdkaUhmwTWnJ4AtyPqZu6HbqkubxrjyHGvhWsIKsi40sdwsk4qi6Fxhr5FGDoK7Kek
kQyF0dJ1uTwB58Y9dg0AHAhRrSKp28OGQuQ8pcdKYlkoDdekQlhmeZ4xJpCFhv79/p0ewCbs/167
eObmmL3nlvvfrEC7rwgC1wEBiHmKRPX4ZT1nE1bsT1P/WeGM36aPyvd3ru4CQhpHvFzAagFTc3Bo
NfA0WRSlCBO1iO7HUJrH5Ayp5OfCP+w5kZUSjOmEj07eqWasSHYlspVDvpO6aaRF6Qj4SOPNejPR
gn8PKcJujJwoPVmajgmA3AGhc44wcoT9dKqLZvRjx69Ps8aHpZpGMqDCCTPLxyqW5xaX2R1C9geY
ioPxW9W8JnypEMHLpvy0T34Mp6xymFfMR6HxILrALwDXhPnm9ESRHPKEXNswtpEDmLAvI/8b0wR1
cUYv6DrE1sfLhxTiLv0B8UqcNDqkmZEZW0oJ/4TmcYVvYDy3g5IHXwLlUERmWwMmJTssETpI9wXy
t9SodnCLSJEeSpbbX5qbfb2am9d+LdZXSJ2+7N2nwbJd0Pv5bNWOvOkXEL4+H/o3orICwr9h5owr
eIr1xl2mjPlR0g/c7NIm/V8bHE/C1HRsmlz/LXD/yJs887W2ObLHBGZK2HVz9YlL0esfhHUs/xUq
FhAGe/gY7I2T16jbV+CKqWx3vIvzrRFUDo73Q41xoSCm7p9e71IGQAbsLNefU3zT/FjXGvxrXP17
j3+oz789Gmp4z2mYfjWTfxGKWUqYyO/Yg7MqNvVqV/Qqz5rh7Xa0mNYAATv6IoLbZ8YscEe0++7N
pXTw0+66VDh1z64hMqS4i7TcEVo/yJI6EgpjPjGpCMrwf+qkwZHhG7BaZL22Jfuo0fijX4S/K3Be
5GAamFmTkzX8Z6FdbMFG9aAKFTrd64OwaYVvw/njDWPx5u09TcOLs4gmSiF2msh2jmBMku1nAYaX
jfN4hRFlBL4xQ19Bkb5H4myqvQv94lY1lhzEmAmR5YFN0hyIatBEug2QZM+01gOMO00hjBIV+q94
0x0VhQXWNssOCTiaZLUm1WgsUFH19Tzeb7EL1rLOtmvxmsGtjSY9BzXOm1B69CJGEQuSXpP18k2H
WauxVDSL9g2i6hVLxtXjRaHysXVCr1Y7PJ+5sNYCOcExsXVvd45r2UthuytRBCBlD1ygk8ircCps
nRKnGtfnSbr1fBJ+DM42n+f5CG0BZA82B229INIESjB3TULvpHtS/XXbCqrPZaRKiDtX2uaJb6K0
vbTa97xb0e1ccR8YN9MLxqGb+FlBCIZCdf8qcftAbyy8SxHT2iJZLrY2Mv4AXKTsgVhYaXJKDlfD
4IQ5S59GRNY3iiN92myV92g9te1UKfvVylBlJ0LTxFshOgBJzfzuHYdU0kKZYbKmwERjYw9BNlYK
XdkcN1/NLjzipq3nwQiT1K9xqEDlMJy2HQTJQvpwFCDQQyj1vHkg0nGjyhMszt+qZjKoSecUGqLb
c7BlbbAAG8p5c7oCkckwa1Qqfa79QSurW4rebRRD15TOCsnXsKc/fDn6j+2tqLQq+NQka0J2t769
pZ5AXXjCpY8Iqxfw//FXyFxJoSCrixyNxgObYyfh5P+A6+vXZ2nyxrBbEIjEn336Tkwto85OqvTm
9BBGsF4XfPr8ReKhAEffsOBbjyFHFp9d+0Yjyq1/MWwWHHe/LzMcpEs1DNx02ZIa8CM+C79jmnFb
bYwvanB1ewJnI4Qv6H2VkUv+Qayqz+eanSrhm9SbbCPkTO2nZeJ8TQ6SvQJgWASAYrq5J8urKWnU
5hmWMe6UicOvtpjK8JbEtXlRN8C27XI4s+QMk7TSbvr4aeMzT+Ke754C+Un1tBAc1AUEbEUqUR8y
aw2GejvN/3TluR3dE4xxo+6o9kZHiGk4wQlMFsbzpyRjrNyEaQF5L6/07VoxKBMRC4U8hqbj6KEd
LRxvCkLf4rrCPiTNl4IWsSo+zpXnlT9NJyYzDeUQvqzNNWrT/pUdhdh5zTkdwcKnNvyTJpDgFrP8
33XCA+8AhHCJIdrEKbllwIksweYPRzKxEDDb0Wq9DTpbJ61HzUhm98Xlreoj2fTrRswfAIKWIhDB
dKR36aaED9uq8L0GVN7tJEIaPvUDHYkGLmNyHPDDYgaf3bdlk38M3QRuXFU7fE+B2HCzf2cNqVAp
cGcVDvdSSOl/JkWlff3r63X85ZTmjQnJiajSd7y9R1RKY23+Hsg2RU/8VJESRiTNVCjp/1IhdIi8
Rlqwe9uXhnO6Eeg/1Q6D63sDyEFcs5QgG9IPCWUL+W3Ozr+G7kRSPOnNMI3efxlKMXhkppPwtB+T
7tJZ54XMJMuSyUat+II8TqoIjJ8F9+rg79ZlOyhNrMWlEM9HNJt+/pzbz3/cpQqkkVxmX/xnWfFq
28lmM9se+OhP/NswEnDoS2MtCeWndONoxDhdiotS9oJ+WWlLdRXltmoMXlZTPQAHxPlsM3Eq+qsd
G4MG2j/c6bMp7jE6Cu0YfrcktsUItz7z0eLG2ayEIYdmsghjGZ+mR9NuitVALRssHBXAbcydh629
51OgWpewH1T5Z8IbgXlsFZFH86wEW+OvwNqP5N4OjSBUYI2/IZYQbP+FNb5BU7sagB2xnbx+rL+h
hwsyjjOE8UkOrRAquV2kVaA1wlqHwnBYnJ2cvnyq9jh9nRlQ2X5Hw0r6Lrx6TsiWJQsOz7FkC3Ss
R/KULDuwMZF5phCEhk4vvKrWjZpE5HLutX+K0zBa/8rLALAOVbI9Q+ZN1lpiET2cH+wWU2U1UVM9
8XNJiJWzzxGAeotKF8BTfc0dW8ebozUGWAvDJnwINr8FWUJ/0koK4wKOZxKQTN6uVOgfZAimnMKb
QCMqcg6SVRP/4mEaWGnbG3P6QCYxjoZE1UPBObv0Mr5j9RY9Hcx+aEX4iH+eMj79PjeRSMPDwYx/
euvAfaKkRairiZKxMWLLlP9tUq7CxhaAcsq5trYFNhXMI4LwwHkMu5wXD1BiIRMNo+lhuSaMu8oZ
R+zWVMt46MG2NOklWh+xvdLqox0Qm0HSm1p+iO7J66QCVXGa5JYGorNAiImvBomoekwSLEitcOlR
9THJS3ckVi47WHoR0upy0RxXUJnhlGRnyfw1+TGQElniNS0JCLaFQi+5L0YWGmVq5N+Lqgt27SKr
5HjsN18OPTMx+6rpq+npXniOLTekJDOXklXZ891rGNtd8sNn4NSpevS7EnRxOEnMFwbt4xySGBvZ
gWVPNj9aTSiVPOuIvfnl162EiDwRvwxjiKtu4S0ruiMSd7IG4c/0Byjq5E/z+LFX/AEjEJwpXp7q
Wv1UTwQDfCDDoCD8CJv7L9731xEH+Gid28T4nerm1/1wUMUXytxRvD9LU2kiDOZax9SJAzoKW9r+
rZtMjLSvuRHdkKk2oWmyUeEupzwUkE5WSNRafrnrJQivZj+ppn1eOSSymivtzp7mPOaDLucJJL60
0xUkfUGmyAmR/b0CczQhMybcuzYp+R+/+3DXDZr7YvT2ULL/j8LTUjjD0Ac+kmKK2IZQ0O6Yd0Yw
SuktPsmgD9MZK14pyxg1KeNizT2l3XPoc51Y++3vn10WqzeEMRbgO6sC/BQ7NF16y7taKA5Crok+
hZ15c43IQUEx2xBvkApZP3BZ1zconqsu5qreAdXyLbNRjfASkBMyCxhCXDjY9gf5Or2ZbXSmDt6R
zxw3K6WuxheQRsoMHEAOxYrqTuR8Fuo3lNcMcpmV1wAb6VuudzfVHujGhAB3pNlyHLE3uFwtuwrx
Hply92t1ZsvFTXFGcGXM+DpPknWPnxR5bUc3omr7xQyPwD1w5Op8PR2Z6QnWc35M20FQexoFBg5H
28ki4gFCn5RsjgwewBszDFfT2Y0srzJTsIqRXBnltCb25KBQq/bmZ/CGZmCz+DvxwwNfkyBpit8A
5Za6fO7bDlobvaHxylF4AfAhm83lIVuaNXQyUhbjdMm+4MmfvcXfItSn57cfYhqNqSu3aPkGdB36
6DZvfZvaTvXOauu7w5jKIpE2L3PxVNajwKHko9XhMCKlYWm89+S073Q8wQDHSM9fpwSYsOBW0joW
V47wPZvqqamCefCVE2aP8N6IPcbKd/FGWlfU3dDqaY7+4fHOnLjJypTzR8nKhLTpWsfK952ObI7O
D8tPNg6S04XfWghtzxDG2IvVbZuW/GzzWMM+UQxgHiplay3jyck57rkfZXKe0iASXvhBZ2h2m5Ef
cL+WsSsUvtG8u/d6DYZWMUzyPDO3rkUPhDykLRYktR8ZvJ7ZycHQrIeye/zu2iyjIhfh/8SoNboZ
5Ek4ygkDeygVU2iPN6m8ZHIrZ7RclHR6Nxb+EKWbPaEBfcZUKm/PhqrEBxXiBUkGdtovgG6I+twT
mdNI4YYu/cPDjQHzVl/VswwTtAIe+nq0Bwe4qbblRWz9gBLzRRX9C0g+3whQ4VacIus0kp2weE7X
giFsOq9iFHn+txMGTpzVxJBsGwcQWtXzaa5ijh78VlRZae3OhKqWsuyyFOnXKrCYBN8o14jkxpyi
5u4FIMz0jjDL6uu8D2+I9V4PwCfMb93vQfPGjuLSAPtkp3YzC9Frewxm6/EX8WAn22a1YI3BjMkB
Ueycw3nqNGtcJ3aiGA8Rz6vZ8yXaGsZeAp7noJVS/NiW0NwOX0lFKJx1Q1UDgCIbjbfTcV+Xd6gb
LgtXaPTvgnkm+MPmgfO56IiifC3f6nQtISkOKBhFXIdDst6mXbaRGqGWwo5o7bvXjvMfVsLV8QN5
oAx63N+qZauH2P7hSkAXO5gcLdL2xAzTmHgpQNSoMyQDauR9cFzoLokDJf4/Qk8CqObFubHo+xJd
H2/1qnSWBvF9priCB4ctxAd1HXk4ttKyPX5EYQBMmTbSci1Rca370432QkeLU0PqT0nuJLclla9c
34C+IUK1IEekxpmNRmCcMgUAUI5ewPHRdczPMYEoj2fdgPCW7bFEzKTiCUUKAu8xz8SVQ3FwJFWq
wnsD4ldRGXFQXnXAmWGkylR6vODWZS+VgoTmOubOorUOOtu54I7JSqxJvRdr9CnRUsYGYl7lHym3
sy0Ria9EoBrFXxFILZ/KK8zEMlJfOJZROg6Cz16JNfJ8jdTkQ9ObHiKl03aioEnF9JwI3Ph7+xGj
Dr00Q7PrvPksNo3Wz6ZAiADBq0i6S9ZHm1TCL9fFbUfD0DAD6yilro/lhMAVFSEslEz4fiC/KSBF
rjBs0N/e/IoPq1jMvSCxz3QbD7wIhrZ2jx+sNUCBc/HMkCdcrWiBdi83GNmAtezz5o5sUfVugtT4
kYSQCjYPFJA9fdAqh5RxlYdVfygmdIt7BzoJ5gqkTpuQVHYG+qE5bENFFHH2Kkn9RqJmUHUNiQ01
WsQuAqbtrh3HK5iFdGWI8QiWw+eFqie8eNIrCUHHWFWldYjnLAymZAgwxBPMbqr7dTKQ+etMKsin
1AAQZziDqhwOgPG2uB5gxmNpgZgZxfb/Hy1g6/+3jmXiX91oWDUZbp5GJ+aKRu5ArrcY0FrKpZDq
yJ/8yAwqBCYUt6nYTkSR1x4fkk8dVletT6i/c24dnfMCH7MuZUoni5UGj9hOAO3D3ZoPzTtRwyS4
LHxK5K04h6DG8I1MACUEvooaDCYE9/a2MMdhntyTu7lFtMXZEL7x2hzsSLmPTAug1OqoSL1qZHPX
OaZ1Or6ggS76PoK+52lKbKuYkwYA0n0Dlh38Kmln+AKxgf2UAyCgDKvvmbxq/6LixAZeIptxCqdD
3+dtiN94WGXySTR/vftakAZz+LZZpY8yccclKPug6d8ZwDhxCZAF0ZxjIimTToLbDTVeBdxTZMSw
NaLtgWwTafc01prLs44L8eT4p5iBjOwNrYZQHO2iTUFvi/mNcT1P0Y7+yHfA0vRl6/FL8SRrTwE8
tedX+jHIbfQVhfrq7xHT5mdO0+MPCjavYU/KikkFm8ni74J8TqtR8B5NNvgKzFDib1zqNmzcyRcn
atz50CK522noqxcap2donM4VIKuOPh93yR9VNTu+maKRlMpQqm5nVvvm6/u3vlLhJiKPLjsLhs33
qpB5yG3NbyIJVwKDHRxwYGH/pIFpke7rOtLeMjALhOWJS0IDmpVWw/3c9BNDoKb5tLux7HLEP8UG
5e/2GBCcFvNwhbUs9pl2VNGnC+CZGV7pAKWhiOiWRNzCltMkyLyS9UmcpDFkVn6vdIymTG3aOCoo
msbQDwxKqb42Qf4ctUBcKz4+leq0J1SVaYWeF2D4c8lni/AvtreaeCQBqq/JYsBlAsw7goiH0Uy7
RJwLaZAaqAUcEL13D2EKuFkPFC1xczd0xNZyjn3N/tsAG5V1fbpn+XtBjpFmp/6DFWqrg2AUJpyO
q0qtk5OaujAMJ7QfWRQWQGg6UGYj8Ifr0vMTqukSPkw24GmrLAAjcvk17HtL8KntemDVeIMtCd/T
wufIvw3RGdlQtoEayRWnjhVWkssPHgq3U8gZne/gvjKh1ceXoo32U60YTGflz+/KDkF636JluALu
svgyLejVH7eCoOc34r9A22SG9zixgY624IVasRxQPh1hOGJ4JlQQxH//laTt+ZE1tX5CQ7Z3zrFc
IzhzoVPJ/qv439yP3S6dwCx+BaPmJHduErj0YkQ/Rb254PsLiCWw6J3V7hMsMt8AFJKMW/m5Fuf6
VSBfmJDl0pAsHw7y7ikhIINg1cefqBo0/So=
`pragma protect end_protected
