// =============================================================================
// Copyright 2016 Amazon.com, Inc. or its affiliates.
// All Rights Reserved Worldwide.
// Amazon Confidential information
// Restricted NDA Material
// =============================================================================


`include "testlist.vh"
//TODO: TEMP`include "sample_tests.vh"
`include "test_defines.vh"
`include "common_tasks.vh"
`include "cl_tests.vh"
`include "test_ddr_go_test.vh"
