`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
QeeOlAKopChjKMhTXwe84WVf9gmZ/vDB7++O3BjFOIlvezF9HNZHaa2l+V+jrCPlbT6tujlnIp7w
z2XYWVe5lgjPPM8nvMEtVM1kyhJOqlrJsw+9mr21utks0uWT+jkSH63812OX47HoBb87HtSRE/i5
hSiHCai8kf4hVTjJiZn90X+Dq27gDnXJCGWgm7JzUZOh74JDWl10eXFGBuRhL2AQg5k1OyMQ2nX7
hsY85TPvUH1DLjO45tQ6/pxUpE4Wa64fWvzdnX7VPMjvFbmeeG3sn57bQzM1oT0tW3meXymWfvj/
b1ihyWG0gg9ShslAue8UCEjFBvv91wr2v2cB0w==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
G0LbhJuY27jJbZLZNTx0slIYxbiMBbAGKxgi8PypQqJNKqeKTrxOoAqNwsyqWQjetjWdf5Drfo4v
Oq4Zqzt3DfModuPw5wSqmWGcT7H0jQVPy/dzzKSj+D0L8YanURoWiNU4K3qEloAiGggvtB2iAjKW
hBzYS9t2OM4hAN+KiHc=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
VtZhWjwignMv4vlskQhE+Nsnaz5CjYf8wqkb/eIN4QAmCG2MfSTkOvbtxJdbq3r4x86ywdx2P06v
Xxz0k6x64vdrHqceA+4igUKtQ3doqm+FpprACvG7/IOvzA67xYhk0FM8qDw1zTWFa6LwFumY4ulF
cTTSj9SczToZkCK7oZc=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12128)
`pragma protect data_block
yqXLqeyf3qWuyfMtI5RjCk3aGif5lxHFlV1oVkZaQ8eQS4Epozd2l19B6Oa3ZgrGhwKoA8rV4iHd
pdytKCANZhC2PxhL8n1iuNGUt5QiPgtwWCdcDTkkwICOIeX745ad7VTPFKiBe2QijKG/ganBOtwF
BC+bbm7Iy5BLAEplDUCNo32IMh5Et64Vl7LIhHX/rLI2ch12/fAiw4ftGEvJrlCv4A1iefP+c4dl
dSBzIBRwt0ZcgvpUMJs4Pz5iYy05wlLkxl0zFHHZJuPohZWU0cJO64eKRMjW2Tex0P0rM1AO4IoH
8MZXpIKB1edgk8vsfWjDDsk+tvyrCcdz2w2zE2JAL/1WbNT977RhjxGJD+wxP1+4ul//S4DbBJz6
16sdKh5+q3tEq3QDRd9ai0Hkrgthzuo9BwcOPnZWxZ4XhImuteyN6C4WQwGRRZCE0pkltEZS921q
SUQ2x6f5U03AMYu+e0TRhS0Xf7+N/VG/2G+fGA7hsZSCdS5sZAAq/j/5Dka6qZa0jdh0/SzBiQyI
rAdVgilT6JeylZdYk37LkZN7SffXAjc5LQHrjyKn61kyMkrEhJeE+Bri0Hzq82BbXSwbu+IG+8Xm
QOzcMaRufxsS19Zw3qsIkx0pcibYu2GGlPLDi5sAc/T/HlCb792Aq0R7VFmUFv7ZZ0XzU5opJ+SI
am4ZLHv/EAMVHrIoqiCm7G0uKPSIToibydN08LesNfPQ7kpYveLTcziChz0KPPCqhXDhD+WSI/5e
PxG8MFQUOTEkg7xxGLBIAuDMXQsulChie6//8wTIx8RcH0eo2cq1xC744MPZss/L+HYmHJENGavV
7CK0WqHGv0QJtjbRLLQ2aA/Tn42Nu9RRB1JtIYfhLncURpw9eCHGFqnDWON8boLJb9hNCDgE/rCo
A5hXoNoC6OWr676DI53+NsGAeVBvvzOJTLHYi9qRkpG2a+UQ5xFATMGpRrfcQK+SYy+jj9SOoiUU
AdgduE4P0XhxhxQ3tneZ2cioScPtaDXTtspl1V0ZYG1jTtF0MTtNWO8yGlAXE9wvF/Wg46HPqUN9
MFq8ueWzBErjGTGkB/SF87TovscvEMN4WoVBhUnMY094jUsUGjsf5XKij7hqW6y1aFbvUbiSAH+N
BjnjHA07vxRWREytXaA9wmKVdEtamJgytJ3mH2bsQHWplt+hqsFfEJrA1HFibiq72Osh1QXnNi/a
91NCh+kw6aq4ZoTjHsudb/tbVq6+x8ASbNwi1K7GS6iMO7/20whY2X1MglC3q2q8F5hAdu/q5KHW
cYHk91712vXdIRxl8SrimHXESu/VWHn96U3Q4sGY/ME+ONrdXnTtqc8nbd50VXgKEdUjurR/nl20
LHKYH0mCkoAIG+yoo3o1NXtmf8yFOUmjzdrFO3bNl1QUsDW9u5hUIkmqrVqFbB/HXJvWsmHvO55B
w/vBpzTvWCeUGqZH3XJhj4bLVi2WgzzwFyun3drlbaqsG506owHciPb0ehY82G2sBe9LG5L+uRZL
pCtn1sBk/A2JPKdOUcHx/RZW3dllCiHptqklAdAMe1cT4lsYIsERbtOzVrVtesWEOqDOIuf+S9Ls
yyuZ661rGIKCsU9xz8MF/i2DDVvWpg8sMZq3IkgxfriYittXQOb8QU6Vsxd63seN1mphq4jsdHYk
EuW8GyMa4S2hB6ztqtk485bMAfUvgZMeaCEMaOAiHX0MbzdQRGH3Pqf3ZHai+5n9dwHN1y5UQIqU
GbY+SkVUTtg+kh7itAT0N9s8L/siZPkTeEjNEXskAOVQZwHAY5RbTF5CeUt3nb9P0gKjolrevqKh
MOWi6q9U98hfSV8yUY/M6/uTkrZissHPqgQ3vrLVIvIQDhGMfu/RggvMUH78QzRLMfwycErTdmv6
eMsrByFS0hdkjSE2EWIpBAV80KP6OfHXdnzyjeZGDjGNSOBIUSXAxMUp1AFVCvTtSGlMIWa+fhjm
JMrJawIBjnOhDJQFW3bRnbq96MIOPiMXQESR7bE0O9ljElyS0dH3Tr6/uD2YA5q7ya9Pw/tewThB
9cgV+/DVWDkXC/nXXorhH91iGeXeGvTnr02sarjRySlU3dVJCbdhxqGKcH18VUz0EAtW2mMfPDEh
Ij/Uq4QiFG2wqlShoTk1+vqOCsbzSPbOoUoCD0dRZDrLl98l8PI9anC8EOEjZmgtI+HGZWE0uTon
no+wuaGQRJMLe1mDGlcYGZJAgcE89A52yOmyBjVOmtQz4uUf/pU+6dbXKQdeZFf7kak49fxkj9rk
P/UVZtOB5j317DF33d+7L3lm1717gRj/sWstN3IJLwiLyPrYtSoJo6BaWyXoKFmFKSl/YJLfXrdc
XsrXvnq+A/Cg59kRMJygNLh1nuF/D3UpMgZmPPtnY0nbrgorsCsYw3LTmbwcPWnLcbeboOyH82LG
LP69nwDaf70s4CIqvG7BVuFhkW5aInqjos1A9Kqg1DdnuOsI6JAJJwF4zYUgIuTSSgdfiL+ADtKj
GFe+AHFYqgFLDZ1T8VNvCOeGbgZwQm/sE4LfwVTDhyCztVBmtIykj712HvxcxQra594M81T+KVjj
/w0FNjB8Aj3Hlvb1fznPiMc0mrNw7Xfzmm+SrHe9xGhQ8OyQGAqTslEo/ZBGFgW6GiUDwG5gMoa8
XpG63cqbImWIrWmz6RLRe050bgGKHucgfshG0RVASyZ5VtKSVgt7KHbqRtlBJe9Jy9CUEneieYq+
q07T6Q5JB9EKfgReCAGG4OHQNdE/yofTgiD/eAS/c+4G7wAQ558/ucRCaxH4atf1Gzh5jNMxDGjY
4L+xSpKmkhpHBZz/X9w2ifupSVPFz9bWgSAS4vcDwBIRlm4sDKtPNIOb4wH1pQQyiLn87AK8blXk
x3AX42ev4NyhtP7M6XXkUJDk4Zx3r2e47lcsjIapXYpZ5qMWjtEC9lqyjftPzL2L7xmyXNTeZctX
vQqzfGdxAHmCxHYzuJ9yGT3lVe8HoYsQFU8na1Etw5hoJbtbS0TvDCQeHsDdv18m0zhkkFcfzTpS
BofRD/qGKoFpLFODyxfU0FuA8td+SC2TWt7GOeec0wOt2g3c0TFPJevPbKGhfKClzTcU87p6whAY
HWZJChyGGRBvP3MduOy7FMtQFKZO/JeebjPGWjbo1tpfh6olFYsJ+5pkxosT/iYtCdwTGFzoz4vD
yBAc14wRs61Lcb36Xv8N7O8mPEL8eAUCMIvCBq9u0tOCcFfJMFBb6udeUIZCa2P+E+D8AT3WhE3I
Tlc41s61FlyrgkDi2nnwtqqfPblXMA8xayl72XEJhhWlIe0gxxX5/QDmPlbD5r3i6ClsGPD4PfDz
Hu9Y8BXp8tNDLeIK0bi6D74eCkNRL3hvMsUJnB7qJo7+IBDyl+xBgdks1HPkvQNP9/0wwjnxNXxm
ELWfyFyZRaQvz4IPNOWEDNXGdSZgxFO/3Ca76lPq0ycwOb0a8tHcmsEmlL2JI4NY2uSgWYZexpVg
RNEHyLHpIoigRW9joOAXjj4CEBC/9vSb5ZErMcU0iSMSfN9YQDJq8PBCKRnHy1FhfB+AzvcTpkX5
ROh8y32oynxe4gtf7HbdMoY2aguaFviis7XhqCnNE1+0xxpGJoV/14HKhuOCQNHYnC2XJR6R2Xp6
9wytLmIJNFUmq3euOtlZf1llzZhC6+XHyI02qdlWeJbQfcRvzUIzLvtIB1LTNHlnVDvgH2U1niRy
o4DIlvc+TiTGJT+nzjKitbaULPuB3MFgrf0HZI2Zhi9kp078t/yS2N+PwAfYTeXMEwdRVLdOQBOY
IncaeY4sRGUjS2eDYaw6HPPc8eupNrjzOPNsMyGGGuep8ff/qI2whNW3LOlMk+RyO1kN0b2wE1Jp
+2Mh99LY82YMtesDuXnTdCIjzDb24t7wsddjkuzdWC2ICWNUJq3Xob9xx48Y51SVlHnq7FyT68R4
jsyjyuCXvcGgH6uXnqSEqqLNJugBhdvZH85fw56hlXnhzh0LTHUiZmq/yqp/+cHVXr1wdsRsAayS
HBcfd2y+FaPFTq1u908M+JCSLrqxiTA19b2AK/zVxvjNUQwpOt08Q/H4K+RTqtC8vBkYLW3z9VOC
U3CcNL2KjWyEa7m6+NlEFdKejCa70Uj7RBl53tXu5grP/Veh5BP7DP2Q8cC74k5e3Iq6PN6nYOBf
utr06BVlZXVpqfE7/CmgWTo4J+nJiY5GSEWn1hBXhbZCW+WbCFgbUHXhfIahDpj6voyqpY35ka2p
qF4d038BWYtvy4xUWEFvrQ/lW9JoN+XNAE3QDOv3YshJtnhX/WShzm0HtrRL63n4Mf5Kq3IL8m8o
LkCJAq0CKaXYZexGrpJiUbNNdc02QeuGbIRmVC8Ne1LxBpqfpjH+ZAYL+7Lj6OTSGRctCeVEumOv
BSGpg5icecDWzoOXtOjnvqrw/MjeIge7V08aehWhycXs28s/XQaS9+w87f34lbVDUU5X6s1cfIfB
saM2/UVjdfdCMM1CjPQ0DYCNNGOXRyO2JhMxpi3L+ob03OCH+KydHN3WDYutIInl+MzKdgDdPqg4
XRGvil7CPMxDMRTyY0vvSgpKZfI/T67N4M7K6WM4uEW6vInoWBjStJkhQab+Z3hf4wDrH5wGnro6
IYbWYtCJz86xv4JZa/QDR30789feStwhEKd0ztnIDLz6nLYV2TnDyrn2JLcOV1h7JHEPfGnuP7bm
woAaXv908VlbMYVxjSuNKL6TLb45Y+aY1acIDFG6iTtLQtmUBHOycO3TZbozWfdBqZ82bd85/IH+
tF1F7/fgJjGkBduR7KDBG2JXb83t+Fyici2jFemZ3/JLcNQhUzemaNTvmOi7t9R+ZvFi+5l8/sBb
STpYHl48SE8UxcSD5Eslo/0IoHfjHNN8VJhYI0iRxAhIBq56Ogsq6++oqWuqww5mBtDmwVc3jKCh
7wgSDQWzGMGkeP3xEfZxBhRjsU+o8FYfIgkrH9y+k+2nzEXbtbDc3C0nGX1rMSoCQIBk5TtYfwEw
PwcQLzPRpGvfkMR1BPznKkxC8D/GyLI79p4XxFKkyOIrYQTjiJnODP+U2uvnFR5XO/dIXjwAdUsC
SjBBFkzxpaKPpdsmeRVfbaB0wOmlZhOIUrPOSbkx4OAXe/sO7Ru7GXQ7tudP/OUzKokrl33ptgLn
wqOrgnE9C1uf5tGjVE0brmQJf+7kJ39QKM0veYgveLXbMhdOzgvYafBccZqh5l4+PIOpP2tvQBiD
PoncEed2gCF1dlBRXvUh2PC9OdTta6NwZYh6E8CRA9ol9ZJqkphaFDIDrhTVNM9cQ3OKIuxUQUoI
LXyWIuzBhPXCMskKz+wKvi5SqdqcECv2qjn9g9a0cRp42bTcUMPlGD9T37dLnQyu3Q23GIC+1Vny
CyfxEpot7zQwmGwbsWtPE+P3oKasz0I8leP7Mepeo5aRW80tNgilt52FAPKP5CwBdPQ9MmAub8lb
xVKk7Uy+B+G2qc/DVool5XQVZbYkegdZDiVRTbIE0U5tUzhsOM3btKF6gM/hwpeSHF9fw6u12hqz
ddRlUMKgy0ACU7lST3dV0nDGNljSlQQPSPsY14Yee252qGpEpO7c66kRy/wRP2uBC0pRbvx+Jeqe
npcT1kwF2UfTj0uHRMQjMyl8LMion5gZPlF2JyAQQXx7bnfcaJqxQBRKceHYjJXKe54PS8WzDfS2
7sLDBq0+eDdhXex5DB5N6qJWtutVLi1vF+xTF920ok9W24xcXXt24JDEnr7qdltP6s00uQk81c7e
xrY8Nhs6U7wgwpzzDsKH21SlCAoVTaUrt2vnJ0pmbEEdGGIDANI90DCLXTXR5JTF8PkleHapESjM
goAXFFmRM2TENa+p+1ouoVUo3BZn4RwbfkZ1p8hLEBy+bGATVcHll0TTv48cPcVug89qoFB6bTrZ
dUe+b2FP8KJNqz71d1dhC+fjVmvBgSfUk22tcVPAFm2v9hBscoO7AbnkFF2vyFI8hEoS0IAdgl6Q
kgiQf2cJnpY4EwnN5fMedGfjKiQPQQWvsCmUEHNqhk97TCnyQJX1SVrnTSTBEnqtmX4jC9KcjOT0
O50CiT7owjAcm67/FHeb8HPRIUyTb4Y7du8HEcwF8xITqO5UZppq2kOrNPl1AmKEiP/tndbnwRvx
XxnAOseUYpLojTRb3En3jivjBgTDC3uJtjKBf3q6NN/VM0PJNvz/CsZEd44ayKaKEbEcAbRjtqmp
mRR6W/yBmB0b3qm1tlYIgqLGthkb2n5Ixt///b0zGKzWVnKoru6Dl6MY7ceG9GNXmnFl835HOz9p
gxuZi7CL0qkfkS8tJUF13ndLWmTmpZclYhbWcZsrgSyDkd1scRJduPeAHwFxlzvj4zcMZNzCoCLA
ZR6Y0CWKukye9QUnSCNCgF1eh+RUhgrXg3Xg9oNgf2QzLHbn/Z28W7C9PunTutAEis9GmIu1swpg
kqQnbZyPzOrLw+haUn7+JOMk1U2zDGVmsSOIrHeeqA9cbN1h/MZV1867UbXSGSuivpiik49UoaKJ
7heqaY1NODOm5KGS9yX9HjLEei0qY7ByUvmdVU6Bgkrp/ZDhO33T14EjdwuVtrbUrTDJGhSd4QxL
Bg3erjYNo3c65LJa329F6HheH4YkyY9Ok5PfMYKhyChIMQkzOUq+Eaf9jurUWsgpXQi/399/8SUm
WdJTEkXIsLMZVNNWRsYGxOoCjHf2XUwqZVn9RQLwwdDzjX9nPxq4XHFigq80ymck/r4Chm7LD3ez
eiu646Xbg0EOxv68jkjpDW+/pRDjn/tn7/qovNxecc+R8B2oH23XD0Ca53JUnM9MIjU1r5Gir+Cb
fEyp+vxatia17bMbEOuscTEfE+cbTYHCf8K8i0EnsA4eLPfiFiXwZW6m6sAmXczzEGLXRxP0ueqk
tdjd8Jup3WLkKYKDpBN8ZrvdMw0RbNvSnmZQChvEWcRdFO0fhjCzp+HMi2BAzsJ6KiWK03A5TRA7
ZjTooBRQJgI+7aqzeY975b3uzz46rkED9krbnO4xsdu6yLa8iM/d2xlfpB9pJ9JTDcuw9gncQq+4
erQDcXUMJuFo28UACETsQTL0LrSIV+TmcZRvi1KA8DQxRswNualKSNFqsjbzi0cpDsrmcLSeA7vO
+Md2ROL9+vhvyEIl0BCP0ykHPNj3X77KZXR5NQ50Qiik681gK9CadPpJLYNJdQ94VYvJGENKhj4Y
lHuk6/7wvTnBBno2s1IFFpAT/wLXoxvXUwjlm2ThtrD+/06cWGMb7VLF9/gPOLSM+iOEELgkZ2d8
ebJsuSMs3eNZP7Fx8tyeddVt14c70axw7CvQD0Uqe1sAFssCwAJh2fuir8qZIXlgOvvufOZHfLkN
kUS0X1lthxvGnbmgirbZdGDB7+6kDHoSiVJXMpcrZV+zB8RmVYwqek8KoUfcDnY6NRWNNVOZ/WSo
MjRCrzfBRKrAG2qNRBzQJtCsqZesD7NXIuyBbLBi/GofAOhtzpwvLK+g0A8HwaGaUEpvTmKnhaGZ
NYUomlmUT6yoBfhQL0+HRUl/mgBL+KdJm7IXqsRmUn2r/6HH0H7QVuZAgUcJKYlnUb3giA4iz6Vt
FHZHoP5nshA61h3ckfLRGHg8a10hC3d1Rs9SNGScdSQSRz4zGTXaiVKVkV2jgjLiJlum6YsbCwFd
HYkTCrv/MBl6kI70+qB6XUrNqjep8IDZAzodG9m9reQAWC6az/0I6YMlSMCuZ5+mO5kIolKLpXxD
OMJ0AGQaNMV7jzK6FddkpMyNNaOrkVnXdlpWpTchZzCjZ19GxsAZqiejVe4XU3OkgZOQUZ/qkoHR
9i4U8KiQDOSbPwcifEqlXw2u1ujbhlNq61MuYXtpfTBoJq4Au03jtKrzid+fgydxTiY7jisp2Dez
eOsz+TJTIJB/GuzOM/8vdDEpcVTDOYp1iwlrATCUwKgCFsdCzwFlPwu06QJGWMmqVovSfFQoLnYv
DJCaHAiEjhEa+4ME7w2yUoCFKKF8lDZKghPAYCtEnA5e4wQaTwx18d/URvMBa9Q18+2JA0ZVNaAm
JwL4jdNpzWYaJKA07G3vbnTc8RIlgSAkXexVq32mBOFKzWzm7L3Q6LqBxhLUR7fVNDQBc2vTqWoM
aCKyRhBf6P1HZys1m3YmyQS/uolk+2rzb0vNBqLuEHMLUEoM8t3FZdANaLbSh+aUnHRQYWEqwmf3
1GwW5LihH28xDrjuTokQ1dB8P62CtpJdW2VJOPPAHaMCXSH4JKI/ioRxZuEBCTZRxnfYJHzWGReJ
MPSQkiRNpod7+oHoV4jFqEg5v6bOfgvFjAOSvEbLjb4jRMnN/BwxPMpNyhlndaIWIR2EjrjvqXWV
dIauq6YKUHFvH2T3zWIQ0NQG5F2E2WoO37f6Ep2FxGJOj2eLaOpqAQVz6P/UushEJXeaK4hvX9sJ
5u+H2EZtwluFPN/T28hv4jGlTV7RS21vYmSpXD8D+gxYnrBchB3OZ7zwm0mrG8/+plP49bI2nd5X
phP26+imHqWnNAouzBFVmR8eYXqKZX/7Ujx5TE7epYURGH0h5f2M62zDWTUzwN96ccK9RMWDJlW4
lDt91Svo+btt0ALnxrI4lUjSsIcrJIrc6GzRnYvhPIjenb6rvJ7rh6oM/68dqrAOAU0ps7ufr5p8
nBlkfl22lGQRzRgdVETH4vFLWX1YWfbcZzKNgZaW/M3c13YZRxIGW21VX1zamBvVmYy1YiM3oMzM
iAKfu8Dt3g8+I13CO+7ux0nGUnHEvTbalxvYK+yJ+y4376AOWDNAfp04FJ10IOSXY012Rejrt2SZ
0BglWys6bqKQoayGCNfS2pAh5vJM2yW8A6K6Na+U6muH2Nec1LwU3eQJhv53x3oPMCBfA1+Dc0rK
5HJQFRpMVb8f3yJecms+Vlepn5YLid5TzcEvimTDGGk0yRX9n9pta/zPQmco41NPvMs4okrH+LoE
lplN8Irl7O3oKK6JLn6YytKMbC43+BGqltrlnoNxOtuM23xmq266uwco2BH56y9cMJI/444x7gu2
ZANQWNbnO3DomEOPQ8QGA3HNKrCBIySXcA2BgldrtgMSobSDWgXgPBsWW3fnU9SIs667U0CK8cCm
NRY88fgCErb+Mb3hbJFXhl31sPKkOImCQ4uhkDaP/geq7yxY2+YhFvy4E2tVuHPw1isouOJ5wEGp
ctBmyMSG1ntKecA6IfGMcuTFacgPBUV9a4zVQin8mFEQDkphiw78v2XR6XUbqXZTiRVIDVm8vgKD
aBQA1v1KRX1qyfMoXjdS1O5meAexhXcwsyHet1aqdDW99GqmwmrVs0zm5UcRJzxEGfCYDgWNXjD7
RQxtFhMNEUth4P9yXKy0O2BaEI44toxiLAgHKdDhBas8BuGoI9qNLr/sPmfw3ASSTr8C3Jzj6N4j
pgqKusD5maQoLBusaOi+9ygLGKw4k7+NMs57ohMtqethzNAop1eVbySEv/0lC5cHKYMKJxtNIMBo
eiinBWR2MeVozuzgTftrespTUiJtuGEE8VGqriRJ3q0pe0HvVlmQ/6p2wfMztj6PG/kTM73HTnVG
dIF3fAY59SPQN0XFI2PJzu+ZXtcsmch8sqvLaDdvZkVrW3Y9eh3qVnAYXzQGfM8UK2wLENtmmkM3
vJmVorvfd67MmoZMzCL+3Zc3pHyM2PnF0B73ElTpO+vMEtyCDu5JfCWpQVdK2omDQ8hpgN0FpxN/
I9qhP+2p6d7Y6YEd0842viK2/fXYNQbKtFTjgoifgqqcFtBxbF1g2U9tOw8wrrq4spTooI2hytH1
znb4swN8x2KDtZoe+x2aB9UgPsnPYnvYdwuVHk87uPP3zPTzdbU9HNH/Iy7dAlutHmkmh3uLYKIc
+QNlpXbxaInmrMYDoCD3Xw4Dm6E0yKSDcKbc6b4C1MicsEJzYZqBQiS9bkVceIrzqONMysm5rq05
qijvyw75NmXWdaUj2kMBR7XCFBxH3X3hKFrUkYhMXNHS0g9tYCGcQA+giB3yyyzo7kxWpbSmkg39
AhqUAJE/I6V8pWvrf5iW/i+s8bJHfkyCpBNX5+GAbPRTJIO7DBkwaEz519A4VDr66LdPXN1SHqGM
a6wMIIKBRuwijHVaBIAfknAaY5lOXU2QeKurds/vEhpbBYmJqEdg69zJmKv7pZ0qY+Z8f7CA9tNi
5y6QOf8wCPYT58iqv5B+m9VWxg5XgTVYDah302F4F4rIRgrE23VYHVEuXyIaToyXGWcSmJGSeFm5
+/+dJBzYdXPq1FeS7zszBGUvhNErSvFK3euRb1g70G6dvhzDHC8u2bakvhD6tRuHnrbGQhZS5f9Z
jROoCIso8SHsvlCny6TmQR4IM+9avYSFsywBGxqjwZ+vBTfV3OvTywqFVONzXSjSxei+eLsYix/s
GEaXHTOsxojRQqZdWL5YQxMVTK4Z7ONZm0lo44u6miixC9BDbxsD/dRdVRfc+zNmgRA40GktzcYT
5blX9HTeYxGGF1WN+ihBMx5w3FMpdXavF+1IWs+8xZco6IE1+KmSHtNcM69ZW3LyBzCxBgrfOzSH
Zks1YaOPw+k3IUrGZrjV5d50sFCeaEHEQ9R+I9ylHanS2iHakMX8T7bN5b+jzjltKFEcB6ltZpu0
CrhV4Mkjsz0PLavIIxunjTVlzJrKBZbXx2cAIJ61GYjoXdkmYHJkL17sJQN/Dul37Ac0/5FH6i2i
Iw+pjJDkq1oX6/+8JCVGfkscKsOpgG99UCL125h7cjxuNzsfT1mo+7XUx2iVZrxdFe8wVyrPvRlE
k+HqS/cVgTZe2v+R831G/8JWNhZ4leUDEQqOeVhkZKc5SPyoXCdPme52liMVHpl2ati20+yzRAbv
u3wPoFlFfyHBpfW1e4zg6WZasgdnBT/5LPK/kawaUDhS2fnHFzSziftvP8Mlv3xtxRVUmetlxqqT
Qj/6k+FT5fkoQYYfHLotz7iSOE9vlbUUF7yo2e+mk02LZLo5TCW2R58vsAweUfCB1Bnr9OcS98ue
KBscZWu7lxXexHL3GOLQeGaBI8vtFNddS3jZO7qg5ayK4feOe/61dowiF7pGSUe80rLUwbb7//NY
iujc3iL8c9twU6/jR1U0KNImuojv4KAknIvzYZRX4MUxTgKYV4vR0vau39GAxl7LRFOIsAy9DTCU
8D1YD9VkBA12F4F7tSp/DwF/6Tn855QAo4HAcyqj7XvLg5tzyWkOjYZ4DQAX85fThA+7huR2mFHE
g+elcFxkPK1CMGlO/G0K54Z91whRSa8jNdoObwYpGG/Qk7Y1xz/Z5TNEPIdWDLOl0TKTWtnwkS6x
H0WL/Sp5SANVr9SRF6dnkwditQpQh1Rc6ZpyqR5kAQLS3nG25ZB+pmjQFvudb7aguXrqxPmiBbvP
5SzX1nMUPw5iRip8gU/tt4dvjOm2kwmFGLXCB/lS2e5NPAotYqudH1qN7KMYN6f1iibBkzJzT2BV
jmOzAvxdmVBgLC//wJFDhAZPIxStLsXM9TXGcgdPEFrzCJu6GfLxG+4tvm3Zx4egmgorrC3ekJjP
VQ6osUapGOWxQgkbO9Pg/mJf91PM7u93cof2PUiZluk6CqKqcK+yycEYqSWlIlwYbt/HlWuz0mpQ
+cQZiiSC7wMjlSLqVGxx5YtLZRlu515xDra54BgjSJrvGOwJE20YGLGkTKq7yS6Zx2yskTjjTPnd
rHYnsNe3k5w1AOyIx5buBgHjTnGIZfjjae7l3x5Ocdqu4RHI+y+t60VoKxIUDWsa18KeyLMYNXfb
qGVxX5wg1dTw3WBiYyQ5B+b7y0MV+nHkqKl9LI5UE8NR/isOcrQdqQUzFWGaw4wJ5Q+P5R3hHPx5
5wYNG+zfofy1NFJWj3KlxObMegNm3QSNM4EZToBgMcGEeDame5ImiB7kK+urIzKjNVBxMjDTgeHG
d9GwMEjzlMVX4xythry+IlA6j03B4nWcr8TpuTwqdnP9kcXrbduDgXq1Tm4jldXczocbxeD87SKm
3yG7hCyPClWRgbr6x3RxnvnHjhEC+vxFL1pCXmmPjDXxdO1q3OE6HUzS6NotL4VJyTjwIE9Nih4v
08AXnVm0zNH0ujCmNCKn2+ZsfmcCdU27ru6cIH/Y54/R8Q+NbAnR+F0G8ESvhCSPfPzKomnrX+Nx
M2pilz5E8bq54DBUMaNUBacY4VLV+rai+W4szmdUXQFufFuVg1RhzfVxFAYcLfRPHLhO2EaAOUq1
cNLCiBIaA5y6OMJS8h6bDkJ/O6k8m/+P7I+obKoYQwFJBCXK/25kE0gLh27odcJfEUweLJS7AHVq
pdMstCM61f8Kyf+NNwD2dUntHBpkVbgecWRK6VSxDZnxd53UaVKPCyJrcT9dsLrwwE+M90rAF6v6
EzJ+sb4V8F0K3cWMCa9JcRFSNlKjV1TpqvJLoBQwGUHqGZ5Ku4A6u8FZ9yZgtlEGf6QVbSsdU3YI
c17yqoVN5x5c9Pe8KA5fPfKbPTezp4/lt9b5YswpLA38U21e7F623iaz06008WKGIRdBovFiZN4Y
QwiKM3/ftz2pCv/yupCzSKoFyS0K6NgHVs6NbBUTv8VnUCSWxTt5UllvceaidkmAraSxk/q0esgW
3pmbjHuN33jVLdvuSrV9Kx0ISzAM2lBkKBCf/uYctH4xRiDgwC4H1N+sftmk3iJFU4T9JksX/3yD
eZq/NHaHVxpzHzjtxz4Yz/QsoJe4TiDIMUpnmyt6hZcIZ+ag/KQMwqUcuVCr0drc9h1iHdAmb4GS
hk2echFS44DmPolhVcVfCyn8kmVPIYNMaNuNS/0sHfqSrqD/82TiGiO/IFhinAGOS4xrlqvTM1Ko
AAbGD0hRTCFu+0qPLNmSKoqOfq/xzYvauwGgU/lDVcqat6lcOAq9xiJgHcZAQReSFNGsItpaie3F
u+0SU/kGRocd1SLIkSNFjI9k75qZbaNo+nmqkKfMYguc2ykhoPapbNHxpMC8S2Rj2Msz6IHg260a
qPoe9fkCE1eNyenqGbEE+ACkuEpJ8dxBmV4Jgf7HFspFyANAKgjlxuRmNf/uNonaeRzolXqhyN3Y
7BjM1HWI2aKVf0rfZCTH11WyWe+jzGnp09eLKsWaWX9YYJ5mTsQxzPBFYLKb6o3fs+jmUmHFcoky
e26VTqhWQATab2cOg08gShwP6/3sZ55jccWnmqdBWt6TFA9rz8U5214fQooFuzcA/YsHtex8IDhd
kebgdHR3YgOgSZusxywe75tWiLzuygyGlGci8k7it7uk6Ojpqin8mLDyZOTy+yyHfvHbpk5AKUtb
lpQROZ++un+kMO9ShhHO60A8DLTWSoW7hmhENQRh1OTKVrCwaBn1Vv46y5hATJdjQ3l4Ox08OodM
CJ7qAEd+olfDJowbLoW6MaGyEu2pYGdIDKiQ1P2dJ2aYAXZ9kz/dahQGRM29fDQFHcmkvFFQNnav
8KCRwTa0KW38R766C6yLk9pSlBsjkmH5Q+gBDmjb/asg906ndti+JkAMcJPEs3/opI25eTRZrnIi
1uA8EqG6J9reM/dwj6/gvy8PCpbnEnFRlHz2q/N1LTRBjkYodNOJfI5mPFW+Dfz+WhtAj+wCnMn+
wNzEFZkr+x6+vKI6cVRTIMGXpmVF73e1HW2w22ivNjKqvHzD9FDCfo20nagrC26XQEQGAe9O1m0y
DQXnWolVK2FoHr04G039Qb10FIP+hbs5LaSTjbLNLMP7idwecTXt7QPFNSHQpGCWD6538eJVvt19
CYa8GSdWAAlLyVVKxRKVJletsy/SmIj9tzjxi24zLRwats8/yVR4OtJf/tbshHFbHPDCGtuQdK2o
Z4bd4ZQ3CJ4+09km8SiwwBjC1HYfMi7LsTQNn/GXT5YlCl3UUAehdATbffRKnhcjlYvhUD2e1s42
5w4K2O+F9kM4mXoT+UqxmWgUxamXx6sPsorN1n+dqlb1r6GetU2LXYeQvjKiKzUEculdqodQfiSj
nhumTRLz7mcZu53ilngvbVI4MhvH13edO+4kNvUE29Vr7Ygq+ZqfR7pF9KSk96iDllP3oy40lLv7
AKJh5dl0QuaLws4YC+zItk+LcOfvRYOXwm4wuuGn3x4yfahBmor6eGqGXb1pbevsDvPGtsEncLmb
odhavr9h8aBlth/9PgtCbjm83uNoyjKTHH/aHud/0rzS9rcViaqd0FSMEXXFjqsqkeZttuD/Xsfn
0J4ESAKS0Irzm0UlbDSNzVl+MURlmCwEgjnRYDtzcs7PH2Sub26EOmcU6+QyZ/+OfN64VqnldfPW
trOYzxN8HAduwJJFOwkrhYPFGTJxr2ErUwbXlAICDgq0d+Ya6zErEyApTnRJxIj8Nv/6lBCGlU2w
GsdpbIJ0lHTx0pjTZp3EPTJkAb2R3cjip7dIrRzKjcmLYJle+W6+HNMdC/aMXHxftH84lRRC32fp
Ir3aH5GmaMaQUVTYoOTsCAsteqMVfc3sidRQZZIhSOsCCYsdNz03vLrKNsA00rcj/DjMNGl1XSxQ
f8Rby1XYA2sSpCgTJY1XyE3rf8TgvrwRTIAlO12tIpwBElcf6pRmlFqE7LfErIdmYXgUVvooL3Is
kwGHYHfwymPwuAl2G1WBWz1IG08K4lzW03Q2cKNaOUhXSN1HfGm1BsFFJ+lhGlNDXlEuL+aWhOby
W8tC0x/Jbw/dA3z8mWBHPRDMxePDVF0xrNGFIJrfjWPa1X1L2+NMHrXyN1RbLLXMYr/LWAtUuN57
g+PTfjO2xo1NbuqnHBwaORojhwtrypiaIb8x0xHwDq2Vb070kZOLrLw996Sxyq8d47EESmLtq7JL
0gcfSAj5sWx5GGXfe7iZkZIgu9RnTiwT4i2E+qkkMsjlxwDPtciePQqxsZYMpz2lBDSicBUS0AHa
QyOR3OksvM4mHKUpwL2uLM0wiK5iYaRwSGMu3+LmNQo5ltj4/7LY2ace7g1Hzf65oHjw8chJq45Q
lzzGYQex14UXL2+P6C8jhwH0fU3cksuKn5hz/62Mi+yz8xYpGuCEXQWDqgrcgbzTYJ7lzsMMfIm4
QV+WyVIwemqc8g4HDbUOEBlAsNQ9Mip0T3/ET/aJLqIHJXPNMD4zeDU/OhvHioncgkfxDN3XjDa+
mK5oI2vOG7Wb6gVkR1CEu9Yf7fmXjzc5LZbOsAgaYHJpLp4HspAF5v9xgsK7Coy0nynQrIo0Z4ws
Ck+4rg0SwGx1tjkZIIOPNPA4tV5lgOkDw/wb06Jzq1o+hy0i5yj79j2Ujr99D8HAXBVySVqc9y9K
nnSgtmktqNO7cYqw9PIrdVEafJm5V1sV4YeVsr+i+SLz7xVl8k9c1xynoi6Mm3gQjQOwHWNVqHCI
iCImBYT7s6NzPDsy+93ACD6YDA46nF2xb5wNZOy3I3VrwsvBLnfpeS0Eaih/8owR7saBgYDOtT4k
zKrABOQbxTHKPDDHxMBytZcmzVnJ5vHQC4GJbAGC3c+45M32yGrCE3j0KtEUVFy87en3Wq0/rNDk
H1wmqyRx+X/7I4K0yfwkC9EH3ZRpHuP5QYLcTR2JTLkf8BtMEYhp0eGFaTjKX8d154VRJUTh9Cw1
Ac70UZvwDF/0NwoyRn3hbrgToMnwfLRrNcGaQvagctnzxmWnaX0zM/gkmtHXOKmTOTg7TZEfgndI
8drpqr4kY9BMU+gYw34EHMPtCO75pXeWXvkdk/PiS8z6wAaVXo+kuW4pr3CSiXCY034u5YLtomLS
sO6Llf7rRfnWCwpD2vlqtXLLVyEdgCqKHWXzT1n2obIZgtZqyl62GKAIqDYnEOWnMKqnZj8On+VL
8Vf+3EA1Dm+0ZzSKz/Rvi4lFBrsJuRrNU+I8bQwhzVDgqYmMMfCAOZ0iC1LIiDuaVIXPCNGjITij
zkrj962XRZ0fgmXOCJlmO8p4PyjBM5h0nmFfJxymNpU3ZD1n5/0/FGEoBqqPXeLTNNrHmulgVCt5
yD5Pq+pJHRjaZYbPQfWyUsW8WGqkqWOGYQXEyJ+oA/FbyaZ3UdFTpu9h3HI4F+j1Ed+qCZFwiaEt
nTcKTA48xQe16D9n1eEx/itd6P9X0F6/d+ktOyL2JZRnjB0tblJTSwYdSNIoJP8FD7JYi4DG6tUE
MVnPNo8PTUEFuNc6VnH5MGm9z75CiPbLmhRTyaaONajXSB6gKaP+iodd0HQ=
`pragma protect end_protected
