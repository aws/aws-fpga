`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
iNHDlOnenizaCpxWQSO9tB9DSZsNDj3R3jayLLrGiprWulaz7oEkFYWW56QEjHpd61lj4qIzy1uQ
fcXI51WrDEAhrig1l58CIY1gD3KNzfkmDD125FmEutx9V/SXIunCq1kXQQW568jcOj34bCT0T3cs
Y4OoBSXYlLpbxSDXG/eb1guyfH1LfnZB+BAh4pYt8ALG11yAjZIx0UGERG5bZVj3dc6CgOvx52TQ
4JP/2NvRfE2+qnHQtr8a3BGlBgPOU01MDyl6Pw0WP2cnfWsbhpBHevqy6z7r2AIUeZk/7zJuoy2y
1M3IAJ3v4EYwSePl6GZF5O0P/Nwf4VyjZvXHPA==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
heBKvkKhInXCDIydBXWOt2kVdqgovYpsPXVJXE7ZXzKp4FN2x+JIe/tue++d4SX6Gr+OScK/qOVR
yciuh5J7WP++qAFf3SnveV//CAkAzZA7kJZWQSrQeU9EB8R1HoMxrOFPRNxomnhuRoD+DDhEXy6x
iBBfEeXXAH8mbxHG8bM=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
mVO7BAGU8v4rw0Pg5zb89jp1yovtKiCU9TjHTJ6Bqz0gJQbxIZi7fEUos1w4H5Aqg9Frx8qzFMJQ
GO3oLZihROsYOrtJPqxj7gL4NgHZ858UTCZEszwz9uKZPLkKYBD9De0203fnJbX+pXCAhGVwsoEf
iBEmBi1uInxdX2XWrkY=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3376)
`pragma protect data_block
/Q0H1A/S42zqz+kCURTsbPEW4YmVo6BLBkkvuhayrIk0CSk77GCTsPk98cwtSzMlbs8FXkhc0Ktc
NcexoMwQlYZgh3seaZwuJxRYlOTTvRcANmRhTgmy9Q9XL6lXS7NZeUXj5GCOoJl+v0h0NMDGSVrY
9BBjMYOzanM9Q7KX8PJDYNAZnwF7ShtTfK5AOnRzGA687bBC75wsALj30Eh/8+jYjiuiR3gqX7bE
92DuRnstXrqfUP36fIiJElsT0cEfzp6SU3UGAT2OSNOMtkHzQdI7xuSxeehl4pSnaIxO//InR/vl
MSEdEO6U5OMZ3H/F5lEpzaFfIOr/M7yI7HK10uVP1G14onvAXSXbNfKOZ+Ri9aDd+RvYjzUxpu8K
YLhMBObQaf9y+E5NyeIHmIGBfj2B833zodZ//4Is0q2iIdRoF35s4rDVK50R5S3D5F4bvSkZbGck
ZLOk70OnMlRuHeSWpdVMBf6ASMnxyjxyfZmI+jcyrSucTE3l6ci6EZ+WWuTMvrrTdzeTnp0xVGS1
BoiZ0kA4iqs1Lc/2enotyXJBpl3PUEMR5dU+hCYfQ99IzoxX2XdIL+gshv4BF4BAINCDrp8OWl8t
dHkjFuka37OiMzUPJZak7FBg2elW3nB3R6wzQgFxc2HOv+2kOFSdS8cCwPz+lLBp0SNTAB/yqT/t
NUEnz3mTiKepNXIuYcVuc9e8VDI7yGtku5v++DGDQKQVKIwvHAKLognC8WmuIND5tsCYt/j2fd1l
za2BBkZWUz1Io43T04Z43Dq2c90/9i014maznIyuLOzZXiHEQvUUMbdz1zbGL+u9Z6fy3TfYLr2J
nP/ww09odjRS6jG1wo5RcbxfROCxApqR5z5nV9sWq0LgasLqwn1TYn/xtMftIG1xP7XckuhFGwHp
aikkMLPhbkWNa7FMzuRlM4LlkbUJJMnWsPt+o2k6ICoBp3+wV27+Cs6CCn/li64WZ8vVBi2BXX8F
rrmPV6lTtify7JaSscrItYCbIUFXJjmdKO7seJdCmrxUjacYY2d+U8+8BKojDPXKn/MiHrRGZ9Yt
F4k+7mgZFjAzCx/Mcp2S/gWexgiUo1+IN306DYewgIQhkqpzMnwJlC1HPJmNKAy7oOEDzQsmQJkO
34Is/Ah9ldLDp+y1f28O2HpHPWjVSSNzUED6QoD0x1eZlj2JOxvfpTVwX8zKpziyeWOSB4rFf9b4
3UnVKn07imqwtlOXLuno1VKEggk7/JiKLfIpP2QgvN2zMQ0zeQYb1R4i7kD/m/X6GeTq8c3ibNFk
JhNJ+vT70tLbJMbtKPVLIEvjBhZnY1I492Yvw8wX653V061D+x1PLoeUHt3aYDPQYKZTDqKHWtxF
KC6iwYAzq+nWEhkmIovjfxFr5byCFLHTkGvV91L5bBee1SIVDXiaOPJoK/O398OGHokzkwDgiVpT
VYnZW+hjrkYGj8h5OGlrp1KgzBN3/w3lToW37S4GU4jf0iOSVg5TrAppLasrE4YzqGn0X7EqDgwA
C4zsDhqgbNWO5rNv8eeWFInqHa9QkBpt/kdzyWacE8ES7+O7cB0aXEfEeVLVtNIFq30v0WYaIRdS
Sbr8qKK9kyFhQD284qimYXjogHFtjUQsMd0aqzrmwS/7BsTFLnsCaexxYHGSGl02tH8xZsCtoWqe
GLIHp+11fgADtuv16GwPLhrFHWmbHO8WoKP9m96Risv/XGP5us8273cRIcY8nCiVQZBV7jfyARm7
BX2Vw0Or3czNtvel9A7KtMUcAI60r1CH7HP29dQ2sMJHkGEhoIPXQGHgwyHoVTJN1nyuTpALvuFT
bDCrj7GeJncVK/eL1WJUI3wNP9M+5nXx8WgBXfwl9iA5BTIRehZjula9r35VlEGNfc3vow/a+88t
qUgqVvXBT1xWmYtpBHwYiV/3/3w3xRoFGSdaQfLUOrE2SX7Xm5iyywtfCQ5KM+wkz+25VpX5++qy
o/sZwpxz8PlFusX4LdnlMWINg7TNljrBh41hGG2Y6XwIZQAf74gJ8zFtdg7KLYGWWoXNoYWp+0Ey
YEw1YqxjsjA6nModEObFKTIkQ2dEzfcg52OfNN3sIICRxRHkt5XsyGUK+9eKiC19ExoHb3+NSW9U
hTbCJO/9M2UkDRfV7zDxsNvgAzW4cuAs9Urk2zi4lgutFy1mIaCnadSvJ2PIoEJrC/9uG7neWugX
AjKHl1Xe4PN5gpcSErj7KL8/HxSAuE+eD7qi4KmsEfJ824q7Arj1BErRubBUjybolHG7lcwJzaUb
k93eMq+Heyfdr/+mX4lnm56VoXTkhi3hEjaP3yMBOChLzLyZ170FCpbJio6fsYZTrnu1CrvwHSXP
6k1n4hT/08PhJothVEv3U629fj7FYS/wfXsB0lDhVUO2ET85WphPIn9duYPQOnf1B4mQUps2tooS
2O4A9ipkpGchruxC7z9BJAZxYWf6nUJrFQPBThScvSsgDhRONbzHDLzNlPbWFV4R3GvytZrWiYqG
o1h4XD9XCLUWNn53LcfEyv0rArkoOf57Qjzs7J7GAJPunD8UlfDUoFELKZUpYVhOL+8rVhLPfiJu
3V5m6g67eARwxx2N9lku2mKfCQZw1xXvnZDOtmvKBaiUHTjc+bN0jc4YbbMkn4S0yexoI1tW+v6t
7oW4OZltzJ3tsdJch5WJdc3r52LnM9zfeZ+8r5NAV7o0u+iLM+076L/Q56fPnooeFYDwXRVAfSl7
EXP8jU7AhKL30w/wYcrwfqdcDbuJg09qBYEtVLlKwdosNf1ODo2+XDRRk3GAOudaP/LW9JZ/Ou5b
RlhLbCah/4VE82g33VtVIQ7G1SVE3OdGtm9Peaobaq4zLD6TzKb6THuWRqP3m0dV/z5dYxQ27dwe
7TU3hIg3uevel6btf809UMjb2S9DQGj76OGQ2HlXsfjIMWihrwepSKKucHL7MoZaGVXUVgXR8UBl
wCnpA9XqteKga9dYTD45byNNW9F+Z7fqQJzPU2bwoxhX2as8+Wc0Kxr8qrNjolYMUM3jDdtY71vZ
hSzQxP3qxaO5o5/mPyzYkyLmhTom86Bvy0aMGO7gQDg9zN5uWPVWYQwRpjKJyfIV9qNR3NMFmRhl
dRFdo1LRGs5GeT3yRUMz7GRfH+y228+PvOaOQL6zZvqgqG4rzBnnQul+MD1QDXikNcDLE7/FiEv7
RBEmCNaebWFN17S6a+9nhAFwug935Q52OYNDjN11wJMa4mfu0iOKrrgk5/Ae6ZQd2X2EV0TpXr2O
qSsdx0ggmkMKVyDJCVaWlgjhC77f5uynF4n/0GzoDb+puddbiepLxGO1XxdpSoCyovxB1t8+fg2C
MRNVoSx37Z1zWXOXT+tiKGGfhXRCXxGnUNNnedIA72Dzsz/F7Yzyb78CR4YXM+nWjqba8mnvI9OP
LqDNzEPtpN6UZB7kO2txJXdHTRrDMWX8IrLdRMph5ztpvQNmKS+BiPoirkGk5X0++5Q6pFiLdDml
5PyeiXLxKaaCv1Okmav5kwGM56NgfsPxUTR/4hSjK5byBR3j6lEiAdRO7Qn72aqAQi9kdQOV0VH1
V8dPK1aObCTkG7D4Uz+l0uhrMRdUfEH8wZBhbuTcwPzqDEgzZHkn8B9dkpUyyUPd5j4QzG5RioMg
CWhKZ3TGLo2ysIBhWvZJtAkdDas7zAAIOisC0DeZ0rLBZG+i1rsUzvTnkFlJsSdsXn7NWa7zaxNv
dMGfkbHmwe4UPuTO6ncjRgQDMnZP2Z7ls5bnK+f6BFag5A2elSF2kLHedwKVUUIlC0WWMi2MGjQt
x6vhrjs5l4uW9xnCDZUQ3DlDwemXdR/o1udX+ZdqHeBsQR3J7ivqk/4F4RwZ7xCCMi7mLa/FpNNt
gn+kW25nzfk3p8yt2L1Xi0DTc0zjezIF5FUkPefZ4lUc6AKVARv7eyxh7EKU+zQpQts+xho95Dnx
yLsUXTxnpJlI/Ezjx1F8aq0R+5k5OxOCgXFEGht+D7iYbw3D8gYmBtbL7f4sfUauRnjQn7eE5hSd
1/oqcWkrlZiQu0xybsCcoK0cMd+sYInoJZtrKCJT3KKHiGh9nkOSSsKZe542cASb65e6Xq9gAp50
uS5B1+1MU8kNIoBFePfyuh9jaQ5Dhdv7t1rsdwlqPOV37fqIJp7eLdPer4kevflqwuzZb4QeITJO
CcZuUvW8DxlG5AGmWvDXKwGZUfwzdqrWuyfko6IfTMqiPJniUoG84QbdhB/aNbiYAviCBxtxQRkZ
45GS4Q/vqlqNECkxmpU1O8jDWC7wUZWg61SYZs269P8De7Fw374vKetEKwJw9oDby7n0YYBkz9E0
O/6lWqpRCr+waS0cK3rHaIdr9rYSllO1u3GQJD/PcwwLUwB7AhIy76pC0dSwSMfnX4WD4/Z/sJ0A
+quT1UtfNpCShWwwnmMOHWG9LarjO0SOLDYYt834l+ZCyE9qkpg2TgBESXi8r6MxiVMvST5UtBvo
/UFm1qJc7ZYDc+3qgw==
`pragma protect end_protected
