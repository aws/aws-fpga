`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
grLspj1HsKFWJGbdHsAmJug0vNShr/R5naUPPzGadn8uKdtywx5VP4iAz1pi3N/KB4UX7VrtZSB0
pgLNbXpyuVpt2wSAIfNrVkCI8CUOmxHOKQ1zpxdfzb1W+WWyLmCEKPSYZZ2ZjN/G7p3WAtg+CaLe
mrarN5jyRYOmyk3wC09By/0Mcn0ZbodNoHWuUyMdFc+7DzeglmTmwfdgkR83xZ2GFee/vDfi8/ec
/LeQbFYzxf3/XRq75tX2wtGhQB8p28qQsL9NSB1N1USqsjuobds5NCdMew9DVU4+SRc6iplWeqoI
FO/rnSkzZiYbo4APw8IHnRvaWyL6uNgxfgZTZA==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
2U/6nBBjJkRLujHgI0aNxDKfSySQbp7ctyLOp4NohuWl/CF2Bi5nxDF2glrCRrwW/nxIGjE2XxHY
cgayo8DPvpJtMAcA70s9yX4UdVNVl94+RfkFkDOARV8iV5NBNXbKUfI2XHa6qes5pV2IHrLPUd7O
utbmnEHaHq/kV3KxcgI=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
H5dlmy9NAbhW4803PK6Lhm9D64n17HBF2dpF7C3acz7sAnLa8BT8QNaPdmWEa+MT1Zk/BA3WXVO/
Vld1AXlBSxJJoVjjzQ1HDN1DN29ERmP+NbUxsZc7mJOhVGW5vkCyrgpCpNXM7gOqqCaxFgGxuJ54
I7w2g30S16AxQ7vqjaw=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3024)
`pragma protect data_block
hZZx+mVl1DIvj2mqC4fzHIrV/ZLkDg1zyFh6aqt104auY9IySYzZ74fwN8A8sWsKuWawlrQbmHvQ
oaPB98+ADCFZnuBzsunv4Q5FUPmnkNi22W7/7GcUJZH00N2wp18kYE/1OntC3IadPVIFPCP2cHG3
Q5X2QlN7Yu0ZSK5ZUaX53MniuR+VgdP/wHFOOgn1PRXOEqlp+rrIsGjH6h8mhL8fQXEFcm/n+mhS
nAlG3NXrva0KcP8uYMWkgtSuVVE0V3r4ymDjaNuJ2yhTQ+m2htw3h+xJtsvM93o6dB9l6wxIOChZ
bbXWGiPmS+7TAuArdINqRxj47WO5MMM4kJ/idQof6bppWWIuJccEZtg5hk7KF+SBBJfYVvoGBSGI
ZphdvmE8AHNCMSgfS0t9weNuVaM89+dMQ4e9DSxYxeyYgTePnYCGtuqrJqG7nNgRfbxkh0kjNJzv
3FS8omjL12ilyuRfmm8HhPBC0AZWmnW8wwGkogJKg1G/q4P3lqBZ3sYYi/SLgZnJL2m3+r8KXLZN
A8SQt71osA2aQ7Y+ia6c0TLEHUgDqYlGXV4mKIoGPHpVjiuI0Ex/GgPwMadUpbs/liizViMKpNRJ
uEiic+vs5mdQGM1FRqGt7D4lHRY/Q0SXUBxuquxM/17Vbza1KIY5N+tpY9irKx9hcxOkoQwxbpYb
fgRoKZViR+bWjPy1FmoXiNO+koPYN9WiG8tPAnv8PhW4xt3CKS8cqglcPDtXgYatmj7hwDUjzbkF
aR5HTAdSEiLn3aIrwbDGePCOC2AZoQL1o3Xzooxl7q9ioDbdXEie1r1k0cCE47znFT9PWxbNfvwx
0iRKn6pvRi7iVgxLC+7ekQiI1ljFbSCkSuA1JmzdDpfrSBRbX6gaPACLKUtSoHqJwHSAsOvTrG6p
SCz9W5xaJTP40/8E1qB0t2su1yuUd4yjyc/OFmWEf6Dm70UVZPGZVi9x4ALcq/bHCFUvyVrL0qQ/
rIHosybcJ1506Qv5Qk0JcGUBafQ7rhLutDAQJoq1GH8J4jIexyl44l39MZ0E6zrZKpCAfHI3+gFI
PfNaoJT2Ez+xHk4znMpuaBOtI3g9h/tQaC/aJUMCRKyptJ6+YkTAsq3n1NcW+Ya0R0DTCWftCJHm
Qqv0PP/kedKIC38oaIVqB2R+zOv6MJe/VA3Mb5neh9SxHCbbzZhVkOuLCwoiJjlUe25If8AYhm5z
6II9MnggvbPGsTihJ7rpVlTVSZ8XrE4NZ/ofF5K1Q3WqIpg/duQ9PoXRrKT9RmTj1YA+ZbIdWezy
TTZS309XVvQarpBbZwJq9VGcHjW0NTCsakS4unKxHKpCjDNe6ZiyLnxC4KkJmxelcXG0ta1pSFPL
hFEtz0YbP4h4ouOYFgAEJbv8cq2FgnzZsr90UzhjUrjogua5PxPu0CVRtYsRpvgD89jh9tnmRX/h
qlmsxlCqhB/0vOi3osW34iosPsezgGrp68LuM4IL0IDNG8cWK+E+lSU5Xu+SZFCt8uFRHTh34NoN
zvikul7G8qqohyIxWZcymc0upn/brUrneka/qrQEroE+prPrWP0ydlatkB0LDumfBlBf3AsgI341
3qesEz1nH8vjBcS9BxYEFaKjJM3YnKEaUoH+0YJitIl/UUI9zQzdvjVtgVWEf2d/6cPinDy+5cAq
OiUcV3CuPZEOLooUcj0f+/WQZWjgXu2LFhKqecRe+YpIbpQlHlAo2MNjj4ub0xV+Xo+kwLss63M+
XdvBFQ4eHu5Gs9JLkRpTGD+n/XyQS1avTWYIBp4FOfZd7nCzXIuzU43sL/Drq3ja/yndHOEbMW5T
zeasYSLhNcV873e3LnhVwkP2ix5PKVCUWhThXg7D1FnxOadegwpzCO/3rQN8eYyLSeO2qzW/UiMD
40AJLMtIY8SJc99R6liDS5lrZUN2L5qc/jwUYk+GdoHisTBVK4RmD4uLP0XwRDuwjhQQpLITZdAL
IMgEF0ZCHb26dby6700lVMOYac/Ge7xPpq4qwk6/DJnf6GXpJXTtkRfPUbKdon5my6PTM2wwZUjP
Gg6PgEw4aOpuIaeKrZ6wMsdywBvXRI5E0OmZ4FRkCgyCfd+2v9ZJ5UVGCAaDAm5zdw0JXIcwqf3C
F3ADkiqmVwA8/vQdlXMWiAJAJLwWAJxijrgRk2lZ0t9SYENjbR0Ds1AWpHN5FYEYpmpCzTRtZ6q7
8xyqJfzUEnGfjpzTVUdJwI0NtW0f6/Zo5rztECMYlzLD02g/wu9uuO3JC8dH5aBThKg2oyUHNjlj
XfzSehwSVeTVvQChbtn7g8jBuuTAw3xXbtIYNqXHPyfqloEvDcySjoCmp5PiI5ncfvfGMnsWdE7i
rQLN2zgicmqmnScZB0cOLKeUNWTtHR6QgI3WQXzZhq0a4T+5I6E7mp6MHeAKutHja18vm4powcAU
QcdeoDdrzM59mokRvnCQySWVA6Fv7IJbt/09O+zjtzJWlzAtvQEkCh8ZLMkXKn8vB+brokzfNouT
PK2MXcsj+b/8JAqnJX/IgN2I+QJGSrd+hMt/DHSxXEFtqTNSEisnRLeovVJvu1O8aE+Gj0dAwDfk
ktZL/ZMlTyPomWwtcP58K8/qjXzgFf4423EmPeCDabdA/4ODH9vV1e0xGP832i64YNNTR7u4XKSJ
1+jvBiL4QggIRWqRuVfa1o/ID2c3dc+wbDVbrDFAtGLrGK4UxQuxjBiiPyNZOu1IH4crPn+uu5zS
U+zZ+NJ3FdHeEOHtPhCY3AkrJzbu4DCBCFCsUcloG8J1EiYn3SSftNBgwOIa0/yYCldBD0t+RHMf
wfh+1qWIVJW6pKiMocTgy1R0iHxodqwhB28N69e53u1ZPYSQhfrWWdbRojd4PEKsVJbUPOHj8gZG
R6BfH/k6PvsOzTqPG5jczX5KGb8+a1INsSbn3hOn1957x1zQ3aFHxzTy9Vk0IE6HlSvX4oikJR7K
j3yJBWR9jqEDM2v/Y0lAs9Dk9tlxVrC1enpph3gsJxZF/U/7XWkNc10kHddyiaFsh6cRmdGW2fke
ko91ZRo1HvXzpS6p6H+W2Ex2YhWySWDH6aqRAUNwaptMEvklI0vAvpR9RuYK/sM0Kctl5T/SFGfd
9ueWjh3SsF+lZNAnB+Qp2W3CFjBEKbWlTlG+3w9BrCyM0+/nbSYCqwNNgV09yZxIMOxIgLjXUa6W
a3i3xvXtbnFs7VNQoVny+ITClrxTFnLjpdtrF+WevaW9QhGJLcSN+cjsfrcAlDPo4fnPLl3gkPlF
3Iszz2Nlym/BWcRVZLqlOLOcTvqMPYu1Ia7TZYG/o8grOBA3s0VZAD2wfpeuYKEcm2XKrBfIEb7u
qTHCyVXPCTGZxPOzyszXY8Ma+cSD28ix90tp4u9GNOwiTSDhVncyKhX36iCtdOmC3kVRXzQ6yscY
qDsFsFU0ZkT0ZZSP5sro2Vwu3/jtIbVZnMckUUpmBuFwOCEp5dL+5a12RmvXwuZoFG3Xqm7pAAYu
TOxb7XVNeyuOxFBQLEs2p6EtwuK/ptRy26XJSxMxPeQtTF+agTBUNDt+MGXTEa6+DTf9z+9yjGCH
Tuzgp/xo7yjLV+zkMZkx22mVvkTzTu9ciZAF7hi/ZDAC6TfkYKQhUH1c7JRgZf0hJsKIN5nrJzrV
GgUDNHRmNQM9K6Xi3gFGckeC4wI05NSxL0BwaXBIy0LrO7feZpJe18Kynb0dy5g2cmAEaH17DAsS
Ijz6Nl8A+AkmXl813x/8k8lfJnmIC8AHv1XG+MFmYOGcgdE3Q4/xbow9Z3lvwqFDOrgZ5H7TQ+4R
msSqVWYZWak/STZyCTzvoD0njhKTpCKSUX1/Zq7Q9vOCo/HGj8zHT2zHskVEPQYK8r3s13yMPaBC
jmWOncgZnwVjgqCEBq6yxHH2mGr4H5WI2HWpEZUERi741gK/LNRYkMyd0pmiWyzUL3HYwVaVF0EV
1R9IdhO9QdjvWOCbe0dFZ4Ye2jDhWqlltn3vPBIJsGlGJZ2G9nND0UisyBNyCGcj+vGl2w0HeyLC
zYyf
`pragma protect end_protected
