`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
TPE1KBn55h8kuuaFzuPYYFOeDUNY/1yaaDFbiCo12ysiIN8hHrdtvU2iPWrhmboducjCOaHyDC2i
aBv/r/RmKSDOM1geVlBy6X1/QldADdVjH5ClghJT4Dgc+5AblKKZyQQPcvPgLXhsXUnRXUO3NYBp
07ymUHn+bYbOURP9yqUhBjcEbCRYgAXEDxyuei4du4sHW/j+pudLv+sJ/tcycSS5apNcWTNTuqP0
4n4h2yl3P/E7CcOwJFJLxi/SL63SoQ43BQwpDWpUlIqZkM+Hs2P5QY9YshwmmQ/qhedLuFlViAue
oTX4+Qjq144jRzmU18c1KH4AnXmGh+sEl6h+nw==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
J5MD9wCBUn3Zdo4ROHtKiJdf1KxvGmqWy60drqkQ05J9zh6JnyB/imSaPw7e09CBnq9CdrN5VFPD
dYjf6/M1zfQRiFDrVjbK3MLifQ3s2ytcu907afkAydweAjNQojsenUEzd0PTUaWHVe3FF9PCZV1o
RonxShvmLIMHXsoptlQ=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
FErVsr5+cKToLCImywQ4bANZF0ceTP5ALVZZttsUjbx/PFtL93sNc8iTFQRuocnKXtIIkeZFhZPL
DggcvLtuDsR8o2LV+qyCj49NGkQaz21WXzKGxA6WWamQ4/VroRREemmKlcdeWwtf11L2JLRCckiX
EM7wBI5/YC8OfUPJx0s=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2704)
`pragma protect data_block
xnz3BRvRE+3Gv3Y2TMB6zXAKi2Nj7BGYNtc0z7IrrQlvBiSLmCH5qa0i/Y3ElxYUl/5s/Z+kqKxR
H1Jc3za40eu3nhuHxYa7jqu04pOC++NZl8X/RtD3apwKrSDBc2WCEFDt293OVL10pyUsWcKkQx7f
1ydHRyJFleF733znuXmsrbKGIX4mmG/5uV7Ta6je9cgoDPjlU4IGHJSDmWj85Sfb8fzxbGF419iq
J4tu18cg73nmCGKHw+sqhTYolPl4TejMZSnwaKmhJaxcc/nsZOTE8qN79BT6Q2Ct2xrW1lkqN5US
NZNsqpg3PStLJBhyAuH7dne0DBd26QR/pqh19Rxv51eIBip5e9ACXILhMOfJBuX3aHm6DKMXMVro
izxcgctj2Qdt/bdIG5Csh2iHTr9Ygins60RPx03aJ4OxDE5BDX5XSiR/ItKg0qMER9RiQji9Pt2N
XacHDDzEEcHw/o4ifVqYPFWZAneHagWgkIxB1EvXv6b1LcmMBUuiIv8QY+3CLmpSZsLHQHnhDpCA
Gd46eq2q6F0EAVmpsVZMXCC6UYvH8CyvKgxK1YQbI/Iyyn20a8S3FKccU6/AqofZv6A0u6g1sDcH
mS41PizJgM4hosn4S3kGa87SO0gigGAwn6HacOPQDaZiiLsc77aHClB2mviVBY3FwBt3/VYQhfen
qZElwA62fngVjgiuztEIqWe5dKLa6zFMOLW1Z+XZ2yndDb36px9lJy2PUn1foI1wvnAACc2sUZo+
UakQQ4Hsf6BN4gr/Agd/OL1RfhqncQucl/hNuFA0/2t8iWL/sxRP9uM3RoYf7R5QsgAmiG3n1sc2
MeGzoui3mObFfkjN9EEB7sMkUtzotYm/nRe9YMLsxOBa6A24A4mtigjDJzcLsLaazOHmn9sfWWPT
I0p5tMIyv0hmlB03Ea+3dhqcuy6K/Lq2CZrMnQ67Eee/iXICtHhFaJhpLYsnd0Y5BUDJKZmHrTSX
ITEjOdMpX4v6W0Dj++qiUM/Q5sbGly9IYuLLQiKumIA26tGte39RiqoWqyRkQcUxKJC5Llo5q6KX
kpeP+y49EkuYO210t0F1C9cjqrTUEbteUhPBCQEm2p9J0z42sAUQfqR+vK43NKtoozQhWD7wUqm5
042X+6Yz55oCBN9w6lrYQFJ/yZ6DosxUmCCstlWDtIRK1Makzh/EHcl9DLuwNE/Mib9xTnv3fBRH
1sXAlCQrz+IVSWskBoTLly5ycEqU7vHLuKChVB2LVpBv0Uh4kqXnMfFqboJpfHUP6La8R29FCNcx
ysK685OT/IQtdiDyyWiy+/f8g0mUroSpF3hl84AfnJIR3+rBUitbUPoAYK9BoZuSAGI2rrAzUCvL
mAgxJA162PRIyVlDbfJ/h/tpYh2FhzjPY72prFHtW8brQuJVTzAqiEyQJUr43JFxV3SRpKHJ20p9
I0MtgoGwgcG9cBR6BgdN9ZXxZLoIOd9daERTBttenlY1SCQb9ddIHFgWWg64oH4AtayohRdIXTlv
QGjM51DJw225TotcEYLCRo/cfAJz6v4/jSL4WzKOnhtiKu6RjWxHvQyn1V+GL7D0aT61gcjUwhCj
D1STfZn0VPhP3WVI67mzWQq9BMIbU+ycUjZd12QgTfykNvFmububQidLVlQTPm2YYANfAqdYgc7d
31ME32Txi3FpvPWfJ9AA1lEOlsohOMb3GJmQCHbzJSXZstjo8NooCwIRWpD14ngLz1tbvu/HzAXM
SvQjfYyrn1xxK6+GIwKu+b99W7UecNtbMuwRI6Rcfat7iPmG85rCFOs0ztA5BpE1JagPaLcyYBXq
3WDSGcQJyf2Wy6RDRSLxSDZgPeV0oNkDDW5S3dIMm4gqZ1xiYDSJM4VVcExTZlr7bxrOuTwS1dHl
LEvSQUVuxXfBcIiQEdwGrjdCd5N0N2cWvm85QktsVDk02XgrotrgV+8jyJwQPcBkG8Xsq/aJpf89
jOO4ai5jUyXHxoHjrr5ToGJC7mI27ITNC/opbvn9q4xRoUZJaOU5fT19dr8pDig3M2GuBi5Q6Tkf
y3Ct1TBz5MxPBbcssGx0q7lJwjNoAghoGgFQs6Wjknp32a2jKhTbDPvmse/CHbVPYHnOLcvKNtll
pAPn2zV3cuzN0bPY276Bl9uIrH2PyJXD9rBN6KLbQlBjZ5IAv/p43GxMOOFOF4kEDShTlkel6C1n
vL4Ezjtfr/VKm5IJ6n7Rztj3X1EObMLbZjUFQxeMYE8RrJrHXF7xU87TVpRJDrIjyN2O+XgnL/vn
DQ3Ra9nIb0GXFkhAWQzo09LCH/ArqQsYVIDxcfFig7IOEPYSzx+4bhX2j8t5OxGI/47ubcpGqep9
4xhVKOIfnNZjKNaZxx2XD1h0buMQmUTQYzKVWAYLXWxC3y8209lJTUfYvG5LVbosH9/jO2c9n0ab
PqVMZiHmDDThfetedRsiOWfz/gOFv6GQkPIeVZn03Vyut2CAZh87x/V+4WjsUo+oyPjABf2bt9Z2
fLqh0276ohyz1BDq2T8XUi1o9MI7zmUTIxGww43Ayr/86eXeEhPAcf+NkGEGYMvssmS2jzSEj7e7
hixauraBLOnk4g/N6PKJNyu/VL+wuaqvzXOgr9pTQGCcADK21spbRy5WXQNgfX8OW8LDzYO+Euxm
JQOLvJibfyIqbc9JcttK0ida+WUDTpB1UyI5uZdGJ+iZAar5Bwx6mq4ss4qIcpYH7AmZOm08HpW4
QOWy4BQlhFFtWfvGK4a5JqnyPHdFceHitVS2jTCfLfQKDGgJ1cBCY3/HhJ/vhbI35QEvOdJBguW+
dW0O5DUXAQa6MffDf/ICCJMP1HsgcoNmiz91KRMqz7EfGP2KBUUPEAW4p1EMS5YTY9NElIMvzNa2
K++OoxiaBJ4fI5tZR03LUZu3oIZgPBEwXMuA1Yg3dNNdZR91GUqHfm9tuXzLWcpv1ll8/yETDyKZ
JfdPYxnIE3dzwWBy4XIkrqkmw5q7DG9OwhQMkSK4CTOshq7SWLuL4SIl39+2vfiJsTEtBDzgQFLK
HlYuQp0HiU/JQVcw9RgU2Y0p2et7SitxmH8zRzNlQ+oLVMOznueYdXRjOS2qb2BybqO3lJoGWI9+
pVWW7oXby0VD96NxxMCVsyuDt/u7rQ/floBHX4NLXJsSwT/MoZ9K0c3ZP3oai0MGA1xTd83pt18O
tF3MEvzxx4jCchvGosPu+59+JoRWxTxN/4BH+sPRBInuxU69PifEt6Fi8ZgDQg3FVWzWbV+o5zoW
Kz8ZXO0pGFVLzHwxE01/36zXGB2XDxXrdFH7uytYRPSepACf3spZ2VxRyODBTRR1JFQnsnAtAEYz
g3aBpGggfU8WPlK0iUdm9a5Oj9wGjtqO4J3OOquuivYzSGAcbGI3NBH99sFMyzNyGZdk5GT0JW2K
j0/9dRyNJATlfrWA5PA2L7P7q7ihO9rSzLMVj3GMfeERnL7iCijjyN1DY9rLq2OBiHBHWcgRqX6v
gKpwIw7tT80vWhUy9x0dYs16mernVUSi6lv4U0lWpvg1gEG0UWh+uwgAz4xZ8C7NoyR6NiAuH4Lf
dRtSySnmgVjzorEcCZeKjtBnsL3tXn+rEg==
`pragma protect end_protected
