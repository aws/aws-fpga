`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
VXv65mcVVIv2opEk5CvOx09HwABaaTskv9jB83GwtVHdyzq58iWr/a54HwlaZ2qpAI5j30ZwQ8N0
LBlETNg5hLzkFe3+7hPZ6J/5dVhS3zc79xeOQ0UzH1Vaj1/La+ivIltAZBnD3X0DKW7yIYzoJD08
m2FvOVg7/Tmqr3nS7vs97pGpL+HkcMrFq3UaGWtuQnQNaBRTn+rdNVyrRZp1daH3qn2Y+Hs5/prr
lchc/+OR24cWecxSsRqU2bVLb5nC535Eskn8SudvPCCK6ihqFj3PqRVVMTBYOJogSgNJ9GGddQ7b
B3yPMezyKmvy4484W11dYQk5jEU+OK5qvMI9lA==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
xhKBdJupAB65ia99VsW+QUQGtBcHxx483QN9iWmxSffDi0AKndjWb/ckZue7EqYyoGQpNvhF/L4n
GvkErEloVp+wjZgHLT5KAObxR9a+6E9dBUKm0Rq81ImNDBBBJBcGA9eDI2Aw4IWLcTHFuhqhxEKt
i62iur9V4XeozfD4+jA=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
cjaaN8jza6FVGPnq2M5upzWrUypo7o+S6SMbz6VVqzOELFLEg3DVaZ/LZvc+/af5aKQukBsbP593
w8uFZX+3kyF5LvzOZNtT+C7VQsZddyJLP4WXSDXz6kWvdTeSXKiTPgsgWsBwy/7kdz0vpTvRqElV
N2ll5uJ17SP7idxKuFI=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2160)
`pragma protect data_block
u15WK37N0mesQ8f8ZEeI25Plo+IpWGXWYQx16WoZT2omN3Vn+hGhZYVhmMpMmEKl9gRPyFRzIW4Q
PKKu/8Y+hN78E/fTnMsYjZEq03n5L3rst1uoaM7iTBM8eut1HlaSl9SRjzcw8t2tFwgFBk8euUzH
y0CPgrs6f94vzGIZs7quYYW7geXUTU/mcrA/LwG6bIGg7LyG0nEFiIQpmpUJKefELqdyDdS6kpHA
qzF/YDCGGqu2Uxt9p4vsayTbV+bnEC1DmQx7idMwcrU0hS+kbiXwCjV1xeKGc2YGnWCRFc22nM+F
zQ5N99QMMRmtjy9lKpurGnLFFP8G2fiZIAdkRnqzJf3VPa1LdpJNHNU16c4jvM13FB/vE6pFpPZY
kyDrgvbwWYL27ZxKfAx9SsXtvLiURFCpOrkqf1VHIk1VUHi8hs8Qj8RBeV3gfeBylXZB4/I7cUdn
CkQR4Fy3Kvsk5m5+BqE5d7vnwQ13sm4royETVDg3gytiq0r9cVHkVKcxVPUYsRpfvrohZNgeddTV
S8mWBzmt2e+Ye7zFymMgK6QGcxsRKqi/itZlWQkdTSoAmBczMX/dJsX12KiQOk2ERY3NIwIh7KAd
2DNIbqb+fzx+vP7UtdN9Qx05aF3/eyYiDLRnanFgFY6TsH5wE9v3rBLgt5+ZhdpGqH3GW6weJL+a
whqwzpQ/Zn0/cKiAaoty/bWiiEBHlX9pOfbPXRdRzNT14eklFV2WKgi6QJd7vsGIvjcs4JYyBcqd
RmVyRLqBAZhh2mz5AB47r2AmluYAfdCl9cohKk11qYwyjIhsa0iKKmsW8Mn1X/tOSUFOP95iV2m5
YHa4JG8QHshAXZIVhb/9qUIu+dCctZMphZzGJYXBMA8sE7guumZ30Jp/IPauv1C6q15di2CRdgCv
CbgshK3/KVnYtzRbObf56JlTjYJ3nMx5HsS5q/tlpTAxriUJvRUsGP4so9fCQhc6RSKqy3EP4fCT
X5GCDSflIHR0GjZ8efbTpb2BMpWZAhpzWzGQI6sqEHZ3NBSV9VLo6yZ3Wb7nAi5Ccl2oLhSVG7LN
zsFYWsJhURKM1KQVdRvV1mbxYs7szjGNzRgfmc48Vj46sb4Qx5m7pQR8yJolf4OfeyTI8h63q4Fa
V6qK0jkbgNa8GlqGZ/E9AsciDUELil0TzK2o8gYDFwdsmReeftXy3vuajRHhrpjpQlnHdfiQmUWh
x7Chbbz/nOfGaA/Fxmfzle2wo53dxUopiS8DcdmqXGsqfC0Z1WYect/lOW9NLgCIPtkivvFOfcja
U+8RrFWAQcW39aKl1XinWl6Li+SVeychd2aGtBrQiF02vlYqkJVHtSykYUaQgZ/OB2VR1/sCvCXL
Wzuah7fdpkk5usb8HAMxwobnmTDuAzNs5K5IHLtzRd8IW8k8O/jBTZyyGllJLpaJDvfPQlR/IxWh
9LI6pQfiaNdeNXbkBktBqorW8/wgrHkTqeugBcWZK14tWmyJgbFEgf1LGG5b7fCSySR/UNST/Mfn
9RjNawG+I+2ZrmjBJ4iWE8QH6H9LoQaa/SUDYgw6/yML/6EqmJOufHFxbbPnHDqoCLvJ3PrchqEh
WFiiowG/zCOh1WeBQKsnnJdXhSKo9hdbri1wZjIQ+HZo8kwHfunIUWVqAp4Dtq/Q7gErNNg1tk5N
fSZvKLvkQzMnD6LlU4uf+tm1ZcFg+3KYEqnKjB8hyEpXnJES+ireqgHn9cOTnjhh7Q6xqFSN0olq
apDYSchlDXG/Cv2YzPcI+OVhifubf/iAFqFB58OJGAAInpecCgukW3QSbHaf3XjywIio846CsPxN
iXVWWn24WlC2eGF+CV/ADFS85xSn3lIKgtYaprTMMIvKKAyKG74carFCUgXYujaqCGU4y0IoJbdv
pU98oJLFOmEpxH3KNF2BAowj+1GjuRS1pkyB7aXdIQ/eVjaLveOM6ZzJ21TPTISJpjHXqcm85Fsy
NYpQfOtt8Pivsy47IsOoUCMq2hHCZxfpKWj1RkS1k9SYuJXMUVTeSizK8i3duL0QOWBhTH4tp/lt
dbR0JV2KBvfkDm+FvtwCsHkGA/scpdvRGGPOLX+Fa3Wtxe5Z1VS/u8eHgk99ra9PsdtbWdg3ok5r
pkhPNeze2ggZ3NakUYFgDP+7O5tLqi2IKbCORMDELL0K+Thwrh7Zhs1tnfQ3cK+NtTfhBCDI6DCU
dgTQ+9PRTYqXCxjF7L1nO6ifQ721g1ny2uwPj4jQrObwaIk8xjxeDTgCr+pa1l590H48Xfm6G8lZ
m4BFPKO0DESSRa+0WSKT+KC9ol/h+4qm30lx+R3IEV1YERgMFVnOr2E3DqBdrGrOjRs0PkyWxGwB
P0Sx73J6RMEGhNgqguXyElZYMCuaaidcJCzvZSoAUUKHiM5EONA70LE+kfj6twOogYB9GgQ5sdgj
xV2MzQjwFjmm5Z0PJth3KQn0naazEGUTLKYIAZis1QH22PbyrXlx89Iv7wcLqBEdKNimv+XpEUKL
7j0+mwHDJd80FG5xwTSYnZ6vCGA6fC+3QOYfkf2f55ukxi7j7nJYvwfany1mUSKfjpIq3m8kCBuM
PxXRDu9ySdeF0XFQwjI36xKMlQfLOXErCoDDGVrhikotYUAsywyZzBZ+FvArop7ifDxQqkf70AMA
L5UDRTGTky9VKt8dhmy4wsKEmU43q7qmI48tualQWoKuuozQ1rNKE9Pf5AkBe9d6oE1wGL+KtyhU
V/0TVQo7Q7pUUJI7cfrNh5M2KhfGys0a+yiTRWS5LV9uv98HNEpha8eJFeRRSpff/hSFGvy5cHFM
37kYOwFb8ng5oehcsGpsPIY9J+u0PhIzlrfvkVGY1bfI5ekXACYFeLYWwU4zpHvYGebv
`pragma protect end_protected
