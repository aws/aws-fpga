`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
TBcMEV4WB2R/PzPkjFMnyj75TXMcJw8Ta6EiT3+X5fDYA7IXp8WkHPaso5lE4oBRoWDmTBO9/mKz
Wxs7tUjhmECJpdOHkxPglIZfRRuTrsLj0MrPhd3ITnHIHOCFITpzq0m0yrQrMlmYg5WcZNECGxH7
Idpu7OjzRINPsISvGDMy/l93Cvpkoe23QFyPC0GmzZ6Kvi5VQhj9m/9VK+2W68DRrSqeVQrD3EgJ
Hlc7nkGYOuFu7ME/B7I//WxZupY/nNj62CXZ71upfgbSzETlKaMJq1txkARoG6pfEmdq7OXULt/6
58Bl4UhvQ72/lDpX/1wwWX+YJaE0XyO6c5GM+Q==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
jaRdDGwS3Xh7TGEl9gsAgLgsePTiDdgIDMUHUz5W8n09fOpgR8RgHoJJo54+sB8SgDv+8JwGsYuu
xRDk2n0iWKxC8J+FqAGOec1vZacYmX2EzbJohBRopJrD0sUII3tqKO21gqFqNXKIl+C/GjZ+bFxb
1VelRh9NZxpvDAo7w1U=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
BilqDW8rq9x2PXSZYl6AL+AUHhL90/oiYriO8LVPRbUpYHb7Ra/rt83fA4ExV52irfGS9zQO9W5j
7G9g9RDOl0KsFhW4jc3WF7MmG23eOCrcyspmCx7+HeO3WxLD3FxFrYqkQO6flHSKtpH4DLEn+ZOW
BClbVLIMIh6O55PZifw=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11184)
`pragma protect data_block
ARMUSqBGYw5H/hARmBxzvPLlmNOvd0xfKeO0diFjbxUHjuzgtUFSFdPda1jDdI/MOJJChgUfGEMU
EA53IlUrRWXHY3Pn0XPYev5mprBfVotuNg55Pkaon4YJVYDwXKl92NWpFy/gCHtci1AhRkJRsoOS
jDJxIyjLwabYKUgYOm+MN3JNHQ1aOTWuIHvajsYuvxa9abhZWqxAHgaMhWB36/zljQm9FH2/tCM5
3sViMzJfplAKv5kJZ9texews+bW81VzLf7S7v6GmAKgfylD/DGSD1uWbsYWQkCxGJN6PWQ2v1QLo
aMmwQ/snOJNa+VzAa8b6v4jrauwPKPebZ/PV/y4KQ6Z7WEAydBvrt8JiCURfXBR7vE8mcpABiMrY
wk4ZkApshvneM4vg2Pg14TRHZq7fAysCnLrjs6NrQEinCQAs7LNq7TO7n8gd6hGMjUfoAycQPry2
iJHjMjg10CLdfUAJZNkJnmP3TfLLc2at73LB1oC12ZFxz6otzr6uGNkcxA3DdkZdniDKVq990A2N
OWy7joPPVpyRWY0m9JGK2Lewqw5ohEy2nn7BPv/Oe+ZMzOpR/Cw1qMFP5ZqusX7EBc4PzP3Cbv1N
ydb4NARU1HDYBVdoi3N7yAwl6GDR0WqYAoQwqJfiPAwD3XbH8PRmMb8UD7DEFSPBgrKc/vBpXXeM
trttNdvaOENWYag7lVVAd41kH0GvkhE0qbKifsiYSfaL27tFXfj+zF1weqN3MnzTIcUQPf6av+U3
2JrGHprXIuQzacvIR5Gyn2K60dOOycDKhBHYEx6z+TV9HzxNS8CJK8w1d2Su6m+c8ngC+MRCVZHD
2NSDE4b3MWphVwJeAa3BMPbM+e0vzt/U9/qW8Hi1a7H0F7xhYsNf93vXHllCYZi3o5hTDlnc1ny7
6rHOyHocvRF0fjyzHP+OM8j2TsyEBOCthFSuDtjnthyMa/G32VCwqLbvyMp7zUJTm4VtLzGN+s7I
XtdJR+3eHpUc7GS4F7QQapg/V0TnhpKqnP9oosn+NhCpTRbL8aO6Bklzqtf4moL5cif9t/3d8VQp
KWUcOMOLgETSYOtnJMbe0GqQZFFCuFdpVd/s7k8x5lWGhZejTqOLSVZSioETdqfwJkv6ekMcyOhR
wBf4q3J4t4XW+ulBrq+wczPeKHkfFDJxcAEqqYXa1qE7LhnL5gzEvgAHZhFjvLAe7k9Yx/r7HQb2
yCB3oeFheAr2nYHWH3xEcM6nz5c6LhIiLyKuoyc/c6QTRfcC+i9NlIW9rnBU3MsMyRHASsJrmnEN
QOsZ1cAA53+LP4Bbjq2Qc7BMcVqGcFq0KBhpMqGemnnb2KRcNA2ihaDDx0aPTKmq8b1TbaIk/isp
b3uVqo2bPp9wxM/ymYBebpRUCamZqA1Xj5RzVc3JNYyOzYM5jhNAw0aCX3YUcURIS5DxFdeeYPdl
OcUmo8G05i6ZCAQokhYZtK+N12vgnZS2gRIMTsFB28HwIcsdZAvO/gPYgwS1QBVJvcjRC76BtHmB
VrthffpjM+uVpz2Ch08NjUUVVxK95cVdaZfOCn/mKQmgqLQKooat1gKOC0rCPla8nEkgGMzX3KFb
mRXF9mEbSSFM2+b0OufRlNLZiSu76eZ4akBX1xiTMCTifEUAEtZxutnfALjQl/w14QKLwDYU7CCa
Mt6iGSrJUEIShoTd7JOx2YYcVLmIGEXE9encichF5oZxN3ezIPgUTgl/sC4kpwkPaopdTEVc6s6o
pJghkaqSK3UeHnedKVvHrsjAO4ptwUNjd42xW2vNFA0lbihl6NQkd3CNaxhgRCu8JkiVfNlAqn7S
ewAv9jazqtblOdOxtBoL9gIOx1T7GJuQiKK9XJK86jijjLO7yNUQ1O0RdDb3pPMch6h4DIa3TiFR
hJfITDGPU1exMeyYOcfOshK/a5nocrhD3okPJrETLNnCZJaLGc6tgByrT4HIK1rlYIQmGOFyHLdS
k9UcvnvJBub+Pi7rJsLv+YRFlENqg013LsgWyJv6venH/8Itgu8a+RNJNnmMSCcO8CdxXsUYFxQ7
NOWs85v7d3c4JZIbwhbW60QEp3iy/zpiz8imLO8xyDWoNR30wtAlQgxX9KKsYCYnDnjtJR/kfzhJ
gXzlwOj1BpPZ8rG0BGQIS+v2/gaRhRoU4L2lOPECVCys6DrYItOLd6vvxLe/esCHtjZzsSZSmO6u
dnTyxkfYGbCDlkJDx04Ztc9mI7xFRGNdCcpW69i7GbNLoqbZ2xsp18RZDEW2G1iXQWQQqgA/P8BX
2KcOMByCRsFD7AMQcBwpnNw3aesIfiXxQg6uFZElnpuxZSud10ScIKmQGGv1HZKqoC1OjgQ1/j7H
ymsaCtdGl/S7/7ygB3YupJIiz64HX1FnXmIBnYiyVE0C1KeegAREjGTw/VxRBf7KUPP8qK9LZXnx
gFYpPcpRhA8g+sY+7mr4zSdvWQP+Tpcw7RCNTKd8G35k/bL8J0xIMt33tkNpYJZq/7vOgzN//kvf
nPeIrj2ANW/m2iltFXw6x0i/ItRRKrnkOOv0c2sPCl0bZgNPBF5P9ORHiedyUpkboH7uxkPxFadb
MTATB8wGC4G5c6pHl5EJWrh1JQ7RaGweP9qmaR1R6hcP+f340dayI75tNYjPGOPx5o6k98ruTYxp
FVCIc50SCCY9j5Z4b9eZk5lxZcB6ABGZ6tvMexhdjXctAXIvhRJ4yErNcrGZDsqOs4ivbAauPBtN
+VO1M2PEyQTCPZY1UKL7yLNlQxD/nwBOWAa+8iiZurRGwEFGPpGZofA6vfdjLw8ZYHtu8cYwxnJl
T0MurIi3fcBzqizx/ekKTBtteEVA1M0SC0citfuhboQeBYuEJoakVqIeHmGxeJGjiUcVzXx8AG8G
ocgk+MH1CdoXIak998QypsK5vR3BBTIqsDnqBFqDEx2t9tHUKcdH0vpWixGvuwnoPfuwYccqAq2G
WbQhwp6TNf+3+UQ4ZFbCi5KmtVJclwcItZU60fFrKLOc0b5+tUSFl2lVMPw3x5313NmVu7VvJ7eK
j+81mEByeyOLELGdpsxkpmFfxtXTuDHe+meBi8CIUdsszsIHxlvG1g7r4W+8+ZxFfNojsy4le0eH
m7V80hD7SW0BmGMNo//rSUoJkJzJe9OIiT6YDPcsecLhyPA47QhSvW0TjNLlMNPTAyi1+mwyCAdZ
TyCas3G0Oyg4TN16c5jlrg0vJfdCsNmAMZxu0IKJDV4lVubYaUeo3tsF8rVe4pymDc4m6eCcNyoc
kQxkmI1SZIuTz9EtJgnLqVoWACF7caoL+pnEvooap9Y2MRbFTiqgMuREHp9aMymJPJ56ZQhCjZLu
TW/XCjrV3s4w9rIcoh9ymt77ZPCwbkODhh+wdn3Qj+RIvpt0gNHQcpkVnieJV05RWQi8MVC7O4b+
KdOkNR1z+mlkZWPUEesXUaux2JYCnT/tt1Y7oQSxWoZTQjCAfkEaE8gF5JXULvFf+nAAUMo3d+h+
aovmhrFWEGROCX7MK5KAc5h15M/LwnBZTqa7Ht7A9v/UF+keS4mKiEVLYo874N+shL2ESkUpD2hz
EgL6kGcGTyJYnnDSOBy9GiGEADxseahjNxMTCGYYxzLUxRjEE1ws09eNosCuLPYNzSfGQWagSska
h1p44EWAICe9wyBdcVoaGfrFrUZJaHS88b0v7pZ8rDeClm7dcsmPkADGcAvWbxtrpGffI5xDriE/
ucKaowhiIZ4gFzEAhFfqkeJb9Idsg2kVWV4QkJkhUegGL/EAeqFjkPhbR37lr9dLInTn5k5hcvZy
MCB3+ffLFR+RnYRBG+R/m+NI56Tvrrb2LozK2DMHNwm2VRICw2PN0jlO8fK0dpeLwPn+fOv8o3Tq
RyvXHoBTLY9O9Lbg+TEC6MJFh7eUuROuJ+Z1bV40RdRmIlU80lcJwybN2essC1+6v9Dqe3roS558
kd4ddBg0OicaVBVduDlx08CR3/f3xVbAeOCDug+cBY6afucx87TEe3H4tAW3jSLCDUfFvhSKnSIa
0T9SWFc+VV3C4uE4261/pDOvo/r+7yZRB2BJ5/oosUCQhS5HNU4NhdP2PPdZEqrcPLPca6TN+8KF
ffhMKBimuKGMJxdpFJchNBWT78Gi7BmW5h7l+kOJB6fz7x9j7HqYvXZEcDbuBtaHCKde2tjGeCIw
TAQmkasCj1G/53YkME9cJwUtki8lW3chy6TusKLoIUYQsHg67HWqOLFakMOzymA9GVsQDNSy9AsD
C/WDx+6+BqM7KzjuD8wvl9dC5CaCPaASkseTuJBXYUrwiXG5kR3jTj/ftaFZ0S0E9GtvT9BLVnnr
b0UguQTxYA1bMXBWROCtih1aJi6OB7aHHXe3k2dHgHqNPtYAE3CPgUGAaiN15/35eN+lo5VJXVF1
2K3jCeYcD5iZS/PUJH2xFvrRBj113NIjr3gBwyP7T0uDB6DA/VOYQ+ljnJ2kzJoC3F/MItaB42Xm
zG9g+i8DPMp3MRT0NzGT5qDf1b/LtAJ86OqoLShgogtq0pw1sNhhFwozUfehkmLiwiNEMPDq2ZjY
ZsR+na4yMT9FkJqMsPM7/KjB+L5YKQqFWhTh/cepvpIcbhyKeGuYP7QVWc0IctBOTdNsshwVl+cv
uI6eAbR60d9REJOm0Si1E/hVWlk6mpWjNdl3FteFbgUUHzMrgzxV7p37j3MGDfHFis408OgOZMdp
/DOqYbqrnoAacxf8i7WcTRSal57l3wiDJr4PyGGjGZGNvNgxTYjrEuBkxLQ27lj2cQOgjh6iC6fl
lCkMK4umHxDHCeA1N+HV1LTHr1MZS+IEdLuSx9QmQZZigiw3jQqztVxRG44i5Afs+8WuE1ejztrK
k3yAeqiNQE5Nu2Cfx5szyQBWIBlAWtjB4Ibl94qPkOQTvnr+3QYf4a3SbQpq/1tYZrPGv68iCJXF
AMtsJ6bAg+y4U4cDsGcQ2MqKKo863bKxQvHjKkf+EVCX1+RFfChIC32hkaFJGwy4KvC9+ULG+jsn
VvUSyFho7G+r6QXQ8MDdWb6R7dGK5f/gRCNtcuoW6X5hwoSV4tsTPBYC3iQFMX4lDq1SkZIfwzJk
cOXb99vAF0j3SeFhVl0fj8dwODIb99G6AL3XYYY1JtUREfcPRPzI+i814nnKDU3K3SX0zANBwe6p
BRnw180c5e6memaMhIj/hL8mtBu8v2H2aEi2alGM42IdFL+fVUN0DqLB2p7zT6cLNPOe7zac5hLL
NgIeMlH6LBvBFaJkU+G4AvEHVMARA5pIGSYg/i29guBrP1m8y6nQsTkcouf5BhGRjlFULrhtc+4x
Fa7caZydpJKm0Yj2gBGhqiMJKKQIeorZh1kgU+cvMd5zDpSGCnLVJxyaaEqB8D6rFHetLEFN5ZoI
pQ7AQQ1N07OrdBs0RwDx2y/8CXehTQkzRT5HZYox504N7O72Jq/vvvcuXJfe4bP2jf89mKMn8uNN
g9RamZZgA6DghHInCa0LrmaCfBoDQZhr552yBl0sYYtRd9pDOocDuYbTOqOpsvDSHdoiSvBDfsln
vhx6SjBClWpZUE/QwSjL+y0DZGYedr0vl6jP6VQaT+uUE9iOXsbEBxJdWWbsNJOEGjorWSXprGFW
4R09uVwJiCyfKhFIraB0zGBh3c6/7WvL6dEdG5Wt9eNDu8C3t6T/ZYmkxoBvJVjl2/EfL1D8xW7M
ymTjzJ4H+ZYqclL3BelAmdiycL7K2BT8C7Q+5ItruY6T/6YcSyg7qb1L4P/lp4gXRT6nETH3VnAA
UBPDo3Hr7Y7SvxURfQ11gOkpIwhsNRbm8kM23CLfeY3NEjMM9hZ+cUfTfaHE/EjSgxI16UiPrHu+
cpBUU2coIZ+h+TEsWPdDPHd8IoYBY/ZL1mtvt37CnFawE43LzVPS05ZNZe6IjqSFS9oYdBlt2vs+
sKbrn/KrLvBobH8pYpjL/iyE+q08OmnotAseFFM1iePxzBeZnfd4g9tV5EzEj2TKfHEkQ8kPfACh
QXGzHjvGpdAa9eliFwktDTHeF/tEaHlJ0nk4FWQxSNYDNhli9ZQPXiu8ZWThAMCqEtaUz86Lvp83
05DgkSv4pXPkuDWxhp7rHnlSyxI8QNKKQuGhSGzVuB2QXN2jmZUSNhs6ltjA/t/ZiQ3Yq+KrFpl6
+lXR5dFz5uSU0q/0uQAzgIoiB9coNvj9HCnosNaE35lOlw23pQMz1KDmNnSaJnF9AuesWtsVnn1L
w5q3pm1QA5Wmi8w1QhJVYcnn42TDqQHrUfXD0ewO495NDpEmV6oPb59nBiJiiJxunpIvvHL4ioDQ
TCUv4hHt1Kpi7fhuze4toZJuNd3WP94d25bUb1PctMqHPqfffzNmJAuTevtCQL1nVDKts0Lnvaez
dnfjoFEy+eW+FC6UY1+SGf01Qmu0LmAPSUhLsmEUyoz6nT0mKK48powxlu1dYVXKYQZOfDoQ1bXG
xtrB+O39gYqfB5SvKTKlhhtGu3bxF6CyE6U7e5XD9AQara0/biyafUb0zMGb7thDXUrwoY4/mAzO
5kajSMPnJy6zIJ/vnifQoXUxY58o7ohjDzZytXoijMt8231jGVVDkUOjtPp7OUO25ajS+usJ9B4N
1GNKwRpyMIfKEetV4wXwFJONhO2EMDMjXmVxEAZ3Leg97h0Z7IxswziWSJ4CcyPgOtf/evpRXpiN
WtvoKbrbMT58vgIH7Av4SBhoHtz8+cMhBmHd5/TRjWRfCnKmwit7VfidT4YSd42dfuvMV8UNfTAs
QyOl9PROhlXWC9xWzZRDWYUOVUwLXLH5FhC61hL7ML4bbMnj5r/oLHqusFT9liqwLJFY1PZfq60P
wQUXc7GW92wGaD+bNMml0+oGxlwls4VFC3igtekO07PB9CO4kuEqHKR9MmP7niD3WuSiiYLkAZvh
Pke6Oid1OFZpK+xpgw0PciN5OnRxEV/TM/uIXUvo5/Mv3QNlAvoYFbnAJPJRLCLXXZp7ZPO6NgPS
kuDa7BmE82k3ck8T5Pa5KNtyjgrg7G/C9sBdsNc2mmEj65xDM7qfCtBkqgGDdUYAxqNw5SvGIbB2
kzR5dMU53dGxXRQ86VZKoWZBU4E7ecISjVRjNJt3Hp/Mwl87Z7oYyhjIl/jYsESmwtqKzXegJqCk
IyzY5kBxpDQ6xsf/Vxc0LQp6brXQ4iUfcHINYltr30dx3KSPCG+tEUaRArC40mMqY3UwZBZaga7l
rL9TrTiL2JULB1z590bPtgV1hdwUt5x0mA39wCaG8g7V+geO9AYErFBydefNjslXNn4SZeSG1gx4
VnN7Y4K1wq31GyYI35QNQnFluw8blizTLYiEUgFZhRiC6AsX9YfY1MwUZ2nne4bGwkk/KX/l/7Vh
HXHuw7NFQ9hjiMTe0diZMTxkZWuNq8URJSmc6JaFJucOhJWi6a8gS2jJFcjKJF75G+fJ8yzfsYf4
D2i6bt4UGFcNFFvLxcZJPst3NUxicf9pDm46H9OZ8aXxxEmiNtD4xRb4kAMAdX9w38Ijo7kNwich
Byr30fhhOgIc4VoVqu7dcfRfbI0XxqjYo/M8jbLbnH6KEUl/edcsq6kKpdDH8M9WyaZ4WXovpfGj
GEyexT8Jd9wEZ2RJEM+GUvw4Cfw8lPR8mFKJbudqJs/4jK7xqIZ0XIjIM/xUQ06Vidj5/cB2zdSE
nDreHoDkqgnDicD+Ns7bkbiZMAvyywIXuhU8JiNiDW8DN51qbeqqDPMYIV6eUh7Vfyqm52aXeJVF
M5y+bUnM9X+O2rl2YjWfCIgPJKfSg4Bp7U7egY6rOElhR98lulpUZ0yVHlI8JZQHyuoJ3aXYQfzO
aasReJTA+FOrT+ES1P+z3RtmFxDz9bi14Rv2AtjvRj8zesUOAAdHwCNXJxguZ8nNwjrAVEX33Ayu
Z0f9OXXtn+ulzZIAN4jwnbVucNvgpVjewPmXZT3e6xlHHgGy7jY1LplpYkPHPPUv9QhIEY96+JSF
3Gx70VTa0wY48a4ymmXx9ql0vSzzoqj7hwPBaYas6mXWob7QYJsHbOLe7kIXq/T3sk9natB5MBye
VqlzDwQ6hWS26iL0LCYbYK+lFbvGVL5Qg8w5ygan2VyitefmkikhVly0fAzgK0xUrKXiFTTJNyxI
uSYUvkGL0GT/IiCtfJGJwe4RIrBilh4Lu75ksjLuCRnpV3fNqT9mdZStFvmR4m+UmHnBzwTLwwCF
iIqow3CbHUmFBs8I2kiKFQaijEAdcp9SrdVlU7HbkPY3QJK4vClvCkHuv20zDl+ynOqeGBCIqg7I
cntqtPdGLGVDbLjmRCypbXK4943Qx+D5taf2Lai6ggbgsL5H7qCetQndfhYxh4bgddlbw0irqabN
2PhZAEi1/ZIcBoY4+eWmJ05BwZeMlJYAST8PJXDQkz/HJTp4O0WmnAWaXH/2bvlf1qiRsd0bjUR4
/64/PO7YUn5+yDdI65UesWASalK5XqMfrYJSUoUtO1PnJyjrOKIqgTNiLC+QgnP/If4rl8Jqx3ZV
6Nboq9vGgkZ8F9aEqo6sPtiJDbIbnFruLCHPCj1/BduqSPGLekhZnEAbM80PtX1kTNFzWwmV7DNV
hzdp3nfQX+0M1yXLWBMqUPWcmNmi9OSfY89lqHyjvHbrf1Prc+fvP6e6iQjU2RGMEH2JklYP9AFX
gNSBzClebxMsujKTrr96ZVPviGLXquGKDQ4zQaCVBq2uVYCeBMdr6j7jPw5Jk1ul2HaRj62KgAr9
DGFNWe4R/ngqOUKXigV6Whdf/WWm0jMGhaYCSrVdpOZgDlphZuHnThoo4u2ibL9ugGrUkzYe8hOM
0DedFl50d+7Oqa3L9OS3eKFFYz4sroJFW+o7SakYnTuw4UjCnxfv6riU394jd70evw154HRi8cX9
DyOUvbHpWMKkqx8yLj2QCXP4jj7wexnwpCccMim/KnKvVj9rpNYrsI8behIbZEE6750UKlyvv0Xh
4bEFCO9SNk2aDqdO05WAptgX1BcKbhY9YSySqQw73c2D8nYkh5XfwfC8LlpCJRdz2UIu5DRFyYIu
hX6NgiCgPoS1XQ9LZoPEtHkObqQwx3MtF36JVxWLfBzqjJrogbJ+zR5l3TZE1t7dSsMDj4Y/f0h0
e/6SEYJ1NQAcOjtGpp533L0UvY5mepoJb4s5uBCitZHSZDK5UwgpnBTk6u775Q1z64/BiXkwaE+R
jTln+54/uojg6/o7EcmccXTyYhmaXVNjTFXrJ8QFngW310xLPfB8y+nIG6eOWpGV0SgRXdtN+fkn
VMFH4oW276afNzq/WxQ24ojWfh3wqG3iY0Cb1KQWtrF96V0zKyUfGuiqJAUCQAtAuS0/QjmY1jBs
RJxBYSl6/lS2Ukh+ACzrOGxP/sjgbOUMdp4m8JiQRc+dfCdwjgUVmCBo1LnfJlpMQfZnbIOMSMAo
rtCfFphJLO5OGHSVm6V5ebVNO66cRW4+W+rRU7t7BV6O5KdTzNGRLxyBNMNORlk64ZUOnD2vbfAE
FlsqSbJ5ZuknnDk5a1odoxKzd/KjWaa8w/npKsxGD1mrFfadI6ZsMLPmKQjZcA5SpfDuDz8NcOqO
IIq4ahVEwrnDSoVXNGwRI9xCgsmseKQYTOU2y7tGtoPDNqcPsYrOFj3fkFHWmvTBSgSnqQGZHVEc
YKg1PbnWcU420jEE2ICQkZxUnmf+FpW9XEn7kZNny2kmGU/MoVzF5/6CjgfpNKpxXUFbIgPJz48S
Jx+5os44HxLVWnvf2a45yIlDHx4ekOKkTTxJeXnOdEvBq4VqIgtNhYQFOugneh/ul3B/9ecdMp1u
fQYJkDt4EPwgtFMBsdfP+6nwZHyDh1ePjP7+gWfyaHVEpxzubirD2z6Vy7avyCCJQ9vor1qpNkko
9t86PqYj7cjnY+EIZ7IM0XVJP3aiuqjY/M5ogCpzU0FnQhJIbJhsAxPj3Nz+a+izotWfuT2tm8fu
ZrrFoLYH3YcXKY5SEmZ1XBobw4ZPARZG9KqShtulhwqLh8NCOuoBfWMiubhEpm5SYy9FIcEYEZuo
uXx3E614fDsO8E+cC4OQtnbLpMDPv8WlqsKmkaGMiFMSkPXkct1KcPOzkfoWNTum+pV2/UsrabgK
GK5JEy1L3Nr9fY8WKvOI8bpYoRWbKnaxiBoTos3qfws6+lNN1xNJACVkGPbhCscrgWhGE/yoaQ1L
/fUKOGs+z9uPYBLjnZgn2VSo/vTRzelQg9BOAjdLxx68HuEN1XMDsZ85wevsYIU72KksvQUG2Gge
H7i9LgLYSEWdNLhH9DR6dnI9aKQYDx1jLTU3KGSjnkKN/eCFuuvKS1wTJPf/9flutuArfms9X/CV
V1+laGkNN1wXdmokW7lqobtrZFZA6YcRXqSBqNP4ijQJkzWjXHpJ2e4oBxP5qRMK6PcKsQ5PVu4a
hX6/xiwnKWUnx+xXXod2EqOhlvu9Kg7whMPS2K1TjFGg46l1b4drTaRJWQGsivxCLEvJ7xr4MPtl
jb38U0gl0jNnD/kQ7gh+iawHQVbMnORj2HwsexUB82x4x2AdOhQ57fgukcjBs9nCR4oAsIqDK49j
yErl6A7DrbktD31CJbcdhxuCDTvbSKCrFA/OufJmvD2HZWWCGHl8icrLrhIsVtFKOvANX2fvl8Za
0MD/qiz85dHMaYth0+1lsQi/cONhf9W4lJGxRDZwBQcy8YfsxJGTwQaMqJzCbmh1DuI+nfId7kbE
B/3S3wiD30NcMxGtKwuPi785bZZvhOlfnl7k3gmykv27IAWy0ZBlMVB9udJsI8prXXMpB+DqAjhj
KK09SXG5AWbORlawJb2/w5QAGaawV+Azk5NICZ0DOnarNBuWDSRjcH9Zt4RcHpK3BDSHL4Z+3lGT
IdLt9rtQRavZnZQyscD04qMfgImlB5VjyUOQ11vkhbH12mVKI9OhPcC6sLO8YZOum17jvonqHomi
qf47E4qPtLxukslMLw+DKoYFLyraTQP/vT68n7z9jOZHAGH6hU6tiRyQ8i55FtP0aSYz3EiJGp/1
CLke2pcvWmE5i0voGKmNt+czmNjCYf7q+7eMedKQLY36FmGsfqVLd9JUXA3NthxoC0twQ/CK5Hf2
bvy5xLkin54AAFWvWxaONXpqD5SIpgjVHGprx2VawDLCw9HLw8D62f33v8v61GYa/ScLGghx5eiQ
krczceHzhZKkn52ax5PVNvT0Sy2SRpeTmRysEwLI1KN68s/6wkAIJNPfaxiFTBLcDcXCOW2hr37R
BXO3gdwZPwlj5HqXckusSp4dpbUEx4yXlE76T5ps1CMezpS3kVe6btF4H3ssDeeEu8JsCH+N4P0t
ln/fZc5OD/skV18dqZSXQSqQPh8Vtk99EA74FsdlfrTeSq3khIpLxPVn/INtGS2CyOA566m3q90X
AH5SjYDDM7BK6LlIvlDn+wTMXPSIVmPtd2zIvD+nQhpQD3NV3VP7YlkSHlkyNBIIUu+Q6Sql6egk
lkNjr9OurHKs/dHJhJgipQoGc1LDrHieP5O7EeyY3F8pcs7Ek+NGZLE/KA02AMKQBqzvT9o1i22X
7/4GuQW+gLVwEJKFzTzbIUxBz/uIw1oZFJYCVRQ4B5Gq4malD/bwCsVgPC4tvnaLyTn9mAsH6G45
6x8Pwkv1zMaBBcTK2FqY+ZhP1G1z9aNwVEz6WKPCkjzR0nm8NYmIR5LexJaXIwy5xGRXZ6gRAa0w
hbbmKW3NZyqlTe2tnxSqs0ouhBT/VfPl6vQo2sVHntXfSWY99/351q6Qa3J5saAwqPJ+k1hJa+Wm
06R5DDWWRNxj8ewcwdzVutXxZvkqxUsNwnYoAv+H4GAiYUPQOMsBQjOi7wiYYSgLZOWqBjK6tErA
+fwULbH2X3PpYqON+u0IPxkFpjBhbg9HI9THYb+VS5c9kRHJqYB/5bdjvRbWFUqFtXgAV3gncDTb
i9mgMvjcl6VLXPi/s4xjMKOuFgvYhACRqdp4lyAYIdst3HZW+H8H0Syx8uV6gArzSKfwNjISOZNI
W5lJmnle+0M4L9liCy+93hRclV/wKPBPPvVctt+d5gKO9ib8yexm6MMJ8VuqQIZIbKFO9tOqzQFR
brrtJQ1B+QcpeGlHHBaUuLyHj7Qui4txj3E0ZTOsXr2XnO+FYhdRoMUM2lP5rxni5uMlkppCvjKg
Y4jq7mz/HJB4D8g8l2oCZHS7+9qsu3mMlGWY7Wu2GjM1kCuo5DANu/j0w6NsR3dNnkSaf9q1fBny
lj2ZUDdGbUPiSswAIoEpifjEyS4xFgrWbQjwgc4hlhFq7N2DuGyttueLMTFZtREfzF6AQSuvq1CA
uL6LOTFU3lZ7rpKNyR0p2I+Rzt7qu6MAOIOtDjy5sWXb8fQwTIBemYuxBX8wBk7hy2cXpX3rhtnv
lxzQd29SO+gcZ2kIvApO83WSlGzgekxi62DbFtdBVfjqumt5lDdMruAcEUmXYzeoOLJFB90W/5DI
Sf8gTE0BwmcQCfZx0GgVgTsh6MFi5NOWpLKvcx754/QOL4K7Ht0JYHEeiACAQtk7/QHTmpHrYPOv
awiGZIC7hnoL3S4rdJY+RlTUM9lLxCio54jaVUJz7AK3y37yhS8XFmngOpTmOUzI0JBe2oAK8Gdc
yU0iuTyY8E0dzkvB8BeLNSk7PDo4kTDoicf9P4tCgx2kSZnCeiZmytxwehyaZwC7GVHrg1b2TJ87
Qwbt8q+OnxLTrYbdLHhDfqXjdU6KU3OL/YpuLfY3e8pyh+94aiczCTJzCjn2x+KKG677vSOZFfg4
056OYtnOquKIAitPHpfpAQ5PVBJk5cHPodycfx0mAh6taOZT2K+TxfxSLyhdXFljjTM/gM6NAuIK
xb4TkEmb4lsdenZWF+nl5DEmtW9mfJ+hYKzdolOX2OIsorhCoh2MeOTX05menf3KfWiS28o8Y4wG
sRAq+ozVWYSotrOzTfeoM1UAKXvyERWh0K49LoVBGOhXlSfiswuNfbYtxxYtdA35cBACUqORmQ1e
pWjPn5aAv4U71YMOejdzWE6qeVUf3OfWoeIj9rNqjc0pFRsqKqhkQ1ThkjZuNUS5uE7cqOm2zJRC
i0zT7tXXc2ChiVrllJ70F0z1a0la81f06myh0iDW3z+HxJAnZZZ0aTTcF/iWEcNxoCcla1v6kLWl
LrATb/OYz70nN4gYSX7T51dWRcaOE4WNbq4PXviyI8BmYs2LhPqMdFjV1nHErT6SrzzVZFe11L8T
2gSNdzvLtKbZE6DWEL3yexaIm/pgJQKNCrziwLeLv+3IkuErSTP4+i8Gfza9VyAVmuGd/uYHUUF8
FNPb/izqXv+MovjrHzkzZ8V5F8+4TA+zscBN59iJTpJW2tJiqmTjynFuVRC/0cwPOM/1hsRpFSit
opDJfeyQG4aMsHouZkmqShRZAHQmdbAgAx8kSkm8nPIgRX1AgQs8xSYmF1xhseshxZ5G+929gajN
cFR+lXlnfQi2Cy2VM75Wt4IFi9hUneRsArwBqxCxx8OHD0Js6vyY1lQggjew2DEa/lObC6nsyQPN
85nQUcvYL8FZ+nPg6apvEsgzRWJI0rT9d6BNjW35hzxzZ1y40nZVjSc2Ti84txwvGmiGb9Ut4yGE
dKpux6v1WeiuNPub232bTzKWaZjaS5sUPtwoRUlGy8dQrDVLTkghJjs5mzJ2SefjY/4f4dJ8YOAQ
O5cjA4RabCApEQBaCD95WbnOXreGMeXhtfzt/XgxgaCndf+36XVusGiSUSbc6U4OD+C0VA3apN0H
PmPSU34Ngm77zOIN3Odh/G6HD97iLaTw57pmYAO288Mjc3qFX6cy9Q2vQbDE/nuBc5KHTF+yi4LS
MeIRWH34YQikxthyP7h7jDZp6D1YSTyfjUGYjRVbMmIrSUboY/bOpYKp1gGD9W7bC6186GNF9H1V
qs3HSYKW0EshqfkYdDWtAks4dol+d/jFNGEqN3RhW/2+a+jLWrDC+lo2Uj+eSTRSdY9drwuZGtGp
bZzT2r9zTPg7c3mY62rC96WiiO5FiYjkYoLQ/n/YyV5Z3y3WR9ZKDzuqnahLnok0l9STMHxocVk+
FtwuFh3ZeZK/tRU7xSTjF/mfRi4drqtROY5gH+GgVy1yb8eGFZGVYyOWCEthMXgWHVpDW6casuze
vmznISRrle8D3RLUXSoSUuGg9/Dp6dYAGOYC7PUyMra5qk413iH8/2i4rxcmca/D/6vp29bn0fhT
A7RwrJGmZwvQCPFoKXkCripeGHSqvOYK+IPGiPr8RF+6fa3L6LqKsjb5XTFCcx0WJUiY0cfd+rVO
/5dGmcWay0Xwk2aRNGFOluBggK6GSadPjfc6zrKacfMXdSW/G0pIJAet9indTWOgaMHtL+wjGa7/
rOV/OqrkzPGRaW+Eqa8QxZZvAocNg75FoSsZgODiHx6CVUWmxRudWmaBHrcIjZj31gNleTEGP20O
gZp4n9/6HCYTfQt8nCSNmMyKJRHv+3gLOH6DcCBf8nkXKwjhPdwJbddc5zjjt3YNmtNyqmM9AtDL
Rw1rDTx2xWJwaxxfGQlVQGo3F1YP029n1GUjEJA4tX0On4gwpQcpeLXg9x/0cyMXhXjQUimdc09K
sFkZgjpIN7EXgR6CyNibdyzlYF8rLpd2mASj3m4bYzVHkwiAgbVqI8W6LYflpx8FOzEWDF6If+4S
3aPXKgyqiXGMjjC9hMPZIAZAasKYb7GJsL+h3YH8BbZv2xfb//hV611Ud2FjnZLbAiKzhFGeQI4E
svKH/A/0g6TnjqKUWI8HtrA9gQiUNjCK8M9mObFOuEsOYCrgKFQaqPEtaX4WWsS+UZUFgHZ1FozA
2N+nKl+m6NU9nt2t+h5K4mkXxETdJVZ+eUyuQOSU0gE58g19jMiGDde+KOou9gZToUyR75l3I/Dr
8nRISEf5rFKJ2hsC
`pragma protect end_protected
