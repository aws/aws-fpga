// =============================================================================
// Copyright 2016 Amazon.com, Inc. or its affiliates.
// All Rights Reserved Worldwide.
// Amazon Confidential information
// Restricted NDA Material
// =============================================================================

//--------------------------------------------------------------------------------
// Stats interface registers
//Register MAP
// 0x00 - GPIO 0 - read/write scratchpad
// 0x04 - GPIO 1 - read/write scratchpad
// 0x08 - DDR is ready status (bit 0)
// 0x0c - DDR reset (bit 0).  Set to drive reset to the DDR core.
// 0x10 - AXI Address - AXI Address for accessing DDR core (refer to Xilinx DDR specification - pg150)
// 0x14 - AXI Data - AXI Data access for accessing DDR core.  Read or write this register
//                   to read or write the Xilinx DDR controller registers.
// 0x20 - Write Words Low - Stats, number of words written (512-bit words).  Write to clear.  note is 64-bit counter
// 0x24 - Write Words High - Note can write either register to clear entire 64-bits
// 0x28 - Read Words Low - Stats, number of read words writen (512-bit words).  Write to clear
// 0x2c - Read Words High
// 0x30 - Self Refresh Request - Request self refresh to the core
// 0x34 - Self Refresh Ack (read only) - Self refresh ack from the core
// 0x38 - Restore/Skip - Drive these signals to the core
//          0 - Restore
//          1 - Skip Mem Init
//          2 - Restore Complete
// 0x3c - DBG Out - Save/restore debug out (??not sure what is on this)
// 0x4c - XSDB Select - Drive select to the core for save/restore operation
// 0x50 - XSDB Addr - Drive  address to core for save/restore operation
// 0x54 - XSDB Data  - Drive data to core for save/restore operation.  Read/write to this register triggers
//                   a save/restore access to the core (with XSDB Addr setup at offset 0x50).
//
// Interrupt Status0 - bit0: AXI-Lite interrupt from DDR core (refer to Xilinx DDR specification - pg150)


//--------------------------------------------------------------------------------

module sh_ddr #( parameter DDR_A_PRESENT = 1,
                 parameter DDR_B_PRESENT = 1,
                 parameter DDR_D_PRESENT = 1,
                 parameter DDR_A_IO = 1,           //When not Present to include IO buffers
                 parameter DDR_D_IO = 1)           //When not Present to include IO buffers
   (

   //---------------------------
   // Main clock/reset
   //---------------------------
   input clk,
   input rst_n,

   input stat_clk,                           //Stats interface clock
   input stat_rst_n,

   //--------------------------
   // DDR Physical Interface
   //--------------------------

// ------------------- DDR4 x72 RDIMM 2100 Interface A ----------------------------------
    input                CLK_300M_DIMM0_DP,
    input                CLK_300M_DIMM0_DN,
    output logic         M_A_ACT_N,
    output logic[16:0]   M_A_MA,
    output logic[1:0]    M_A_BA,
    output logic[1:0]    M_A_BG,
    output logic[0:0]    M_A_CKE,
    output logic[0:0]    M_A_ODT,
    output logic[0:0]    M_A_CS_N,
    output logic[0:0]    M_A_CLK_DN,
    output logic[0:0]    M_A_CLK_DP,
    output logic         RST_DIMM_A_N,
    output logic         M_A_PAR,
    inout  [63:0]        M_A_DQ,
    inout  [7:0]         M_A_ECC,
    inout  [17:0]        M_A_DQS_DP,
    inout  [17:0]        M_A_DQS_DN,
    output logic cl_RST_DIMM_A_N,

// ------------------- DDR4 x72 RDIMM 2100 Interface B ----------------------------------
    input                CLK_300M_DIMM1_DP,
    input                CLK_300M_DIMM1_DN,
    output logic         M_B_ACT_N,
    output logic[16:0]   M_B_MA,
    output logic[1:0]    M_B_BA,
    output logic[1:0]    M_B_BG,
    output logic[0:0]    M_B_CKE,
    output logic[0:0]    M_B_ODT,
    output logic[0:0]    M_B_CS_N,
    output logic[0:0]    M_B_CLK_DN,
    output logic[0:0]    M_B_CLK_DP,
    output logic         RST_DIMM_B_N,
    output logic         M_B_PAR,
    inout  [63:0]        M_B_DQ,
    inout  [7:0]         M_B_ECC,
    inout  [17:0]        M_B_DQS_DP,
    inout  [17:0]        M_B_DQS_DN,
    output logic cl_RST_DIMM_B_N,

// ------------------- DDR4 x72 RDIMM 2100 Interface D ----------------------------------
    input                CLK_300M_DIMM3_DP,
    input                CLK_300M_DIMM3_DN,
    output logic         M_D_ACT_N,
    output logic[16:0]   M_D_MA,
    output logic[1:0]    M_D_BA,
    output logic[1:0]    M_D_BG,
    output logic[0:0]    M_D_CKE,
    output logic[0:0]    M_D_ODT,
    output logic[0:0]    M_D_CS_N,
    output logic[0:0]    M_D_CLK_DN,
    output logic[0:0]    M_D_CLK_DP,
    output logic         RST_DIMM_D_N,
    output logic         M_D_PAR,
    inout  [63:0]        M_D_DQ,
    inout  [7:0]         M_D_ECC,
    inout  [17:0]        M_D_DQS_DP,
    inout  [17:0]        M_D_DQS_DN,
    output logic cl_RST_DIMM_D_N,


   //------------------------------------------------------
   // DDR-4 Interface from CL (AXI-4)
   //------------------------------------------------------
   input[15:0] cl_sh_ddr_awid[2:0],
   input[63:0] cl_sh_ddr_awaddr[2:0],
   input[7:0] cl_sh_ddr_awlen[2:0],
   //input[10:0] cl_sh_ddr_awuser[2:0],
   input cl_sh_ddr_awvalid[2:0],
   output logic[2:0] sh_cl_ddr_awready,

   input[15:0] cl_sh_ddr_wid[2:0],
   input[511:0] cl_sh_ddr_wdata[2:0],
   input[63:0] cl_sh_ddr_wstrb[2:0],
   input[2:0] cl_sh_ddr_wlast,
   input[2:0] cl_sh_ddr_wvalid,
   output logic[2:0] sh_cl_ddr_wready,

   output logic[15:0] sh_cl_ddr_bid[2:0],
   output logic[1:0] sh_cl_ddr_bresp[2:0],
   output logic[2:0] sh_cl_ddr_bvalid,
   input[2:0] cl_sh_ddr_bready,

   input[15:0] cl_sh_ddr_arid[2:0],
   input[63:0] cl_sh_ddr_araddr[2:0],
   input[7:0] cl_sh_ddr_arlen[2:0],
   //input[10:0] cl_sh_ddr_aruser[2:0],
   input[2:0] cl_sh_ddr_arvalid,
   output logic[2:0] sh_cl_ddr_arready,

   output logic[15:0] sh_cl_ddr_rid[2:0],
   output logic[511:0] sh_cl_ddr_rdata[2:0],
   output logic[1:0] sh_cl_ddr_rresp[2:0],
   output logic[2:0] sh_cl_ddr_rlast,
   output logic[2:0] sh_cl_ddr_rvalid,
   input[2:0] cl_sh_ddr_rready,

   output logic[2:0] sh_cl_ddr_is_ready,

   input[7:0] sh_ddr_stat_addr[2:0],
   input[2:0] sh_ddr_stat_wr,
   input[2:0] sh_ddr_stat_rd,
   input[31:0] sh_ddr_stat_wdata[2:0],

   output logic[2:0] ddr_sh_stat_ack,
   output logic[31:0] ddr_sh_stat_rdata[2:0],
   output logic[7:0] ddr_sh_stat_int[2:0]
   );


`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Z6uhfLwj729rYpSb/F4AmCSJYOWIPaMexRYhlWJBdDcmINccAs3p8zBFPfzqnkPjKsy4/XsFeCU4
6xNcuUopswg3f7VfI7Wx1bDt/mi2Ul0hod5Bt+9lxxhOavcwZicnFI2hx0n4TBJCh/7UryFJ+gDf
lxgmDSQlp56CCncGkWSeVgUmYdGqPWGHH5ERP7ZYqAJ607rEDqTeouAefY+aZrYz/nGh2TGGO50E
FltnlLlIdxKAFbtgFhlTQ02MkjZfPdOyap1d0KE24f0TUZIEvp9bvJLqPqT6lgEN0Btftptuy51a
3Zbh5Vt/RlPOPnMPnPsy8bSb4Pc1uD3DZJo29g==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
zE6zreo2tMNYLFuzkqBniDNKKgRrVvdL1AsTE8AY0YgtaUVdeAIlSWFYz1P7EzmJvPEJajIUHXHp
aDcDDW9vjLl9f19FM/JOcjo6EGaIyf9aZjGoc+ddmcl5XYNOokRGDETYkSB6cWGC8QRgq77hRRZ3
DQ89sEJg8D2QfRhm8WU=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
RWpl9t3Nkv5l7Wpp0BTpdnQVlzUwtqqmnIzCvWN7buMLEe7As3dGqCoHwG+rsLrPDTjSDSuk/mjT
Xx2jWZ1EnEk3ZTCKNyXql2MkXJ/HWwD+cKzhoLqLNz1A7QxsvuE1rlmdLNKS/q2lXfhwha58rslo
oBvSxSMLR+XjfRAo09o=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 46672)
`pragma protect data_block
qchxvd/IVapFTGqLFY9jDliqLdJMqHyONzrJ1e4NGh7Z3TDRhZwb3A2lZxnj8ilPBIvJUDOc+sLx
yGryPwLG+ZYRl6U1t+ofKhZI1fxPeIkFYpsBsrG8qdjyyyup2xG6q2tnIgrBig775YQLMkWe4fih
0bWt7a7ogsN2GFTlyQmze39L8bcvDA/78vlAtVFNFCN7juJV59Vku9WCNNcvFYQA5lUT/t/iZC1y
vd7jP2bzAddyRlFobukYxX+ghsx/yaEwsygUyiwzoWpoukjtHIppLgIXas2ixA1oaBX3HyVmvlpn
/4nAKj+1YSqOd61z91eFPnAC0/93VDpYBspSHBJbKBuO1lU/5iReE1Qmf3gzoFQiebA2w4EMLjxT
kw5djTaxUa+TW25Aax7d7HR6GIo+3erXBVMZZCDVm5JwFGSysIHyqprOgwdChcfY++9hSX5Cyd/A
R7naxCIpTPrv2P8eo/BDh9Bd++cnkJYTi4mAIU0amEDZEczuNN2t4ypAKq6nt4X74mfLJrDZOiJM
FSkq3dEVRJNJneYbnMxHz96T08aIiSbtSV0MeDiDtX+hB3dp9IKkk2kkoZkhauDZ5xR+jhxtmdjt
DTyj+sXsOb6HOZ6/QByYMuTpKUrBua/6vizpWhfu3vQoJx0gNlwMmbiqaXBsSsIaqdJDBc0K2DL7
XIA9/T1gy6TN75GuxsN7UyVu9YZZe80iFhAiI/eok3n7E5Sl7YHY3Cdut0n8yPfUnEivrYlU3p7x
hASNKKUavYpgGIpbDjFHsYkyK0NKfgDRel+Y9qDGN6Yl391L8OrIh3GfiTYX2i//6fWHvgIzS17o
uurhdLlyuUGvMlatO8QQ7FG+GwRNFzJY3QddyAB5V4a1SwJ3yLgdKXNjn3nsyl1yEKDsKiPE0QUi
UuRpXY37mgFaDfMuqojjPnt0c40rQA7Av3oGLsb60Lxa/DJHkBblM5R+e9+yBnoeni0OMtkoTVgb
fMX0yzeYYTD5lQlrDqx53UznLY6hlCech3cuVUUrlRXRsn+WFJUPm8ar3TMyPmaipZEd3z14gQT+
DvMtLTHCdaX+hfNdmvR5qxlB5aDXnupP9/+r6G8pE77oV4JkWCcLrU9ZpkA8MG0SHqPNxr8tsJj2
BQkFXr7+cFjyL7NfS0T4w6Cqv6APisO/dK4CsXMPGG+femfylGAWOBh3o626AuuelJQqcUflyq53
qJgL3B1YHgvkxs+nINJnxLfIdi9Dzr/2qSjUgFlBxktQqI2PAKZ85SEcO/s2fk1kU9ttNfzE7pEI
fN+JS2372Yw51XymW26khEEA6dH5Z5OhsaveBrMP5CbbTvn1cECWWsIlPPQWLq1VATnBZ7cNEdCv
T6iRntAXRt2VdeiYhM8ulf3bMfhYWsa7LnHiTQFQrX+cG72dTfU6IdGihFwHopxjZ/o1zR78dNZd
dgw1QPO5ceL/bxXo16bvZDxfdzg1ph5khN2p7DuiXLZ8mkpEyIR6ISYH3YpVISlekGiL7clB6oku
+pz70N1GsG5yHyuoxL+9XK53aaxXdbn83DdtcDe2P4Ol4X6rttt6a05NKpTV4gWBGvs0ZZEAd4Ji
8ywk8Rw306EE/44dxNqTg/x5UvjxDqeGgNxvZykJ8CV8OxVh+kWYyAz71gz7C98vvMyoGvWvvFbH
yuazZS4JGD+LNY+zsIoGAZG+Gx1CUOIfIBCesaLF2URurUcergc+35toaqcvtueqTVP59QZvWD+R
BxPKfclv4rRLZ5Rp6S3Q0RKRLJZ9rOPsfMd7AN3aLkWqeBA0237JhN/r6IrGah0QrgRP9Ag6F88r
b9WSkDuApKbfps6Dwaa748R+D/GTUsUNlL8JJaW6p8WA+qsyYzoj3oJnEjzvZf4EMC1AP4VDxaXx
4PB94YQkKZe+XDmmTPkdB22WTPNodlWAz10sMbgJBu++qBdTPtxoVuzGxvWpgg5VSriprAPgPQJH
w+Q/OOAKuV7Y4D5I71S8bGfIsqmF14VPvVH5A9KHzr7U09e+LqOLDBtnZBZd9vck1O1CMpOSGHV2
X5YTVVdrFnSAXoCH2PSnsqSQNh8NzbYcBg5IxmO+tOoIldgLYXo6ANOWFQCs/B/UQAcHXvKDnTg/
drVA9OdBdcd1ETPNimcz8lwMp6YRFMjlSF49oGlB+iq8zyttPHVRdlAnwno+qLMDVMoRHo5nApDR
J8AAEf0LE/Tb1DHkfxmt51EtyCirvewkPnVHAD+KUBqWC6O2J2sefJswK12q4wAhGlJO9MIDyxMQ
H5YzeGShKfF6KgAWIYRTaF562PTJs5CZFpnRib4dYKRkN1b+ntCtCDXIrQyUSN3KxCPE6hE8/bjx
6wHpXdNYV7fZXMPi+nFAtqTQlXVCMQednseCjBBYA8sGICwf5puCpl3hKceYMf+mh/3N2c2Vvnm2
4LJp5wJoT4RALi3Yjzkz4v0/LwBp0vnFbpMvVTwKJIxNmz2MuUf80jQ6JPNpa0IIfI+Bk+NvUwiU
TMshh1uZnBlpz4KXP/kaPA72K78SbYwJsZYHafb6GVjSckhevZtpQpn26Sfnkaly4wJmxXQ14G9p
1w4Ju23/K52YpEYCWZuRwToDoQb6uDVm01KD7ixF9oEw0RsmvhYsQ03+3MVeNprHSKDd1yVwvUh3
ZzLPA7NT/hCOd6rPG8VSxFYOVAYi8+RcNWHPS8K6OiqY9TcG4SNwVsEJvc75nlbcR9Sm9PLc76Hp
WxgYtNcq9UUPK6j0T/R9J9GNzhpZ09joU4lImTQkWsvKGodtteDRFSFQa1pXRMCZ1K6lZTRBqbmK
f1gk+B5IMbmOxTK35BVIYbzUTo9qbIZbquzxwaDL8eKobxgC5b5ascmnPwdeumYdzO8XEiTKRZfx
54wso4owsSxKXTIGpVguKHl/0mLgqCTvXAnSxbVbFaiDEEMREVFmKC6+Rfsv9cBcJs4yuxpr1xUw
UE6qSkw252xHCUOiTht3uu4ZpOGnxMGL7FvAwxfGp263Ro0yJvOBLROM6rt3RhwXdjFBJyHoRpBn
V7EtyE7886MTg9shkHS+Aeo6FNY3nuzVCDUQOYFHgGgNYDxPolZIy92I973gg0M3vxPzfPq8IHsk
zEY4+l2D4LGJKGrSQdT7d4AItLBgNOygLYXefZCtw6UIyndxs+SIXzk6A8nzToxsznN3me5wBfbB
EI6IBJIEud7TGHTH6qeKFOSKjWfgbT8PrNR5dHB9SDUlnvApa9GM9QK24Rx+lWwBhjJUKUzAGaYA
ATcjUYXMWwqyd0tdh5QKwNgh9kplTi8b90OllumYRkFIxE0OFABExJNzfr6FP1nQfaH+VvqMM2dr
NWhWsG4oZAQ5adyTGjHAWzJuVrXVAje3ebG5PhDrBQ6PLEoi5TUks8bIOSeseMmdCXii7eMfcjI7
odqHWttpxNbyXyJPlYbdPaVeU9ZbnWLThUgcmV30Uy73gDoNZfdcRHbIHhrqkypgrGGrNQQkkgUk
T2P8Lg4jiKS2rYHA+E874uDkFSTfCbbr9Hmlp14glxTrBufRF/NuiN+baAoOzV/bl8vEds2udE8G
5nkEB44TbI2aQfRT4qkKd3U0dUx+TgW6VnBoLHwlGY6A7NvdouOruvlAAOjADuIf3bo+5fpAuIfq
r0IYbNtRfmiY/8LJga1bBOJEzk7vo2icxPdsZbz2oVXlRKyX+5IkQ7E7/3sO3xLlQEZVEIHl0+DJ
FhxnTo6boLJvrAn51upNYd0d3FYn+o619tjmOscUavuk2YAnjvm3FQMFHPlnliXkz1MJgpG2bdge
56nABiXyY+dxnJEn9VWh4y1A9QZ1PgO4rtwx+7coaNca2r5+S3KCxBM75irQt84AbUUTh8sKDjUf
nnCCix3tyW5uAUeASfDBmIvLlglidAAXo3rmOzBppQifwV81YDly2Gy2J0IU/a5l6b54nHrmYWdO
vN97xTAma4tMo9t0sS8cBb4FcpciKaa8u7FJeE72UYhR/zlVgRjnHVZcoivsLAy/fx2PWFujccv5
DZH9Ha5Ceb+K1IQ/2XA2eRuuNMjqMDpgYXxJTZ9fK4Xn+vPmTqBgnqA5M4vEv95UeDSCqPTY5uUT
TAhZ6v20uM0xxvZeC5OjAu4cklvFvFZ987R7IBommPHlZKMXtEA2HFRmbYkdBXUJJGrsp1IoKsc2
bPnXuEhecQ6oilgG52HSfXjwGgyZD8eQ7aWBZ+pjfEsn3psN9QchUKldHlft9geUAVh1v7nousi5
6DYUi02iqLB6RoWB1xJnb3UIYAYhXfSkXTtch15QJpZ0PdEe0Nyn10ZmYgBIp5lHFoA1Nvo5VS7E
hr577UWO4k+m3qUW1d1TNNOznAfOYfbqIHmEHLxrCauPF1bSwpcmeH36ck+dmqxrj+K6NwJcWTme
BMQKJQ2eb+RijWt0seSn5Q0a4uljsVIo3D0lACskBXpzW4urNq6fcSm/jO28BK+ODhRx4I8xnh74
vH4wAla/X8eNDPMkr7BDFWShj4dWDGXGJoUYwmdhVcXTJZgLU7KWe//KCZJOSfdV1ZAcH2roj1jW
bTro8+ysZfl8d+DWwlW+LbwUpoxZt0zmFkie8AIr2+O6AeW+D+Hz4TwAe5WQlu4XaS2wFjo7EVJz
D+fyleBPh5QxduFEC7mbn3qcuJa9MEFSm2iPs2U+Kp2OIfvf1HQlJ5hvp/PhoHz98D1bjEKBjkFX
R3oDfBS2GLDxWEqLg0Diu/neiLdpUVOEOv4jVKYfEogEO1oYNxK2625gFueEopS4955h++QH8NEd
nGngevm7TJBjQNYW4ztpFAdAVDuwYIQbXIgJbJRUZlyfxDQUrzlPtrJ8HjGetnOGg0SWx5w6fzIN
a89s3vb5xukqgNnVtfvz76VcqQZ47HnEWD/f6540vzIEKmuZw4gSRKEKVfKxsZ9jw4GpR0Z5PBt1
0bIhI7QrbIlB8hdTWTTyXyPk3b3dVXkjEVOfBmthAuYkcskUPDgNSIrTRk4Sth1W0j+zuTtWQ4yK
/aAutEKZ408m3eajJdLhqluUctwjfGQJ2iMDJXsUeIvRTtMYLp66nPEf/icwA6WmixAVdpUVQdS0
ikGqHiy0t2LJ1SS3HGUiJ7NqFZn/tO7OUKQ3KXK/HVIWFusb9SNLGCuVRJloaDa/qC1jUdGKCB6u
NDtTsb14RkojH41j6SOHKiuGtW7lQ/lbb0wmaGyuTLa2MTEGRreh6MHM9rNBeKyY1plmrlwyLTp1
3l3sRDxnUL/t9sLSAFTqT+75Fajz9lnh3umCFdfLcuQ/PK4m3h2SKAVl+3LrR2EHj6m0OyV6kGzW
qsi5iwNfX34lwM1BQzYhiQi8ITZCF91hbtx6DgRBs+2/K0MqOky+L5i06WV+PZdy4iY1VJmeyxhS
oy0A6FekX1Y37ELhqEHqkVbZzl+A4yNh0lQ6FCQT0tSr8XAfGBk0gAxqwFZH+G71kzuDJHSzgTwO
15oTzTkTqdN3vT6ITsk0NJGatmmaRLkQPnzONrxF0B1Hhbcoh07Gj2FSDAo1k0eWHJMnZPSzrK1u
vBauaJs0sSFM6sYodD2tPNccPg10hmP3gqYP/jrLa8QBwqDWncEdJZ+wA0mvKCHmEPzr6hUOPnzh
Gq8o/vmQOW8F0lPBpm790OQGvZF5IlH3LCc4dgYwEZLGZ25Kcdgo+xNYqtFQUMx7189P8Iq2OsI9
2FfKRZzXblxkH6yplPsGEjhipnvIxIGMX2/LdTI26jNcJxNLalP6XpyOZWgvxS/mnbzUazSyNJDa
4lPMfCODC31tzmeNTCch7KgZHcoERt0VSic4XtEQihKrDFh4dB9vp8Jzw48LRp37zqD3L6ugOm06
4NMONHZpBAY4b0JoB97Je+AzwWEBW3x4tgc28qCLOkQOOT8Jv2JIo6/yY2YSwDqPcvXkNwsdrs9K
ITxzf8xARqIYWOa0tTu+7kkTXY+xq2Wk7Cs1NizsOcjFnw3nL369/oI5LSjmACHaEieBaKmLFteL
8DwaazwpgzPPYOGCJDUS92+hqwpkDYMZQMNAglL6j539EPqLSaZ9ZiUPdL+ITV6AmFCnPDH4N1TM
+lz7di75cN1K3jetkFtQxVNECei4oHjl/CDvbqqOUQC3tkDxNUHaP8V6DnHR/FERVjFBMxwQWnSw
zhaXWm5lenyHFtgTECczjW0TzUlV9BcGsdSQXjxtuTwArB7Jqf2LCfY2qSKpjJ3NlH5ZD2bgVQkn
z2z4D6fCbVbzfoFc0KN8O3mdNgYKZi1Dnc6u5yNupM7iLaKCyzeCsXatCJGmvW/xHHIFV+FjUS2T
1amtLj2ScntsPPnjUodvBJ0TUbCJLegixqgs3v0NdfbexQXFJV2bpfIWUxWOTCKK3YoL2Tv94Kss
8XvEpYo3/KNJ/I2U/zLbsN6Oql/acINq9pCSO1oozdg6Q19PBuWwQRLwKpmcE34MpU3iGsdqbDNO
qAJTOMTB5uit6UfybsKS5u4e7H1L4c4TudgBBqU9akqqAKNBZamfzpQ2GNvG1rxVWtL+NJt1viRE
JfVXaiv3eYQuK1jG81uUa9THKEUhkx7WJLVa7UQ7hZIfm5z036uGAktYgueQ3TkUzTp/fZIL6Ud2
zEaEqqFALwjJr44tku12VtRZii52yahkFT646IWDjAkmygdpZv/1txwwGmWs6BQ3R8PlbXFOdt2b
PV20jCsGmrBlMaM61JAvellblsVXWAtEjgCSkkwLYj00F0wk3eazKm7Q+AVzD4FPjnUMUwwZaCHR
Yn0+93BilQFVIgd5jcCpgw6BJfED1ANjvrI+pcLwwv8Z+KdGSLX2Qw3ZWLV3vJZZ5ezGmeubXb1p
XTMtW1uCzzNYX81lpQ3GtLxdgoTuzDl7pGAuHrPVBGx0J9df2wEUa0g3QFbox2I4t136S+lTSzLS
RaviQ6dsDGjLZuEoweaAOHJwoiOG+AFyd1Sc2GhQVfBe4EJFvcQWj/v/a5XnFc4Pa19g/KEnHP6e
HiySfCF/ZXejE1/pOztEl3/d4giY1/O/1yUjP+u5nrRN+kDIDbxjQ6+e8G3iFuhlKG8Fkcvyi3JX
qT2b8vhzXWqdnsCtieKfPm1ZhYmxLBbNLNriAlyJ4TgPfRgo/pDV2grvMX2Dy9oZ3yZyzo0+EzsZ
nqwa7WmBDSQ8xXfiEYJ3BoLY7uE722KQBqTfzw8Z+9tCFsZcgs6fjQDNnljWW/2hAFJOKT+Ic7ZZ
41FtruA3C3S0pyCCJktSBnlF4gWSH7pUopfNw4vcaG7Gzc10DP7PLfTQ4A3jQnPVbm8BYzYOBZN+
CkFuExN6Fq+nbjrUChO6u9LXrDzxLGDMWldsTRqiVsJ5nnbx2XU8zpluOpkBSlcdEP+JT2LWIkzk
z0EuoJ7kvETHcu1IBZ+3O9UfpNerZ9xmXgGnJy+AilTrriQk3NwIUDfQe+oXuj9SZ6k55w/5iBYs
ASkpjHz4hpAt30VTzXarB8qN4V8drYXPGPT9dOGR/yUO0La0UviUTRTB9sidvmypaXcrmmk/sNlG
Br/atInOlJ4iOZ9fdRAhVTfBdq67DvmCxHcgULVQoq8AgbD5DWpIYJKg3+Y/AZphWcKM+NirbM+7
+SGJ+lHKnOLfRO/TrcRqIRhxALmTPFyRxwxVhLgAGvSf6+g//cJEX1s8IC4IYD2wT8/BOFibEwTp
K7IkQU/wGRpn5j3pXssuCVzB7nKg0fzmVRFiIVVtZhWMfisYbrsTCxGullstgNICETakUYqfEwqS
+ieP27sW+3uafNsW09LbNtdItce0NFZCMP5xxnDtKE+JqJw8Lm23F1/cx+qlMgr1NYg36rrW02o6
7hsa41swe20nuIIk7YY6dWiKmAn8SkRsDHf/E+2HXFJLMWA6q1yyi5TwTkt0Lf3JqkRzCzCOHpkk
kJd/90LiQPQlkdnZnHpzdrIHZnW5Tpvmx/nbDac+sUf8zr6Hz00VClkEEVHAw6bL1dPjcVjQcFPS
skJDyxSE79DWX7KYaA3LfIzCI4SZ4CG9fshCwIbGkoHS94n6ADU+OOApC0BLyoHY5z7gCSNLgx/i
1W4lEaX4qxRnXyvUf+7ZES8kWa7PKJVU3KwuLBnO7AEyyhJadpx4hy9vl177XZd4ipfi/jL6y0aE
fEIXy2Y7wJvtOPqxzOXXu8/4mLRhusDzJJbe7yMeFJ9vCs72sK/UYPqwOcIjDCl5Mg/gii7e47fe
4cgNxD3WzSS5N1/REirBjljq/B/w+tBdMjSjgRXVehYNPy8rA9uCsfMFiRYMtGuN6uWaUl4eTq45
p56J1UTyauF9WysnqCWZHQVwSZXCwBsYQLnB9r5jEAEx4YiTV8zA0Xu74KgtzPHz0/dfhn6P2/of
OjjR+q5kfISD8dWH1JKHCyJvqW404NkrA9Fe0eqFqVIhqcDTS0YsHi6CM0YWJbiHgukv3hlWrvwS
yV+c9yozCqYxo6RSBRPQEHsRliBWkAuf56N4iNgICbU6bLuEglKVA24g/0GiIZenfyfiOG3UJzjt
G6OrDhKDWbCBosOKQLT/QIw0YOc/r5xagTYh6fguINMUwbAP2+JO7WMBsird0AyL6vZoIP8gh4r9
AqI31XB0pJVtG3aGloFfjgN10vhuyFsiz0Jz0n1WRxVjCzcXCHrXYEo0ApjASlbpbGCYQHAzWtaO
yplsR3+W0y6u2TE9tuD2Bgm2RUuavogD1KijugAlkf8fVwXXpM7SjMNUWjXMVLmb1P2skGqsjcxA
2GPu52HhgfXay4ad4E4jQsBB8SRd3nwALeeRjrgZWufDG2aS+tqhxrW31IZAvmHXKaKJ6R7BqGik
v5kftdDWwifuUoqI08U3xrNvaRvYTfFajuThd36tpOkvJriFr/m+Im0V55xOshE669iEA1McCm4Z
DqaGVCPzbYqT8pmRY73x5upgnD3t4/2vdxPyKoW6XKCvXG14Uf9xlJMhvQZhGkHLoTLrcotucWNI
8FocOi8Z7CPfOcXQd1qbtA1b2V/MGfmZ7wqJiuM/mwskxJUwd1k4Wwz/J94H/Po3P5CVmsqupfND
cE+OHC/McmGd0ulJJkVdKKWFwsEGCdAkY37syBxcet4CFJF//+sEc9t8m0ZELdBSYJc50EakLwLv
kUUqjLrWFQVLNe0xgOri82dS32GoXD+BwPWx0DFh2mzIYD20WQOAEYt6Q5EuggMb45rDm+t17tDv
a5LY5b25B1DYVngQxhzjabIIwBavY1lxeySy2RIGTEhSPJZZpA2Oo0qvwUlSu9k0+OkQt0rOsGW/
ooRE5mGe/SA3PweB6sPBFyIInvPdczLxn/Y2wjMOahzjvM8togPIHpk+9dUgG11YaHunmfcTJaOv
vkcAOot7WGPTuZvLf02yfZAKDEsAbp8rfaBlAE0TwQcKpMpUDrX0025iuP/bKNuZqNc0AvY1ARr4
izweIjY87lubsWSaqvG2Px2Fow867nNnTx2MYtU/YDgUFaOT2saYq2oDb9N+vYRiwX0HKuPJNKWG
rqZdrnDsgSIotAodBRTiTX4Bzx6vbeyKf85dvaaEMf++aQLtGhQDUQ/TzgpKlipL10OUhDRPep8X
w4+1/qCADa27TkLn2ANFv7JkRyIw7/naO1v7BtfkHhkXRDteGqBR+xLQImYuNeVt7jwGM4ahymSw
nx5zwVkpL34Mx7Us81TsDgTtrTmGDQGascV+nc6bHIh3DispsmO2ug56T5o2vOmzhK0zXWqJddBQ
YAGJkwwTtzYOHeA4vFZu7qNuF46TcTEarD9xnpzHZeO+SEXBc9xlBGu/LuUyHEa1KLNV1YKUOH0C
sOY+e6USu9bza3ujD00O2oUt5Ep3VdQm0s+QBaLKB/fr9XotZRMliYI3VGXwQAT7ROV9rzTfFWLt
OWUrQH/9UMg+PHGibp5d0dBeQmpXYzgsMYczt32zPfHObFQio1hpHOTv3T7G+Xck2qpwuKdC2jKT
tX6z/GXhyfXdvMvEViK7HpySs5AohcHB7CODQuRgAi2wVuejrwTGlDAJi2eb8dft9SII9OwS0Ffq
VrPqTicBMCDAWnOQEC7wIDoSHNBImQfPHaq64/3y1q8eQ4tugLkC5gx9p7jstupa+NE9p9QvVx0O
G7gvSU5IpywBi1PfDtMEdozesW1+H0SuhgBv3YRo2hHKJQZzvKR702AfKSNe8IQayI2Hcl26j1vW
cAC24DuJiZYQBbbmhFZc33CD4pEs/RxTKg/g0OmCS//C9qWFJRkzDL4VxNUkRHlfQFPUTYESxGRe
Kay7WmjwdMyIZodxEfmUOTNiLCmmKvXilE09e1dOeanUffpshWL57mN+AGvE9hIizYC5DqLKtAM+
pdJ10PSlqMRS4tMnXw8hF1cgBsL8YaGpP1AQLZ0rhXBzLtsmvqYJ2F/2s8yRu1ciR+SWZITdnWvx
vs707vKRyBXFmNdInuF8d0B9KlNJbXfVStmpMLAfbSD4lbxX3iP8BQvgYYJGmCq9/I+jh4QJH1Hf
CswlE4ftxpMNKRlIM+pXiMmva1jAkHknB5AYBOEGdcdZzb0mpFCfsbyiTxoYRkUmeOCM6TBXKqi2
RBNtXhqARHSXhuSflKEBQ0bBdBfokK64XG78XxpCJyo3+MGNoUAGkvrmdAhmGBoe7y7p7a2mys5d
9rzA2Myk3KGqVuLH2caVF0aysRDneCkPkXYZZ2+nTEOxizNe0ucPKY7I7IR0lcDO63RewP9PjScE
s/yx5DKlJnSMg8vk830GeyuLJJbI2yrqmj1tTGqHa/MW0BM3Lj1lR11ePwU+WIQyOdw1ZAdnzYxG
yuzFj8XeL7U0Df0qHRmPkA+6XQQLUqNcIn66/tAcuMr3QwQMH55/aZtGRIjTY6zw0tqGEUKmEMwF
ctj6deYlISXVadU/Tsj0jHaApflUSjaGdlX/PE/uoB8D2MAtD/TukMR7lWUv+m7n2PwJ+yQjIRjp
CTI20HJAfbE9cm95Z3UUf6mkEuAL8fOdRByUrxI1fWMdnE4dUceOsYQr/aSnvro4BOpO8wfpib51
d22l5Tkp8bUPcd0VVBAK6xwh1pYWwsI13ip1UdEtHYrip1paAzy/Q3N3VRGNszJ5BoL3W2YHx3g6
4HmDhVj5BThyxEYDVnTuCg4y0ZO0oLQ1EsT0U5eS6gnljw5k9BCdxCFMzE1fBBHZ7BXz+xa3lKN8
mDtHLafxQqGh6rY0SHA+sVwwPLfp1ackHW3ZW+wtFeyRET/xzPpQudi/wilXHDnjfhpymFInGytr
adXnimNCb6qWYIVlkOMoj/53M4aFN4opPCqBb7UKchCZE12keIXTDVoCBF+vqS5uqn0Adc5IgbpX
7lYm1VMVpN4zg/sqrBtN1ATymFBZ8xRuLAVLU7SBm35hFV8efeqfmtf7xoEIByvUtY4/B0w4h/61
a7cHvqb7qRPeFS+LUmw+SouzSoMadPlzt5VYWmbchxwZH9QvE9gmpeojmNuQnpjl9n6LeOGvSVGu
CxCmSKkzZjveukMzAxeVsCgUpQ/sZx3aehhAfJ4S13PKOq0xekRgNGJXSSRki7vUNScMtW+Ss5SL
zSVYUNXmwSVwJ4anKP5NllPPrQaPP/Sqf7R3XgExduWqbKVAUAMnbWqQGfNKVuxO6ZTvah/EGlBH
yGjaf48ECBJXzzULOcRQQC9hEyqV1C8VX0e4WheV7BSzMFTQp9d3HiITs708N0zTGfKS8bki9kFP
8S7Ch6TL43Vy6ZgKDSapTrPB/lcuC7vIw5ePuJaG2jAm4rohrkFZg8EWcyMB8q7dD7gW5qBPgxQ6
2+1rj5IGlNWOgvLnHzeyNa0VIw0hLinYalwgiVcw8rXoTFHVtEO5Pho14cONhrt47JV815g4BaZo
7mkwCBTQi29VnFk4qCpi8DxNhck2LUtLD/wsHSSrX3gcZd0tMozhrs+ovRnk2dIZ+f1ECZilzHb5
iOBlnThR3jmwnYhCJh6aCRCNDM8ZWcNLeFQbxR1Rk6ixcqDugubW24sgvmuD7Jo/gAeQ5b23VIri
UZS0hG1MrOArwddG3jktmoEmXLdWq8hjrHjp5QWC9Bj9PPPjMhGQn8k1ZtCQc3uW+6Za9hgnZ/Es
MceXoQqlB+hzITY5OUh5o+ZM9Smot0BC8FazAuaf3dGP44AtaK/9zQIEP6QmyK0FEr7Rnv3jiHnu
2A0QH/7jJPOijEr81cUaI7jn71HYBbRJ+vFSiA6Xghg87ht+/tnX/tSd/6u286jlKVcjD+6Iyml4
xekt+bEaAYM8Fzyk/YCo5MgD65kCsCFlwKcTscQnkoyYzhDvbDEPI1hQolZMhuYMz+rBaPea9tsT
nHFx3OyPzA01wN3mcihavEmqbEFz61+syksn4OkUdLv6ovHD4YZq2Os2aIqid6KGFoYHqhXILZ1F
pkZC1Zjv32RLPpsvdgOSU5CtAB9b0v6lacAzrHB/x1R19+Tpyg+crwFaaQLM5dHUGZSgSsPvoygt
BDOWiTffhBpfS/Ml6d9DYkq0+h3zeyUXBsSgqEYo13E7VZ8NMkb1Bpj+S8TJ6uCO4vxAlyGDzD68
rYPWlHxwHy5aO8XqaebozjqlEoC90kvivz/DShtnJgD8XbtJQKZ/OJr/lcG8C8WkARbV8LDAH2Cs
/B/PSmNp26ZAOgQp9ypZi6XiH+WHIS6rT57mzXruO8CjHNmmhkbOdmTe5i/16HRTi3SML3AqkQgn
/kCwhpV4un8J6sVW71DuOKv+UUiVDvMzQd3HUbiuw1T4hElwmgxpIW1fbCyMpPyx3j/4TYmAU3qu
qup2CNOIk9ek6M9qwXTOz5uatTqmuKmpRGCvmCex/P3jPLh3QyiltH6o4rVb/bKf54DeZykR6Dk9
JCzYiiLNh8CvEOlquNzMkvxEgoaiIbmL+me5ooz6PM1q771DV4Xs0tj0uUWE9l5jd5o5KsWF/Ika
FXT0bGxj9PvZQOo8fQlwuIDR5wt2o+/i0zhdqRnZfh/+7P0Qz8+ojtuyb+fmYcFldxTmsz4IKVio
zLFQDrg3HiDXnftlPZ1YOIg0ruynrR89Fu8UqorahwUwYEpkOHKDQTb0av40C7l56jSSv8RndbP6
PLyafL8INTov9EXoprY0XOvJdjkMlDtATRXxdM8PV97PVtQPzdb2kZh2DVyWbVntMcKWfScxo/E1
pHTyq+GRBJvGcheS3iu+nYgAyFuIU/d7ky3pVAOGeT0AdHui3Ya0/J64t+9V56FKQ+22pkIIcEis
kR4oMC1muHuL8vSYkzNZuSMZfuEp0XcxMwn4sf24d3oyqGDln3M5aZYfp7KjvtRqCqRJXaV6USmD
o9LfKgL/Q39Ex6G3J1vzigBAyZpjqC+QkqIlBto+rSkZ/cbw9cth3V+ARPq24CAgr4R8CVPi2Fqd
J8dBWIbs9qCBy+yOKsvtQINR3pUC465ParkpEopbAeDPn/Lpdn+0IvtVgd+w+lP3hXheePKE4kDY
nhq5L/PajK4nuiE9WFxWyY/s3RkkG5NYyev9F5LTDtPwdiNYPbMH+XiBaepnga28r91TLNAMZarJ
7FxfOsMtdfgU+166kHTVHtlktQbMBAj4jnnsCeUn7anCiT+IRD4GSlt7Der+2PQOPKSTAPjipHsq
EbWRSCrQ0TO0221ZMhH1gr305HNYHe7uZOIKLyRuHMlTyeSrV6RWV/ct49OhzAwdjvT3RyfIwhuq
Y3t/KVSFykudsBGMr2aTELbLeDXcQYe5mxKwcxKeiUlq7sTtSubEB2I2YTaq3t3mwv9PkuvVtLl8
Ja6Lhgm1udjzSfQmpsd0yShDbIb1x+LCv8cc6u/YtYYv/f6Pet/tGspTM8X5Cio4uUNp0Xlp0Okg
Kx8qJ3llQThTK75pqs71VmWJaWHDf2TmU9AG0NNawqrtRHZpu38K0UEbHUUzQibglNbDV5uTIwvR
HInIlfvBQjvbFFaoz3MFHxKGof+lTP2KFi/GNiW/VGPAtsJX7M1GgmNgWGRUOC4nIkgdhR/S9/tv
abznVopxa7NL1l1PGGh3vly7k8TR3a2LnW3Yqa7VRgViYC9yjsao58vDQ+mJpQSQbs5p7TkxYDxZ
1AwlV6b85oi8tgGawKVDKbrT3G/wUlBlllCbK+FLV2HWtKsZkGOk/ca8Ph6Ems9wusLk9pqwLEpb
V1sr3YKzlIeiCVEeTOh2U4hU+cmwsX6PSfk9MZ2SekS+fhGlDw+hhC5eHvvCnakjxgrWzoAvBNRZ
awv8Mg8qeCND5B0GoJOy36gq46j0sOgi2AATtuUs9foLIkCyZ9h2c2VpwL5axJavqXP9aTFm2pdo
PxwXKecRsRbLX9g0sBhTeqbYpFElOSpmo2VSFKbdPmZ8OgjM176HzZ6ilvRDUJaeBmBZXzwSROWv
xKrlHnYq6ZLJg3x3qi63+0rvBqTrElknUqMiXDRMFxhZ24bKrUrymAjc8oe556C10uYXEoZwdTt+
FE2Av1isygQBEAxh02X8E3wOAuvQ0GNbhD4uquj0Lrks69n5HMTbxwTrygHST11uCwXT9PhRbAs6
JQVUClY9paO7xSFK1FUNGo7qGuZXnj6LDSljzUdrAh94LGPMqOZHuw2aRITi1zHfvTnXr7zEOTzo
aW7uCSZthMiB9o0pHiGkNcn6kYJK4Ah+QCYmJGApkEpYR+QGa7v0dkfOt8P2q6oAL1OLfwnPBTYN
F8U8Ip8QmUF2pF4op65f1ui+QVXy7BB4xLuGyHNbvQbywT8TbgvPWRJL4Lqj8UEsYnpKlbtnFEBY
gman7YJTGEZxtOf4ISwpcX88AUd6VeXQQ2wux+m4BOWIAQtCpIRRkSE2feqfa8sIQN8WuvCHhmO9
ppaA/npPRRF3FGkh3RE2G7B22VB1rlsaBQsfHhAv//lAtuQrJUW4zjWCUfSM91AOUHOzhlD4SsHF
3dgZLxnORu0fMurd1TxQEyPhyYVPzxFfa0B1GaOfszwTSs0dw3oUQg924q3mv50Ic9r+VRoJPZ50
GXB/RoNeNBlevBI7VB+a9n6KuPzfjd7ZHDViglefhrKNeDxsX+lZOq1qDYfWpBN1Io4LGgDb5mHy
BxaYPurzUKXulGbYaP8HCYDpZe+hjAN/osVd0rIauE1ooedOGh5+fiW9ewmUDzU90AMSDQoYphdY
esWCNB4C2vdx+yzc2e21d1f9xCj1qwy1zHd5RlK36/Tu8lGAhmCDBuj+/kdVCDce2aZmBWKndD6O
WIqZrQT6xHXZIvIpXI5DJDznLPjacGVI05sAx9nELne1lKN4Ra/TmxrMEtMaGEV4J6YSLmqYjV24
3CczTq3yAogXSvC9W6oSnohOSXAfzrzzWj+A5WCdwqgw4aRKzNQ7ZdSl1wlznoHIo/TqksnLFix1
ifjMCv3tz9jSJrb+BmdWTdA7gnzYus7fLfbeRIa1yAbR+97MPUqcHDGisLiM9VNKUO3Ukv2oXJ2R
46jkeni8YC0VQ0LgrAWgVuL9xnRXVG5pDWldl6omxga7Soz/QSxqOc5sexNmmYqyHdM0KlPJCHhS
/2Rpq7TRkCENrqExKhvBP0cu8aFbTbzVhezFvHu62gEE8vm6xSB3vpVXYr0ME7lQ/x0Z1rkuG1Yf
J4yy8i6ufmUQUDVhjWZ201d6/EbmTxAEUSIxs7D3B6GJ25jZWRrc9lwnN04icAstkjejYy9cks2j
DyYqoW7TU3qUbg5QMo8M4nHPAdhvJYhefDoEwHi8r98Baz+7pjHLiiC7BZk4LGgVVkFfhkyduzQH
Oisrx482a9V6cR2xsCZJN21uYFrtLIhE3O8lPha57RrYUCl8dPhagWQGpcUFm5rPZFIt9p0j8rkY
JOYPYEw/dEcpZVt6JtAZLMUHaWoy7pGw/tjY6r/AK0HFc50RA3lz3bv+zeRBVFtTDWba7ZrOf4js
ijo+MpG5RJCJwJ1veegL0O74D2GVhFPutFnJLv5CzUV1yJPCpNoacXvrB3EKIThhhuuwpjQ/yDfv
VPBLuzAAwbxtIxBa2Md+bMYtJnEkx3dn7falUTO0zgUCL5NOsyzulPFGYlcPzmJ4s9/4SLsbPVvD
hniTuU0eoQycQgxBDtgJysbI9DS9+oKCNw31lEyqSTYA3suVEOTdTwBjYzAlvCwEwaECT4mWtPkz
gpaVKmVBtKK12snL4Kh8JLRjXIRqYsg0wCEJZLEvl41VHsyY4XFBjpfga5W0lxNjC13p7xEIQn2D
esuCU4uWt7QsoSthdMLNb2znrsmpHjkcCd3fQGx1mOQyjqO5sX33gYpgRek48lmQAWE/l4uwCx90
S/A3Pl4SouxqFHWq4uQ5AWl5WEwGaVhjhazxmRaaR15G+DiTA6l4KYi7xMKMEKsy8S1vAQn65B3M
T6m12zL8NV9dUk235hkIIZP7BX51BfNnA7hxFTKEVN3qud68CYCzTNhLXaa07wmbr2DkdCzcaOrB
CI6gT7jZwF057HQOCj4K2ucnxFsIvom/3jTXyJfF5SIcoLNPQT+SLljxN3bCgFMb9Ad0Ng8F8bWa
t2CFcGMYwdGkuVYn8c9xXTQAc/kyEZafYBdRAJfRvesvvuj53NTe9oSCJMtph9iz7au9djXd+eDe
BXOT1/RhhECEXxkI4YF9dqOQk070rRFMG52XdWawQbLVb6RtmdxmHev/udwMvCnrjF0uQftLJncQ
w3ip3m8gqy3KVdPZxIQ5fYeyxz8itr7SP0kH0f9V6rKTT1Ppar3jPonFRQ49u/QbIBNcrKZ2RMXA
lzGMYb3thdAIC9K9zYJl9M8lUJQRv3yvuP+Lf1PdD0oqJp7FWYKFEiG06ekDKhk4rqGxzo+ImW9X
1GFeiLxwXAcAblpV9aSyTO+RzWHwM1urlpRPgNWhVoL2bE2+n6uXc0mqq6XCCg5BwqlM4DEroFP3
15Ps30J9Wy34/m/NqDbxNkva+5KbLgdm5Jih7dA1OdXyCwxsMGCiu707dzdmmy/C3t+RRL0T84oB
PTNoZh6zdWMBw7sdO8euACCR91nMLN9bKTb9vKa/ED5Av52Sl4klSIcdbGcAXKiI+qtlW30uAsjm
MrXR0NwVyNCaGS3OgDFBswjbqtDYBhefOZJpV9XXDeIc97gFdtJusp3dzxewRboMzT+pH54Dylfj
uzoeQgG05BbIbv4m1NSQOQGGLLzLruI1gPaaX63JdPC3OGiwmm6gRphnNQaBguLJsUbKaFDleMpL
6Ncdny90Ik6ln9ctMWkZZ/xJx/3pjT0+oXn3/epN0Q54yJbZweUMLavVdgYoKd6zCVvdJSe94GoH
cZJARi+rz/pZhKtfsWEzMIn/Xa/kc8yddVtNQ6uakyT5AE8jf+SFvaDOqAERrEipRRia+jnZNEXE
BN6rSD51ey0XQE4Hwde39GFuVN/H3Yv3LmySNeJgjhN4/tVuhXcPagcrHKIOzsXQs/y2nT06hLPO
hZSTaiyLTc9TJrOLB/60QDrFrKjnZemrKlF9SZJtQd80pAjWDO0J+gkvO4FlLoSKZfr/A5cxyeRp
LENCRXuUCwJRceieUS2RoH7icgNfz2h+wW7mb9cicz3aibeiMGk+/gMoIpfNAAB8oZRChhQ98woF
uQKl/Y0h5wxZ6C6Uv4fdoXaUJCvrVReNJ2a4boZt7jDwwXwQS7n6ij1/fpWDfRnB1ZdNAWlMmnqg
mzY8mjVePRPeHLLO/83R3ZumwyCVUcvI+qT+S5Zdnu3/1McewJw7dTo92uzoeysAL6l645S+VRt9
KRr4TJSg8+55hs0MlvWdsuW0zEduw+AnQJqtbMZ6zWWFOk727gOTYN2622xF/mWrUU7s/rfkCx2P
VJOvP18FjfWLQOAiqI0SkOwEjPBmWt7fY/CcGgQBYqbokiz1gIATCNpQR2Ccimsx7sRtlTIFXIzd
7GCcThnQ3AqhubNyhaXsfHTIIGloRQKjvnEokILtuwrvQ1QG8FfkaFM8R54jyhTNXDJvtkJF8ViX
9lRWKLHXjNrGO1jbbiM39IOIiFXk92Gkiswrcg4jJOq7TsyIarhwBdCJ5pNZqbViHAXIzzGNxQ00
7xum4uqrXr/xkuEqQvvsKtdfNercQbfrAA/rgyTEb4Q+dzS8g4itaq6wEyAJt/GkCH6Ww+dTvgGK
RBgVoMLZ5LN27ggmaVsKJE/8Bq7kek6QK79lH4U8v9KLPewbuxvw3DTijc9YasDDJ8I2NQ30U5oH
BhiLFf2BM6XOUExy4l8+FgxhdEQW9nfySvby5dZS8EXH9tGYENxYE8ik5lqqRrrS25XpX5ThcoXB
K568tlHcqC73KGbJoYTF3TpqsFvHZM6YHbh8+AiBZB42tvlbJ9UCxEmWDD/BxPkGIOQLt4pQcY65
QcEBFScEA+a1EdOy+TrcnU4tUxGdseWwWSol6OCtTGNiDoE4WNkhMazjmuHat8vwWiHPHt0WgJhp
LArvIirx9ENSeWtNBUDvHC9kJaaEe4saa/veUn1DsuEII8KXqkk+1AqqdPwFSC5E5zHMJlwTf9rU
zHkoVd6enjSyae23OsEjjl+RUHdM/UIP5bBqbVd9+kQUrEEXntVwpboIQxpmgepp3UYoMNxYdMXA
EXVQ+U2DJCAwtOX7PGsGmhY42MXIozaGmf+CzHi0GZTdMoVAS7k0n68xGn/GUKwG9v4vDfNGW2bJ
i+2RoakGiAbGhF3DPp9s5USkGzfafyjRq1R0dgNlidyKOienehmGkGX6IadKURYrhLl9hM2O1mrF
MixAy4ltrzI6g3eO/KZUB9QwKXjodkphqLVKj6ZYvhKyCsdsxF052Z1HaVqODvAw9JUONH4h3Rt5
se1DFHOj94Rhd7IpzlAyiiiEpqZjn7/a98EME7Q9jYJeGWRK5DaYF+WoBo44rzrm00mNTszIVVrf
8HqvsIWk9+FbvahseT4G76ceENhu21v+fm+leUEuaeVbD6di8lfo+9YfxFcYtRwydyrChUuTYr/X
asPhK0o/1Re17HDMFMEseRKVkNJSpJNdHWaMR7Mi3BtZ6QZFogFU16cy+ekXDCqSluKoN+FhzXKw
yGMPfKFv95SHVxM2CQfwJiKhLeWIAdcPtx6QbJIkFQwxNwh+a1G7RVKxqh7D/qC6v8G+9wiM69pc
0Ldu/iLJlFVTXsv8E2JZe4ws2w1Kobn5AAC5B0BaZXjBnKXu/EiudFFt5qwX81/tmBTYO5mftJaa
aA2pCu/IH7kyREsEeB2CbeUAK4DYCXXgGl70YKCubVO/nOmpPwXyzWyoQvREI0u+tpS8Hl4j9a/B
MAn+nGxLocqcTb79ZzLP78PsY36nFLmrtlItuoWsIlbd8OUlfF3wgPqt0vqPp9GdyPEV0bfir5b7
/eTT4hRPPDfqNW1AxeCJxcPCa1axGD2XrkG01ph89K0nQcZYFgXyZLZh0oNkkVsgpHUGxNJuAPt+
IwSEfKUw8yImwOH3bG8DSI0Re6B8XGSwNouHOz7JD8viAapF0QACdDyFAsdBMdcY8fXRTBvC6LIK
zxRRiTged+SP4wG6ky9h3sCsLYBL2TScTebgn+2/oaPVAa4ILlzrQ4T9p52s0KGiR3yNkk93l/J6
wyt5WH6BKTOwFb1iGZ8kJA8OKYJIK+GwlpOLu/SLMA6ItMln34N1oCIEMWWcCEN9JVvcRPp3GFtj
YvBztTI73DIf2jP8MoyckSTAC2PlQeggZjD7Gbevp3gHfuan+kJDffZZhr2iVzOaNnX2c7i3JcGY
QcrhIc2ECZjivvdH2u2dlI49SiU7J5B0Fd8oaHixGdmK0VM3gzrT/d5CIwPIlK9BhUjr6RSoMVNU
1ieYkDcAhFPTPaQxnwnU+z92yNmNr3vOEROTJ8yKC3X2Ntw5mNaNxLyfetHZgiJ4RfdLiBBSZREO
hdpbOu3BgWanvMBHA+g9xs3GUD7ZmG9epMOT2de+SsofMkq4YQcrefEdqh++t9BdU0OuEKLOvyGM
yx2CckQ+X7sQdiffwQ8AsiTUE4p8DUs3B/M07T+qJWlN7qxANYzg6Op9UjbyQU9zIrzYDiT5jvBh
bN0B2wSKOQg7DsEHDhNJv1unuOdrWdyBG4wnlRP5fhceF8+1ijitu7xDthgJ3QdmRDegFfsflukP
Na2P1+Lr8uQpgKsvt1oWhx6fsjgq5HzQY/W8gjmj848BQqVIeYLk3kI8zJooZXq2gtou6zNAe2bs
Ya5fy4uJ6ll+J5WZ7uorTGlbjqU3hpljFGG1xlzp+sGtPuUczgmVjohXR2ZxiOeQz7zsj6902wXn
2OdNO37GfdxmV7xogZDBzQYCGiJRLhwIbde0HXw2nok2FYJeX701L3UcS5BGlM/VO4OZFgA5uq9j
SFvZkE+uIPZJDWP7z/3WHmDZ5AdIKtaTDfk1h68gu2oki6+9K4wrgjqVGFVOoA5L2dEzv0PgkNKN
I3EA2luytHCVeNMuzuGAqEkpKfC42oDLADxaUWa/nrdSIzYBqAeJcZOUTDI3nw9upWtR2ELp57j/
rUvXBdEtB27RN81mInTkQepUugAHlgMi9SqA3RSPanUr6Kh0Cs0xBhlWtnf1GvgwALKTu2wY5K+0
ixw3WOq4xaSpf1fNvwHPd45kDMlgHZ1t9Kab1CHKZehp28SWu1k+HMnAwVKEEfB6kc1omfCjOUS0
tHevhV9u8nC0bh3xpU9QTrAIYLDCI3wB0LQ+1bIkFrX8X3QF39HjxvVxosLdoGS656TdUDQePafr
hRcwFjCSVxOgAs5/OaAhoVlPbyLtFkI387sM96rO+8kW6+ztXtuhjW/bctD9QAyFu327j4M8SMMe
/BiQxn2U6qzzgLoYjmfJKKFGOHp59fM9XPISvLa2cpHB+iqrIVjikAVldOopkIRUnFJAysFgRlji
0fEdp3EbUeDObyabcDY/eaEdrnvypwSxlIIu+3ZBnJtDNk76LoC4LNJBFodOdLtiLyopIuP9j1Ed
k4f4CzZjki5/xGWlAHFoi1H4nlTl3P8SsuGeatfcZW+DYuuVLq3I7gyKuCFrBOlnnKhESr3TsxIf
v96AuVxZaKIBu4WWMIP4zIzFWg23Xz8vFb3sDDg/4w8FcdyYWTM9BD7cWMpCFqp3BHZDOb8LIwAb
qaW0IC6pU4Xyr8DRrvc1+U6v5LHl7lx9IehvdpeSkd0yhHx94yKXeO50O3y7S3fXbFXM2H+sXazk
EvRFdm//jcmDKVrPQA7jPCL3k18zmc2kcqcXe8nNKydrr52Z/CnmAs/A55PwBY01lgmH3A71ZlUJ
V4TTW2Q3a03YYzA4/uS29DWYacefETwIhlp6JQasYdvSbcfxoWK9HNqffi0xiq4AwieimlH/w56+
cyrCzGC5yKdk0YXIkxgF7vs+3JP8J3KcHXJ5A40LuAJF1KVCdGxYj6k7305N5KjdSYPh1G38WSOr
qtoIy641t+2hCLTh659ZvdU+lUNRmKKqdV1gLxXuDWQDv/MS0bcMTPPH60j7huhDWSJ+wro03hFX
2HK7/dnaaSBxL/+N2w4QaQF7qEUWE3rFUC5S8wVDotybFXJP23MN7a9Nndjmkgjp2k0iXdvMApKC
7viBHSDJLdvN2D7H7KVA/nE950fUys4uuU1c7oFRa5g/ve8Jh63QLfkKEfY3OL5i4Jev/E2F8qJB
SR000emNcAOppXHm7+uo1GFZaCh8oI1Sf2HxvEQ+U4340ZGgq7amDx8vE8bAuFKu231XxsijnBu4
FCqPRA79zflYbFjRSjCnR8Fzxf1c75Hkmmr7x/Px6bUDZgeL7Lm7yV31gacDwoqktOw6k3qbSLUH
Mf17nzokHouqcPgl0oHaq2PlfqYHeQ3dZ7ZOZZo+m71iZdZDY7gJ8Y/EpFd7ettysGwigVsPU4F5
EBedxUN/OSPOIKU055zUeDxFHzndo25CUyk0Ubott2GShzzQmBcHlbUzENhjEaFrhr5k2PvUEisD
Ji3t2gP6z+8begXmVygkXXRWPy+FOEhpBgfqmnPqkOS5IZtWbgRc82HW9x+V9+qppzPiesd8rp2P
9hw6sECIm58U476dwlypH9KLl1ibJHPIxc7aG7s1F3T+amFnlC62tW5A+2Jw5muEWfoeqi+fwsbU
k3tJz6yCkinrpwJ8aAsX8ckSDW3p0w5iFQQZyXrXjutTker/xnNaW8FWr7x4HUEyyc9xAz4/h4z8
T7ExbHbtIO2xd+0dvZuH48GjmwyL7rwSkzo6ZlvfXVqnOtAmQJJ3RhvQcg/Vd5BegXQ2PPL3YiMO
C8yNOOVw+Gv4b0rXuNt6nyAibDuVJjODVOAX1YJzYrKZlxhAPynwbbka8HyqTOYUHNrqgX99Mc7H
7ByuAhbDMiP2HzUZTVA8GzuM3t09X5E6fNIUqjMnLWcK/np07ruAK/eNT9SIMHvCH6r/R6kLpmh1
P5IsRe7pM+3274m6T1AKFoY2aQx9po40TU0EKy7+Ma/ROsroPuBFl+PSrqv4q6MzsXptuQx/u2Sn
U2pMl1K7idUKaMDESBrhQ/suFl5c9fyoVSqcKULabICfLXAkqCMIeK57xUd4brjbfm4FBBmQxfW0
vNA0an9Sq/ossvwi44d546AZfxNsqICP9x1wIqhZZzAAEV3FTxDDMvzea+x+iRjJKncMLL7KLwJf
KdwhLhMktEtPqyEdwf/2ihX54SEfyUZmI0KiOHsiSWATkx2yNLDf8xVDnQENBFXJoWH3UKVaZkXs
R6Bnv2RYonYxafkILfO9oRrell9uzd59B36U+RuCxonAhJgEZW8Aps8TIjOvKPLz8R0PQ1jFqZ0O
+xtgsjCrGE2CnNMfXlHnhcTWSWweyqveHWjsQcRdOdrev8wvKqa48Awbj0MgUWIvrnxep3pTZ6k5
O+lC36o+dzVPi9YiNy+kG+ovKYK+7anJ9ODoK1ETnznspV1KTNNX7FfPUpbNMhfnstSTXrvZrOqz
ZZkoHVoBT9BY53bdX6D9WB5cj1LPEMVi2Yzy/hzqfdBPVCZdHeOfaoLzws4P6MmC/1m8VDIvaF+A
l+M4ey78+0SRVdBhOi35bheKDvZAAhCLzre6x2YKQDN/N/c17K0qSf5sBaoWPhtghnkiQ0E+ncjR
GLnqb8p8JBzRef/15qr8rfBcU084KMurtlzxntPuCY0044xq/ymHQi99CoeNezAXy6EWujKi0dSa
dyo8ukVxanHkL+wmAIuJKbvpj97NR8s3NTi/uIDazv0eea0zYEKeEmOpTUV0KySuUydsWs6AODk4
5pGxmivfNKiu1B1DN9P4XsfVpqi5Fyt9XWX96BUCAcCjbEYiw117GOxu5Bktxspi2Ppo+GFC6nSS
ExgBShouf11pTCY3AQA/Q8OnYxHlcgX0ZiUAVUHwOZaTnHxsP3dKE6myHwhg7dNTpMlKi24zGa2W
ebd4CEFyRbjQxVYF89zptF+d8nHWN6SpbcWs+Xch/BbMZpj/lacutRcudDOPmSRhMCp9qbT0O4bO
C4oqlgJjUA4APesDURU+1refyXfi/UwniQnEbPLTp98rjCJv1f1AVSEMWci0xeYnLucOIvzhegPs
MjT7p6Aw+CyGXJ/u6LE42k1YQz/q3bvpx1moeAQHp9RLGhRh27dOrW5nluE3SIHHQUEBmbbDgcAF
6ApltaW4UYf3jVLnoPX2KgXThr1E75AfgaVCW9McQoH3PgTL/iend8YicpX6OzRPwlahq2dLTEFS
TKI7r5zuIgINSkYXDggAPYcfjyAkgA60I+1EVmrluPXDhEJaRY3J9SllBqlf0oKBg7r+6kKpk+Ng
rVAxV3L5RE6WJMRK2wOSSJ7tcyF9s13DpFCnGp6TEZ+ZFSFUrrZ7+Ehm56g+MCIqAvrQn4nRAUHs
964E57TJY9VrXv5KbWGyCFsXBogDWQx4/Cmd6runeqlNqhmfEdQrO3Fg1ajzBdIGlWghKogK4VGB
EQ0zBvnxv3z/XRuMqMxBzrVTw2wgJwtLD0kkFhAcx4mShmetHmL1j9t2hjt2e1iV/NJjd75phFJE
FtadxBmEavsGiKWnyOKgzz1LpeNbdP9MpLK73MkeAKGCjCuG5MH4GArHiadnU/MW0IMzJmqP0YMk
JwPxF1N1ACX4hDntlAa9/gf1EJMmAGGwJBnBcEzf3YhzmkO2ajVmxVvh5GyJFBroO6c2e1sA0IWG
LM8enbT1nzX+AEkT4MTBNUBOgQ0kaGgQSGmSHdaTJyUoT/G+EWnaXTv/kzJJaZ6aE7knn77lj90C
Y79VVJ/pHy+E3OyG9u6n9mP3V1IRItfTcM5BzF+VQZb0aB8W9HLRSxXtvt2m7oL1zPVhcdYSiijW
xzHoawwCrvotooCvLAKNeM4Gy9TvQc9ve7z98T9gFoq2YYYNVEaFuWgKecRd2NI4od9QOA0/mUmk
LJTGAtusBKs9N/wRmeOkouQqHrUuPUDWJebsqAXaSdiZeQOfqrcYQ9JS9iXx890cPeU1dBrYjTCK
5KMb/65vuBV70p6kJILwrmwsg/cxeDUjp4TxzUtpa4GUbR8xucjy38IJ+0H9w7WfJnSZr8Ib9Z3a
ab+6aPY83S77ESTJ3pdpTCJgQBCwPpu9JAXHlJ3dTLTtAid16OHnGsGtEHi3bl5/H28Dq7w4G46y
qknW0KlHEbheyvUD+tgWJNIzKL7+zZcG5FkZdaf18g6rpAUG5pMufvFnXCuqh/oVbiNFcZ6vsTaD
JPr8MDrPDqm99c1wrgzFRvlLzOK+ooS5BYGezi0U481Y01EThRuSbQab/Ld8zxH//K8EsH7kB3B1
LHJvAdiJUkjvJqbIqI9ie6P/VCThVvEzGbsO93jf+q2S27FnYaCoSfBE4K0UFPgRpOkeO3jBQDms
UBMLHSqEF+PivmYvWiDj1XlKa0QNPbW8AKOnaflT7PfSLswVBRfcF/FNcOolmGkx6+PEqFTUI/oK
ZvgBjeO/IMNChMb2tb2ltAqe9rw0IKuGkQoLSQrLR7SFuMDQSnnSzy0i6sHmiDAHrnRn+/zLj45w
ZDC0/XXzerR+Jbde6deUFsOZ/kCmoT+Q0DXVp73h9WbuzHr4JlTu4FoE9KoCI+o+RZaRDPegZM36
qLDada+6C71G2DJ4AsgqW2GzE8RZZdptRu8bdW6mSsnNeoVw2nSsAk26NuCOeAwrGpKXEO49RlVc
PqgWHeD5xWdsiY07+X42TsdAjUwVbzb+sPEm9V/55c0WAB9xALFheme2Y5bhbSXytXB//RWuVx4v
BjE5eGyImgVc2w6zdrDiEUY10hzfVUiSCpH98sYD56I/JAOY1XzIfotZMso6TVAu7C4VjBTJVi+G
d00oYb2FK2+lNDsubDhr9nLNwoBWbLiBrCc5cDcXa7A2/apVATOrElwK5OXAMkCLBv8BY74yVYy5
2JovkwtKMxGbuTejTOcnIeUZ+JjBN95Yhxzpc/32gGPmhy5B+NkDWrpprfDGb1J+ZzF8PNCJa8zB
DmBH9tyMD/TubdtZHTpe1NA+tcLFk8PLJOwB6x5xgZKLN/+flAwNgCbdc1COc0sZXlrIF7LD2ThE
aRCmzgoVoDRM8jIW5Sy+ujK35+8I5Pr8pMiFYUjhs3IYaTfxbSEsJC3VeIxGBgACnUX3JtQFG97a
EuMW0G1cTYdsJOL8KCmt42A2ooRGqcw2AlGK5hQfQHVehpakSZ8MohDgDHaZNhHPNk/tOPAR5YJS
+luDKlZ4I4gO8V6o+43Jqrh0xDSoVlngS4kegfxkTTFa2Q4Yc683nE60fnF6CkQYfoMuC2Aq8f5C
RQesavXSi2YbQHZX7p5NtMHPRw8AOxWyqWs5noTHchqVf31r1e/QQ6eMIJyc4vBbcFXr4F0c9bI5
9bQ79ZQeMgn0mbUBMua2MWCGFLu5qZ9qtIphnSWMpshD+CvoM+pH6WJrqTdNUyCAciDYQeltA0fn
8C8gcR5dfEvKYZneluEzD7a7CAvxYoRTIy2AWRrIxHnL2fsuTLbiWpH6wJF5Kbym2xQ9F27RNjDF
yZ2tOi2tudsm19A/7xbX6noiKLeepLX4e5kx56+T3Q1L7Hpsmn8ak3L/2vylpfwb3z6VmCKiW6sA
1bSP8oNxDcXwwLoBuTLKOTs6kzUnIlABNSYHrIxntGGAiZ8PUJwxntI3eS1WNd/afcAArWTutGzi
msriWJEJsloXxwsXY8M1XH1VplTDcIOrXf2iPSQX1uR0tVLgWr+KzscycgZee9z735K3P+eLyTyn
ZuG2m0IuLECS9GlXqRtkkgypeP1YSXOg/UqmrbOQsQny3BzhopC4HYHwqfHNk9SWTXvT0mwy9vw0
+G5orSCuERwG6HohCHQDoOcGm316yhlHC8kR3pOf6ecDltRHk9egIEokrnLrAunXDF1wYAF9uk14
CipSvT4wdYOnHBQx1ukVfne7LsMwqseM63V3Eww8cAvDTeXF4jy4mDOmxEEnlyHLeLELir3V8+v8
f3hptvF8mUVx6xCvCIaHVTQvc+ylcZN4UPAnZ6H64jgSeMOwTMd23pAshQaVsJkODyzxKwLzX8+r
XVrCUbQl+YamQLcK0gGKZ9LWPavWiQl1wFRyN98BWVPbeMKca4jKkgaXUcVv16S3Vg4WJiS6eUX9
BAa6/Ywe2eQzEEwV1IBAGErxw6Mt3URtZ08LFadHK7fh+GdNClj/O04bzjTHJ2B6/6MMZkk1lo1T
us3Voz/zasaAlpXtHTMpgNgDxM44ozGPdRETWTe+NSLNpKWGJnXfhu6Mf/UuWzhvPckSQlJPJspL
3sVrtk64R9Mh4BhtCpGhrF4bzuA6xrafQJY+XNeciXBVsz+WRiCU0xgcyqHrtU5Z2MuZXXKHumf7
4LfS050ZSUfvqBUAK0/7Y9ZWzf/gj4CjIC4sZ8g7xdYG/WAOI+Rv2EAlNtrYROFFvXwVjp/G45iQ
Uu69IgKuKIDULCDEOu9pcPTlGcyr7gFa5fnHhtAJ9cS999jCm/XNNNC/T+xbWBwAvW+VLIUlIJZV
zJdig7GiEfMUF+/06BUOX1gv21aYp4rd02vXXiM0Vz4ncatSGzX0uGDefmnPlXW26KgJK4+8pQsX
azgV2O4qXFyWruHP0U5Su6oFwwVPq1fJleJ02IWxblXJzeq9qgr4EilV4ZXClr/9MfaAX4dRH79e
QrL/WpjiA+iKXrtbeg4YlfPhvIrc3zqCgpe+Mwi5ma9NHfw2juQurWla2x7zI5uIww0WvD5p5ESK
cckS491LT5Th2iDanDhaCsKc8+ECpbqXTr2vIEKB5Q598zgVKoUQDGho4PYHoSV3BT/GhpWjgIs/
a5sTlfZ8N9Mtt2VVF68395FrVIctVURKN5RCYPWGepqBOrIWfmJhAcREeeapdZicS52zwBghSsP9
0ULGeqWBgSWFpk92UKUgbBkOXkqEWz9PJEd/cCRsPM5SdFSBjXn1BUBO4GrOYD0i4mIQZDH90by+
DvpbiPc3NMOvgLnBy/C2k4jDgmbJ9T0Gvn2sObJGH8pcg+v5w+gT0jJXpqIkvcl3r2UtVk2+UiF7
uenKYKyY5M5YesvYKJkLXy8GAnxe6WGdnhG84SqW9AaET9lsV/XnyKcCLuBqeltK4xJY5xYeLEc0
wBVvXDE6sdNgbE5g24DgBGbBtPVotp0ET0fxiDfzEqcID/HwL2S8VYbiP68nP1x4jdZzPlB7VWBf
r5R2byr7kiqmGOht4eA0CJ1UvUR2eHk0n8LuoBbvd/Oqy1LHV8vnmM049kL3LhHy7Nd4l2QXQxRY
AxvptbS69VeK7E9QogkMRu8OQ3dxwXkBpYM9+UkcG1xUhTzomEj2Wf/bmFLH5uphbaz5DEN6c2VK
mdnWeTn/A8mTBY81SIyIg0fw2V5Rjc4TKWTO/21FW6yeXGZWnxU2SPaEZJHHehY6pAEhed8X/Ohv
BMkVLxT+UFv70JN298K8HK858xpKA7Xjc9Oi3m6R5ggrcrAYPp7cX/i/9Pf8YltpLwcvpOaKfKBh
BK4X2PKr2KFO02CHrS+dU9j+6Uiol/fnoSUr1Qg2fNAryEeNdO8fD3KqqHbsgiAN74zL2iP+KsN0
qL4tGD5jP+Yv6BPNpm3r2GDyUTGG5BPu4UQBQTvE9/ELS1EIcdp9/mgsFrLDiCu79WL2LEHGKOmf
K/fI9oZg+O7OyrEP74sHWGbGp1FlAlLCjwYsynuYlFMUiPkzJp0hZN/7HrmQNVTOaau6MwhiBFPn
Plv7v5x8V8d0afFBhn0Moc3vXfzQ6p3KLmUryLtZfs5iPPWiW312pAaNRigSWUXhd29A/iUwuAeH
Bf61d3DtGtblmmLyfXgJw+Ogm159AtrmC2qhPkzGdShmuLD2abgPhlifIr5U19ySB18M3y9E6oJj
ETHmZi6BcDwsla9l8rMcwCykZVkSEaUknLEG7Akx6sZhzVKJdzoNqcH7Kvj7H7q956uJQ/UR63vm
LJcdj2tjUug6z5cn6BqxgPnFGAI503SXqczdsVPwo62z4KVVKdRacxSZxBUbqW4SiSnz5FOf8Cx1
yQK2nOAbNn05WZgoSQo/oz7mcGkmtLJ57cLQmEPIHf3pjeEp3yoO6iPhiwiNWrODyNWu/5PIxf+5
/SYsQ46OxgT9SPix+edP7v4pxCbDkgcQWRtfJmxNgTPAU1wZs4mF+tHqs8zPJfuV0aVHux6pbxcq
88w1BqN/iR37pfE88ktHARV6O4Kj42AjAVqgVjVbQZMQ1WgTmII3Bn6QFM4E/6PRloMTxMLkD/T0
ACu5s56LBpVuWDlHQMPmXtP8D/rkaHRYAqLNPmhCIvBN69aspoQyZ3vohFGHsKerkSoupv+Bwti0
t0rZJFR+/9Jr1h3Ria/ATHKOAGlC2f0v/8mCG2Vrs7VbskpdEtMv6IGpjVAkDHuF4AfgrIwDbt6h
V9giFv259IGE92pTVyRNIB4aLz5W9bL47wuiEUgDfwErWtKbNeH2PYDN/ks5rXNxfLtJV+0Aa9oM
VZlMUGRZpp3d2O5++vBndoRZZZ4ywIUkaG9ATfMo4O04mwAxvzdpizRtMp2FYf7NENLFNEtBnRfw
5VVvVhDGNaS8+dFigwuvUdJzOriA5Yt7mn4hOdEUwLuHrYsUgOW0Ot2cy2MLgcYI9U0YNT95nUai
ZJGZIbCXJbETcAA/aYel67r0mY/276w0nQQqXPjod6XtMKLJKMasCuu784V46vYOND5UGeByJ06D
3+iAVxyiLiXqubGonyZA3wRvkIiJk50nveFHleSUUfSrQ0zYo/+jiFS6TpHo+JI7d2e4249AIRgs
MTaDYhmYBBwlRK1ZgvQaI3rBVyfu17QOvqUM+F3l2ly5+XRHgJOO0skdLOFwn55UTNN7ALR86kud
TqzvR7NgxNrij6xwJjAavYI8Sy9PwGlANd6o53B73iOfLC9rJQWzkaIF0knYbgtugRvgLzSlyYgF
wgzRqfUTz88tiEg/ZTo8pJr1ziEIewfnsh6HkFX/FcqVyz4Z2szlw9kqBctXcy4CMbr7E/fCxfJ9
H2DRdXUOCysPhUSO1JKi1zXW+VG6DPPCit537m4nIq92gHWL4lQGJ81cMS6pIco9vjJ/HsasXRjO
wgC5iQTAdhcZgFpjya0dQRtqU/Sn6XdixtvftNZPfYSAZIJj+vMNCm9af8vwoSu9iJ9aQ/Q3kiBl
LKMPbmXOckgOE7wF+f8o1XsX4os2KNIpP7RUe2j1P2DWtpYyVmUy6X7Xi1+AERsFtVIyZ+8lQL4d
PfG9tJcXd5PE/NF4+dd1yPYVM8OK9hJCQAwQnw/9SRRKwMDCTE9RtaXNSiG2yE6lOxaiie0tddvC
S6fOltjeyFY5ngNafvpaYmY6Ok0aVHk9DVuSH99kegScWDKnpEkfrv7D7ezeTYsZjSeOAyI8x9Am
L1+eZYITgQ+SiLs7DsPtuSKHqfvwNbc/lD7V87si0VrIe2ei7SJwZQJPnsm1zyDYLCinbqBcXUnk
iN6S3eFq5v0mvIpJ5Rx6p8Oh8bwNaYzskyw8MTqt/YUGHFcS7q/gcIhe3YYBpXl2DZGjl/b3itmR
HrBKbrzxLWp9nrVxqw7hGY8Jh+G/Gym7is1zzoNomf5Sd3qw9euwxzLHMdplS+5o0TrDLD0liL1p
ZuMIYMLXn3LupkaMCss3TGATLJEOKdO3mpc+tWRLhn7v9EgOHJJ3Ufid/1Nzf91SS4Rl0+VjDh+W
TdaBlzYmMq2eCZCcgHWZsWUPVLUmX3kBYfQBjMtRIVwBahBaqAtk1p5TWFR3YezFzD429KGo2rdt
KKfWCgQMw/ZnNQ0ByzWHtNVmCXihBhzr6gZfB4hL4H1EfmtBYOs9OPRExWCm7QAYk4N885qQc2i/
0h7YLW4tWGN/awGWXtbLB0M7D8XVmz7ojzGBXk2G5WZd+UCCPDMIIuHm6RLJ14AxbVH8xKSVY78I
NXvYBErYCRS4Tctz1i9hCpiMNVH0CL1PBpZrTsaTDXf8yZNqbvPBTY0GzvtFMOs7XDPwdwOQBpbp
gez3g/nVxToEcprAAsXVne/A8KGWXp6+WIzroxnmzjFGXRMwTEwjS5Jfj1ME27eIkqZNGbAOLP3l
grH3vpH8NocK2c/4451DtjsvCXL+0SBBMwA8iyBbqoCL9uKnA88bFDKCUKSPWyOWTVlck05wMsdK
6tR3jxxU+wxcBPoouSYENFNgvdJINQ5/fPflBbnE+8m8IRRGUNbyIADbMrcMx4h1ayNtRTGOHi1j
6KT/Laimykuy38GhazPZhHLYNIjS6aI5x0bcgJRarRFfyRsQOS4OTpzq8dgVUmS4XaK4cjIgaksg
noQFF0sp6D2QhBLmTmTQvQAc96JodxJPxWDjgipwpIrBQDZZ6pgO1NWZ3/2bl6DNA+bJ8DEaR4Cy
wiYjBk0P8sUiILjQUlcdLg6f90B1pJ8KkBcs0ui82me3bR+eDxXsg6eusPNKoenP+nWIoQsnZDQl
R2K8EMYr+QNLVCDdDuqh/62GT1MduLoFP0Ujp9xBCHWGVaLUMrkZuNFJgS1Zw6hWjgvw/MfTtvey
48hppGp3jZ7SD7+5pKR73VoRLimXil3TB71OXQDVOBxN3mk7kYp+sBBxZWYzmtxHd6cjVOmxjiRg
0Mn9U9ph1U0SD2kY0gWI3gi/JZDG8Woo+3bSN9Y8oaxZ8Ex+9aCbtb8rkSNK+cw1750KVemQWMSo
g3NY218uTsksaXYdOXYkaKUsx8SOH5bczn+htkyvF67wX8zNM2wlPN4m4YctgKkEr2iehr7FOC5B
Qrnx1PXJ1cfYgo78UWBmTvKI7Mr1cibeNoPc3y/nTg19AgwYh3a02Lt+3dhGLyPv7h1oneTJwleZ
CNSoc4XnVzduo8gzQvSCqf8hi1wq4AA/sQERqlxdjSoZ93jP8nOG6BCcA5TjvYh4JGcq6S0WQmI2
sswODwUChn/FRJJkKCzItRgffr/TbJrcKLWQM9910mv9v7B0Z2dZm4Juws8hbYFIiDHE/6FGiZGS
9kdoTsuDGuY/zzqanXjaXkf8D/ZCCNvm5L3Y9XLTz6eRR/nQoznzexlVA8stz384Ok6zG3A0MogN
yGFEytachQOCw2werBkpYJJer9CcHPdlGsALaicVIubz/b6adqIeHkIZum2PUsT1ik3AZKgzlTf3
ZUZgGjC5BLoDifw7e//aOFLQrP/qdX67jYzD0T5/yvhPjxvKdmqRfUK6K7FnBmadp3jYGpuq31lQ
NapPXvk03lmjmEqlhaMN+BubuEy/DcFkYOWUyuEjfwac5PZy29Dq5xMtadJ8rBxv7gJ1fMLgD2V+
VVGK98qH5P+VSv/+5J9j88oJTU2SymI4l5OXE6KehVYEc1nwMVKWNgJPwaHPuRQ05aUdeSmCphOj
cufVREKEfla+26uYQXZNCDEe+sELcNeJHxTc9mBBgdRUlIQapPhMUujanB8/hsnnoPFIjk/NHQpB
VJa0/sMEOXbaVAmnXQYab+b0KcFx8YG8jBRujCo4qLOXwZNESjdhvahRupmAUX07X5WHXjZY4pGf
KRGQVMbQsJ+FFDuqhylh1+6F2Lm1Mf4+vxg0fbvfC7WLOnHb0NJ3ZdBnOGTvBplm0ydH1NaBdxNx
Au9I2vn7WDfWUeMJwAvVFuCAdQIOmVC9gB5luYvuM8H5F/Dvqygp4X0RpItSBXBXzp0xBC2PScpg
8cnbQX6pEkmVCEVhQ9Vn+kfgh1rzKGmm/VXkrzN6hqii2EEPHzlvCFkJ50gHHcoWIWkPOeR9pYht
Oar+vSWpZKw4udsCIZR73zk1axZo2xYgtymRbzQTgeRXMqi57lzlt57vCTT4oJBzItnImymYba6c
90pbp9gcoe+OEqXNk6aUOkcPkuXESEkXWcf+ozk1y2nAMjTjPG6Kv218L+ZnDYIkT7Kgeq48XlLq
gzcWscYEToI3PrXJs5HxPDgUon70KhnuKN1Owu+ymnNCLB7rlqllqy5dbPy2PWmWq/AKwSRS5PDE
iCTqMGe71JSiVLgR+wwNXJ9PXhbFVvSY4aABmPk6wSdUuEvNlnN4wKaFRCcWM5t78Gs1RSQkILMi
tM64rPhdn7SWNr+7bGGRX5X4GtKzfyWw0A0vftwwUD57fWLEL/hFQrPCeo7mKr+7UAnEHyJqrQep
DuC2BLpcpKd85JSYgk8toCTWPKEsfCq7JHoORLjG8G/KKOUa7Y0E1TYWzzhsGxt3gYMNhaxfE1w2
KE3B/8m5AgVZLTrG9FFRb6FpZO7MINM4wG0vP/EYRKDTkIMNQqxNy3P44zI8anTErvuGcaMDd5r4
Jo6pUHX4kL1d3BPPAPEsKzRqd5K6rt1KRc2968lgJp9kfBluSEYthoOXwFseSYJIdU8zK+gnjpT4
0jSxg2vqYcEWuVKIFc9L7iZ3B67nuQWpd9m3GLvIjOVtk5QWW+FrgxH/4qa6aW0wkZ7zPtqL8Wxy
VBlKp7xVitoYu5I3epLVO/p+rTKzw7Coa469lLBlcKfK/8Ay9FReFi2DiINWh2DZE5st+ilOuWqq
fvU1havWWk2KBWNL5//LEkuWY+sQ40jlG4OdFaO2TZ/Ha2BQkmf0YwsO2YtitjFakskncGVlt5cR
N28lZaUPJAxfWdUoYJoNfnpwZGvjOOby/5IQK1162dAX8yeRxEDolPqknBA/O8gaQBdQjc2mG8g1
nPZiAybD2R1Vm2NFMtM7vBWSehGdJnKwetDssDBEkC/yusRo4/J0ETr6E71nNzcOsgdSWrREPvAH
tx0IRNfhNC89hOdWN7ManMZZGttKEYpLeVYKIt6C5RtKCE1Tw5RcyWZEWf6qknHozIom6PlXfSWU
qLyoou47sDjzls2IlTOAzIVsAFjYNaLgthZPB/81iQ2IrJ10aPijrAJkGXzxy7alqzupdxFougLy
QCwzredjDp132TTBZG043x8sknDnU1VNnFzXU4CTNvA0T4IuQsnbLpnQZRYxHmmQnadg5kNQj5l7
Yk72UE94BO4MWGoKgAgFMdZmBvjWjM0aSFuKxtaDy2H2QjHFDV3R7Fb3Jp8jnC+Jin2tWVhhpQ41
zmg5CJUN/XqlfXLYwFukzyGZP0k/lB39K/RT7QG/nfbYw7rF3LiaGR6J1wSpuVaeK1Q9ts/0vTuS
cJSsdalbnr8E5Y9Q+4GET1PQI6Ww3UGNJHpC9zb7jSyaIQBhiO8ZCpiPiO+7XpOY6eM8ZDZQFlt/
XMx/pG7SX2ZCwbQIxbFA+dUj2cDZxZcEQnyB89IOvmzCKn4UpFqbJO1KXH+R6CICs/bO30N4Ohn9
6XCz/RfVh3viJsI7isVH5BGU516a5CW+1MMJiRnmsB7bww5TIh9A2wRqXnM+VaR6gkgSGzpk3/xR
IJGS6grnVdK77/kaPYPHb17BG2iPZK/Pvh5rPxpLrQvtg0Je+7bCWOViY8EAIteNOTawompe1oCZ
3lGxNFBd5Q/v7zf+xy+rx00BSsMhcSRxm02U7MNhKlvAKP3jBL3/SMsBuLGnDNXvxKm3+mXKbDG+
gf4wot122DufzjsY6ZIf5+b0Vr4v2jMShscYHELAIfYDOkSqKDIEdxShN+QUjVcA7fQ8Sq1InsVs
3fE+0fpnFfdjLvud33kqxc5Yf47jSS21JFnmTRdXFdGrAdY+Z12dvFProF7yrBrOOHg5vlNlPDy9
knH5r2Jlv9VFtkX4i9C/Rkxp5LUyLuSnzuDmPBgo/7yB3j1p2FAtKEGQZd/053S9DKG7IbJMhwIt
b01dcmbs99jG+0KTYere4VYa5w0jxuiQ+P5CK8Vv+ajd3l8iuynksyspj4Hp86NWXLzfB3wiMlnk
4b6RvayU1mL1USxluvBjuAJzgW1+nSUmoS4pcL1uBKMUl38Pd8bf1zj1QW6UMP1W7v1gQZ8s9Hr4
0QoCcaSIu8tayyOhezOnLM6GCTUBBybwmvdasZXuOkqCOrsZWe2NapOvL48/hisSR6NwhrYYpjJO
+UU1cmoThGUn0xhhlgP97ffLUmT9spP36tgpKwwxDHp5pCBqxotr+tS0e0YPivMGrBnyUIpAxEyl
/1XVxgSNFOZ9vEf/GCv1jM/FNztmKhKCb9l60zRUCeNvmFXVTWXOue3Yhzwix8uFfNoH5wrISMWF
OqIzW7m0Rrc9q+HESFe5LaqCv+9PglxaxBnprwDV64ONhUxsT3vEQNJ6wHEoxCN5kcj4XPbgukOj
euCsk6n6jSD2hxtD/5oq3T6zg3GzFHNLZY+9ucsoELcM7SsR7aSxEVZDYhK9u+8O7aVRC4fFx98P
6Oc9edyJ5+lBWtwLw7sU/ohoQcgVGj2hdd1m8C6QYV8C9nrA7BEGu0o0TPDSOuvTdGnFC2/vHuGu
4y9YMoWeQkftyYPhq3GIQ/dVDwAoeaLIPIUY6ZCm113H9LRoVjwOPljDSx6Htv9kP/JFeN703Bg5
AUv3r0GgNKAFEQsGZdPv6U/at3iuGxRsfs8sZsHX0ESaC3ZhkuhgUFo6ECqQqqDZypQr7K1foK7w
kuk8pscVXR+SRXmFoHksEbFoCUMyVyL+UZGz60jCBCTyBpKsuePa0+SazcEfzxassUQDtVh95ygU
PW2lt3nOkrkZKkTKUxGJlsC5L8BrHxdf91baTFilaKUImdCR0lrIUlNG6IKkHRwJsDQ9PyPL6tdV
7xGwZ9hL7pol8mol7G3+sGG1+Q+EhiWoqLfuLLhfcKaDRqsxay/ZxU3PX7lu+F3ml/XwIQnDmccY
F+9Vk9vE9l05M8qpX1nYGQqlmqNxVUx46owD0kIpFSVuMG04lDv477qPuplzWgIKggjTX9Tnnngr
/JiMmwlRKK0xYeMQmRBKuu1BGcyOCZcMHa+vIResjTS8sWbkhXdzKJ85Hlot/wIKV6poBMHAASg/
iibu8vcieej9fkn+VvLKLJrb4MNir4fDC3j27NjEebXp2LT6+bhvTM44ZRZwrWOad7RkRiybyWKo
6oHU4zaRRuYbC+X1qvJ2DMhtyRghuwXLkrvNDT851akgp7CDg3BXOgDlKH3SRR8FC8FtTQ4tWVNR
zf+VvIpNeWw40sR9Vg7P3y32wQqw948n31t/hmRQGi6uu0Jsc9+Z38UzuVuwyUMpa/qZy3A9B/L3
11ksCAFiZzo7HGdakUKmFi/euoglK6XV9zEGWpcyRVFr2nq2oENBAfg2vzxXbaeltImaMgfq0Bja
12BXEIqq7G0K3wIZmVRpw+NADPAYby+CAaWZiGulaeCNl0K8HbyoozmineGfB/r024R409k7sljx
WtfJwA+95+/7NUqtVNx1fjPmvhUjcKlZjwbHdlydaK4ONdEdININm2v32UyXLwWDy6DmCavOeYu4
4/M6a9nl2u2/pKjg5K0pMim6gSe9qtaoPliGPsHFrYC8winQxE47FqfymecXoQJBgp4BuvLsPuvi
nK1M6IqslHYBPNvAaz2LS8gu3ldo38GxyXCmzjVjpTwKBG/F5WPcx0Dcfrbk2HTTvOMHhGzmT1Wz
2Gm9K2EjDpqZqi0I8jVNrgXvXvSlJEdihNdB6AI0H0TXqntLJxQ4HMag+BjJ6UuBbvZBzoUdh9V0
feZQO1GgP3wqe65h1dtkTXmRnx0iG2CRPM9pp6dZ662Ohqg2kPATiM9+iAEtNIgopq5sXBn7u+WQ
0ITPXt5XQpE5bTQYAMFs2GUmLYM95SkSB5YWfdv/EQ76zJ6FF0CF6nkeqtPRIpy9fAjIbV4IQlxy
bXILRUMcchmz3mfs3exGzUt695NJBxShBKmdrcVENrgtugwgu4N0OMpTc9AHC3+zJlWO5a4gp1Zt
arFdSIYO2AuwHBSqAqwNQur7Ebnt7BpGAXn+y0qB1mA5ntAZOi4cUK+t0tQSKmY3Ql1TOJx3zi90
EK/Xm22WpoAVcDyD6xi395Xb5/djtH7zRt8CS8yDiDWqheTHDFr1vYGLtqxJBvB+uLpHvax1qIFy
VBJGC4tVH4PH4k3SPt56CWgM8Ld4D6/+qLW6ZrcQICDYvz2/H5/V4pdSEsiHr2J+EzWP5Pir5OLM
y5gk+YLeignDAPDopjPaw42/n3oO24QvDbEQ43FVV2G4RAZcyk7/Zn0L7GsMnWM1fjKV2yKD+UzM
1PgjOxE7Ua2ov/N5S8Kn5EsmndyWh+5Fg0YKxDkSBeeOt4+Zinel8S52vPnalIxhBeQgRiaRjDi1
dwOe3g34AAAeZJtYrBF/Ud4yNo9uHO0e3s3WC4upqccviWBJn9i6hjpkavE2YEnpBECpIoP3OAJ1
EaxgqLZGGpOBnriSi247GahJ+qijShDoIsQVhdZQv7hMuLUd9tZGZGvDGtyYwR7knKoC//HwaPXq
AsJndol/2Q9miyhWxraXpHgQ+yFXNExckPmMPmpO9hXMZxQG2UlCk5j4OD5twneK6m+bm5c5dWfo
sVpjXeGpvRzAuCad9nU9/1sgKzkEeYFOzlwcclZscBQ9VrVnI3idV1P4ndm2fuR5fC583ZWqpCMo
qQmzKQp3QXZoDaX8MTixL3tPJeXnu/gh1aAtbrZDpvBQpXbW7Ni9M3RCIUarkorHYvbXBQ0j2/4w
R5+jG1c4BhU7yC1CcUwAZm1hec76Tj9W0iJLiyY2xmSc+hTLNmK+ITTp79sXfHzlH2fBPTtokdFl
mgvONatTCfsuIcagBWhW6wgrO4aQtN9o8DchW0HgL5lW30kZshpp4mf4tBSGVI/aIhQfVkUQitCI
9E/GCi2ZwnSyAJgnXPqIWVHh/HlL2qOADqvXsdXmLkF1VRTDYLlwLBTglI5y1OHJibfkjM6IZHOQ
RE8Y4IZb/+2Y1WAotUst+nMQFwISZmNDMCBczvVhYG9aCRO8Nw4PUgCvv+X71JlN28JWCfcpZdls
HNoEX5KXctyuH41yXSIHgpqUboWnlW9JJ+LwUHnT+18n8z2HKhabUeFIoTT876BxYYl+0/Dg6dXS
c796XrE6lyZ95b/4Nu32XfIKOuGzINzNkWECvnYexBUJdCW/KBAwvsT4Dq/Q7TO73L85WNPr90Ho
v9xK3kjfq51KUDMP0aYKeXLdXZbrbmROTgevVDMzlar27/32EN4ncDCJqN8w6Sp9i8eVwRloWPsO
ZUjY780JsDDcQNO74awQC2cSbq1uzrXWE++KzKwJVLiEBb3CgEhKWwila5Ti4z0Anll/1k31smoR
8c0xDxn87eeVcIDg7XySTVf68qk8lU9uRW8r0ktsgAHtuQU1o2343ej/camWdMc+4dtXnmNhEyiw
2yn8j5JmZKnhlTd0fqdnrZXoBJIfVzobDo54yOyXzdgf3ihJ2Xmn419bhKlqOt6TP8GYiV9V/1om
M7dd5t2oQk0hvLajRbvwPTdNYg6fXAV4QCWzbJeYky9sWw9QVkTjOhPxCkumEL7gPH0Xzh9K4bbU
6pkrDxcdqpIEtq70GqA4dPLzc+DqL0qTDHrE/+hc8h9x2PwUi55vg+BRM5ecA866orzyhAPsv9Zl
SSTdm0AROr4Qd2QrWUsONK6E9ezW8I/oj+urcN3J216Jrzba7Bd3iLEpTg3ubly76x8S74rtiB9D
sYxxuqrUTumKbptHdLAvhz64TB1HuVUhLGVeoZdbhK2QUKzJK1iIURF1bp/CGWrRvAbsZS4GN7C5
zi5buvVeLQujEsrsZbrIHA2VRb/6Cu9w3sJ8mGkdy2u/5pImA7MCMq3mhCJswWxiAuUblN33Ckii
82/uW1jQSLlwcPJ+lWGNVcZiiu4RrvT23HkWbMdKifxdl/R0ez4zVGO/z/48W71RtwNf7iMz6RM/
DAXK3PHpN0kEATqNZRTlMKB6uIr0lYdde3vYw2C5u8xaeLEuQohiPGEQ7Ly/ZuE0qZMYgKVabhKU
x11feFXFQxeuB+dYHy1SPU4JEyX33Iqyn1MNjmgaPeMjdnswPlj/GcZR01H9NjO0r2xjOZl8TCDT
8kTMC4NPhMc0FMgOUg2Z9yR6ka9qIqqkYFkHRagonprCbem3XRlY/LWvBsQlaWRvjO39exhiZ7Ll
O3wup+eL2J+3MJcGRZdhfn3mKYfli7PVEMexh8ea2NPIQngqR5fUzroVCaGIMII4HfJjadBquBjY
7rqbQ85XmywaFFcF/ea93tXvj+4YHtSsns/mmNgLs8WoX9isDmL7nGdQEbFQLCfbOC667++blRlr
IyN2/vRGMy085ayhE4KHUJXVGbFP97w2A2Ai0zFpOlKVPKUymB10+8+W8dAicVjsHJVzNoq7meJ4
j3WF2t9l8KgUQLdc0R5hS0RAez3z3XfPqkXogMZaAemSS9qQSrcIsvs1bp2LSCplzltH2usH3W37
HKQiD6R49DqSMHYnyjLGIRYTUnhI8qgL/a8IMToqcQRz9FFJJsXA6/SWSlshkzyE7gjPtkpsQtqS
R4D5mGZbExSUtAKl/UcUw+q8igBtrbc45krho0OyjKn9tc95Rhxrvg0JZRhPX7ygnXgbLIT0YER3
WcEO/Z7zH4qDlNrRW4+4ut+uvbt0Hu22i46zLzRWiZLaSRRJ42sv6u6WdLj6bzp0AD7BbfWmfD43
LhCOJ9H4XCLw01y8rPW5UGlgFpPMZWOkaRNVrZWgwt+HI97VCd/UZnH19I4aubC2Nes0wCkVrpJu
zdEXOnpU5MqIOgDsLP+Vhw9XHpU8BqITFWQ3BpyzQSitXXNRcss6paFSiogUsqzL7/Iuoz0jY6SC
sR2mZ8/I031bpO1B1rqHad96IxNP5VZmSvRjn+4lB4Za5+GSHZY5MVI1NAg/UclOxB2PCyaeREEX
AJfeiWrXF7pOjP1Ve+g1+AznxCjbTuFABaAmIK9o8uq0I4AXrQ2yqE8t5ZE4Fvjn3DpDrLW6r5Cz
fMfvebs2/mEpzmFKot+N/qyS2mJKBlKfOEzdb41FzTR5t/xQlp9vdWI8UwRRw4AEQQOMNoBfVgKY
0ZnWnV+8+ZyXM1tyhKbnwo6NurQU5ycFMqqOmbphdVUDaezrZsZmQ4e1bGtu5vCeLMbG7SQIad9h
ecovHaE+fNG9xHyt4nbCXei+ty+OnilkSXVaYadjlXt7zNEIcMD7YWiHbasVaLrkt3QJhcxwecj/
PSkGm3YTQNYfiAvSghcJ1hcoxDvxIRvMc9UBbDBABAxY2IO6d9n0Fu7ditzmEczv6FDDIOfr4aF2
g9BakqGFPR3Sy75pvUmp+qvmkborblSH67uEU7jHAA8yRZPm7cdr9qbKubrEosYkorCvnGLNIngI
70C1DbGBz+9PatKrF1va/hK2778vmTPoAZ4u+aNmsifN1BWwt7AdGVG1ltnt5O6OaRLP0iZ/r9DO
LU9zb9paESWXmCnlFo00SqXTnH0VxYxmzsdMkV1Scl2XfJ8b7eQrDeytTtv8Q9ww7dfILhN39Get
JrryVZDr7rvXNH7/WNl0AUbnlX6ftPegOdqLlB4+/INlkEtCK7oY5j9NZtHznelbw9xkWi3dZ9Ny
XTCORvF9SO7gGA8V9xdFaaH4aQP+PARosZQ6qaSwvWUkkEFTZshBwTjkcwh6oUEac0QQVl7Yz8Qw
4tvN/FPEvQG8oLwSFldSCjrWeKafQkdonuJlGvIZrtBVu2/G3yOK9CibUmKMTaXNCwKv+s5XSDg6
rJC7lgXUrCneuUVnbMjPr2pIiwB/oivDYnX1zyxV26yjS8WOYwWbYUMIboVVd0hGEtnkS8W12y1K
pVXVN2eDSsyo2cDtQOG4Buepw3rETYAABrHsyho1mDQqaQ8RC8LDAY1A1CcXNzTrXx4Hxvc3d0T0
aQSnl6Q0RLcIY4cQEtG+aQt4KlbFY4HYMzfPRqeTVKcTKqdFf7v8IluEDM0tU7EZoui77QhMqGvS
ndeZ1+d2gDAsLhLzr9wflro4In3ZzV1KLfwVThG1I3lNPbjBh0pK8xenw/Ht3vx+UgMb5ez/55dk
DyutImv8oJF9+zPtxackYLjSZ/A12ICmpSF1/G7ehn730au9mGsrmrOPbr9/S+SnEyhH5A889SFv
4Q6Yx9D3B1hN/5TEdPcuf2TFKldw1BsNwMXobnoWZVN7jk7SzbYB43mMISTp3Ni13YLTfbAWftgK
bSFaAH+/F+9HJV0NVcAMbHGjbswYA3BmdMxQ0LbeNdJYn88XzzM8ZzYMaX++Oid6ap6S9d6rlcsd
g+Zgk98bn8S0Ni+hP1/bnRSR96JELfxLpA+4eWysOp2/vqtk/CMNkJFZD9aK7EpgGjbQl+ekN4to
i8d0IkfOfRpMjyfOVIduk+ERRWOcDkyLtXPNRxu9hIqNYMOQx9jfQn6czIdI4xlGfPlKcVJb8x7b
7vDFmd7KqXol1VUPnXMQvrHBLJoFPGDXErXCPgSS0uMNIsZJK0Nl4BQRY4LlS94mPLQqPF7uHHOE
tvSlmlUuo9dcjQx6THGyyt6uo2+Be6gr5rpnYokP6LdrPhNHapapkjQemuJW6ZeiOxvilE3r5mY8
yuBnMtZaoH0W4Hb14cR1sER9855JnF801yr4hXccXf1NmTVo0Qwv8lf3jIkm+EBpuRbSbvpTxI1F
1FdltC7PH5uOeCoU+uR7y2IE9LI/4ZTY5IQY1ZtZvWA9S1LQcDyG5UsupnfRm9gP9iDRc/hV4Ffc
95lS4WFXqChQQgOzuVGB3RK1jPcrXQ/4N3S8w3/3qoDDxU9l6eXsJFOdHTmRpnh8sPbq5eEpZJzu
9btU/k41lsjSOu57Vv8w2gIcBpWwlC72t0b+OFCsIJzOQezvb4ZOHi/aIkeXCnXxkm9+PWrHYYRl
Ah2a7JK8gg6Lhr1FiMf7tOnGAXUnKxfhQjksxCoJniyRRasIclRyAVXEZEDtRbv0ZI8t7owmpAl+
/HvSAjDl8UtKn2xLXHYhJmNhGVxa99/92I1YWii/IvneasQ8q3Eiyc6kIC6b3ZhxjAsMgrdi+p49
f3PRWSaBPfEEoQzTI6xPWWjArn77ybfwJMbYN8UGPPcwxpdLkS9urq+k/ak/6gQfJFPIypJvZ0la
4751Y3niuTobSMjshdt3CYDRtzrNPNRIwsd7zRb6YGt2nsTS7k9C/R/+pe96Bh9RbwisQ+aTqQKN
jCVbP0zumBRQTjVzOySbbaZ8X41P9v8hrR7cpsPEB/EKMH/wuyxK+8jMI5lMm11ZnRln2QCiiw4l
ygDA7+xWmZaVzm9GuCPKZBKMGrEnycQ6kY+pfOIu0k4j0XOY0T0f4AcTYR9wbTKaY0QX/2N8JD0c
iFSbRxuq1+yifFsz/Yq1Rc8B5NsDYJtFQ0pJMEurAaBIJzyjIK547sVW+7ocvsuKsG7Hd6s7vrzw
6IcnQP59svtGOTfS46TldLpw3H4JsMp213+aMklWICUmXEFcsjkVSdbftLdZaDf9KGc7MnonlTeK
cAgRuaWyQRPyQzQBfLoEy2Q/23eUBVyepI4hs9SbLMQAaaESD7ZTsNfCC3TDtCzU+FMUvNMWEQRV
+4qx3T/3CchTILoGcv/wNCViL/+GXCit2Yn7H8jlSTwM+RQ6QXZAFfNUCXbpwWvYx0WMWMpUxV6O
KCurUyJhqpNS7E6OK47+xeSZf2VKdm6n755BUIOlnhjLAKc3yt5HuuKHvWgpN1re/S80Eivh9uKj
y89Lh+YdewmTOzxMAYpOuhWzT+UZnTdWqtgKF4ouLKXCykHRseIp5l6sJVYPJgQRqZA3j+f1WetL
xYQ46xa5zN8oirNz3ldHzbYnSs+4ogGtYWeh12YV+u7hXuT9zRQFa10+ZikrAyRmeCjJFBRV8K1L
bUSZ/2VmDJmm0Ld6iDGzb0Gf2OVwzvRXW4NxIrPjB0y+0H8qBhLTBAmjtLCRrWHlhgQMP9p1Aqq2
QiMh/C9mkzmujwFEC+EG4MGoOdpvwSETe55MCUcX5XTTT7eTIpsdpH4Ky5VdZ26LHjre87W1i51E
VlL1ALUAjkcTBfX6jv7bGdNFRkftmQ5sJ44RGTQuS+yhfVLGwgq54/HbLeN2kus8zHx080XTE4BV
LZMzgKSgIPzvNy4L1QUxO+jQOxEd+RoQo2GFc44wrg+xppWQKPaVjvDW1toeCyeS8EkRyqtbYhxA
z19cHKKNDnMUoG9S2GSf97a0lhzYYTHO4cDz6JrKDNp7rP1drkatDnwNaFpUt9XM7oQZeubh6uOu
C//zUDZfq4a1Ca6s+LuNRoO845hEFME4DLNrliJT7Xj3iF0T5SZMKByw3wzlHvy/ErgC+8VhNt2P
JhPMJxqS3n19UUnCRAUkNS3eYDW1SD3ynaSpXBRSGO5RVo4G0NhH0YPmmFCmXSyByGy4z10pAXpn
aa2shLmeL2MeEt+nBi5uRJpc6wfei6ENcHvBaqcoJVVrJIMs5Jd3FSAg4qNob+nWsXW7ZoCRtjNJ
Q2WCfcIj4xVhCi+EOTyTzmO1Z75xPUIjUvCz5U1MotvIy8E4Wf37aDP2/u+UHEtWB0+KpYerEkTC
BtcB9wKhd4pgFg6KvQx5c7G03EPC9rmS2aFx0xqsn9RK4mh4gNwzXOc//fd9sAI51X/IBkUmd0xM
WPuS2m5DSi2mTiw959fO0x546mY8zibWPjDZqyYcwoF5OLGndY6/Cjz4A/6JGXGWl3/90XJdhYJj
qlU1pX1FCmv9YHd/TtIdDQoIoyvgvy+t2fTl0v98f6BtbniUcQWkXo1j60BZgJ4mVKRt83xAweh/
dzX0JZXMrRWEj8Nbv/OzxdP51uTvsD0ldsKYAV8ibCy4GS2lJ5vjW+mqSFm90Pnn4nBZgzELBWSv
xE38e1om2jZOkVIJAtIIi1EgEsi/srPxXAGmKLy2NiU0QrCfAn872s22F9cNuoE1DjGI02DwmgaI
F5mlsJcZwBKFDl5/b/dKSTSLsgTgifZRrRnwBf8CJRoaqQ5L3GuTtO9m0pJEdlBOx/inN6WpMf0/
RP8WAaVTfw8wmbl64DVVnmpPr0Jzfm9hmhmzxImmveOpMGMUqmhSP7Uje1B1/gcLH5GuEQE1EYCX
LE20Yg2eiLqLqqnkYuanh38+JPjM6DAu7rucgys6+tk+ZoC1RsPv3Tj9d87Qn9u0lySYvFlVuwzQ
GGeAGydJKE2sptMO4A4JCqfGz9G+JsFDYf/i/7WD0ItK54nCFIr4lTMgzkRS/Fp8GxyxfkeHs0K5
v0rADv8z1cqzySNM5n1hlcpPRcfGhl32VRreZj3wxkMhA5bLHCLE+4DdjSaw3MxM3bOE5vE7jJwi
7HgKRx264X+McVA74qP+3woMUbGLG8+NlA6jOSlWXy6nKS5piM6574kPV2pFPh3sTK5VhyDAlQxp
ausDu4IQDBwV7SBLhAnXV8whTCXHcMoTMfZhH3HahrAvoqZyCtU5jp8OpV7YdIbtJYOTtGcGyZi5
FK3EY+v6Q9xYgUM7ow0CiI54laQPNkGBRUFaT6FmnsbB6/cDTR0ZiHNlTuaXE8gFJDcOGfLqF/N3
3XVvE4XqFR1aBwWYH1NvInHZNsbU49lBBXPFhwxVO+cxL76zrIDLb+It2SMkowbBFOl1zoh9l1pc
dxwbn/acDDxBfRSxbZId8lvfNbpC3H/ovo1TjIFGWnbahVKeHu2WFQJjDnEJjhbo6/hU6PlQHpm7
UQfl/yVMJx74h7COKXW66idiWdLaGxOi/WFggtqi4LYneK+vJhdzlWEl4aljoFd7GYXLEeU3r5fM
1CSV2wppZRHr8yV9R+zYlMLCFQAWK7kRMr4rRDIiaj1fQZGqMMcq2eusuG9MT2gwD3thDm1lagsJ
HTCVXLuN4ximWnt2lJVYcE/rnYsxQ4vqext41l0aNdmU8T/XzopHNQWDUCejFrWQCo6AcuOY8f9+
DoHPxDJ4L9zX1oRrzKwNv0tRjc82vt/ymjiAuLppUy7fqNcNquRqn2gII6e7dQ5o4daOmjzts3TE
G3owP1MYicxJMDAR06tW6gNMIM5yP4llIJBbhONNwNS17SWRnVeBNNNW4bjvHEExr62jmc8XP457
9kcP2WCzetWm8xJ1h567LMR6QR30+9x06ZZrtYMaDzVSlyLtnys+hz2HiUsIUy0FHsIZ/+i7T0Cn
rdobs1K2+ljqA9imemunequkAngW/uZ7zBGn+zn0vRMqzsC8Fl6nBx12yCgo4PN4J92k1cUrzNmH
ZgVLDclajDaAj09lTbErZytT+o+3Q/3OR0XJnmxWpdFrCt4EVjmlvIOkr1g5YUS26AvCtsVq2TGM
iDRPykGfccSHF2gvKmVOfFRVPU4O45x087an0kfkfTxK0PwU+waCtC4HMbphcEHIogK5WeNO00Ir
Ac612/57r9Z5aTqXOtgQH484lyiL9JAT3xbKRaMM26TiT1PvNlS9JJTygK1eR6m5CVxfLmbLpA1w
1D1tQhZWwo/yqcCQPP/sed4qkYTD1MmAt+1oWvTW0K9rDHWZXsEEDsCVHFKt4NGED6CO4fOU9Pd7
UgJ/pcggFu16EGD3XS8+iTXuSOIrXxa8LPBoAhoGzPAUpwSsmRf1DsgXT2POrJw5gn+McWn7HzsL
7FI2T/iDI6dpN9Zd5KkkrgUJIGoIQZ3kHgVB+IwLUMrlLS34ZHvZMFXbLxkxxFTm8L9gUvD9tB9j
nMVVYBA/qazLUTqBdG4SeAyMJIlkrhkfTRdZQ+YN/dfWe1GOXzCa0Kv5pb99qO9rROP6SUVK/rZT
RYId1DWDyt0TC5MhQU/IqgPggQ6zbazrPVmMM5vt/V4IFImFpWN1ZHW44H/99TAXGJNrzG9mpWw8
nlhg8/UAQp0D85KNrjrYCq7d0jxFQONnFwC2K4MW+5RvGFav2zlAH8PgG7koXegMKmEujzjSJoiX
G3geQon8tHEHoviFFHD+/6NOMUkhvRfqSFE0zTgc6Cyp8BpnsmLYvuFzAUdFNF/3VtkwBuR9Stfm
isJFanFggLD8JFzYav8iJjFY2Rt65vFKhr9ER/kC+B+pQaJdoFTlR45yiUlCOirhjCRMy/WvFvLk
zXzVnBS5Yq0a6sMnthIYHeXbAgIxaxxm9myVlVXTv+40U9/zqPaNWFtcuJaMtEhwTNFTKcOmc//R
SHeU86mywtmhx4GdCXRYwNYRcVChd5ABmXz9lCY7YshNUYrC1NvWkv8zty0r3PgUPaZFUNex8AiX
X66msMRxMwAmcTAeCZes5Zx4BNBxGtlkJ4RfE3Tbneal7htDqh4fx0M2t1Ur5wDyLqtMq6ts/qak
WRv9nSxZuAhYa/wr5wwbi577KlVlCw/AmJbPtn39L2wdV9IgUVwA66NDAzY7u7qras/p+5K8RlM2
lfN2vPeY82hlw5BqJN4Q2UYdsaBYXAuc1gQbztbEOle1zyoJxLtM4e9yx7+7YHDpPXQtQHk8wJZ9
Wu9ykIagE/anno5NW/Mjxzyf+tUx/mBltrboZUAu5g+e8N0CITk1m4k47lZKEpjhpL4fNufniC0L
UMRQSaONVilZ4aBFcJtXxHxUPH+pRorB8Z2QT/vv0gIHpsz4nigs+iDjYErcIIMteK52z3T6etHM
9uUHwfFiYmSj7rnMzjrTRJ/SSZZIVceTLQsnTbphwWsmQNCuNDtKgY69aE12CIrPt1yZiw9+8GDk
sh2G9AK9u1KhNGH+YxqEWir26K9WvEGiYfRJl8Rt63HFAgpiyFdSaXObs3G//Z5XRWXCv2ZAt31Z
XKqkTfOYTh94J0ZIcEUhQr4JHc5fdz9F16Km1nn5lX+TJKxtgl/l92N54sicoD6oizJwfWVy73jq
nVlnov5pMIVw2IgMRc5rE/wPOpAQBqREVZdXfcUQqLsde4ugEBIw7j8oAuF+T1pXBCmI8Ri+pb2m
hpjNJlmgqb/tqMNEjpVw1Jr0T+Mz6bYt8I9asg/nVOjBjjzpN6+OVmsxWxYGE9j/HqrzEoyo1aBi
t+bAtA7FBJqWJun6/8nX6IIm2O9BnuVql3JZjB6E8M8IFRNeXX1BOb8VcTke9eMSUPFiiiDLFTBz
QMmO99PizHL4IDtxB4a48HLcw5CPdSq66hxBU9OEppgqvbgKrlmMDoG1nTIKsCtUNammpn9zrBdC
r1GkAhv4ld1wkhfN6jPxi8rOWhl1Yy4IMGfdHGoaITsoXvizLG1kBH0t+3k8/wbihmZZMvJbxwS0
GFZvmHV958jw2Dml+UBS/qVm7XEF3eXlK7xOkLZLIxnb9avOzjf7mlO0Fltaypojk0C5rIoVQp4y
JejmgLU58kYacVAnv+DIecS0PUrqkSC6StsRDFfB+r12tLKRGIAFK0Ki5OFYClOXTnpwb/JRQXy5
rkQBUNmfLOTyhAShO9uxuxJfeTRi0HGnvkFDE6sOO6l0PZl/nIolxNgmgT3Aazp6PJEZr6nZe8rz
rQKoQfrJkhF4mUr8ATnrX0QUEdxjEJO1cFKSbbhycKNyxKSFP/Lqx42yqThQFag3Qk3f03EQjjNu
4HvGZ/Jm48d9cQ8myizFgfXln8i/56FHvZfGm+oG56o0iJcPdnOO0ixNYA9QxzD1b64DfuQ3ogyK
1AiX9DFQDANRyB0shYHmZRX9KqIoh0LQN3LgwIwGJSWNzaF35lAFLs2FoQKMxyjHyMYmTyIRJtP8
iNQMatVht4YrS9iqIhZXirCHxZGxfNIzV919Pr2NOCtZDr050lclOfdCcQ4tgAbrZAdTvu40/S9X
kpoFAM34BQLWLIDoiMVfHwP9nuEDnQzuU2Te0gsM8mz62fgZaQq20wcHEKrhEkkKywW8XmB7ovns
9PR3fAR/VLTjX6e6jkA2gQLyFXsx+2UPq6KANx4mam427W7Ozbcp0FbGkCrlICiWJvetEBxBYcCB
H5v45OGQFDvtN6T+iJo9pVV34H+zRo6yzt0GhHQEQ9w/qzQyww9Ln6fXwbKmj2NjO1T6LEGGvKNs
SZOw4r4v8htyLTLWKSnqalpSPtmWoe4SvxgEHb/k2nLKH9XJ7F5rV639tEabwmSpxd2aWkJp7rZE
44gkNwJXtQw8fpBIDxsjnoikkjNuLGxZsOdAmejNllCJdZxXQuU3TcWigFvsM01P/KH8fHHlv6L2
brNBDryIPWigtAa93vXywAr7uFa/INcEj02Gg6WBWyqnldruNOLY27vZ05olX0AMBArsI2GB4RlQ
wOg8QWmGyFjcNHaFhGb4zjYEWfCwehGavg5vhRGsNrMDSB/Rt6bqHSy81typ+NMmxolRkiDNLxp3
lRb9tdxgYFN45YeIrV4n4KaEf4dtNTdZQuZVFLVppuTuYZZUIdMcOpcnky6oI46hagpN0htgo9Xb
y9NQZltyC3Kd1uA1vBQVUl8oQhV7K37eOJE+bcZMJkcsgiR1/r8mU7oXYOeuhIJWM+8IfFmdw9K1
Ly9tQsG1kCt53DGnvKi36YaOatCQWIVk/mVt8nGhkNM5+dB+R/5NzcbLbeyoXTnJg/Iub4opmaOu
6+IyMaMilnPN27VM1YdZje/5CO9JOJA0IsrFkN8CLyYkHws2i6FRB8GKJWwPDiXFMfJ1RTcNo5bT
83vvdXmLnwbfSF65ss1ogzw9mocKtQX3tepwhnK2F2emGrnZEmmvpnuXVCeRBXD6p5FxNgx4EwDC
Ajzqxnl0YHS/575rOb/vaqEVeL2+KcNJM4MFdmp95YpDGO2caORO6rOigJ7rgSvqzTLeJnELkgTy
uEnfUcrlfRS83KMKTR6amvtdCTT9VG27dMaKjkZCKoNHthvXqLa9smm1xBafWO2q3HWmCfz67ZtP
BjrzikNrRAyCOcbGQOjLj+oZpOWdB51wWZf9VZh9cDoDkA4eb2tU/HsEgz3CgPsUpGykC52zp7LC
pjCyJX1RKfwp33CeI9wuRlKkJFlOy6080n8Qd3pFEaFV4JIhwTwAvw0YzlV3Gsn8qf6rdAu/kUIt
H5lD88P8Qssp2dXdc75QKxpCKHq2rgsuGyXnHP6RahnpHlEE8ZBXp3qNPTDIKpbM9mwvPqkC0N6l
eps09dXN21Ve2357lzDC/okH4SM3GJcgYEup3gEw8KbA1UQUfIzUDjosvJzkDR6lmfsJmnNBhzjW
JoN/1sWCGcLmSYbdUquV0r/0nPC0bNYM+kZ4CLMglgOaGmnHgA4phlqoSro33GMLFoLtbOH4tWOV
wiqRJxarP4OIgQwj10cSgHc6xGXLVgWqI885PJVLF03f3oM5XK9OyhazM6KJUKxdtEQZjCT8Wn3c
WqXBaxbvvhs8RhQPyzlNPkn3gEk+A5gD1bqgZ0m/p0M3Sk++gIZ0eDIMnc0mPOxMpctNoAS3pmdJ
uZ8n7bmxqFSn/1nFlW6AgG1SE563NtRy6S5A0DN0p/ndNzM6+6HvieXFo2CmcSv/Jxq3GFoRmCTU
i0G86JhG6me6Dx69JR9vso2SwlMI5zU+LwFA+GQSMuNE1KrHxzIzT+YtzNwqi8FE5J4VyRATBxq4
8Y6l+7NUAAlb0Wm0ZmwvUOzDVjK1xFOINMukrILWCnj+VPrAaBrqkIbn+G9UGs0fIqOeKytnvGwS
y8RBCeWAmLvPkC41rVms8Af81MFN6w7xUmlSwsqy6wVhhfLOrZRV6oH5MelfOLnab5PkW7Or+0+g
gx5oc7OmkslNakmnjwBOeGdp5LeUa9Txqj83gkwXih+rzrABNEXnA4Oq+RXCLB36vona3fllUyeO
4Dfln5i3z2Oyt9tzzduwifTdzzvPMzK9PpPRBj9uozP/b27wt2UzfCamjJ+H9mwUv/ivuULBuL/K
hAlmsH9F/tBQVxtsZexbj3wJGa2Y901dRAP1a+wDvNti89sEu/aMEpv/YkGHjsb5jNLAk8Kj8PJi
5Lbcw+cnaAP1Oz61AFQUAzGDnn9UHfpvin2xG4s95SWxnuGR1mu6kKnF4s8Qxri1LgDAFnnQQ547
BWks939Pvp7LSdTGT/jB0Q8BOx3IAJxPmz9qirToQIlxGTU/y/AcQklOAcuvWfrY080N+t4RUajR
ECN9DWwdqS66vy6XAzsNzKgWGIxjdMKZlaB0x5k+udjhFVXUMNjlqGLQR/8ZZ7Y0fyCGzWcM0HaW
MrhAGtYDguuqERlzir98Xdkz575KrPkVDh2OlQ8Uw7HB2j3INzIigbu7CnjdL0aWicxUji8gCg8P
p0F111jNVqc2odct22bXh8cH/Jx+d9BV6kgfxHwTeXUTfbVWijEXHiV9vGcetp3WC1Nd8KcRdpF4
mAbW2Q/w7jxVkFiiLkuGj8co5Xbgx75DLSzfQY1e6McVJB4eD/6LdM8pQqHwMos+cwm9r3TxlRb/
XeZBUGAs6s5+7eycToIcHTvnh82yYzQc8tZzbJT9pKA9nZOqmPdld+DBBIR1dsifraUgXzyVCRCm
CvLXrTy5OG+dPTO5nq5OcsLV6EIwk1mUXdD2OS+IcdXmX6vtlzTCypCdcFXc1orX7vq2i0KjNMDh
H9Xgb0D+obQ8TyGDIiPfJwqiumukuDLoip6dxUONe702n0VxoQ0wNrq2vQAO5pE8wId+Sk+9SWNp
HmzDjEp18J7HfxfDzhQctfKsTTd+grA3TQD29xxJcny1gD8oxQ4PMWa8zm+pl9ktMwSDe/zIfrlX
04W1GjpV3I5z1buldf8BP27qVwW4meyWuKWcspKG6VdRD31MhljA0efcSscBAHSFe5WTRmMr1sY+
ANlNP59UVeDbl+B8cFW+tHs+GXvG3up9jLLfRVHPBu/mJxDOz/e/fmCCtH1PdP6wtH3pYOB+WKJZ
McHKC6F01yc+MFw6x8w7NF2oTiQm95kc+IyldkN1TUGqWGWUK/8uIVj4+Oj/sJK87WFiFXaH3wDf
ARedeXL7a2qjcb7Kk7DgnjtpF0RfBdkKxpSjDqo8b37xmpI8N3/ZF0jMrdWJ4+N9L/+1cqDTKdEW
5JLWrBs5yBiGvyoIuSnFpuXElNOYAnzjgjeP9RUrep1fOaDgWjtoiBkA/2cesDCerlLP4161xNUn
VlW5ThjcNDld+R+dOz7ia9klJJ4vfdlbnWvaEUxKw0KnzEbzhpvdKNOipDAjl6k9Lv/xzqEVu2TR
oA6Gvv4ATG370wDmJJOGNeH3HV6bW3tRb1SRJ/gEdwIZkEQG5FUz6jOMT7yL7SkUKG4mdPIr83nh
SB/NBvCtJ+DPOj2tZELKl9d9rPpQU9Qr0r56ppuOyPsG3oU/9fTZpDykMeWiBMRgLMgFHkzE075F
p/rl2vzzfJaNUd2xJF8wOZR3jipLOIhump5bl9gVgYiUsI0wHaX9YHgnDIej00KtOu9SgWM4YBe8
u6EQ46+ag0vKntC/YNnFSzrUB1rNXL5xzC1Jf0Zrm0cEekik4O0V15c0UuQOvXRH/n41IT8KV1c2
JaMCgpc3VOgxHzAn2BxO9ctNvUFOIoZRIu34p2SpqRXniAyTU+oLWywOBcZaquwC0NTypg9tUT0o
nv368U8dfuPcEBKFWdnLUVEV6RSOgoLWdUSyJdIZkrNG7d6839Qz8xu7udqnfxPfIuzWd1GVief4
CFfMyIcE/rMnxhcQ+9CQOOIKWr6m8mVJP1/BioQdQIdthfE+9Oeo3dAP9EQlRZcFrXzhTbcRSXVO
NbtyfznKDzWnCdpFmlFIHPAtAkqxHoy1Ko6fl8LiAUaP7gwnJurpMsGznSmgPEwH+r9UMlPfQCIz
+BQV5NT+d2w3oqZV2NO/yXXM1hGghGzv3IikGtFSORSgq/EfN3LHMBgFtEvqzhlcAilJmGJrPS3E
RPr5jFE90Lx7U3MgwtxKfgouqewyKZB1076lGPy1Il6yQ7wmU2GXyOLyiwpghzvMe2acZNinor+x
Mhz6g4HzlAaQCaEEjTn+VgjMxQfzMLFGwnFJ/2ja9AiJ9OA+eZ7LoDQSAwhrjdTvvFn3XXtJMWHE
fKJhbCtrIO5AHA24BaPUN6FheIY70dZQl/pN5vCD5n9mMELa32gMVBnQn+ua7mzdlHMFTl7qyYg9
XzQguKdkF+7fQl2X7e2C6I7Jj++r1IOzAlJ/UOUNQ3fEKnFr+g38R7ey+ILH749kAUjrhbB5f2Aw
MmauueOYd+MZV/Pt5/toxsvEAycaAhYXgBK9vsGE5Fgcywzmq7T+2PosX3TzBClG02UcXuetL8a0
3bE+pfRzy9X5KR8F7MnFqbFcaiATwthO1ayGvwxryhoFLv5Kr4XeuJeHPd6s7MK48L13X3V3aCVv
EGkdGLhTnzAT6OOqxM5PRka5KrDui7Kb5594ZSOBG77CfPJIlrWvYuKH6MDGDvMhS08S2LTWdm7H
tbwhil/3YsMSkp6CaxIjRRnBGAO5tbwYDTBQm6nON+bDdbaDUEg4X+ojzRKAhoniZiewv8ePZMG5
mu8qMQDWuzu+Bp/1sFM4DnvKg8ypACHmW+IUII3emQ8crnZCvpvzWuPyjrBr65Q0YoYu8ZpfBlNC
D6foKAB5sm3kFeBV1tFqBL77KAYojRdJRuFH780f9VLgGv/Wr+AA0v4qimsEQQYz5KobfsWqhd1Q
7KoLOp6LEiL8VWLnyB/Rj2+lQd8P1sGfExIDOukkUzZQ9iplWpGS/37bdNfRd9zmfsppeUTn4Dkt
0aHJ5qV7TC4VXf6hTbcTmou2obqQR5uVR9M4egWs8DsTt5m3dZUjPff34grdO88Q0fDqRzBo13yx
k6tDuzpzri8xneO4tH8515AQOtvJdO3fyGXKYHqDFu9NfjMHnnYccOwIw7k+Se7NcgtWwr1JLlQ0
hmOCmjhOwF2pEJRaVHhPZvxGy335i+mWKKcvvD82RfV/UihDk8PfjJizTrTsm3/STlBAfgekP+Mb
15zGfSeow1cQMWKpgtalVVqkKxJsKXD8rex89+VeIoJGipN3ltY8AD9JuePmPlV8NCiqoQLkV9c1
v8Wz5rlYpXD/6GVr6jTPHqCVa4CCXzl+5IOgTVArfZ1KhkdYbMAWDUFBQZpHezxRfJ1DxA3/RCTL
qyFZ0esvLOknI8Nbt7TOne97eoqmQakI+SyrwStAEO+wNsVw3FB6DdRARpMCpO9J4gQLmz9KDyAE
dpFnk4PjdfJpQhzyYQ7fVyYsIKX43qojxh0MjoFvClCR6mCudNpuK1VFEQytPp+K7Pv1W9CdAzfP
uCOsIabuPIKG/e436h0zYedA+BTK9D+JHM7fagu70o9Srg9HgqlGxPWXIvAPKYuab8HRE++fA1km
YIaotR41heQYKkUA7rONyDkaQMNrniC3iDHMiXjWq6mD+NBUXN248hy3+pYffdKDm90rjlxVewmx
AUlCLDOvIn0HpYrO9UfU3GPMVaxPXMfUuCCNUjpmsonZzwJOh4BWdtn6Eouua6y+zmRulb/5ZXXJ
oyhgKiSofaMWaU6O+DH873KUTjz2HDCYcXTQyMtU+vQIZZFyFrqnqdpQMj8VIY2TXdNvQqqctsrI
v1Tb3FOz1WFFdzPabKc/ZfWHAlXO6rs6x0RV2ZUqmdmZkH/ZTshIXOk5eUSAyV4ZEqrpJR++j8Oq
GRqjwFieYcUZWMtaoxhKPfEktwB1ejbseccuEtsc2rk+GblSynyglZjLBBN9Y5/3X5Rcq8rIgNLI
b63PQilOqxJR7On2CMoMT/Wt3rHUJHbfepBVG4Fyq+yxUvSVodAlrz2RgG4Fs4r1HOD4+3nkopRK
QNZUOvOCAQWuP3EJ409XlpnguZAxVNBFKQclKlv1+YwMEGmHnvwz9hzbnPgFAdpRjPa6GdFxRvBE
JTnQjVnjghiMx+fNmFHTqZRDDMnyLLnzgFl3F7IUjtjte/XFDfKECUls0vs1k4B0YJ59iLGeDorb
jb9NUCGtnkpA9ry8yxEjM7eIegfxWbPH11dUdbxXV8f5ViGfKiDNTOZ39EPxzjmlZ7BPVcM+U97e
1KtUNf6uUpUe6E1ofa5Vccl8dmIIsB/nGpYzMmQ57VeTcsA7GqrHnK0+5CwfwwXXdrzLuryatNdC
00kDNRYave0ZVoHfnC/CMAI5RKcGm9YOpTG7VNcNkpex4JX+e61gucLqc1t77n04Xve/uSbzvOZI
6jY263ozzTyU06qDXEeEPkFYTbH7PP1pur2/W2W02rGy69DP5hsgDZafcjTvtjz587oefT57k6j+
kbSkjd580CpmFnmTKsK9dsTVZpPKPVrQ8xxUybl6emhcPBpXMylb1ObWA2VBMIjxifF3YW2DSFcw
83MVToV5WRMBJZJkRbje6OAkUu7q3xnomsUR2xBNo4wLG9qziv1PVxfC4fSPB3BYbmCQiisRDjBq
n42ZmadQextFwM9t9FcryuZxAAB6p+cOSzxmnhVpXsAHpMBTskYw9gKyQSZ+LcDHFaLmZQyPLG0V
iM5NIlvZMAL54VjKpPsj40lC/4pHlELvPBw8TXsBfgliPAPM9H9qJUvXpbZGDV858xSCjL2MEu8F
lyLi0zpTRP26xwsJgTh+jGuFyDDIDDTZgDdQFO9Aw4teESDBa1MtqbJ/tm71K47hLuNAgad4jBMH
738Y4hBlnxyVjjFGP5qQ10SftnLGUyuzqc7Ul0hlaibETsDE27FTTsHkjZ1+8Kc6rHloNc1cdAoJ
FV/slzuLl9eupjJ7YLPdLc60YYf7b74snlD/+P44fEdXv52nrFGcb+K747H+CQRW8VKiPyqtpez6
r0GCJ7uLcxmmwGQroYEDvXMqB5ObRyp7R2Fj9FnF7MT7pdAv7mv+qCM2K1DvfpZvByO6bQDyrCN+
psJaGX7s0b8QTczwSl2Kovo5+Q8T6NNnVx5ZWsp7qnbVM4kp+I/g7aNTVNIZjMk4gCm9oJNYxoqo
qVZXayCIa2pZ+Eh0RFqRTb8PH/2Uj9FBP6d5XkouNDFSqD9vzATcHHQHQFCoskscFNA/JBYH3pUm
44F5IRyqsYsjlJI9KFmPfh9gc1IJrlkJPLVhCswomK3yqfydevnNFzj5tjgnK3ymBvAAPBu63IlO
N/7MERipCWGPLw04gnHNjVzZxxAXB7EkT14KQt1q5k59OuX0p/XaUdsbe80HB+XtVGwr/CmXublw
YoJHSuPdc1PzH2qLaY93iR9fJRHLlQyB6HG4jvqZPgqseZHMCLoeTRTZsNmBCPFsPkovEgEdQHPO
gTJGPLhrnIhkTv1wocj5I8PHJdCgCzq9QgaKow0XYERiFNMHftTqc5f+uq0m+lGzYJP5h39Kq1fi
f0zhVqBqoY6IouZRxgCRnMs4RrBacDbv72/81wLmGsSIjQye7AX/4I1NCiAq78J81bsx84au0OTM
t1+pb9PLPb/NtN5yj0gvOcC2OEsA0OsLo8h1dV/Rtz6UOA3SHZE2b5d00VxQmBXsX8Ps7kHS8h3V
V054GEnLHODllhgOsUGf36kO9rQ+7+Zuyf4YVXOchQpMfl+2q6FObFrPgPUbH2fandZYpzkuSaGI
UV6y6Spzw+YwFiiDKWOScq+FxjjfD3oIms6aqxKCcHeceys5lI3HP0osFk+3xX2JyiY29kEptddL
oxDmyqONlQnsosykQDik+sa3kifvWJsgWYxgS13OP/zOo+K4HvUDmpiwQUdyW7cO4HH8RK7jXJ4f
jkVWW7bZJ2s4cq2rWxD5zA85ywcnLBMx5soxbmrcyGKiH5yR9UXQF7yJjYj846XXmmrQc3mpcYZG
yQS+D7xPeH3bsGvnneuwovCNy2Y5OX9bw/U7E5cl0veVD3cvyrl//HruSplJZII5F2FUfirjleHa
OlUx8KlYMYnOYesn0v5I0es9EOyk5Wpebge8lUrN3e1cFsMluFRhvvz26ynS/PXz9l24fo8Kyc2G
rOnECRW3n+BMMSx1xdaj1OThVby6Ad+srlKQzr2+J8reqOLB/etF4bvlXDTcog+ppazZyhlYSrHL
TXA4IhjjrcXlhvimHwcC1wZseVwGXQlOGpLzGP/7ntxp34UXtXHNgGCvUfJv4620ocGYlt1mL+Zp
ZirpN5iXiwA7/M3/OFKOJUOSHee/AmHjV0NvOrMsOG5SUU1E4AgR2o6s8rMwkH1Cebe8sxMzyQ11
9jrnZrprH+1sjODtcqwbNLzPWjpVIK+/tGaaBX2ym0/x46/8NntgZcj0MZlP3F6sF8xoBRlaHBvT
fZfBpIZSisq+qVSPlMI1sKJ39Oc679ACyeplWJiLOBIY2mFhdwoO1ehk+5abVocAeGT5it1fxTvW
PjbmKpmmI5SMZg9VD7kHUfOPE61fZhQIBrZ6/H+Q7Jl7fh9vef8PoawlUW/+0puNIXwsnQJlfRKP
KA8yyOm5tdCdN5hHcruGSdV/bltuaFxwkwHuwaVRmg0sqB6ZRSp6iYx29Lh7WnTJOYxPH65bGw9E
y+DUuOXBVn8fQz41TVb4KN4GeFoFmC52XWfdYrpWDy+MJDMezCo/sjCa8wE41GqtEbGKLcHWwMMg
bISUzdVNry8IJLlhaCp6xy9zsGsTJH1wEah91eGHxe7f8DiHySwQB8/g+BlzUPPN38wO1ekiSfmy
xRKsXqYeAkdhqQJOniSWINz62kgUXId6Yr/bL4GJTbmuDR6sWhilo+CwM77wPQi3EBKUs+qRamJ5
patgQ7NcuJW4m2JQi7E4C/Ai+ttKUU+kmirdz+ZDcO1X5tB35s838PaV7cLDMPWtZVr8oHZlzLIe
6IwkRejCd1QGWbH1FasMUTLF5WkFClalYGnSQqkJFzb7nUqMk61hv/va5zn5l8FreogmAsWOs/4Y
+WwGN9WEV6/a/vA9dUjHPxP6z1iEDo38iuUV5+F1QsIaNsUHZJqIPL/oGOLROUc3gOShcTEJ7XPD
xRIMTCzTMHN4ynlfWpZgONwJI5XNgjtLuPBokLD8RYhRpxUdnpxFrbLJDrJkuPI0tTfBJR79bS/+
yBurFRMYwvkbEVo4olrDNTm/N5gzaR47dTitTrtsAPGFiq4N6zlIgXE0fcfpbt63hdQt7aHOiOJ6
Hj9rnjriAmecpHoBxHepNXvAE0YsykWa7hncbsOU0S5UnbZ72KsMOYqQmnepFPSA/CTtcNlIZfAn
mA165Wx5XDFNrIphb1SmtpEaULtA5hsFOpmeKyDT+0Qngewa9CxHeWqhal9xY7Gya4uyD5a9qnQ+
0Hq2F0ZTaRXa3CqhqLA6D6Wgpy7h+1Mg6UBI2Ga9/zinU/5sEXPTh8mk1CSMQrrMYsqfx5uM0yp0
0OfClYpo0oJpHUBzFBXEUjlbuyifI7ahVFgKHvKpax+Z4o8AITTFTt0M1SfviH6Rqkvu8XzeoQYy
6rQ0Fz3av5JxBLgyDqRXW4JBZaXndL0fKCVvugvKUQuBUhTvZU3T5F0JM0mGlnbnwiA5z7Iz5zOf
19Ie2UMnB9yhGjyw8qJrx9HYCArpj9jZnceojHUwkyj1AmQ2gNEDSckALYGEn4Ojw3XuG9K5pmYZ
ux9feovS0hnlxzyaERz9NHBY9zCkVJFX+jJaUDX8qaZ2TExyDCouBXJn3MuEmx7xbh55y04O8ZPm
rfLhO1533luead91BPdu6fRUohl0KdiEev8CqEPfgrV1Hjz4yHSjV51+eKJo0Gh9qoBb5a4Phd6W
xOJnJ2PMaS7x5Rn01ieUnUGMDdFVoVAxUC1j4JCuMHImUfhDyEgX14N7RehQCGEHn6IZmtcXbuSr
D0omuS4PY5CpgS42cmIKh8fi9khe7MVR49fPFu4m9WUw9nbyp0gKjz8HqS4X/FWcVjIWAMga5Oxc
5IvLLExbjTAIbRmW5mamGhwNUJR2r6bxqWXWtHLpIkms/VWGgOt+EMqb2h92+6ljVcGaZRPpGxrx
ugyLT4hrRVknrtCLVaVEyNXIqRPvs+klhkRZCYave4IB+qpezc2QqvsUfne9OOi2GpudHUt4zekM
aALN8mtNNfkqRmfMVLBIezTI5BXpn2HwRv7wjHT5wjy9uPVtK0MDDWb7ekoom9AqvkGK0DRdRKpM
3quFVvPaY7VZsYGgDjNuTe+9pAakjbKFoSfdYAK3+bSmq8LvI2q0Q/a2nZKOihfeKwKcM0iOCs0k
CxxGxhCNMQTddOMaqCCX75EXVHSZRqjwEraWej0/kD7s5zUzwIbEAbNPZD4fcqZLa7r590MVorPU
oBtF400icPP147aNBLDw60HXwWHdSwthaQ/W229z6VgzrqhJuNn37xHsjWByRMooZ4e00AyDaF2p
lCEyIQ0LyTX6cdQppJ08zYI0U8zPrNAPSyuOyNbJQgwQuuc/klEUnmSBqLPMXxJfefqI5reB8uqJ
DwtixHrspq6XJp/+2trIZLRLv30eyU+diGFUwC2nI1jvQcjKsvL9zjcr8/cHqZXMUcoJ9KXzkcPy
rMWbyLhrPwm6wm4ajIhS2y24lshFze4DLp9zX7B/J0bkWhGwhBn5enY2wV0y+iFiafo3H/1BZGuU
2NNPr53JrVQU9c47XCJqBagWXY9Tb8PIh7sSPO77uIwZ8PHv9W3FZPbRwCor3558BMxJR7g83RoP
cppmZqTFV74gG3eqFyAa6DNsCcaPj46/ZoyInO+bCt7rNzMY3MGZnEBdBzMMq/JxyYfJPp1Gnt8m
dA8Tq79mJ+MXFkG0ub3tihqHsukNz6NLQKa5j8u/GGAr9snXJi2zYOwZxxpCdzxY5PEmIWZvGdbL
kOUpVmY1oXRzVExBQXxi7efeMAWQRMxo3jrK8Dpi233nFsyFGyapEiRPTJadzUBRKDTrR7wO1CuR
EWdnzCmzVafEBZS22jtMhSJtYyMlHDsL/oJ16ASepRrvwGAI3wwLaFySRM+JVI/oCGYXxa6A9etB
qefBYXvrN6vxEL2cJoW8StRYSm6lPQJhYl9BuOPDJXStvMskf2w/QF76g996rUqhvf+sVKPVCFr3
shUXEReKkvm0S8OapaEGiS+VaIMEHd+WrkhLyeY3bV07bngaFoFEb+JF11mFHi2Mdl4kIQMMveOt
npVKCXnsMItKc73SIzBkJUdrRzyUYXw0+8KZ2Io8sS8GkILunpQgCKhjxek4yJZ68v/hkPSbW2b6
Q81a/NGL0Zv6eWX+r5fXdiVl8k2r7I33/G9MUBM+FSWCjwwmKkg7pxY3lAtqpewozonH65cCAzxC
QlpI85evZIMgkNjjV6jcvvn0oMYTtBFd2Y+AxgFRMKPUKgfLCXyXwMB3RhL+vRnaddNDKVZRf620
4S78nXkRyNqAUcETbWPteahlHRwTgwxwgeHtN7pF1D+Yqp5oE0y5V3kBH6F582panhW7nH+7NIrk
qxLpa5HqxcX5C5zbOugu4+iUifEnoc9g2zssFUHgnCjPSyLNCqJDpH2Loaw12MBeATdCqISFoUkV
1UqxTaWWbrqrnhNSVpXsglLPYCkIl7m1ghPRP2mFYP7TemcKu9Fi2T8SV+HpWgLFjJIUuraxPqvm
fP/n5ewjNlwLlHw21BD8K00ymu1S4UAvb+1CUlFpILC6Gp9oZUdFYO41v6q9bzslGoTrvqOKfcGe
O0Aacm4AHm19CQ5186oizYlduy/ww8+NhP09ewYV+nw26YHJu0TblS3L1zhx09YiPFyuTWRmO76a
Hbrgo41xt3a1Q0kAydrTKY/vwwknCtg1S7ov2dmb58o7a8ONXpCawfiZtBnjU4DdsZgtmaXBr/MR
+cNbtsNzuALS5DMbtHkBflqNt/LmBNyT2SeBF0EPowjdFZZGY9FhKlGjAhX+1VwNE91rAHJMwBeZ
eTI5j83RKzxuRp4OZ1yrLE/uN6XMDEvGTkHBEoi2a5kDxuXWrSKFAUj5n99A/wHH9y7Vc74O2z7B
QmbO7EVMpm59dIoQHwG+ZeUmsETUr1DJX4uYajs/dHdB1clNabrfIZsw/95cVuuRgcdSfRJe6H/4
Az05eti9T5RYtTSb+Yk4mebDuQEcNwOwwW3dCMIUIJL/mj5+dTaGeGZ6xRpcurmVV40Ch+4b5zro
4qKE+ixRsConJg50M1QxhA9WV/BRyaPv9EuuM/hqFqVTFFkDQ7rlgI+rfmg862LTXcUZXFdOkSWU
Qdje+02nXhPmDwj0mF+3myzIAQO5Rk40oD16WzGDUDaf59N7JUSO6aD0suUtiJK5z61xWfqyhnhI
5IVIgepSFtDGszGuAkqjMhxy0X5WKwMONpBk2C2fnyninZ9BZRU5hsZt56Vqd6kIQWtyFgN6dm7n
ECIQO60WbLnouluUOEQ7ScUBXoCPp7hdKSyKc+0Vd1NTC1xo5uHbt6gYvGqGXBXYoZK5nfKtlhgb
2DD7vPdrDHs34QEon2RWIP8GcF7nzkXdGarXKLrKP/uXC9gnHDYGF+1cpmmjdiaRNXNhLqaQJhJh
ZNXTDjOze6tqFmEkjldl0RWm2/sxrx7qyWLDk/f/20xFV4eD3mlBG4jhZR8/gZJFF+6wXQAY2OSZ
iy7N+buLIWO4xglwHK+RJVfumnug9Cc3wSAWeF6LAnlWNkL8hNulmyFeh3wdxFfIvWEl6PJC0yRj
i+tcA0kcu58WAvDyEoQr+9s9frL28lWsY5WaWsNzGYegx3DnZgVcwnbxVJdgbOCUBAm0IgDeioVi
GY2TWGEtftKvrUW5Hf1CfY+D5dpV7bQty/lipP0Djw8d79gd7H2F+yF/wfWGRxAh9ozF4vhZxTxh
trAtA1vEj6LE0k1rvAUDvFMLsyFD3f6VhcqDAGnuQkivtHMMGlGAba9gzSoWv4a1I8mQ0fLwjrDI
O2PiSL9jB2wOSVbEY6rkB0oDOO5T7Dbak4g8VAslmVcFRFM5G0Pb8iqC+EHuy5sorqszSDk0vGL1
Big4z6HJrIxvViqEvXvR/BIcaHorbEp6Mq9pdcYIO0SNS7NmKQjO1nMbxRerbCmlQEdrR7HHC34n
mBw8h4ypjV7OIOq5iGB88M8o2JnFIAL7IDdj/1JqmTCn/CxVQP0/+12hOznDRuRXWkGgHfSE2oyU
zRvMj4fYsKt2xzDoPM6B1qg4VtnFO/jxygqDc5XLCnhmrRFZ1zJQXiMiifkLkycNc15T2RA9Ig+b
u/J6DULp52dnvncyi54u2tZFIOOBG34S/ndUDrq6OyjrCuL8dD8+gWeP1T13XaqofDIId8/cmiMs
AAb9swRSm5Hl4IPZCyb7g7rm/TmiwQxPyBLNJujs1pd1Ss1DQAcK2v5XcNDyheisGocNTGzQsX4u
f5UCS+JdpV6AbcJYoS8EUcTN9+EOr9cm5kfe/FQnBdpQ9uLfhAWgjK4U0LTm1DIMgMJBeINyPpaS
c4IAqsjmpQG90Cj7KS3h8ucxDXrGqRwJY/ZQBK55hOaxFJMfL8yTLfAfq7ed2KQ+a4alCO5VNRhh
0CYDXkKd5ycNiiav/O2fgfGaMvueD1v6ceLIn+aCRuCq83gNspTwSfZ5SVDhJ+k6sOuegUJmbeKU
d11nlRBoXPBtfQh6+8lcd/3jbkYFl/ZW278RgThD97FqZoN239W7dqYevM/Th/Dc/S5xj6rarT0l
9tUy2DfDVQNQG3wpEy+id6WaG53p5MYzWKzTdxLkYmskDZ9VtUQzsM4YT0/UnAB1V5EHF7UO/Ng9
jkyVCWio/gNfWytd/yIF68bK2azKtvGIrU2Spd4xvCuKHoWJBjc6KlVC3g885YDWf/2YxstELdIF
f5Y8sx7eg//02xDzGkjiLH0HW3jDljMR2KioIxD1KUjyAopYL/TA0bZUEU8lvMxafqqWRNo5lLU9
RoSB9nksq6VNj2PVBn8N9Z58e+z58gp6BIlnncaQEd9m+d84aYIGQ5fnd4SnImeFF2+oJKdUsF0t
kCmjbX0hkxJREPnIMIzY0VOrvVJt28JAiN204SE7iweD6C0/FIF7fDz2TNexVDsOLKO8+cfjKIIh
0Z92TaakBHRIAQnbragbHcdK/CQyn0KffhtgcFIve6SVbosEV3WwhflPAA4GsCxnk1PraZrambIO
uIrvGXmhjhKOxW8yuCySM7J4b/2ghBaB043bCpGe3n/mG++0WlegyoyjuI8JXBlzGgU/7LNbvy16
cd6r65vkJwi+SjbdWnE5Sl9a2l0a7qNU+ShtThwz2ps2k/R/gy76lZM760VsuYpQ3Hz347ubaAnO
JaPcW6zSBcz2GmkvZks4B46vy/TMblBZnxzEfcxFt4XYF2WpNVz80LZcEZK3CzQJ4zCH7oiMd3Hh
6HPdfwzWXN/+YhSvqbbb5XSo3EYx0CZ89NceTSZgOaNx6OoG5NrDV8ernGNlq3R6zWFcvurts89i
vxJUihNkQN42fSt8C895rQcCbdPriPyrYZHFnbuBSW4edqgRrgpjKe6Gk1jn9KBk2uLxYwPh/+5C
jJ8Y44qz5sYAwzPV0sOzMbufla62xNJCHOduIQcfWxiLfLqjwQ4gw8oHpaBdsn4k7qlam8qAqTLx
3wv0zHEgeOpRTfzPcsJS5Gmyoaf3oNZO6zOGg78HJ8atvAf4xW2qKRRl6T/dmWtQFLfe6X38ybyw
bRKrHkdUbkEyi0v79yJI7/mYZ676Ul19E+XloP4PQEEe4ND1U/4ZlfWktwdVUu+JlCalT3IRDNkE
ae+u5wSUmmwCDZV1Y2VRbJBMqrE7ZRauDdDY3gCTvpz12Lf+qt3DDeKh0Ov7ngzZpvBTtEsR8ZgB
q44tiOMA3j9byoqIFrAtc+jjmNJFhL0wiLq6Rnbs/PXaTdhbO/jIH+o0PWzf19JWI9eghzo3YvnA
TKDo6gjiy4Le19XxyK2RvBZdPNzsgkcN/wnDkmEM240+0g+yVHPNEmrtZ5VPB3jr5G/8nkKFAhgO
0LUBFkyOk8k6+wyhxa2efarXm63vw1HpkbV6RVMlKeamlXpclYRLgLbERwQ2amLhcjz2qXdFZWzh
Qe4n8Iu9DnqAok0ZF6RoIV6aN00wrS+m6SNkT1Vt6H6Be8DEdRoPcO8nAE/wNyF6E7Vn7CahWsGN
ifD0M6JwflKjNgBurqgAJ1vHvqQvyPnnGPEIfGS0Mw6AV3dzjrkyQk6+AN54qK2JEnjISsgENkdI
U0/4XIvPCCuOnF0+iR1xuWi4iIygt9QVQUQSv6UhYF2L+2XAtqFA7CQNFZXdeA==
`pragma protect end_protected


endmodule
