`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
pHHsWlZiMDuZXgp/om2LD4crIA0Eb5LR97V0D358l4tNQX2/Kw9tSGDgFf7XRl63NZ4OpuYrERBG
k8UhFA6NzaT0us7QJMZlT+Yo7j7yBYgMG3QZucGNEK08UiEE3l7A96QUlSiIJg+MhJ9RQpEDHE3B
3rmxP2Soy5j4yN5niwfzKoAz2pMtdMdXHxBlnXG9W2oHUkc9QE4mr5A40TUc0thBpVsjiS6iY1kP
mUGYJcDj5rgnFOVaG1xApFQ26fDtU0hekFk1Wssb+bQITr4zvEhkjLmy14YM+aY6awLFz1ynsdak
gJ/LaW7mJa7Nj3e72Uh3cOelf6DfZat2CVkWBQ==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
hF9i18QX4o4Eq4JDjRc0pQvAICDaXt+y6V3rDkv+JupQrmnO8MQtclwdN8p29OXU8HeMzX5IP7ew
nEHhEJKtcbrHSDGpJwC1vXqhFMy5vgMjGNWwG91pqX66dmiGoj+67lWfd6YNY3NVLuBKHxsJUXBE
naJHHYtlevjXLB7YfQo=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
abVfOzcXAnvp+2gENAh5Z/AGszntCdJi8FOPWrGZ9HNBx1bgvmhggYA8OrAmYLK9XObHSOQv6/Nu
TnjuBvdw/rqLN28tQHuC9wdjyDkVhLZfwHjs7SFGemYaOV72LuyPIiNodPOpDpNzYsGI2Wr3/XKR
400Tuk86OwVH5wm8SuY=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2704)
`pragma protect data_block
moEs1rATZQs3upgSHnO1TdYL33Qb/+w96ICLv4X19b/8iNtYEow1Bci+O+kTfz0sd2vO3VMG3Wv5
+XXZ4lhDpSUY7KTh/eGImbRinv8sHle8YN6R28nLvdcVXdISLgHQdjgopEBRbWqtzgwAZk6ZHqdB
fCrsq2ZpYFrKWLnOuViyyHrpPMe4yBU8DMrArUrMdoN/VSBt+78rRmJzmIxpy/dZSLYPj388C+dy
wRsFmaKHF3h22mmveRj9ZDmEBDfDheEIs4HzscvHSCSVMMWZzbC/9P6prgzhmAyFKGIKa5dqRAnh
EpSWPyTDPMBB4R9ZkDxT+TbphVAp6sgYB3zSugkPTH7hMTr74HgEiIbgavNGGkwPdLPpiPiv0Pph
jAUPMx88ZbEDid4ksUzH0ixHej4Rq/4B6GP5h6lXbEiedKdoiN7EC+XXq7lKghLSxSdP6lm/q5xM
OpSwYMB2j3OvRJ1PHgocGR3Qhc3r/ZDElDkg+DqyFbYAh2Xc+gkFDpKaz1lz+b8fHUluAn8NwWSd
GE7Oi5U4JzPNDc96mXOL1jws2f26sfFvMjhd23FaCGVJdQ92FE0koSpjhapzhmLY+uLarJylQVkA
KLlooia1/BJ6djDtmduA+V3mDaQ0bVsRPDXfBwfuAH0rKzMwXCJ5ubh3uyRW57Dht7/L9BB/+B98
YTx/MS+mdc77rUtC8dyzm1dP+4Y8qzl0hR9GgV6zzBXy3pjo8OBbTJdj+FAuK1/onBKfvWatE+Yk
UdQBdz3RSdqEVI+PqLBBQooE+Jue8XmdNEcRi3y2ooFmuhU0EWwD4FMmkoGjR4di+JLHaYfWn37l
9qqcSZWkOQicnY91kaGGXI9p4rksi8L6m1TTDtNqf5/THN9mizWqUm9l8R8A8hibbdfBFfY5Tkw8
Ih4cV7dCf3oaUZGCOYHJCBmcVsT1xUbRWvDrvFDYz0JmAvkS9Vh9KSPjgWpo0UrMP4F6Dpq4h7AQ
0lhGUYFhztya+xErJuG4qN/1x6+45G5FbYhjGxv3HpI+2mXqGI/hCFMLeWyuCfY8cuqgihKHd3ed
v5gEZ9qPXFUFtHOE+4SWQ7afIgYRENA52Mblu93KDtxNzdIM6zmFsTCvYrPvmNtDh2EWu2lTKzJK
/iJjHhVf4KCgHxyv4HwM62eL65Cbl99rtR+E6SWyoWIPCIqPMEV0kV7Kir/SzstRBSjsIl/Lj5Rc
IKBvsu7VhMx/9uVhC3QzyfIDelfZAstxC8JsrgiMte1UR/T4bUOd4aikT3itgeLVCAafQqQpmMvp
7gBGvt0GBrpi7oqOYPfpVLxJy0d/HJVij5IzvBvoAPbM7VR2yVbu5XvolbJyzpktq6zVdxtTukya
v9eJmn1SHGtgqSMxwrVou4h+oE12SjxNmn4uuB3uQpt1kfyxac3YTVyTulwdpYNUHXAjKNmxZLSZ
H8yTHENkKL3UIC5q5Vo8xZf6+Oy/L1RtuTSVwRLx1rmGTtOwxHTYoIyp5IQ+IqhAwYGa92cQj0qG
N4ul/wXBE6Zj7et8V5bV7/ReH+yxla9D5VfKsFzG2FH6jXci4Na1PeufN/zMl9ltRGYw2hIjvokS
zZPuRQhmPPytQZZA6rIbQ7YvzoPfi5vErRxClBm7XVM8Lf1Gt1On/O4jS4IUpwyUfqHhC+RP/wbS
vYSHOcoyRtYN7lzXEpYdsctvoA4R7xqvFbSyYuopW+QgASW+v4sI26C8OPLw4ACEEsDnle/jqXSK
RMKq1LGA0y+HYeD9AQqjVeE8JLZCqESmumOWOtvwz0Bb1xUYe1isQ6YgBwb81+Poiqyew0uYtLGP
K3XtcsNWE8r2bQZdwmSYczgBi8wj8hxAyC9nS/qVyL43pUd+lDwsmHibpSFW9a/o/AafUq2Y0fou
W2HzgnUmSvf0/7pEmbOyaSRbomY4pvaSNgA/R8G7iN0zZJLenMGfHnya+Uv3Hj3hKM9Yravw+v6p
MQGVO33nLp4eqzkbNOsP04Gn8/S87UrE9ZGR6sDCq24h/mkAJl0yiXgrVPQQnmRg9HZL6S2JtMuk
anp7j3UEEnCIxDL0f58lHADorDi1A4kyxtm9T8t7R9RMHdl7X0nhkC1im9xFnffFBbULJbhqS+J1
iF58y5pARt3/K5xMt6Jo8HgZf+t0mhrB25de7Yv2g5aN/Tj6okAc4W7Uu7gQ3fb6DcSRjw+xke8Y
RxMV7I7TYhKVZqp05S4SgEciVlntHmO36nnK+z5N67hrR5/Jr6pjOzE7Nuk9MMhs/k7GhjD80Nsb
MVgkiewInII/L49LGTqCaXnyBv/CxII5l2d0onzSRN73iNtG2N0hFEfnecLvHE1rcUtSJKezd3Wm
mmiBkLTkIqc8xl6FPP0uuCSth+HM2Od4xZ+1IxNuAf8yDPqbeQHaB8FMbwjqgHvpKiV+pOTPKapn
Us99T0/FHK2ZRKVKe7IXr4e6Th8iaH8nf/86vTbJmi15QN5uy5XRqEV5elk04rAHrwcqbgBN8B3b
v6jexnXOyMor0FDnKwv91tSMkU8sAhjUWUEhZEKtiedOe84Gxm2mtix66hUdbMQcpTrzZbBxZ74M
/HZHY5Dq5MjI8C4+ARtaEwFmhKrj9a7gx/oHaXKcK2kxqFNU3quq5GkqDuwA896u2LQ9UAuaRs5W
IK92uX09kkXakSOlEicL8eDi//1bvSEMkkbuCPSbL8GagcsvXR/Hkb2gp43nTUMjAZNAqDtXKy5o
9WHyT1v4XD18NYWRp3l4R0BKZTXegdHMMp2vSUUhFZ/UDyasw+vYkiSUucUkaPKHW7HeLsFc5eaE
8erT22gF5PSA/+uCZSjMSuv1FMEIZ5eQFRf2bGdhJmBUcQlxhD+EN+ZCpomR0N37XE/LwqH1BMuk
A+1JanjlwfF+WjC5IfZ6IEPOVnJC57KXRc1G0+Qc3s/COeHiccY0i3vGZuur+DK655VEjveYmeQF
h1GHrSj8Ya4Gaa90ilVA1kExX7+kiaW1YEgPOplGVhTLkDCE6HoERMDqtTRFHuU1eP65b/LT0Ij8
pVs0lGRZmIKAqFRPQhtnc90+LXLIjJ2Rei+31i1NhRUiV08Ypmhqc9+pg1fqNrrvjR6068YCscT/
ancahqIS4/mMA/eNkpzMK54+opcUOzJjRf11WP7dui7b8M2SuaVvzR51vX2ndNC1Hvup3xNtkhG1
9bFw49lNlpencvIWJMewu2bx4SE9bEfav/f4tK2ManyOMdYcD9m2kyJr7CCYAD/D5XcBQYap6rig
N5BWm+QI9OqNrMjI3CZbH+64P/8c2zRSqDvM0egcfFt9wh2773WWqZT43W4qLa5RiDtU0fbrGCy5
lSWhxR6qqe9yUQs2TdNjzyOq5kevYf+tYKxiEwkX501vB4yNwcb4LXXaX59N/5hEk3YiHZwaYuv8
wgUu5rjtJNx+HCMORxu+mxv9YGf+U/61JxIcIlFDMmE8raVMWB31vEmfJp20iCVye8gpvKc+7Pho
gz1x69XobWsmjmMzxSGOPRNwMnNwmtTBeuWcSDR+dVamN/tV7tLLz6T62YnDNks9GzGXEpsC6+QQ
eeQGBCh/Mkt8pAJUJRPbu1YMX7BuqogUwg==
`pragma protect end_protected
