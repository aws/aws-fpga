`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
drZ3AxBUT2RdaVGKvgFr6OwxjUzV1BvNAHiDiuKvo5hBxGE40Q/jtOzfODzCMi6GgD0YndGI0xPc
SXWv4f+4u3KnP2I9HVzg2lYdM0lvVqoDV0ZEEbwJxOpsDn9rIHjOSNqbzr+YtUnkMviTauRRyWlt
eeA9UDwzAxp2z4qp9+O330B8iNyGVCq2l71Nzojz4s68kUlSFJKYYE7kl+XrYNVPw8vpRDcZiPY0
u94KWVaaBonI+sTNr1EI6kBh+x4Rxbex5dm3+Prd+EE6cqlQ9wN9xbmnWjNvebOUDMOtXzlTtMyD
eFdaMLm88AwFzpHkOeY15y3ggMyTl8kcSbhK9Q==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
C2AT9kDB6MRhX1NlSW764ucT/9AjuBNPTbyWrmhHvfMA9cYnQdgXklEEgMrFWfmFBCB5yjTOLQb4
sBMZZt3ak9rrf4QWG+Y80F4MnZfGgGVTTZbefR/fkPQ9u1VrrN70OQPBlWhVHictsPXc8uCATmQZ
RG6eYRCqQUewtX+okqw=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
iDkCSwFh2VBGegsQbJ/8z3X8/5crUIh5/YFrow68YgyyHUhBsQzTNfzNAYavWGh+DzsbHiNVn49H
acd1K3DdoFcGnnmFQJ8X8UshIh3xVhqNVSMEHuBGOvWLBTFhUqadUh8leO9Y3lRTDsiMDEXpw+7i
TPIH4TbAGFG0QolJRD8=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3488)
`pragma protect data_block
s0rEN74PkdQnFT9wCHgBDyy1ikISWQAGc/PCpJbFv1pEzpc2gYyyeM3biks0mRfH8TKY+G+dduOb
8QvkzDir08Ro+K8mq8Whgo4ReQvt/1Fh8qvJBjwKxJMarHk54WiAauDXWDLCfsADkXJrxyG9w6Qv
yTHTzEcl0JX1VIzIu8V8d+hXkYdg5Y26491+WJnkJMiNwwlhvFmtZjZ882IAog+thhNyjaS4o51C
bIJag1SOIJHGqQKjF8GNZqCkfbD83Hy/zLUCeL/mLQczg/yKEkRmVJcV4Kyz5xI/PLljzEBdxp5d
+7Y1F6B9yWQRKaT/IsGCWXai5Mw67H0a6TjwCNlj3Ypv2OIEH9kuDaZ4hFSGL3gZJE0VGjBlEuRL
K0uAr8dRGY+UFGeskl9U8POJGkq7oOLDXPY1Ibsqck0zRBwo5YDgK+cQ8I4zv6W0T9R6ObXRZEh9
yuW89lBwPO5JCmcPevr+jtRuoIqecwZwjZxs+pNZ4xQJa9jBJnpQzmcdR40w1BikRpZa4OWH4c8k
r49MblYonWvrm135gsCRGv8COFYh/vjp6xYJ73uhDjPIrgeXm2oUd5MAynuFLiDgksMmBYW8YgC4
pyLKHDC/q8xvcf4YYdO6g4qoG613EMjOPBtlWhDjgHk21o/+NI9Sb+NNe1WmNOTWpLrD8AUvVVZb
+EOXhrZnpPh8oW+aOvKj5ezIrJPjZ/TPMB/aVQv5dzjy7ieBYTafQrD7e5jElLWpX4KP4g/nrHv2
F7ZW449wMOI4/4otvcHyh3xT0dAVmpSNw8RyEtuGFz54Ws3tYuK7Ac2SYJlUB8A0hPHqClUnunZN
SkseUb29JV1YYjWxiOe2k9IDhIOcEwP0gxEb8Ht6nvL8U4CZkf9RXvFOrvcF5Gxw93dCntWGdqgQ
Halgp0GdXRkVkHW58FLe6Kdq0BXZOxBnMl0UJZZ7y/aTkNgrsfjWC5hBBBmrobvcEOdXjr+4pNuH
wfUa/vgoz7NFHHKnhAO5YmVw/dJ7IsrW00u32/rwtieNc/byG78MboGP+24tMQbJHVejoKpKmkna
BeRbJ+fHBvboAh54Vu2748aOpydskUmn/FL21zKt3Vmmr9I95HIkvXicYqz9JtyAjvtJLqR/25Te
TS5+tOS1S7gt2xqaR2ozksyHJC3kHq7idmfzKquihDOeO76+RB7rSoMfAtT2//Aj7i0GTX21DCsD
xFXmKPWORV7ISY2cmj1O/VeO+cy5M9/I/Wr3/37GCuM5DTdMS/nUE2Ya7hZtuw3IrUGvuuVWWiNu
/mWDcmeHmV0Xc8SCV6zoqZ2PSch3kaWk6f9FWxL6hV7Yhi6JVVe9WGRmqa8u0nROlcHoe6MvHf7F
doxyHEyJ2Gap9CxElhjD+cheWJuEEsLWb+sPDd+WcCebRO+v/cu5yumNWjrGjsIJo/6SAQ3vAaYK
d450dePOEdUf7IX4fNsLO3Wicu6KbL+HjUJ3P6utAYKI/T7hBYNQMnpenDb+JepYBp5ACCB2tDQC
WuSvAXN0rtd8OD3oTB7vC0pWvOO+qsRrZd3GaF5JSfrd4I7xd9ZndUXBJhMZrwZbAGDK6orFChyu
6szX8OnSrYOQa3u/J45IzWE+7yPjGEznp3cxiqvXEkY6QWAcdpaBNcnZYcsjk+aAty10bjO69y4x
i2S/zmjf9JP138Vo+bPl52JMWzCSlu3fGGBG5XghhOtW7goiSybMPV+bF9LiLBCeCEaMqerV/0Hv
/L06fVpVOnl90myfzVHiyyLp0bXul3m61bBXWQ1xp35NYbRh6i3v+gs9WEnEcNZaF62wQ532aJeK
2QgLb05G0UkYDNtw2Bbo2mAxspLDoffeRzXnUjvGWpITi7lYIafvnroPULhRhUphTfZeHdvoHzyk
3+h4wgdBbPPKEhxttd7xJTQXsVQHrvXZmanLO8dQd96PxRmNt4UVAvNAHgoTf6uYGFb9gkduUZW0
InTcneuhFTEwLqq++uWzzmvPNN01eaWKrFhiZNwluG2cbzhmyg+MCjeGBT46xU0WklEcKWXS8s1/
Ck+S7opgIIdZ7Yj4jwYfKAAzHuggi7EPnxc6n5cGWqs43seG46mNFemDCupvYlovs3zPA+O9ET1E
PqQ1U7sV7eAeJ6m1hfq1BBBVTUHO286LduwBMLm94YBkrQIVMPOnwH7IZ6teN3pozsIyBviFQfcj
KD6szjQF4Cn9XyFZGz244oOloX1HTE9X+XWoK4aVUl2NLbvoRffD+wkZ1Y1NVh7FqSL44dRilDla
6Xo46iIP6cX0oLgeisSTNkZl6tzIvdqE+8LGoD69a4SPk+AvD3WBHg7rJXIDbSGilFeL1aury2GM
Rzcz4K22DWKjueWl4j+1c809xETcEzJeeptKP0mPx4fk5/rz7Wyk97czeiMJ0agZ7bzXtodM2o0J
piwe2Nk605zKyzUjs6MTlfKjPDY4k1KRtZyPDky/Z89DTPIbhweE8IksSs20P9krChk4IRrud8AN
ADFCGWjiVQJNcmaL5J9UqzqTZR1OquSIV77pFxsYiui9yQ5RL0kYDnw7824QWqJj4lAhOJg7kKrq
osMyrFsFK9BzZsKivrFkrs/yEUmJvly8LWlzIWLjwKWDjI3BbYdeedH0v9kO9T2DTAbJgN0y2UwP
BFSvO3l/nVZ7eK7wcFpqSgd5tr7EL5VAWU44Mv8ahUrXtjewbcVP1BRBc5kuwzHcoo8xh83Uk5rG
H+Uzx2mzK4ebZkf1gpILIkZZ6oflOQi59z2A7/fjY4i9LkZODRGVnMncnJOn7s9jcdZWhBWqfUYm
1HMNQZa2eej3c4ygovG4lsucJofEFBODsMLzqmeCsD/3SyTYCzB5VaXQTwBeRfGKLGvGMogv9p5d
zAv28KUbxMPAlVL1qSZ8RuynkJiJz2e5TMQhqb9eztt0SizED4sYrS/IcLA72AeDEQCLu2p/v+i6
acxewIBBcVxi7rtWMrg5yJjV9oaNzNPvh0UAvdr/qQOba6pEmKJRYHOH4HUp5z3Gp/TsmXiI623r
kpRHVCCu+twfUrQxj8I1F0szc0gFhzDD7+1tkK3/cipc1xdyo2S0rU5zDHFd7ztRN+6NiODeBmmh
067c3xgCLiKOSKlkIkPt7xer9fGwJgXvQzp5p29d60LphxHX3HSG/TlQEtOhk2jusK/WvX5AHYFL
uYNe+fnwI+ryXgcXo1kKQZTIkWt9+wwZuM3U0EMc949wHPjOREvCYBz/mekkMfoUJx0OnghFwPaH
ZUcx59GkgV81fRWpgVE2gjHoICYzyE8vqo/q2ixiC2SzzspgyoC/e89eIDy2cjY8Up98sv5MLP8B
5u69GfgczlHVfdRmWTJuzqGwG+zbM2LOBjV8Dh595nVin+dZ08MpSHQO2iR66cqv+UeZ+dA7jo3+
Spmkzn66PoUI/pLDGGStSA4PzPQ98iy/ePrBP7xJKQrbF5/9zjtjv5m8suqO2NMPR5KQQjjOiRaZ
NpFkKTpq0leu8hU3epaUNqrrviquY+sh1Qn7b67PzS5GJrFHIjoZ+TgYbtk4oyRoCBlHJqva1Jpb
qk3jKpkIWBn4W0BwFwqppEKnXDZZGToSvICAx5tCPL0iPWRLVULH1WCig4+fUn58K6Ry8mHGu6Wq
JroSJcK+6UtI4V5J/KDTblP1yV2/8iciteJOjdyy6hrJvexyBG28k/pSWdZU9SsI3qT5pHQ8+y73
WP+QzkUewCdICcMCYfBC64DDjGRS6I8PGRTwqsTKzXmAuqgorCv47K1uZcmllIKF0agsSzA7xhPf
62DoJCrbnGsioAtQb/JHcEKwOdcMM5VdAEKrcmIpRzfLNAitzB1pT3zlFgYHKKMDHY8h/35wgi36
Orogs8ogRumGwYkeBDKaNDzepERtlyw1cTiqGe21u46RhPsm1RjqRpXw8z9lYYimU6C2qz1AiKT1
c9ekk/cKnwRXw/VZca3QHlgzvmcVoqIE9Nb98iWQ/cadRKUmlsiiYwI1Oruwo1gCev0jYdLS8XX/
6mjYII7YVcUQb7Vg/qI0VCKSLKHXI+9VhHL5LX5oX35PjdZG7Sw3waT9dlyA7It9CetZrDxowWUh
TJYqgPc/QJqrmH6LQFYwUS5nbasa6EJ0JJacMq1v3xcyRIGUTVBJRgGWuW+Pz9ssslMNBH+7/00m
Ym1baCTVvu+JxMBKrc54guheC6HdkIhrt0CI5X8h1ruxwUKsCP1B4nUJQYj9qyY3WUUmhj6nQ1lw
nWIZUUEx4yctXpSk/nzJgJjC3YpZRauJba0l8BN+0nFjIk6RWdMI4DiLXPp5jefDO+qev2iJ76c6
nnZK6oOPSvjLCLzI3hpeo3E1lyK+X9cyYe2XYghPiAPcC1FgmehwBt7tDiUd8chcmawgV5/wDxXQ
X+32uqVNoc6Pn34pg0qjMocYCof/p+YOGGL8UaQDmgxmF6u+eQCT5gRxpztJoiBDlUQ4WwmjLqzH
7AjLc1kynctFD0aRq2Cih2gRkIcRlzoqzOvtjNedIFLPKMNj4SOgsl/hygfLQqmjLZKSzMTitU2X
KwkqzU5yVaU77b5YuHtJagfeCabgcwG4zTf7DNNg830/3tecirORGtbnjvEwYTsys5EypFGiRc+l
++1FCNNhxRjbZgo=
`pragma protect end_protected
