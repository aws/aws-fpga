`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Vlb1+jzAJkdpYoo+9Ef8nRDJW7vEaeXyk6updoKJgXO5c9VRCdznjETTfqdBVoZnAIuc+Zf348F5
cwgHbYNLKREWB/WCxyvannb3WBrFtGKEx31J78qI9OiFPXNnmIeFNKN5QdxTkUCUhQ3vZs2G8uYb
Rb6cwL5wwK/dhxOmMxFJbWallTLB97g1WP9JXwRKRvGbE1pOv+9wIbTrUUoWXQM9l2IM6sGf2LuE
7pb+2eQ7jrRFsTJJKHh6ry4BoXqyDHzeGBi40iaLDP1a84GALIlpeN2hxlFdRVpeNsiQ/0rLa+Fr
69Tz5Bv00BxJ5yK37Fbh9kvmfw9vh547HvkcHQ==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
qRe2HWSp9V89a4wQiGXcBscE0+d0JrAWsudQz8Ko5pOuCPqrIOkX2/SuNfbBMFi6vglA+wqKLx89
G+YJ5/xKp0O5mbiLqojXcPwsm77MaPny8HdJlTDBb2ozjgwp5kQjlKwh9joFfJgMkUncSlkCm+Ex
qzby6NDgPhJGYLazeog=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
O+jVfy3F7v+Xx7RJ6m4kmoHIzo7Tt9AXXgciMUtq67m1C3pSfJtv9olMS4LQJfTWGUnakruG5cf4
6r7P4jgxY3kGfEyFw8Kj5iO7Ad0q1XSLrlHUCr9nomOWd9JyJbDgPZQshAZHmxTCxradKkEJmkzx
MpdkPYPOVvl7O7EiVY4=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2672)
`pragma protect data_block
01hN0dqP5ViR17eqI0pgMc2LJhhywWGZd9iuU1ASxeHDeFTl25eXkdhjCdcyC1jKZ8O32VC9NB9C
UIU4bZQ0AGG5j1MXsW+84Qp4PEdBsC/KWeyEhWjPYjqWXeC6jyQommQyAwC4WrxdKz0t6sHW8KHx
/pCyrKKDVdi3p2VD15eNSGpY7jhALyHjngpBcoD0QzxGY7KWaJsCmg0nZYKlmwP1iGB9WPR6CK/C
LkcFISD/3PxMamlmnr48tsWwCVsV+mrH3HzHi3AIe5a9FhROqiCp7/n5fTYDqpAMi55CTknDGnho
0i+XQK/zpDs4MS+FCxiYMzJpa62Z9N8VD/j7F7ro/934WlnrHgPxZrvR58FdmwLSfoXq0ZgY/RiU
rYkpu0T/LoScqn8EAcIq8X1Aagzvkm2ifsgPLzcViBAPig6W2D6l4PPCSSh47wDjoL52Aj6n2C8W
OumHLmMYWOYT6r8V7y/Cw+iXo6H0yCASLZ8pVO4zkl31b2zOnrivfDg9rBqVLAv1UGm8yjQ638BG
qq23fknZ8E90HMeEhXan/JSX4Te5EtI45ryWAMT5OnBscZOUY26DVHWok17NjJnHoXsF7sqiT9AT
3MUfJL7vpn4HYgWQC9ymst4vY4JnB1hFix/v521HG7w1Sn1iQ0oKJRCDkhECOv8c8l5bvX0G5qkL
DiOKDkbzyB5RbVeJRXq3Lqoem//EOefSiR8Rpe3nEBKedgxXWn2vq09Kwgc96TTQh1p6IwJDoN48
vvzxAhIsvjRZQMRrcEUXRSdCRWvmdrp1u+TOA7FkJ6uRlYfrfD+DnGrQt0s6PPH5BrmohVgY2WcG
s8MeiK3Gd4KH8+mt96ty5GjM096AYAUtjNR1or+5d7QU2IDumrs+Zpmm0pZ2v8YFBMQKog+J3y4L
na/Fasw+OgKhRl3Tu9z6plJ14iOSwCVVZt5CBVk6zukFaXpXlkzqQ/qA6oSX+xUQWDHUcsC7jbdw
JIGATdM6WZEVCFbPT+rUwgAvU96AVPf4TjI6iS3W9Zf+jEQ8ISd9ZWkqCYWy3f4rjH47bo+qKRZS
xRZNjpJgOzBl72H7LBtisNdndsCthsXKb5eyUQzdx1gftG0N7nUOpQ1WDmq29H4CRPSGxYLOrTAZ
x4DaIJRz2XWmKF0yzD8b1aVJib6PtlLrFX5Y+LRLU8S/LvxGg2Ble+dbG1QU+yyKjUFLjoYSE0r2
IsQZHqQhVv/JDWf5MRqftoaKNcelA385sMQ0EmvBj6gC4ki2L3A5cJS9Xfz7EUn4kbV0OEEQ3sn3
IogevWCDzfNhUHKxZowdBI8WZ+NepuXBjrH7bT2yokKcCObEt+urc9DOYLefThfMETHwxFouGu8I
MbnQkxAPwYfoPXW8BWELKSK6iXdrkiOWR5M9bLdz8gKS0p6HqzYpBzimLspCzbiTtaDa/oectpip
FlQ3TXrpsO1ZjEw/f5BqqiI99/28zXeSozF1idQXCoava6ahr2MeBJvwyYOaWvxi6OSoeOJZkdsh
E686CLcff3e9cQIpkSujT7uJX3OUoQS3OJIv/nZtqWyJV8VY/Yzlw8t8/f9n0ANS13DShqsP66cJ
wHqiFaumQclNShGDSvjUEpKceJYi/TO7gcF0bapY5pluC5XTeltrxFRrfQgmnJw7+gDD6vo3jrce
Enh7x3zQS8BGVItgrUoK41aoom+N/rhiQG5IRFH3/8XF2qCyjqMMRmXdSmh2qFp1JlATUUF8gGvv
3XG8FAx1h0++XRMF/ofBbfWg9YdCsYYBLLoPukznq2uM+e8j8u9ni5yoMTD1bOxelN6RDI9rQFO7
uwx3U+S1lltVokikLlw+R+MhrXgXRZTdIjnmbx6w98YJj/mgTPB71EvM+FY0PP16XxS4JS3RFRGO
4Ghc7X3viDmNes0RxrhcWcKtCSqR4SJ+thw/7IYzuHelCrDBtI8pWThhhpSfTScZlmOzgyshGNZp
onuLl+/bVWcYUbNYC6dIXxYXed3yaNpBYJHGS/kFKmARK3zrja4KZcTyDjdd/kY07NXTPd/0OU64
dU2tTe7II6NYAUpMgbwHX3uMfvCLB3wPI4r3NWndsTXL95XETgQFDQB51FpIWbbi/TYdweA3+Fvn
qxMpg+OLVjBWb4LGX5IIGkX0/+Jh9SWtMXLp53j2A7FvDcqh0tx0FSDioMpaqy9WXgWEJuSyU3DZ
FcAMIqPaCkDJnx6El5Cd4YdI2zWvOguDSulhsRwaBKvF4OycfEshw/jpsQUuHBIv5Bpsoafs+ZlM
+3bj5Hy9tPQzL9VRTbCfnOZfjPEDodLZCdxtB2t4abJCCkRzblg/x1176oA7MwI3aol/wJ+56pnG
GG+JRyGfBT+byVseminHh2gN/tcxmqZ2bVJvOq62EWMvq5n8LIvx00AHoB3HIGBdVJJ8Mov1R0iM
Wl7bxq0l8KhCGK1TadxLVk+PD8nK9RbdktR5G74rGiF0yCcq353hgAdLZi1+sbXU1mbed5Qsf2AD
6OOGFubdjy59FYt2qSJpUDqkZ4qc97BmX4/geBraGE6gnNnMtP67EYcIHdqokvf0JQEZegvw4Y0a
DoL1ke/ZrsCPyIRi1ZRFWs5nL46wItwReDFESfNzwMH/+SzFoq0u/hf5MptGwFacXB10I13RGjkZ
j46F3pgyfJyROq9S/cFcSKPSMfSV45DYSXPu/LODILx3fyVLZk3bAaEtpl3Nq1NbXEjI4r5cUH2F
sq3ooOTsopNwQM1j9gF9h40w1YcD4XZz/95zBkg4Q/cTcsU6uh1sKxvdCirpQosQeZm93cjgoXsV
ucgY9zQwKMewafH3cwZ3UyeJeViPfxfR/7CaBoSH2siRgBOE2LUEaJq34jzDdBMmZSLohm6x5Gi4
AyDx6r3MkilPAlLLAHSD05twCzcl6tqxhCUxR8aAyhsyqB0BvtE6BK0StUFP5AeYtbh3VTFKWtn3
6i3KqR7Qze/F3cCTzWj+tbZ3lAD76VjtEGUJoFccpIQGgWbzcHNLOXDlv8Q0a1WfZzw4ttsmzE54
87bhCETjRF/k3kSHkc+T+fk4lZ82li4pdaEODUoSLSQjxY1XgQwdd8sjnvQ4/3kY3lmnSmCfBYDl
4qxBGmGgWEu9lxmIU47bBiY2PgmF4UBeI9KL4w/+qcE0lyi+Qj63jOtAkOisENc+v//04XKJjHJF
yXknS/8yUSaiA+8Iy6CL8Tx4tMdVEzEuiX4Oag/x9KeB/hRYRoWOZiQ9UG9ydViX8abUoge3lodx
BmyyKMy9l/jQjP4bp/yWTATovvtLK3ziZeM03CXg7Al+eb6F83Ahtl9LG+i05tOPSFOwgY1RZ8FP
GRkSbJDUW4+0doPY0UAGDd0Z0Mk9Eh4/7rpcErj0h4FnHFT4yKemBQOQD1a4O23DftV5fODpK+2r
EhXzeWq50tTnY4KnimsBu0Y/4MvtC7J5pJVqytqlJ8hZU2Qf+5U9Kej96S9NKoILhyNybcv3Lfol
UIuG/So/7OYqqKuUfTY82LmHw2oNU+6l7MxH8uEfUaGTMMwOc8jjlnZqqQrD0eSmiXM=
`pragma protect end_protected
