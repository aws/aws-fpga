`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
hHXkOGIxReJr8t+4zQ+Mkk0ZKJC/pM22YiJXNhJHF19H0dn0mwfVL86TtnM/l3EvBoNkH4VVAJcS
gIH0eHKc3b7hVTrgZ83XWSD16eIGHTKDEwjEI0AbyyJitBOUrn9T50JvvIkO9tWPyIq+gfS1cHcD
3owazRC8Fc9uExNljO86esGwREuBsc6KKZNuh/y/9X0ebHeDV4ZfnUUpWwxcj2K8RuUCcHIWGfow
8dkIwiCPiMDZc8HlujshlS+GU43sM0WsuYyWu0yCFNR9hMKbq+kueuz/qrktMEurCO/sI2j7CK8a
rLcnFSucQQGZj+4NrCQZWHUf7YiGTfkD26Clhg==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
PvIPBcVbKdrAUdrADsQSyj0mW4nqC+8bZRUQS+2Xf/K8jfqfyQcj+gYxfvRGh+jn4RzzB14jOdBL
10unaiw4l+/dGf/rHtMOBQQnhc25e1ETRtUDqCu/5CjkhjyNZnRHBAxJ3YMsaJFf03wTt+wFVx0K
P+vhuoBiiySty/xDVn0=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
eZkZEMeZFqqvETAWU7A9KN78imim7OvrolNxeuzj8MRqhiP3VwSpn3w3tVIlRKMb4Ss3ys56A8XP
qYzEQuT1pjhvzwAG4z7FiV2R23xLlU0V4Gk+vB3OrMdOxEPuKT7OYCzy7FqjHasbQDW71OVJ5kga
yiY4ZJT3fmYyEsWFXeU=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 21712)
`pragma protect data_block
FxojBAdhJgxxTIsNQIi2GWCdvlqSJ/N5MPUar7aZ0E1einPsnR9+OZCimZIAHe1WnWyk3Im4qifO
p85xVZWgjowxj0fqIiQVwVlyPKYWsrVVMiMCvSbTRBqdLhXqcK9k+t2kHk7ttqN32/LOPniNwvzE
pbALVFxRW+Dd8yViG3EvEnguZM15s3F5jrJMZcdG2JG9Po9ufYMtj0IwBsdyRftoGli+7wNZMt4H
RYac09N3CIRUR06xkDW994DnfNnZ+840vRYHmK8mBHZXBeHwUW0rPAvMl/g2XsXLrrPHLrXyksLb
M+rdFuKuQOEnUQfNiZSCAxddqQquend6ZHOSPZqORoiuYyINBZZ9X9SR7pP0lFaAkrq/PmxboP4z
5qX2Ypq/BThU6DGuhrL9mgGgEZB5A0yqUaSw0GpuqnFk3Ylyw0kx7P2nggYyyXnTRGVhWdulWLAv
JU4jvZwjTdfbZTQRD3oDJ5I1PLCVU09sAtgCx7UL53Eo7UM17bmAMukeaIL2SZTMYXnoz2ed6dPp
Z086SpoYsB/VzRv7wUAy0X3vejaez2NTNA4Dt3eArRvK/kR9p2cPcePS+K8JWl+HFZkXB7su5Fkg
sXlxGhx+xVi6qWsm5nO/F947N+Z3cVjPn911hv482+9EFaGaJVkvXJYwe7TIvexcY0tTsyYT2mVZ
pThqHLSj99xklj7ahCpWKDCB6eagmBa5faGyvZ3Uz22Hgn8o/XkKkx36wJAYc/zEWYOALp0lyzM4
9CRraGtu2lfMNS+U8m9NU2KshtbrK1WKSOBoHe2hSj/bwD88EZ8TGw75PvJjRGoGoIGMHevofwnJ
C0eYSyooYA7GVakK/lUq0o1QDf5MxACc58JkSZON/CZzYpS/uSh3mkQh3FyWV+/COQ8RkuQK0jit
ZQWfrBgo5xBUSCmrvUok1siahwSiLSzSUgXsRgi8Bd5JPxTaLGc8Txqb09Q4oG8YgGziSQkiXYtA
j5Tzn5VAW0JUZLn6aSpshW3sd6N5rKy4AC8/fPWDd+LB8G4E5Lh5eOSVmR3nuBHJ2U+jyVnoDVIW
7wEshfX+8H91Jy7jkg8Z+3e7fjT13OCxPy219RC3uQQGfla/8Smdm9nhi5k7ACW64kH1WIT7XrPT
O9aynWwW6VWjHHX7E2ayDCPQ/l167tcWm0ee5S6KbqW+QHMAoCgY4uMgTb+5uJbpTkSIsosOG5Xt
FwLYJtR4V+LsFxNI4qPhbxKqQxcCuaV02R2c9dDYuQjO98UM34VCz4CkFwGzCl0OFbjdVYawqmke
cqs/WCa8vhanf1kGAof/Z+/6irQTvT8bOHPB5YJDXUj5FOF6n11oNX+PdUk/z9H7lf1EzL9sdonf
+8LMcLvwB3JVwHFoiuoIeb/yua0Y/fE3DxFB+lqlqCsi+eajrwbWDfzBZMvtB6k6Nkzjp6UFZOGC
1b0cNLUt5UtZUYpzJql7PDgXLDmM02CfjcZcGjDuw8jF01F/kLBw7nDbjkt2TCHQ6Qk4DQ9kCGyS
CTbL6PCSFoUeiaVEJMP5K9p+RfgLgGaDsWZfqCP2AyvDZcW66ETWSCLq+qBHUEdlvojCQ6nWBdEr
dV6ldkQ5B405+DVSOmK0eGSqj1acijMnU45RYpp868keHrSN1mJU2Ng+vt9swpCoteRuAgNwj8vn
AyWDju4+PcUwJYPbsseyyazyIgiksfaR0hlJaab21Dt4cYIHJF5/P0ezOFiNPesftttzbdXZ96Kd
H62WbqcG2FHHf+S5cR0LvLKgedRXxQgTFdtZa+aQYHpRw/FHQApjrP/WETzBgoDDNt8L7o4Cb8zw
Yjv8o5MsUItsDK58LR951SJeKlIwFO82ReDn/+Nncq8KBnCl/DWTg/PAvP0YmNxRGQSSoo8SPjPZ
fCcB9Y0F2WJgM9DYiEBG7xLM3xew+K82IblAJq2byWHlTHC/pVGTAak5CWoQ0HlchnKapRlx75Rp
BP+jg+8rhhL+Yq2CYCX6guriYrXtNTZOpLG4jzwrnvBzvhX+k8wnJXzvX4oD3YFYl34y0v83ktEv
J3w4MwnmXZmJFWTxy+sM4FbehZ41SmRn56B17J+HyubEfVK1iZFqeqps2gN7W9Qa7ycQBl65l2ds
1uuC5Br0dL6gghwbfAzhJBD/30qXMul8qWW6vBuHqRI//VX0maiAV2cKb/rnN3icyksx1Gq7NqeF
ZcRClEx02qyfNFBHoGiTAZy3rfI0eRNFhotm5KdvAMsBrZEVB5J+WWmN3Ueu1yJ90wZKf6UwIMCc
GdJLtPHnoHFJ6WOm88lxtqDbUvG/DO3cOS59gYw+goy7xTfVxeZhiWB7tPoO3VPrrYXjzZS0qPpV
DYpEQwiG1HnzKTirhtzwyNpCgi4LFIBl7cVf+X9Yw2GZrxC8ZF04RbTtRuPKzbBbYfJHYJC10cbe
pPD/ylyDpYfZbRey/fqbZI03544yDJ6GAbhhzs1VU2+TgkerJw28+m/vFWU0l4oChIY/jz2+Oib9
QQ9UmRuJQ6XpywjO9zZzWVqxsEsUp7DeE0Su3rirqhA4Z9J+hmJXeUSC1NtuO/Q3aNvunZcyVhY0
rJBM6i66QixfS2Y/BDZK5OOK6NRXkXivXkdum34niyikuAVfdjp7C/C3VZJ8UdqSYkBoOMcsHJva
jLsZIYIwkFsRu6f6z17TQgmpuecljv0ikigUldM5EvUH0D8krd9Klfdd2fGVbxV1gToEUTUHn099
OZAqfxdk54HsiXa5ffFx24uRBNPin562hPgbyp5aoh+ZUT24TYnAJHKY5A9GeeX6ussi6YJ2oSTF
B8U0HSJ0VZ0Y+jFg80caJg5Q+ucJ/wIZU146R1EgOw4xYFQjFC53GbmcscAtREYTybOQvTBXln3v
Aqj9c2VhQtPOA7xzwFNln4AcHeiaIxidSGaUtgGq3DMVxI/G65PNi9kZktVVBcW98sa2wC9ixSm/
00etDHfpZSLN6QqSYnRGFRNJlws2XFvGA1SLZauVChON1YkKSLse3QEx+OMnniShW/Ma6RvzUW7b
ZJx+qegrdabtwuohaC03ziNj+zhWk4FKKsbOrzMtFDDskPhR4aWpR1dSzM219syt9Tucxf32Lrca
wP5mYvCOYltIy5Ce/NQ2C9ox+08mVlH2J/k79qrLT3fBp7T6cFGiq0EiOCN52FRehtNUZltjs+Cn
uaN5kkjcIJXIZYiSJFCGZZEN5KxgoYGfKtYeAPeSN7JtNpCP0wyLzhQIB+LDWTMKKeJIyCyB0e9p
7eorTfgCouSwauYC9oNt4HFvVrhwyHRTf5bDZTkhBFyxVefcjUhZ9WuTw+yK64PaHuQph6mSdaaA
wxfCVkbdmoRYe6dwCntpmC+wpY5s0z7WFqy718GX0Sr2zTTtUL80/p4+zljtVmWxEMbNYnYSlKkv
ugUUpE54UT3/Sl8gPOUeGi6lip7HahFUwrQQjQ9BXbej1Z/PohF/7Xo+mZInQ76Jg889EHEBQedc
8epG8CH2vStAFlIkxLraVOUtUhzSlNuZ6g6oWMooqnHVnIrv63SpgK6VkPte+YcUO1vvBCj0oVFX
PSIFcyqnQ6/XTJ7+vz4JiXnWNB6We9voWZ38IdHf32AxEAJg+q2L7HhgQn2lgZULUrmo3FfI/BlC
9WLZURfpZ5uJGj4GFPvNv7SkAMYKdpSY1PUPuJCzH2uAOcNwsMUG8uACx1iEdNVawBmXP479YI39
ocaHfqhwDa4sRUgMRkpiQbMmJraaNkJ+n/yuDrmOAVB5/w0Gh0YqbihjuTKzXt8/gE3MvHod8+gR
ZhqmTXyiJ2s5DrKo6xMkn4ulSG3csf1tE5jWkPc0Ov6hLjXRlYGZwhlbznf38G2bUeJJZZtdkhWm
yd7/XY1x3M5ZGSE/HFfk5V8KJ2a7bTXWzH2QxaHKIm9PntxOOLUxlp9zScGXrs/ER4ipPQNOfxvl
HyJVFN8kytKSGjkDaRlSKLPOphmZEHnUzUPlu70Ep3b+QwJXxk/b63hriK2eIyT8z0obks78QWdK
DpEE6ePNaBNF1NhKyS/kSx1LGGnC9nia5c1y9udbCt030BqBrRS+FBuCHrPYLBX84di1j/tNP9pC
4BRcY+GVKJXavwozfk6TthkFeOV7PbnCWmNKa2dy1kcrBXqJdADrRE57zeu+WNO6GiOqsEJ3rzYo
Tx43VY2dYx7HpHDyO/5aCRyMPZ+GMAgM0MRsGmxSUe8+VSsNEgCi6o25RSM02BRGPBudH+2h0m30
dRiXs+abH/3tW/vGzBq63W9D4tq9hEP0JUlN1EQ40ea7+J2RasEYuGEfBRASUdqPqXgDivEfdZda
ihx380guTRKCB/iCTZH2NvnqobO7YBNQm4oUOsg/rTxKP6XKxMeKM3ZD97ZmWJi3zRakm3W45zWV
gJf/kogQ5g6AoSiG3cR8hB5WyiJBvk18knJlGN7Eo5/ACcmz2mVfIjgsFqUFS75GdNDVKXip6Rvn
fQK/74RRqOyg8UC1j3bWxqEXRVeTIptJGyhAUUTQ9u1uRbkZggV7IuhLtzlTk4shLvkR7szpppn4
v/DDkrApAgdzoIDSBf0cAJSmMywS8wTjc5u043jRYWAaQK0LrfiNW7HE1SaXDF/oWivVQUd4JJkF
WsKbXxTdUfY6wvxtL1EgKY6WTcfsJGFBhjqddgSpBBFoJP0oncwPzw7vSmQcYUN10Mkyp/240Je/
BDXd5EBfKJ8Zq+WM0+aUzKx9gU5loky024TMco+L9MzeBWGrL/s4KFn8tnIiqPKcHdGPI9S0/TZW
laPCGijytiAzvUtYtNphHL9nOYMKEqlLwninwpyuHxShFzS4BPp8mK0Vz1OJMAV9z1oVvW7SXiFX
xccVPrj5mq+99iZc3sFh/QuY1uZjrcNd379xB2Kv9hmy4xFFN+DVAavVxf0GQANP0pDCEUB9JknH
PvO/ssvecmkRLSvErgoFqicVh4esSL/W3XcJWgZis1epRDl3vIWcNIRCdoO9oR7BrYTWeiIE0UfQ
fmmiuonsWUpV18R2wJPv6eKPWqpeUD6SAqA8aIg62HqIxe/RWBBhczIBkJHhJPzcP4yVIh6+uM3O
mA/fD0EzeikrA5x7Vpg6enZR0aqoTEwDGmcFGZsP/adIl3A6QauBgxHMDkPhfp7YZO/hnWgw9+qM
nInGH+DhJTajqxuyOIUjZXxsP+5z56wfQjqZzrmfB9ZV+itzTdKd8mRA3e8yFDNAKfMCLLpqNBLJ
qW6DPp3GF5itz+jrha0AKtBQjL9Heahge/F1WOZ8g3focue7T/6aGfmbeWPZTM234gZZbF/l2iv4
/3lD5bMWZYHs0jO66nDHwOcKdaF6ZjIkL40Sc9pIYzlFPqpEq/Y57ych1MjlzKvHt+8Kp5GKo48B
1QbmXVqGXcVGCJjHuTAfujkTnZRUovADaZjcLccXaFp1eZfAnoZyZxvCX0qHFPvmpD5J08X7ulHy
FQq/S7GleTs+tVt4xpQ3zpQSOlSuTLLK7B5XKASmbiBPm2cxpAd1w89BTpIC+eI+U8UWK76PhsJQ
lTxP7dpVEJg9yxPJpbURTy3SCIjbE3YVNynXz9d1dvluihZ++OfoP7SEx4M6qwYQVf+LsKLASSSU
s9XU6gvNcNNA3YZTL9Spa8XhcgLWIZ9ILMAZJRaxrOJiPQW9T0cxgqQqbZn+lfYPsBmSYqWmLtME
cIMTKFHeIORdIelQllWG9vJ56/KglHell8sqRdWAirHn6A8HHvblttLjyKzLftRYTGWJLTLHDWgZ
vsndxQujQkQiQ/aiYidgDSHfmHDTZ5ULn4+jbW5+Tvmdju4F6k8oh7yXGyvz0B6qTFcrp5tCHm2c
vmviFswBH1AYQbTcGcEZcR3Yly98wydnBo1VzrYto3ubzHZUVUwSbV/+EZiTrD78d3F9Ec/3BJ7x
i60D0NrMMmvzkDNwRmUokttV6Tu4zLV3scloLCDsz2gt3yyTbjfrDetQTCqc1pU8WLGPi9+4OVPZ
gguuCepDkOLvjeOtFgx8txQ/wXYOPwvHmMLMilfDoVwIFFkt0qZu7ouhQkBLA1sZLaCXqKUa+WSU
w7ewLnHrS9fJwUTS0yZD/HgbDsNQ0ioq6CAXL0pwq3m5/a8bbeHqlL+q1viz61wf+iBsplWa0SvE
l0Mw6Gxa40h/QC52jKlC6kfIaAaj6ENDxVn1BQY7HpKfkZIqASz5xgh89i8GHC0vamPTYQeCDxcC
aKKh2cNsa5xSg54t+TX1BNkZbdlDyofwWss2AwV8lx+Ibht5ib7sqE0V/8p4J7+XWAo1jXW1DrJB
QdQVDRPqtiqvvozvUlR9gKzkH98YyFzfX34nWn04IPMcjRUB3p4gMOgavCpeIzbRZGxVi2hJ0Jp2
DDVIMx2CvkRHcjHvMkIu3EAmm+3dF6OPB2rVDfkrQIqrduNpN8RShbTgArcauSF+nvQDkC0k6vOz
hLg/JrxV2BguinFuahP7+a5ZDaHwCi2N820kVp/0Tcz6djaGYmNtEIU/SZkKkhmFh7I94QUv06/k
L3IB9Z3hL8RFKN6q68xQANFraXnr6IiIZMSxnC6Xm4qRAggxGRJjtpnx7/VXR5Y42asjS8lc5btE
VWA3t001zE3AOQ9SmP92X35VHAf2yGNmN3WkBw3y/L1XaqceE5Dqn2HgGFffh/A4av4yMN/OFx88
a5dQrTedbWQSsoMkZwx09Pwwd6mnURRJipd7dW3rnSKzhKgmTaOSYjx6+M5T/ieKyVWDFLlTswHL
ag11WnNT08d7Aat0ciyFcvxDmNpPVASTrXSw5fkq6KSP5lwJnj8+Kn36RztBY3BrGs8IWjMdV11x
AwNwZQVXTHz9frW73cJDrYCLfOui0+LSkw8RvtXggqRV4g0XIrb2N1BYFos8zHnDlZpDNvKuXUrH
BcJUHQdDKaOA2StmtFARK74AzBCQ1367guuHKgvICge2FMg3ovb1xAhEM2WWoCCqooRe/UQvNwdr
2gS2zeY/6iB/CK/gpLVOpN9w03AfBzZMvlugWCQV3OE4z6u/t5gklSmqZICgEAmwfRxLYiYTaH5T
4HlZclfJ9cNRVYx0jT2SZZMom34ITgIXoYMeQU48aWjXpQCWEGPCmOWE+V/GEoCoI3CytlN2hoxr
bnc/BDE9lK46VNm/eD2PSsfYtsgqe99shPYYJqJDHbFXVD6tGpuRL764s9F25GjgMWd7c9YIJwls
II+th7DWfFkXU5W8Jv5vbtffzmJFBZNt70AN7X/cbTDcI1R6BXfuxQtZboGRET3vI9aBj9FlsgcX
JcC/wdamMIDwfSd8v+8DC+5BaRTgPA/kF3NXxr1sAXFauz2XpeDqdDK/LlhjgWoGrdIB2i3N9cZW
27S/XVfZAWCXMBlohxB8ukEn4PgDSpcSezM4I/Ye8pIL9Y8MuRbpQBkO/TEuzJTVFs++4UXIMg8C
B8RsOVxhyXX1IRjKm8Ms3VNIdvM5zHz+ABAisVIjRIL0v16ItnXkFwE7DTjanBc8aiOGLgXAUxl9
TG+bigUQTBjEVxljz7L3V46WssTR7vv71iSOm5vqfBvSbVYu1eUWh8vt5nh2cXluc6bggr+qE3j6
6vixFjGlcNbfLZUjFneGzqIGGhlaU9Pj90v+81NXrEvrvol8X8/tQ9h1fkYXsH+fBKIHrERCz8fC
EX6iNTknVROwSsZhjBI9iMRx9jL7DKIxuOQa/9/c8HeqKJx+Dv+VpwBDhkGc8DwvHmscf/RNhghZ
MNEz1k07NgFasF0GH6vckeAI5OHF89xtxdKORtGMpj40zZ1d+5/EE9vD2Rpf0sCIEgD90uEj94o4
z3sktmjHJ5MM3Il0uAgDZkxCduVPnpZSEZxkhR4cFDewVciLUnBmbXzm9gdJjyTLCzQMOWv0ncSw
0faxaP2n0WHrVsxDy+A5Q76fyliLR4gQM7XbCuSTD8Tki5uRAtyJMCtQrOtalX6KgRRvK7wlfL/m
sAFD699n5o30jf01MLJ03c+S6kWpz8EYiN693vFJ70jzvdlG1B31859fNOhpZz4X1M0CVwxh5tff
X5bK26Dk93XZ4IDh/2d7uCucSqAMUosy0cepIe5xwKzhPw5F+hqQ37famPEjTyr6uTXv9cd2jglw
wt0tKaqScZxdPCyBVyYPJneCdcTd7UmcahMVXv9xXV63Vtn41yDCmPhzw4gsPtlk0gofHocv6V9A
qkFvobTvPpx/f/zpaW00PZte+rA7kiWPw7OwebD2oTNYqsSVCmMbgllYlfYrVky79X2I6mAc0R2T
JSQ4LTM5Id49dBcHfgLXLxjy7YSbvIlBJ9GtuGGuDJ3YBF2o7UARCIjdrDyLeRY6FDN0mf1bWPWl
z07aeHpuIxHRBbxBoFpZ3ng1pH6VGPa+ieNFt8IL47KWg4AQX1TofU93V3IZio5WQ5r8BjsxUroY
pSHvoS0qhHHDHSSQl5AWGSLhYyxiS4MImhS2J307XOHUH7lX3eunCZMja2+XRDy/uEXSsOUCWL7v
Ci0w+9qjny3T/F39Qm/wAsaDfOvQBUAWkPGCsXjWEIkQ48sZbi1tvHeIBqZ2fori6x8q9uk0VF0R
Dicl5orgYfbSlPf9KxbWDKNCjrcmdCH3QsMhsmXaRuoeFtrMpO0sN4hFszv4LBOHPYDi3jync20F
Kf6R8zjKQH6h8iiH6+WCRHT4Ehwz5QF0vuspXT3sV5Yiv1TgQKLy2iiWLp3urDlkj3xutCEaRiQV
/pTYl7xSGnoKxYeQg6GDy9tMxq+hSfkyTA7baNq1q5IcGw14f4u72eh8REaCIM69clovxSJeRJNc
308zvxlCLMc7aStB9Q4FnsQGsS9d0hM90dXM7Lv0O+WgvPlJRSI2t0rZF+ndVsUv5BYd9dWOGcVa
GdtoovsvuF53bRsFpndUXXquynOjiqVUG8qITpOYxcH4T3sK/jP90zcOL3nd9Z/0jY6LDUABpwv8
mADDvOB42FDqHZN6DKIfANewP5e2ZKlYtsbicbqHrEDSH06gUCRiF5+Q35fzrqq2DEks+DN8Nib4
ptrSDoey6gQoyisHifrxif3lcDKOFChrowH5tXWK7jPMy9hZ/A+mJHF4DHtDPl1WJMhICTDJl0Og
dd8qdkBh/D6d4ubp+cT9c7OZuNd/jAcWWoDHSShM6nnvY7vVb3ADWtrq8SuVFM9XzVqB9LBbXCrk
1mCXAsywPVKXHL7v4xLz49gqT3tYLdHWZKo4Acj9rcl5IRxulBtmtW7/Kg07DvqBuxFaKfBvXu7z
q6BPcZaf3zx1CRSTMZiP1bQ4derSJ3SiIKzobS4OPkNFo5AerrVhatRQ9n/yO+naVuQuw+s9Ku+f
7s9WzQwW9fA74upYFcLruKau/1GLCp1/Qy5dZJYUVQvN7OJO9VWlIddoAKLxjxeBINo8LLc9GlJk
koWT2S3nBl+9v3eOkXHuK53WKtboYrjuyQ3d/Ah0Pw+39Y+MOG5P+/kaP2ACwGbJ/+IB3AV5aAvE
98wa8POaCa2dmOiuQp+L3miXadIOVrcjakk82o7DrMz+wi++v3r+D0OTBT4G6CqrJGQKYFcZSG4D
4yPVuhrEd2RRu1aofUeZq9eeJ8Sn4PVZKftjOCPqoCp8r4lbxemuvOvL8dokg2jrkwQcYX8sutCi
ez3cSJvyLkAo3MCC1tVuWgcnOsvVc/02yWSPbN8U6DBHb+cMEwuzgzjqcnSJA8jkiUrsLxvStC62
NdwFXVrFKfcOhay0umpvvzmYrvjAVkYEqSMVxoCS+wLN9ix32hLTUqlekmH5uiq3OBS3OSmwcDyM
LgAq9iXkdGc0eB+MXLVZ8KlfGD0tPx0VyWTk8lWIGj6U/TreY3JVWo1K+DUU9qQ5It8DKS+5Kl9L
4+/xamSt2t+29WRIK+ywvGVCOHKDVMy8tNyR2hZk+9oQSMBNfqggZHrOyoQDkTWjdbuajE/ogjOg
DTmoT6Gir/Eym0HSOD7XiRyG0E6EHl8HJ4hYsvoCSss6PFbd/Z1hQBd1tIjKxL5xaj86q6Ku6ZjF
cMVPH3cNNg5Eig9FAqnFC1ZkvXmM/sxjatrFIlXjCmyQMnpjUn2ARx4qF81vQfPArmp6/w4vKOnv
Mmf0cFaQil2159a7bY7w5wg3sr/UmdVTd7BwoH3/ItJFN28yRjbnU8HDwcw7fpXvbVumrSmAnf3R
GsJb4YPA/rE0OlJDBXtQPjxljhdgxwkFNkwB48ftXFOSQnCfoBEJifF/5zEOpGWqqlrAMW9DyNJR
I0HP6JgchGqvvltbbci//cPO3TZX6lDRxFAmAqTdsnFDhgjsrWWdDEcZt8J8xMc8tVkrRlesUD70
jxHI26Dja0w1U02Ou4CFK3trju4kkPWIhXqhBe5F9D59jxlC0traB+5bodsQau1weWotOKW4/3pK
huVJpr/h9ajmUHvNllpcBIM+LUBT7Sm9c+GSvMrUP5anYJStHAtLtP0PDF3IjtH0pV5SRipCRmyj
ewb2v7vsnBlPmyKRQnrt31Vf9F9c5VHLQc6K0mKHSJF8rtok/zAy6oOz+46CSoMazp6EpP95q7vC
5Qkg3d+H7unseCaYG5V3EBlBp/TIWoHzoSRlj2thLjove5VbLguGRWhUjccwq4strHhj6t22LLNT
OWV0P8hoOY6KrtJ19vJxIdGRYmZGYnzzSEytL1qfpIh3jR12hNQTDzgm2Vs5PFbK1M2KDsJb5bzX
zoLMVSGQv2T10IP0AM0FIjYvZaU9RjHgXK1o17mA+n6NSrNOOEFsvQvu7/MQ9+lHQLnDF5xS7MkP
LubtrCF7HsISFxpfXrRCMalbirlZhyE7WfCDsnyB9CiTxvCkt+f5WdocE9T8pKkkeKoTZfDLo9YW
mBADZWZU/EPUaxZdUN6ldy0mnN2lTMu8SiW2VBXOA2HJzG1umdBGjAVAp5SsLGstlu/dLrthAtqL
zpcuqpKfuDsoCRyC04BNWXoeG3n3cgau48gLGIdYoPE3BVCEbHoNTOtXpaGtSnbUH8qWs00fBWZq
jvCJh8HUB3CqNjunQHe9QcrK68/FK0saKj5lPXTw1WTeonwQzJ/Uqz6BR5oXR5fkaA0Cs9J2mslM
hiPHSaShWr1cgfz7/0JPFGXuTvNpldFRJHmVb60Qn0qO1Gdn01Z22HpmmOcpDRd+MveIBjnoqruq
h4sUQrRTBndyB6bkIfCyAKZk4PIdGV+VcoEoAtntdYPFRiPMAMglue/N+SpqZCcgVkqRkzuaB8c3
TqbX4Ri7jfShuiDlcS8/GgC9L3McPKZDnADC/OKKomit5iOXCQImmSptNEiMmPqlP/rqflZOI606
h0homoVe4FRlf5G+SxVGz68As7Mbog97YbO/pgL9mRxM0KE3D5+cKCO+LHLdd1qEwBMOoaQ5eziW
2XlPGhfXNXWJqsd+LeUmsr14OEDDeCgPtB1uixP0PbZj9wHSYeBSCiTQ3HFw5+OzDIUdRk7YZskg
PMymIOMpwBYxrlNKXMdJ7FuRNimsC/oIHaR60DaCNfugifG5M/nKzdvW31bU0xaX1HZ32a76WamE
hH+khYtryaOJEwkTo+W9DueN/uthCSVgV0u1iu6y+UBDjtktQsP6BLSoylozuv51UJGNlWyI/ZYQ
FZjC9XxkI3od/ei31ngRhUVP3T5YUx2I2AR3EfYqSGlsQteCFKKuqZpHbU5rWkYwzNgTofnLP1uV
35iOCo+h9UgajxtB+YjxYR+gglzz0rZTN6N4drFsTa+RLpHFPFuSv23w2C3dGRd19I/UKuaGbcQD
20AhPaP1U/RwtfV7/5H8+JoztiD7PK/TQFCWgMl5VrXKQrX+RYfZ4cR12KWC3mbZd/1/OOGiO7we
hMHtWU7zg8O4+DgUkNk4ba87TDb/BDxEQGHMHd+zR7gL3yo9ljy4mdWrZuD1BTN1MlLjDxbMNei3
/XXsdcEL0NODlWFU+AiEk//45zgUQO9CYeQe6ie9wyTamYz6AjCUjAfMWzcJK4jvVQ2vrWuvG1NN
r8daU38pQF47nmaBGW+E/f2E4uKxbmkaTC5VKdMfOEBjbTUTthJTk5hZyzZJumBkwwUWMo3bG4hH
1JuCO1E/6EXlsilO25eH7Gy3HgR03pWJfAcOI9tJieQTSETzhILAZdjlt+84Xv/UD4+Sepbi3m+F
9Gbgv9WFpSBYsF+3qohpyCohc4EjC92HD2Nm5HnygF0r1GWTdZDNXj/wETK5PKGR8DBTMijcDdgF
PXsttGaUQ/wx5+bo9E233c5Na3GPZMMdYRqJz9Rlz61Omw4tcEE+DlEQwWKw6G6wbDPKbv6T5cyS
bHRyq1bry/nRarcwMw/PzYjgHUQV9cT3wGqjrZcUVP8DY+cGhR5RXJoqmlzz2KG1n9uQvPDecaXE
MxiZ/vACqrC7bvHxhaj2KD8HVwF08RDjil8HdY3m6dcMTTynBJrz7Mr1d0CGxi5M5MeINf+szsP3
EeS90V1Q/kF+PMq8vNBuXBr4CBkJ0IK4QQ418KvL0iEIeoI9lVeYRg/kt9QeuuAbojJav/anIZNl
xqmkToNEjkRos622dJpg7L5qxtdOmAiVQrKhEGHYOpFWlyVsQsJiOKMIlU5BVwH4tWyVkzeBklIw
qqbfs+y9oqpaCAnX+cJunv7HnmaCp0txAqNuAjSPvECbODpsnjYV2ttVEaTvNbmistVkLQ83JdnL
rqa7zsb6UYhFzYq55QS1SDsVQvWNwuJH9NUe0JuHXLw1w56zUgQWeTvbmZX2hPFwPwYqAtR0StYT
jhqiDroDscN+EHWk5q2eidmV2T6SlACHTZj2VPeHugwnF3g0i2uz2AvAYbNWGAU845C8TMn055aA
WKmBBPUjPwJ2A74JFBuJS3olPBD1WVgZ7dMD41ZI4fTQw8sRCQ06V89ei3bcfsufOEQRIhSIq8qC
/51doVneXMuBybwyfwe/+AZeX9eWWpvGlkq4N75nWgRLcKco0pTTScXcvmJ8B6wxZ1+UstAce2SD
V04Hf7ztcwhVnR2L+kmQmfTBPyXY33VgdKUYtKf4bClQZulP+BZgYPZBSyUfVAQNw0Xeb2OxGhb1
atNd/NqeN97j7ueivr+QcK2lvIMqWbQBsGaZIlIAQAt2kB/lMkW1cRSVXPfOLSly10SbtL5DQaFe
Cvhvk5ZPKRT7gIi87mLpHaw2nT8iFoMzVAEmaobT648JPTbVdbcTTFxxW/OiNPZt1BM5ARYrlRDv
4pcWtG6oHrAPprgTYE3NWjHY6KuS14XCwEKiR+CAH9nzNtrbpPEwRnVfjTTVSi2CpUO1GVqleVGe
Lj/doRohV60qdXVyl8p8WI9yeokQbGODyz3QoThvALpr/JZted1ryHSbT0eg+m11NrXfkshmhf/c
kDomb9uaapUAv/G7K7nULuCGbAta4F9Mte5+dg9A51lawy+rfBBNTngGv/zKr+myaygK7UqnIoqz
C/nYUY/ljYijIadKW0e3DHQvYfQTVdQUKeeyw51b043WGrCruT1QekQAYOoV2Y8nqX6WUb/TidHe
xE9zOM1FLrd0J10yZNehons81tjU99BUKpF4G4gpGQLCwwqIL8srHk9Mkj/KLOL2HkocG+DR2LCh
wqNEa4qLEmkmfvbdn7TKiZkRGJxWlLoY+DexVZ6Qa7AUsG/oyhkzLNU6/peOe6/kip8amTltFy/w
e2YHcqVcByRdCbNG08XqXxgCtAKIIU6+RVtmolh3Jyra3wwdY0dnj6ydm/GQD0hjwArkwmkYWjy8
416E35AqQknp0pAm8e24PjOdf2vJ1msbidxFzxcMI3/69/z9g1uLmZurTe35dL0DahV+Cji94gtY
y44TFnXAeeMiejBNaZ+hDEKmaUKxIVKuMH2UffkWJMTh3CmcQZyF6E+ZsfuFNxatgR45Jsp6jwu1
PdAOAgKVNFa6/wOElSWdW4lxN4gZn96NsYgJcUAPknJP8zLb+UEEuhP0S3fuXyQjFGyOo2htm0c7
LecqdbVvsbQNFrlxX1JDTrW76g0T418Q+c9AnawuLzSP1wvqHupFTDL1/PZlAYICEph48k5+FtZa
GbqtiBX5Kryl+iG/TIigJ/q7vRsiZG1hFhwF1d4kMHO8W+/UOtTgL6O0kFX87HCGlXshVtwzOL1s
4EumXkebF3pN7RNY47y1VbLaImzRQA46kjLXt2KlgJrhmUr5LdVrlAVv7HHwYKHqni0LJQVmkWsy
W3Twn3RU8N5JUIWlWcdmEXoqdk9eHrvyVYgKq1qiPAEEec4UCFVgFkChtlZ1M8zzOYkDUWXa1YcG
dZ9gUAu4l+Qt/3MathtpEdJb9umHacpESVnjiYS5pB53dQcNODFe28y77p8Nnjz98HROFutMdqng
N1qXE0aZcSChkQ7cwwAalODwqEJraeLNuKA/JUScK/ISNRW+cd0MGwA/AECiOvElPn3mPdqT1US+
/wB3XD44qDsqe+zyMwJDHUE3zpinb8abUJZyxUEJ+s6hq5qBOiT4vE11PL/6ZbskdLrt6NpkL8Wk
Q7ASnCZeI83gIJAafzg7pj3pNGuSaqRJExW1F5O0BYoax1ifSMf9X7Et4z6A9bA+jeUJA7qX0U0o
e7K7iasxVP5aRVdklXLVVYad3Wn3D0MGMdQ2gjAPGNv7y1ValalvtpmXkVDOss854UYbvhgnMKBk
OqVHr4BIYIbd88K92pMqN8nvhDHdSF8yDbVOGBoCMhD85Zt4e7RXaK3QFjK07lt+bmcQ+W9NuMcU
YcPA2Ctl9gQYeh8Kz/vN1HmOTwsmV5NUhH2bMdEJgOkRUqxcxSbHP/cR5fOL6GH9MmgSSPvLlLFt
q72Us9MbZSHOI0fslMiHf8lfVnYaI45V26O1t/ST7afPXyd5kWt6RfITsVZ8VVMSrnXeHxG0z8Vw
/Sy1+PZqlit18rOqPIT7DLkRrLZFwAlVlKpR1qq//4Xi+bwY3J+snq0Gc2vFwxEeIXfGvtqXSj1M
RyJsdkwCobC8d515J/wK1l0mV1DbW6TrdzFo1ZD4yibgMJH1gS+ygkrX3Ees9x6ZWK+5NERrmseA
MYuzG1WtL85lK3v9a0YM//my1bAkTKfIER/rtJVlkg8HKRrzJOX7caJFRCC5y34vV+vjf1lFmctW
4ALv+oBEaxwzTglyjziH50aRItP7Pnp8X6U+d9Q75YQ/iQDXfq/YEizIuOZlsxeAsnXC0o7zPpGr
poq2da8wQr2YISPwMsGhceILYAWxFOcOhD0xn9YB89dV5dKk8v53HZmlMvgSMn4R8k8bOB5YO4lB
0Z78LINEbmszr0BojrXjjUWP9xCyt8YUbETQZH///PTO7tswvbgNA1eCoFKJTIbDSFbgCSrqoTAx
vJ7QgB1sk6XN3RJEq2ievpom5B76UsM3o/8MMx0SRXA41daBaGXlMB2XnFsGRNDTx+rYffXIk8ON
SYAVzFwJphebHl1qYQrTpKgOuUD3qcsuWo3MDCDAkOYrx3U2dkJkg23JGP8VsCmIcJ0uAHTh8cIQ
zAcs7pvXweddOCdT/N6D6VmUhHp0YKRHw9Hc1h3ftKLPxpsrtOiYa2uESYTc5j1SUCNyl6Mk/ksa
NiVqFfQZb1ANKIFLZScuIq88GBYHJLQZ5pYwXozBjvI0ni6GlO1QKkNFpUz2/ziRcZa8PZX9owQr
fZLr+lRA9jt3+Tf87YUKaDoAesMTQsKT9xIM2cIkry1pqNYtoIMBsc990OyxaNl2kAAY0fZQJ3NA
3evmjsitG4zXDWP1It/KrjwuLMIQahae+DxhTv3LVB5ShDg9J43j237Sxt58IuRQtmtQ/7yf1AdH
ATC0wia3HgOjIh83ZZMKmuved5OKzHnh8DTED8b143pcvPc1EqrIUTTeVlZvxpaFtcgrY1+etesv
c5/mV6HqdRBbvifA3PW9wRUjUmXguU2jxfchC/ZBQIoOLqHoz4oUlnTLHYMvvmxz7vES8x6tVu5G
GNXZfKkShfVUizKQ1vnBDDjpuYyZLuWZ59guyOK1SuL4takSkDntLNOuYwk2o0ln/yx9If4iT+oh
n/SxrrYKSwP+kJlQUIFoBXacSqXOYigwHFbKvZolK8S1xPcuvgGbYPJF4nMOCof63ah7e9X2xvQM
sN0reETATKQw6bF5gAqyX3LE/vyu2xlHvobw/xQYpT6jMK0d1S2jJpvPLp+OTWtKCnI3rSwOi2/Q
KzjxSpSFipcU33KSfAjDttrVxd/EkiR6e5PXA/xitySeKn/MXOhHApNna+EzkYg49+OGmiqKO67y
oscZLJqq2Rf7OVIPgKdY5bdEl5UZ4AWL7dBrg3sG3DmUi0QQYZ/dUwerhUhpXmhX/Rpg3mNfP4A0
ks4+AShI5P13A1K2w/l7MA/1VkqnwU0c7U5WNsX74Bv1i51Pb0G/ZORlUN+bZCoh/B4skBPT+vrH
n4IJoLd6GU67qJMNX4iedmj+EAjTjKOl4pK0T1RO4D21SNYUn5C+g/Ks0wLtRs0ixDJq9JB67SxK
blvQGz85jKr+t1F2fxCTJObh5xt7O6UiaeSQXyImJcieUN9mpMp4hBbBNqWXMM/poxcxRjbrF9mx
zFZU+ZMrIIJ3uO0HBJunaoHgn4D6+0Uav/Pe/Y5/rh9NcmUBFMFXbJ6wmelB7uqVis1Z34SpDTaN
lyXu08sc6icbptmZ2gXvcuhW/45DFRqIHvLFuUczNGci9MTBYeqXfH7XilWLoQxJzF27weANqReZ
A1ZsR1743KXDk1mA2wPTIolmROxZ/ZAHn1bt7hgFyDjQNOVgzKFQCvSqL3wxy0Mg/BT8LkeSaVmX
6CUx9WiEkbfuXu2j/7nevwDOImUfyFXsBsM/l5FP0FIk2EW5JYP8C+X6aA7pipFBom22LetX9ncs
xdWTS1+nE6Nz+Eeo++6JGiotXnyln5XCyyuXO/5yDjlDlm0M+HHJOHLLSx7DZVOrRW9TDWq5ckYu
Biqv8pOuZ0yf/5+ZxfieeF3DiabGr93NlbtsF6cMGyZoat52rY4jUPObOvCobmaf0U98QYv4B8wk
kD7g3oVERhCoAuyb6S2FEMQVr3EvPMwF5jDYoAa+PFmi8JVeJhA7aECanhb6FCWwadXDkn7v1dGf
j/jB1S0WQ+XOAbEbUJEixe4BD6MpDjeAWa5xaWZUm5yNY+Xhy8Dh0yVIjd0Yt44SrSJxDI4+NqbB
IFWhpnrK4mwecIB4irEpVOELWf3bNy7Jiuz0hXWem3NLKfZ+57lrL1D4KmUltnOAtVAJegxue5io
0jDEfhWE1wuqSz8hCffd7+ZLHst+dRnz7/x+9y2j22VQ+UAbzwQflFaGtk93+G7KmByVzepC19lr
CYdgN00RHquUe6lM1zmcjhLyhYanBcvG+tBS2hCTH6j2OOXgZk9qJmGpQwNaPFAjfS0k6o2SziEy
8BD35RP/YD+61hkVSRVW5aXchco7S1GBrmvBCwI250N4HEjvVXVGYHTKOMUsazFALDkLmfzRB+wD
6gXQ4bBfgccwZBDIO7sRoY17lmW+uqUNE3/Gl+svEcDIKFvQXK11DE23qDiuzp60L5LXNxgF21QV
Wa2LaAT5uMweTgMEmKQTILakYsMnSogwFZii66LqS7v2TBwsUEIKytWeU9RIcX1TuurfxT8iSTtK
2hOz8ccacIspt4xkd1z1zLf/E6ttXKMTYtml0XWgvlcgrW9rki7SycE/Dx2U0qcp5o0DgZS5RB7U
JQ8WibA6YAfwSF495WvQ3vCpbs47MezMda33phYjNcudhRcuZXdeUNNt6tzaHg+r52eO5RuAdA0v
/nvILxZFRe3Y6uI2gHZYYjJlj1laYCCkvJdZyHjBLCka6JWafgKJEmYxizZJOR0RLY6PpLjN3oum
iiOkmncLTswG8iPwlEMBqbSsYK3rZWOUooMKxFdOIB0XIqBD/nSKhZTB+f3kQgb2KxeRVUArVKBv
VtktWymOEawuAg7IdbmU7YN3CYYYcS4Hbr8HTsL/1IS15AT3UNR4MEQvv5X5VIBGGmiDNBiiwARK
srtcWfSIOjlwx3Fc1grBUw1v4asgshMUMhE4l5az2OAX33Znp7UTNxOh+texEh4dr51vOhls9lNy
7gCShZbMo5os8RX6STOvl52M0HO9pyLekGFSdqaFNUx3G2tj7kII1J9mFQkxBZDqbJQ07lgpmhMV
/RVGnNFNDuxhzji8Tm7MZpBkkss272o9i01RVcdQrZMupPJdBP0Vbr4TQfETa+Ct9OW/GMHtLbjM
+1H+clQmBCxO/qN+btKow9UQOWitG4gfNbe8JjuMYIR8W1LyM6ZQR7zX4MfYjJWTme2plYoS5C7R
Ws5+DMTRkJ8qnCM8aN1gOVccDLmy4O6Jon621fAZMM/IbNkX8gDR2lJbiyUWUQcvqgdWPHlGyMVV
DSzdL1JC+lxA+dkyeCrn2w2QCGHWhkJ+9rnk/2fb8l6KyoFVlL4XPB8POoibT7TR7iWurlh3UN9e
9TBiHMUL3PIcjU8WGqWwzzRd29ViFyFUgf1d2uko+Qmgzd28WFHtYyenmthznTE84PC1BaMxcL3V
nhXhpBb2oCEw0HcT2dC9b6onMU/Mjun8jH2sGZK7YZb2iVDjHU901c4QwLskDbAgea93WfdYisYk
F4w9bNvxdGBZ2Jd2MlqV5yJKYo8CeWxeipwW+J4jQFuvRM/1cOc8ZTTyF9tPRgVO/9JRKkgTSD79
JLa1Z5XAYxH2QJVJnZXhy5ZmsapWm9jdug7K822DaozVq8heJucpgo4xNBDdkTynYsawDKWq1pkD
6r21AUOv1ABjVReCCi2Sw9hPMccBQjHSHRDJn28PMjK+h+VLA+Y5jgL4djfmzoAC4ML+I+YLwhyx
OcYzc1clopmVgvSc//tZof/Vm0rupxMMIqffP5DXxTPve3L0B4OE4hUuqJdHrIObWDTIc1TLsM8/
4dZ96o5x3bGb71s9TJBbuQYHdGR87Ezhj2fSNB4lcgddXgB7MbkOfO06Nq8PBfGeHNfhY4KH1JSz
U9r+OtPy/zSLQZHYm4VmQlHuj+R7OyPD3Vsfi95vhOyiXa6fMeP31DSmjdPgBybIISf/mcZRdItx
nq9GUBkLZF8GCI0K6ufYUtDkBmmZTmaOGDa1IILXrKNlnC4HLmODY++/MocDmD/b62QPEIqIp03S
eZyiJ7OG00eTpTvHZS+jPXczoN8hogLhr7soGGBeoHNgKuuK3/jtOr7RJ01QQwMwS2Ohb/xfEQsK
xdxwknB7MCdoN4EC9O2Ht66hLBkTeBf4yTjlUg4TOrWIJHAY5N2Nj1MIan/93opj43U/3y9SbJXR
gLkEV86ActCf/Ql9JGioSCNzbg9NeeJYo3M8MCmF5O+ibZd/LY8rBDVhYkkUNjI/twPp/a5F8H2R
A1DwnRgKE5YH6ptlmi9KoOJZM4gkk64l9bYyzJiDiD6Upkx43LRpO/k+hKlj8JkCrMVUUBUKQrZN
gLFDcO5iH7zKnf1cJCldw3R7uERi88NtDzNDuMmPMldV+N09B7cljIf/a+nIweF6F9555WIvSfBH
f+LiV/bz/Osz32vIh+4HoXDHjend64h0jNNh6ej80T8RegcMSUqRySEZxqQxPH5+d+wW56cEe2Gk
/On8z0+aTrcpVRsnPwtQ7Of++pGaU7qMPNrMuVsXSl3TQgQ0tRw4WIz0AC7d9pFmfYdJECIaF3EB
snimsglWT6KafnAk/n7Z515nj+USjmiHbc6IldM5IkcHUWSyXsH4ttANzqtyytEAfheU6SWg9+HR
3HUWh0oY+3G3s59xkp2r57exICHr/HF6LaQLCrdfYpcMPy4rSY2yb40igKSmZ0nOQQbv6DmqmXyY
vp52pV/uO/o3IIVa2ybnTgkgljWCsG5xVNOcX4R3whfXyxW8/4DaFJWkbKHiwGDz33VaHLO5Vbiz
DpzTbmRrN58SFxBZihoLrcWSBCqjsNnzL57tWEP5J5llY7IJVI7es6Ndl3U/HiYMBrRysfWZRQhT
YsYLjwLCosBedbfs4M4LU88+G+z+eR5t9TwXorzfqetWY03yJ70Cgw666uIX0LfWeqtYrNCAyw4w
jbOlXlnEgXdLnzqXjo68Jrre1vys3Lyep5Du/OUuMw5HC3kJfBDitQZBav+1ftjLLX8c+Gy4dMKC
FFhrLIW6AJVAbiFr2MoRwH62fDRTkXzTb5dtjY1f62Ubrd24ElKWYUcwzUNibJz6DbVCE9l4eRwW
rYIQxJerqI/ZRcqhOkp/gj3hR8FXKoVHhYKYlFPeZ6iCKt3huCTVLV6DEg+gajP5fHXvcCLdx3DV
Y61sSkRzk4Z7qypcNOWVsRC+pIT1K7T6nZoeP3yQsTDSEbdgMCKLjh+l3tPmSwcehdjppOH1tGA2
EMxSpOz1A0pIdB54LRTH2udVHyp/z915BY7rcCtRZtcXPXi+mdYPUHDrVZTaNiwowwQNwBlMX/My
/KPXkxzVr4conZhqRH5fU2W1RMwDRn9dK+y0ciCfv9VvlWxjBThqdH1p7qV9lKYxp7LDd39Gup0T
O/ItVSsKnN6eMcGEMZ1q1jwBInrywSKQiCGwcrNxlEzEjvpsgK3sWbVGU53S0VeBcZpX5wPZYrOq
uXYR31Kh5D1sUBv1Y8tfSsU9eQZ0c5v9udg4S7APprVVvAmpf3ebUJ7KJQ7JKHe1HFPP0kvgrORb
79riTMKaSqzFnor6XzC42PbxFnp91oPsc7nkar5fKNmGkQ23QWuREN8OGItAmpMyRQJRnfzI7enr
+kUULa4YzrJxLFqRLyI521jn5M6eukAuvYqij7dfBeUs+a1kN/1hdJGFGl/PdPZ5mVk6Jv9TaugL
rCh5EKuRRyO8Ruxxl2fw+RIAcVsN48eP4SrL1HWYVbDAgbO2whwsyGH0QQIdH+4fCXrWFI2XAwOt
91tauvopJbF5CBHYav4F3CsxsQdmC+Ny2yqsMuDGZiT1yJq83OYqXwhqWx0kiJzBXGIXaaCWvdHE
DsQSNXzCHNt2IJWBc4RmEQG4zcM1/PVrzmzIMDSCOQQ/kgu+f7HKZ2FB4QXoHMEfCu8yB7kNDKHI
hCUvXmypWsKB6+HFvZjIxLd7GWmgOBLnMalVjnkojHkkkDbORLCfY3O63jx7m3+jY9h44jmS5H9B
KQF8ba3+ScImyFdrSS0/N5edglUrVe50i7Ax7wVH8H4eMcx56jucqmpsYmmDt2pFAIsBHnU6uDx9
MSfNNSj5iNMDcMWPxmpW3n04kG6W4uE7Vi4zr2yVj5BS0U0pJvuuUcIc07Z/q3t38Sv6FVy4Yavh
3JsIxP8rYdVfJWrrCE1DUKsWTubXgMjwxhjB/YQOci7xecK1dMK+uBMhtk1I9GgLdU/xtJQUSrFW
eeUn0VVA4UIo9spzkyg1crGvtVVcb5GNEMoLqBscRVznItkrC8XyyPt+T2KXniBdtXK9Zgzo6bWo
hD9D1hofaV6YDYzZwfS0+J6If9wzWplIJp8caw2n/Qi7qkV/bi2AKDx9tTYe53TN9TtkldX9vfSD
XcKm3omhMfSkMsgPekooIvPAfDzrktA4rJ9FBye21x5/7XLXIQAuMnWUU2XzvHPcW8nD+tYrQt4h
19WXL8YzbBOXJqRMzkAZNHhY68l1CjIwm5tZsthJKnxFfP7EXiNWZlsA00OZXtr3m8TAyuLw2J/4
ESXYc4hl3YutNMExhf3Ok75FQPJU9m3BTT1nq6Z74AMLCa+MahPO8D0zr1mLN+GlApxyrBwb6bOD
1ZW6lyVZEIYtk+V76Ds9onuYjn4avUtZabfmLDloQw7cukUmFeMD4qBd7S1aG9DFtd0LrzC7KZ8l
QEibOXQ4HiLAC3sT/hjxMdt5PXZMQ0Sp0fiFDUorXVLxaBcjCFu7WKbVp1Jv0sN9pEEL4yvRIGrj
GPW4PHADg3wTncoT/q682aBevJgxTI5/eUgA1R2qgJXQ2LvxPLSEGw+3KPPo4iwT9heMq2fwIuHp
vXPfkwTqqyASNhEQEHOxxGDUon6m6s1yFSSg79bR0kUqk0T2ed0BN4VHSYyf0a99Cpiz5swIlegf
slcNObUOPVq3CQzPYFxzRMAzQd4qvp7Sq1yKI5mZba1f+Kp9hGPnSmSl7bz8W33ymDvC+zQQgHBJ
9I7czMj2xI/8ajLuIXdwPMwrC3NqFqfQ3J0NV/xIR8MvLWEE5hZ0oYstGN+3jIvSIWkJdM+0sgi2
tCI0ba23/Zs3fpkJA3ENU7OuSfQ+zDOr1y2NztQkzafwDtpmtuG7rq4Vomd0x5Ck5i5QvPJRZqCW
tlIc3KXgHnopTtYArySbtTxjg7Gi14JyefaCiZxiy1nu97JmsuqQZGWvhan86j7CAjuWmw5hfyzt
OFdiQd5+idmQ5FA2ZsMCkW4gFPTL8tCUG99xAkR0Rydkph/h+H/w4Z/JuhReIsGeb+BNB6LlwIaH
GZBTdoi4705o0/83Kf9QwQ7iQ7UUCYDmgX8yyiSi9ZVotlui7rBw2nW8XFCPe9HPabRYl5THfRnJ
9R7MLiq+ERw1MZCslN9M2DZDIAjmcsA4vW/EG7jGvLWB+R9iDdSYZv5jpyM8X6t3w9M5mvusaBV6
ggdFKKuhSF7NAzglRy/mrJnIkc8icDDc9w2qztrlpzDZjs583xeKNtliDA05E7LJWwcimSyPxxMM
zHi1ODXZ1rZ4BBCPCeNShvjhd4E2Dkla0F/RXzqZJK4cLIpHG/yktd7vloAfU9p8G7Dq3TbNBn2p
otEdUBhzcpo0E4nqJ+qfLYI06VRtE6IsIoMEverFmRKZG5xyQUG6e15fofd8hvgnGNNbaii+o1HT
RoaKV30xHrhLLW4jSRY5Wxw7hwmiKdgMaubtQLYj51AiZy4ksZMfKEjNdMfgGDbTPO1PCFOjVMj7
cq35r+Zd2QiS6uLTSQV+HXkKWzBndSyVe4JxA2IUvHo4xwEIZyw6E/uTZUEoaLdP07Ch0U/UT1jD
DzWzvRqYlOEJaJ7fCRqtvIV7xy/QIB3a0R/P4IKJUEOi6E5PTbUAUZsFmHF4DXkTvqC6I60lOSzs
rLspxAXkroJ/6nw/ehhK06xrOnG/L4rj3l5OD7HlBQjJgsEoCMTfSgaxMDqU7zAr97Cd9f8pizRN
vlDr9ZnRP7710Xsw18Lwwh1E3u8+CFPOh8NGgbjb2p7f6vu/lpf5LUTzOID3dp1crFg34Ff2yAcq
NFda0L/KASQgvmED/UCT1+VbQS+7iuGxQgkl98yt6R2KdQKiTD1SdYRLL5klWso0kVUYTEXGY10V
jMrqVYSHLi7ymnVU2bfQ+yaez7g3R4kzuZkECdP+6Yp4mWD3rrv4M/8YjhN9KVAoXsv6jXE/Oer0
8Ox7NVeaofeqegiNIycmuQyAIAQ065TVHigLvvHymvWR7vHUz6+uijusCW0tpFrSZkZA2rdc/6BE
HBXU7kqAA9ByidWIes+Z3fr1KchPx9M7qEtc9iiv5NM3KZAmn7vp/PC+oRYJE3yhakOouWWA3ZSR
oVkaO/ORCsJdAqchKb/fV5U42fw11If8FgQJrJCVaWYPR/YUM9saVpT9xme6kb9TafkvincpcgX+
lsusfsPvHlD+Bs46wUkNWBtTlNMna16dp4tDwMC26iiiKM/VYkSJowedU1/pK6HaGKkWyD6UNGIF
8rjLPUalg3v6hevCeikYcrsuHJ8l3wlSEl/LU7AuraZgavqBD5c+hV0HIBQHqdJhAgjSiZcSuaE3
Hqv1SOvGfJbSGY0yY8lA2GMMzeX6sQO+MO+o6wpkNz5qk82TZY4cR1bqlSeXzjq9V0cK1+F9cvOy
IKM7XfRZ3jpf4sza55XJpypUuiJ7eU1ZrnpAj7NNlVlBR3zlRaPSSFDMeojc0XjUklvkI/DJxBMb
nkHEGk9Rt6c21onWM2E55DV0Ln6PPY0o4clnBOnJ5DITQ9a4k03/UrTQoTXtTdH7oCLbI074n2ea
i7juCZzqi85EgEuHq2ZroRde0cy8Hgni3Ms+PblNQU09Ro146UVSIHoYvByVvoBw2R5Vi3vzhY5g
bxZ7CbdASqPjNX2Tpg5/So6yqU3V5FolwRNlFPslKAFWw5ITQy+M9XGvwxAV54g2QndSLBBOok8q
QpYVJzrHDegMHb/nb46aCRbvbggk5X35OTYnZLPdN39/gc1oCDnHn2+Fe+jkS2Yejmd9Jr4pXbby
IEl78DnkxPeAwqpAx2/t2p/R0eG9FBE7Ftk6CUWEM/sFwEs8cHE+rP2BH+3KANQwlcWRS8uwgc6b
S8I/dcqAtjvpNoiGc81F4XVIUpqoyVdS8NIi+n5CSLfJb1xNYspujWBlFWiL73u6cspG0ZOLDfHq
/4r3Kf+oquWL2hafxWinEfVY1wbA8Gmw0+AQ8tjkjCkZ6rwcDZjkRdbrD5UsnBYRfPalbkT1jV2n
UA6/OFXBbFBR9ZLa/y4e1bWK786B1E7JHnXcr+LJMJVYi1X28MBQlCNR8reniFmXxZsmFu/Z8Pml
B4r/yYaxd2Q6dgZgc/Fgkt5FQknl3b7dKdk0yyDKHuxk0bWbLgBFY/HQvvqfJjHP9I4ovgZCCs16
Dkf3zuIKph6KRGWTziD0OxwtbVyOptpD4ErcyK9zdMX8KRhtKwQEESLGfGmKX7pcvalfwIbC95vV
OEc0MXIsb3auQX44qgoYsNQKQm2Xc+Cm0QgSe3+01Q1ju6WjTG9+n38JVWG3qJVLXbJNxDyK2g2c
NyN9JWyHT/RjTdetatmHXpiy9KRwAW8z3LPyHI+VgNmN5H9wVapkQLdfI5xBD1oJGdFZYuiApDVu
mag4CAj3ayZYlJme3tPiAX9Oe4jhScDuE8e8zizdvHc7B7Qj37yVhWUg2WJaymCuBgOodWAjo2ki
GLl5SWJ3bPvZfzWfbGY/4SJZgh9oMdpkyEdlLATVWQKZaklwOk9rVvDop/Qf/+R2W1+gK5uVgx14
Z5D4Yzk+9rW9a2cPezkp2Pcs1LcrnRBCqAwJE3HBYZRvPG4YNy4R3UB77Oo1DClhNmg8+fZXxErp
FkfwZZnL1Mb7jluN58KK+UFgz5xPV1Exfg6MpIvSv1bxzPUxQKDIF4jpRwipLU8NcDAWw1xcLJbr
VJ7imAsUILMdekOKewh9bdqgAJLW2SfadLQv3YRuJRcaZvviAgrqrlYIWZYu+bARNafO377NyIix
OOIHUWhGnZxc6iHeYW0+ES4ehXsUjxA27qG4EESqN1eIpDhXesokaZoTfBvzsGzaGfi3UwB4MAIi
sIPVaMCKnekYvthkVg7OGu4xIaJnyiN4/Z0md1+i+6hyisB+e+F1pwewwL39h9wuKfaeRdzWQUS7
Ecy+BBgDHZV8030jcQVVyNFtwVGJgbBm3zcg7Egk4cAgCAqfFxMu5aHEcH4SYm2B6BT834UWY3tN
Y5Tf5GSmEGA18owEiIt5EM3xyDQJJofTCprYTcnFtYnKEDMU4iZ7RpZHH8YmZUexbQ/MCyUwrGlt
7WAs30a2VzMTv64NwNsC8UFICSyJzoKNbK9zAOw6EPzahAVS7+NU7C3EIzBnA7lJV8KylI17MhOT
ckJpx6v6L2/71zguHAj8JPyDlz/g3m9azcbrdvMp7LvTYBZG1FBOO6KSpY+z+xGossb+aJcWhSEs
FxynFn+K8+Lfwkk4bgR7cpWVyeabnEeu2MSp65heAPdj2yykQ/l+0BudBjGtJ098Dknef6f6TnYX
zUr6lkKK5Cd2JTHmqW/OROMXwA962ckagsTdf75Ftd9s+n4D/jdfK85BU8CpkK4Bl/1l2b2OW0oR
ll5EFrQen328Al0vFDsaVyHO5PcbIRBpSFuMYjuT7d0ohnJgIoYuAMCllgizWC03EUe9ND/R1368
3gNtK8XO0KLwAA2BAcJxnrgHng/10+JFW5rdF/doC+gaXTtNNfIKtDuc6Llft4Gqfe4/IX2s18SS
4EjrDGhYRr9c4DeetZaN/Udj4vRgrWUesxCJrfXYHNnZBzElDy6VR/zXZ0QEZxpEpDqzl+CzIYRX
In2BsQ10vAYGq1j9oxfvwyck+kHhVvkVhw65TTSiJytzm1/2Et6MV2D5LBAuAQ7cKXnzQ6pRc/Cz
uX5hqub3pZiRc+TSNRtKMGGPh4srILZMXNOPaOyhpiZziiNgXZeKd/LI1w6RGl+mUimfecZYJsiF
9O70IHekS2uSv9403OdHFwZ09Q+2Qet6SFM1Muc11+kwgvK0u+5s41k5j7cjvZEuZEZl9cZHf+EZ
a93GPPZIalu4dWy0eszluaQjX/+S125qx8yp5/Spv2CKdHcn5ht4rLPqLJ2J16y7H7L5iVI0ebej
9Jm/TNwA23GVaeEZrW0hJk0dFua+PKFGGIEoLkDPNcE6CO8KzPs8lVIh5N1H0xfV/vd1pqlor+4B
nCapkxNUuc10H0sgnUF+qu9jLM4/7IHGOf2571NT2/8UkQB2IxDKBh5CVXDIgPXOvNHjiChGJVD5
cVvhWpLdncqs6gknDVqHd8VXzIlEHmr5+EM3d0mvzR2IpBNTK2m7Vy/trTPq23nuiMZjuNp+AjR6
bVT0+K4eoOYtxW4z23naS4/liLjM13kJ5/G0Ni3wWZk2xD/FW5uHse0hMoyAReYXfT6RPlO+pA9u
njjLZxEQo8SCtIG8WqhZbszhStblLxszSFmlsgnqrrfigsG1DRB+G+0/B4gY2SoPGUJJnJGMVoKZ
7XfhnwP+OUOQYviAZOc0084in2H+LhbHqPga9uWtjcBwl2C80j0akORAr8VkCNiznvLktS748MCF
O5RUJRLe6Omo2LO2JjSnWxQuc0TqFQSxpXfN5jpCjXfsJPiWx4ZHRmm2Vbastqt0Syc6C2ht8t3R
heOdn/WMC0bPFDChBHbJtM4tvGJzRZiPsorIJQrqLi8XgpbyMFZ45yVoZGKVQ/USx1dR0b5IT5ng
eY0imf8xZP3Q3QTnn5lyYQWkQTQzxLv0zNnaU3ek52mPxz7lVE/N4PDZPaQWK9DGkIJ3bvp/7Ahh
glQzWMzCbKg4vKt4kcyZF856fUI4R9ziavD8omDFj31wAUf5y27K93sr5Lg1wSsJTJRi73CrGoVo
2AS/a5iK8oZqUhL/5Zu8+X1+6QdPCWXKRq95c9YRlv4sELMam+TZzoRZK590tHnoN87D6FnPDjmO
uptpx3Yc1q2woR5qrBhKTtYajgzj09FBTZ0P1NMIM9KnBpk9PiwISUUBXg6k0cZ6RL4mPwt15dCc
wTIVafmxycGDB22j8CmjsoFcLbw0bb+yD+bdcEsJwerQM7xjSVX3Vy3FUFp/R3EXdaHicL4gFwap
0MvqId9q6zCxS9Jpm/cEb0PFdvd0IIwZ+uFYY4WWFfu+2JmKiOh1aCOoe9DeX2SbphWQgWDf/zdw
FOwhF9t29UvB6WTzuvfHBs6VtcGb0LIRLerMjsR9NpGj2V3wSLoW7vLV4t/1AEeiV63EYeSvoKsv
hvUVXTuXZybMpm9AA8bHUbvNK6ud8BQjO5SmOoMRkyHZkpNnY0MueoMma9nICXerytT2prZBLjGe
K8X7H6Kd+3w6UxuUac8637Rl3LhOX3tLgZSouvEIpNpYIIecPCq3bJaPu2rwVREg2LocFq+mGLPW
o0d/RBqrBvPxxb4l9yhEcP0oZ3c1TlC1ffxmSOTFdwEXm+y3MWp6pNx71VnOKOlyIq0Nxilc4dE+
rdKW+EzK/f8wPYa/kQx90rI75eXZfHxvUe7Gfqac4rdgcNJI4qPzhlU337ZMjSXXqVsjB/GiVylu
mBwvwPQ/9mMYTmKUAI78NJk/VA7G+daRj0ABKOdPy0t/LGSs5GxeQe10UtmJnXd0FVtfb3JwO56D
yl01FnpmVlXBEzwgAB4fPAz6neT2sOvyWsKMcDrfCyV6OZxSyoRY/H4mMF+53QIE33xZJQ1eaFqS
gi7+fUIIIeRmn26gV65+9jgko/Po+KItSmg56qYLVFxIqlCSX38RIjtwwaZyF/L8jhxUMteEWB7t
Y5IpIkoDyBbVeDJ2gTFVGN+3ELJI08Gm0FIdCzsabpVjx30QxGv1vAAVjGoD8/XBTYB1JqJ4T/Z9
ZH/SAXXyWrxZW+MO7Pyo6C+wtREOekosCayO+ERHaiDD7nnfFN1g29xnOzXFvWXjZJL9jUwDpN+f
jnMVTA/lFRuBfUSNduuFEiktqJnkK2yBT3Yo1vT7OR7hb5QxiLCp9JP2gCmds2X6hqoDOKatv1ep
Q0hZ0V+2mGYeWUYHPnd3yjwzp3/juf731wNP8BjG67cc3zioZuIkMfMuJmNWYnLFGQrdIIqjqsvh
RGVBCIovU4XDiILU4OtQvRItsx+PtDkAlOIcOsqGyEWnQCtnbqdDOCPjdos6OZwCEBctUiTWyy+l
C/hPI332uSmXmP8jEUfC1YAKlIcW2FpHMjTB3YGCI9iAxzaJlOb7ld5Fxm4OeSgf00EH11t0KmJE
4BupdM716MjMtlX3frlnpWnFrDGjTPiw9Dz6wXqPWe8dze68JRRfKmLH0l/eZnU9uS6WAFCj7fK5
Vg7ElvTQyp97Hit46hugIDD+vPNNia9VYHrCkPSruX0VyjzSXbRKT+ckoEhqJ4+V6fQtHzFb8Pau
oNeqFveKLVeDoY8Ps4aI89DBmk+EsTRKcjpg1VGMZ1BRUPjKyfpcEGuWRhHaKb5L54FYWn2WfAOI
JDQVw9YmkN5c0BI4M7AYvcngn7rEBmwnv+UK6lX6XvMqkqTevzMSZkpY5bGRSm0j8x5dLugCbLqa
veIuuQMm2py5X2VyJryB92g144Qj1rmT6w8zgegI2LUtfoNSCbFp2MWzLs7Nt93dtBIkrUwyT3Xs
W4M7+fFNmNxYLak/KlZhx2k8YxJ2ysOQhXACdUzOA5hA+JL0k/Q/L5W0CGP6LQEcmmWBLP8YmASE
D4SQbANBhobSsmnhpeu0QAMgFTRmh/c31cbhBR1jog+XJZLCtK2ryNS7ZtjgRuK5vvlA2g==
`pragma protect end_protected
