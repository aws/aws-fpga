`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
ktiwXDLjlRh61+YzhAUMNj3bubIus0Ldin30PEy8L9dZGpoj1cc8WYjIRlqE5YX6HvCx/qVAQvHj
BxV9lBOSSHx/a5QADuXPcIXZC+c0rjqGwXylRD4otBKWPvDwNqiZZ5VdbQm3a0bmHZsN3M6hZvFa
01n/UB4uKYN7ZJcmSeOf56tCrUxnB/CVw/rCmO2IcjrzAVNAWEw9qDGVGwlquJ8C4kwmc2JvPNGQ
1UzGhH/dCNgpTYgt2O01Gi4qlpUEYBajVFcNmbUyPBGOPudmiDBeIURyDCHtP5gYdPVFVNlFd9oP
vmjjOQ/ZBl2jCltbqLeuPE5C/nw6zfc+zm0kkQ==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
YxKD8XU1FkzWaKjaSBfYqBl1EAVsaWDJ1VBe9Mm1v5N43k68HE3tgAHanybvL6wYOxwoWAzpK2oF
JQU5nDydy4jQxPghElz+gqFMprSb0Yp2iumR+fQhyo0RzCkD31ytnouSN7EZMxsGkqMN+XJmvoQH
h2yge1HWa3dh+7NpZ1U=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
VRUsd/sKiUuuw3WE95oU3H7Sk+WBpqirL4nvgIOUw5EhnoZK/AK8V1UuR5e/lN1x5medPHdwZqJA
EEIOlNcEHOxLYoPDtB+MxMYdXZcyNs8f0X8b0x96JSOCiX3Ioh2QesjZ+TZuI0u6ifLK8OYfPlG0
QKgaSbzASLN+F5v9kac=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4080)
`pragma protect data_block
az3bR2GadHOYzmPwturDBJvjOWfCOmDjTMw3jb5IYvvaXv+Nolwb+RxeYQgHzkJbGPbnvUWccWDH
OvNEeBpZKnltKOYkcpP+xz2LWU45PcimwNNkbqqZJKTxahn0AO4Uu/IM+hDItArRB5cveMRuiIy6
ZL22Djmxg1zoCJdyXCs4pv/9qpvGF1B2uObxnPn912rd66RCZvReyQXBFUUoanBHDkc7VFGmvxyv
kERpkip6GMs00y8vTEx1DJGm8r6BTJXO9NbK5T5A6iIePpsnbsI9H5rL/rF1NIbUTXdqgyH1h7RM
crAboEgui7px2Rar3TNVO0RCVqSnbB0imyThgtW1juwmo3XVRlgWqF7B92/EFkNjJ71M7qbTIxbJ
w6OY0+PXhRxltMtcteHv3MOekk1I02quP8Yu4+Ckjv8TeKCkQLL5pFL6/hdc0Qke9Kawi8vF2YUh
X1i3ViSCID5lHC5P4MYjEp6v+efdFdCVWrgvQpKzUuONwrxg6rgt2JIRNU+oTqs63rnO084JwNDi
QJcCyh82owbeWn0TM3Z8NKbUd4zwK+vQ5g5l4EPzOBRYeac3mOMcl3df4zRoq7/GLQUq7GqBePbE
Bk0ZSM8sIT9M61IE4/iWdiAj/XkIoR/go/bI4RP1vhHOjTfePfQ3reJpnUA2skTVReWLvDzdFryi
MaaOpBOjODfREls1YmiQisa0h+jPK5KojHjhJKXKX9Fittdc6sccmHFVyMq2Vj3c20fdHTtAxwbx
pdnmEWLVNzH5MZKTpzOBh/Yqk/BAUOCY1CqWfn/z2tDBCZgTQXu+TvB06f0bGMWoGMcpZ4ChGCfp
l+pZCLq6yib7aia5KMSkL94HG7IUB4pMmJjazaLt+lQcOQk51rjLUboqYlnKCQnxdB/1NoLZG+cB
CNsCcVoTOUpKCVXxM6GMscTM47N+u76QJpO/i0q1Tk8IHjcKrh4KPs3IPIyhURn7cO+3/ornWzJW
d41CEAK5s6SHutN8zp/kJ+zVa145k0w6JEXlzsKXWIBHJ/CWs0C3NzEhCLJnAvZ9DHBAD0zo4skn
pXg9zIEKjCz3GRpcFO87hYDQNTDR8FNQbdtWsDI+lmC4IbwkdCq3LxrsU1ftdkPkxy7SpvDVeVLM
nNWBIP1GLoN7YdhTvXEQaLBOlcM/mEQ1PE/ItXjtHZlh5QrGJBxME5t4lK1SW6pePo+quPbKYsKk
sbU+uOyBdqhr/AQKC+9Ofr9yDynp9zqqxendSkdnRHm0OJFC41Sz91edXnvlsAPaJEvkBUFkfFZh
V/Sk9iTERtpoP+UEbyxW5vUwtC/aOieGN7FHzcde2Ao6MH7Ite32+WENUkvlENkDv6i1x7egtiFy
YNxf/rGZ0oYyI6fIMFn9nhP8VS3o7LTeM/GxjEjsDAek84QKmShHjQ9LLy/jx05vyefFr8VcY47o
lKBOHuiii6XH151aQKpxOvvm0BU0gAwHwZg/JMp9uHt//UhqPMaj/+er49qslRzYbJtWGGCIyTXB
UHV5sGs3wHyRAubegfTWItEMBjNMdwAYoNtcB3dSFlFt74eaZzbYkOxASqjS1XlRMvKBb9ZuN79z
h+lPymCyBKNgpAArsp4AUSdSSMJmDIZLL+FgIAMyHRcNiHOKr3PtUPlmUM6LGcHgcjCt65Vz6p2C
4w4GyBxjJESbZ8HKPGVmhU6o9iuAYBNjMldmR4ZRHRZDQ9k2UsiZvW/3Pgk2X17jekjIX1TMHNHG
2Zq3dt2mtdf9vuoD5VrqwYtMPk6soVdHHr+G+vFwun+zV1dgevinL0ETdOPT/VbUPdi2Od7M/q58
EhmzoepctBjwEwVkpIysHII4l2CEGWRL+cWezKiR9XcOF250ftWZwicNOxshvEXrc+UkMCH6mN7M
wRdf0LwrYzdjv5BKSbKQugS7wDA0MKDew7aqxtFw2UKiZToZlJz4YxSUdhE2w4kRMmHK99P98+Uu
WxXFGZZqJVepzbyc0N2K02mY1FuAeazRiWJ1psvxzAQ0lBIEfe2HK3WvaERcxexaNfZ1utjqcS3A
ZaJwXmR/g9W4J2xiYPMWbblr8OFkOh8533vEDCXFoeSzmh3ZvTEzWHJ+1ZgZVtTapbMaVrGNaQOQ
VKgEyWmdXLGp0ZoITHx6jacjqgHEX7DYXttO5MBQQOs5UuT7oV2DdymSqsoQ360IsG2lRD2BrCPh
s52FHFVzi+NUdUIIN7LTYaqFtQROXvCo5BpD/9UbC08kX/W0JPOGQSv/yQ8fTbLXZXN4lP+C3vNK
bizXGdKN2F1TAj7NfZz3tgdqP4WoxyxTGjyuVGjEH0shra1I5Oz1xX5/lOo4Rh/eJfB3fH3r1lhs
DF4tJ2mqHZeelI8OCVkwi7NTslmgh5Xr1Jh3bUjOzvKtXDoMlq59TYiNP2iQeLtuRSDdGE6M85vE
g3QlwH5hEhB9DD3KutVhkb/rzPuqCaRiToSdpf4iNcjasXqfWn8iUbv8eoeO5mbPubWbk2SNlqDs
sDhdkjZ9aW2zMWxJVCORInnxKpUkhk3Aed6g1gyHKimgwoIjk6iQgoLxQ0cAf+dZWxnQj9LOQSB0
49ItnvD0jJZf2QFaJia6e/pDGSPOTStwmFTAgi885kn905Bm3W32jkUvRUSOlmwS8X8KDbcpBiG7
3iDgIhAJLLQ+rP3zqx/qZ/9CzlZTX5CxlrdiqZh9W7Qg2AdLTJhQgWUOmMUsPFU1pHK85xak25ZH
CupH4YYMvnmmisAbt8vgyQjuOdUX3rL+WEqJBGm6MZRl+s9dqngUl9nm6S+XwM+lkUMoTnX05gHz
G4JfNvcP4Qd94C0bWkQkb+L1Y68ua/Syu8r++CWVsAVRyq8CdUz4utFDQxA3bzaJoD5hEakolAny
gDkgCLkimNMtA8RjfNlKHX1gfn5rsOdAIYTB10tsvyaVelxcKGpglP+9LnorW3atbSPJoBfdsPFW
nHL6ijUGaBBqawNjZzxxUqnez+w+B6YBHWdGCHyBxiKrAfAZc2LFI7HqKGsykbjdLHONdpmFE6on
GMXq5oVcTRwcpEbtJxRJyb5WVHcZ8+LmWSGe+0dfwKBbG+0dfOfsVR4XD6BBF955BQwCfCd5+tZ2
OsQur2uSFqiJBG5i59hXnB0jxO8Lg+JcOLLrst+pDh4JF6ghIWF+6Wx+pfbj5zlTlGu4GiiA7UBU
OBeiVDfZMVXRkfdBPEDKAwvZV5KmmN4M5c0p6r6c/9QgUZezWViXyyLipPlM5sh9KKm99K7Tiivy
nbTRnW+sBBJtNfKqDdREXPIboQouJjs3+3uC/epvw2AGOydLwSvuFV02v7CilzXFFZIYwKR+oykq
xnnN8KFETD2blm2Swf7ssTxEchIPWhPylrDsBGvnGkzr7riUGC6na7cKF0DcqfDxF3DpFhTYJeKw
MJJxLHH1z6nEN5O7XkD8oRPGjdrOhAYikWamKLzEOYHEg4YgocvYmglnuqqqGIlhixKUCP6EzTBH
oVZdaC4BKznYG7Wbxj6uSCZyrv7VMWsnYz94V4QQnv0lAXJYjSI60AjPzP2fthyGujd3gDy7itgr
bNrOVKsTMcSNb7Q7QSOSeGu8AJYnn+asJuMdm3ALraJHAzeVSHtqeLUjnptSkkndP5Rxxfbkm+nt
IAF6kPI4Ex9dpiU0/7CvhqE19Rj2ObnCUSpenell0AnV1EZZU1N1ehuZgcIzhqnz9NE99iJrhBqe
xJX/6O4tSaT/eZTcsLPJ8s2H0b79EcHbnlYqVTcipIkCVj2Rw7FkWIBoW+T+8bSbLa+dALUx7ay9
BOwTvgtII5yxEHLp0DdYthcJ8pd6ftcyH+VyCGgKTWC8CoM2FfH9miLa07OHp7/vvwJiQ8Cnf38P
VQXegkn7VYLGSg4nAMghSk/zY1q2a8iJ7mRv6ZqyEPHu6BfIrVXN5M+mZd4aGORJr1c796qRssYV
B0RU3YnUhWsvovxscCVniPefm3i7F451w1lTYFztX2G440QIxBVav4JkzyDChCXaWtpGaFahh1xH
sDCAcJXUuTQxCSpA5D0L+OflXcS5jzAcC0kNeQR/YiNb+GnYxObClknmjULaIxqOShtKpVJlA4Sy
HXhVsV8ZacH5HbQ8pwjK4h+gS6/p709wVECMI/uLmw7tAtOBROZbe4jsMMvmZIq33P+gznzUKOAO
5H9hncFR9XppiQLRdmo8IxCtfPyv5q2feRP8kwrI3AwBE8sjjRUBmoMCzL/hUgDlV2RaG/Skdu14
SmIX/z+Vgw1ZmtPKOj4I2yFFI4zk0hh3O1br7g26Xg0qkMpcw02iuYmAs60QQnhGooN5Anxd/XLy
bKJIjZwbpcb/FPxjFLPSmbou3MOA+0VH8xuD4bv7NJnJqNbkRwzOVCN5u+TnQOrmK/dBVEtxC2d0
PvxUnuRkqvRg6eS58DAsTn32K8VyUCvwk22J1W6oDTziCmAYlvaDNiXKLyEHZLAvVNor7Pa4jEyr
5+qVzoy3nrKhQ09rwLEcv3eqngNoxW8L0ue6/W1fUguQCAwKqH7HQXuA6jmGeYWwpJEz23kIPfad
R0DxwbNssjmzGpg65kVdMyvx+iZtZ0vGlz3hyPj+GEBtbc09hQ0AbFfnWdhuBDJCQB2ZQV/RUsh1
5NL+pXdDOvAKJS27OZy2qm+GneilgGA9LcxnXvK1juuFWseZkpms48rmMGwYYeSCikVt3uva7aRG
ogoCX8Yo7UUw8N/Yk3HLE06nqQKA9+NbcUT4J7C/Csv9ytz0M7Ulrq06W4iTWIoCMdb4DEnZ8LHk
7sdAc6hjRtHRKPhgD3SJtODj/VxE5hIK/LlWETJJsmd9qXg84pZVd7bsexRMG56RTm/KTftMPb5L
WC6lsdtPD8GvyoT9c8kT5SqjAYbMgLLRzUKQWKm8k+nqBdjZ0lwRBa/KdNuw/AT5oXOFgEWEdf+W
RLS01bD7milKtnfNdsjRgcB480sce5KKpZtP5q/RXUR0T3/hnzfzSw8PDadaRdrSheoufMPKYtrA
cK7RmfJ2xd8HrC5NfJjvx963C8FVMVqj/g8sjHMLTfDbUF2uOg5aiZ87R12haKIDWNqd3yZrSG0f
7m+tb1Mj9PYj3j6WkOSgmHeXQa8ENNvuVoTzXrlsxFb3BXGz84b8ClARd/bJMBD2kKhTYwSpQtTA
TZAr+1P1Xfvcr6Wiy3YS+OTtGGttldYZM/WYwCoJsaBD5RmIQA9iSzFiC3Nouj+hdZTjvY0Ev63s
x+ToJOkge7iBuCkouxLsthkguG1vEK1n8FTStEXgehjVScX87m8o8w/slarTmqWXR7Zq3W+Bz8Kl
FvNIBe4KBVl9Cp8ehWjwnvdQDEBj+5zG29Y0iSlOsEDjgMFVj32TMEGlnfYnwv/6YSic62KODXTv
1whqZo0wK5cnoZQ5bKvwvHRATQLV/fIycpDqCZhwiwFM
`pragma protect end_protected
