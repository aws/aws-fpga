`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
pl1HYXi/oNiYYe0zg+gyDjfei5wcEIEmZUtSWWYDmBTfFbovttfIaCuS/tmGGcU8lvsJH0RvH/+k
RfUpMEyIYDNwebtf9fTTteZqtv7+oemOFuF6N0cSCQgTblZ/z6UxyHfUxc7ncQ8G8uA71iIs57/R
PsrTMwlZ4GNDazIYvOgD6ZOGSvfN815L9Xa6KLKvZ8VnH5yMqoYrOEJr7iWBbuHdi33mH+J/qawi
YE5KZWMUzCSk/Jrohs9C3cPAAF/R/dPT/3sLeIUIRIZR9fBgW9twe8ZhR2hifwkw0BwCjKL3rJq9
bBbUfChXqGHuc5yiDqzreGCM4IRsi5Ngz+OxYQ==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
gw/7TASz4aZQmQhHDU85zbYc8CaKqNd+akN4YJhweOtAJ6KFp0uOC4gJYHcsC1jWfZri2E3W3oD3
UmLZice1pYMbjTupi1fivtaU6WOGQ/EQ3lLZ5PGHjUrS2R1EC8Y54FjW7j04NiILQEBfW23N0lPv
uxRUQhQ3WRbo8sYrx2k=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
T3q4RlrQdNPwa91pn49cim2pYiG6lSzWmxM14IoJW5zhJKP6c8EBl0q8I8fDUoZwzXWFOZW7gDd4
LVzydiuVso9ab5lkkxjD52iIiRCUEZ2azux/1RjVeRX0ZBMAaujzl0TvXW4AbBaF6WcbQfVhIhaS
7XzpHEp5czpJAo645UQ=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 45184)
`pragma protect data_block
lENwy0CyV92O9JAFE3D+Dzxp7m4H8CcAh0xPwmq/uss19drOQCj3gwHvJoBngmJYuanqMFM+oz+H
ewuZ0WsUBfiK/S+0RWHja++3PBhd+d6thhU9FrYOQS69qZukclIAgroh1bs75zb1GcISjn+Fk7LU
1GdwOUnfgDawfcNpxkjEActhXwhObqg9Jj6NkHlrhaSOk/NRrreNR6YwyC12kOcZa2K6BJg0IR1d
mrzbRkLStNTxNF5AKPUbw1KyO7aMHl8YGfi0TBx0V1xeBpOdaW2iXktgBt8JQLOIVhkkZCR4Yjpl
M4Cbdm9+w1ipgPl/aoWnBWrR2he32qm2c/IjwclIJVzsKkmDO0VjUhTaOfMlCcTRs9KytCsJauw4
zIegnbM0TYesbooRKgfbc74wwbDyFq14ZWBA9Qv8w0iEoB1pyIlG442pJ+9nZN3WcGOB3xtUsD20
PJTNEH9dWcd+iCD4eF9qbDK7tJszaxnSerr/nau0xXPw26t3CcbJPHxnblsGhQUGEN0I2vDIxr/C
gMlPQ97u93OVxzjhKzHWbFJwHlJFH1oZRMFDuzqIfrz1pMlYj4n+zdcsBJl31Uc0jNZLlUv5iRm0
AlW+18jD7zI/TTL7k5UeCSjImPPQOfamGZjUP7HHSCA1YumlF4JlzF6Q40UrqdoSiYxNZ6QL+jXG
/LINybBhjZDQ1YV3k2Z762PqXuEmnkpurRSNOhSMPIzqjSeLZvrjuwREx+7UT9en/CJ1OYzdqNyh
tce+U0EPhrqcFM6FtmTSg+ltQiTkjhtkxGk9wRibcago7Go/pfkyrC3F/kn9sE33gJ2YWKbWcfXr
lX8q6PotUhPhwx9NDR+HmnHtDDW0aWCfbF+yUJmFbOyew7o4Df6j+K92tfLZnI4pcKOPDl2ns5Yu
hkZKAG8LPJV1Do3oj2iTKPrxtONHfKkBfumHV5Ws5ccsx/MwstF5CksuOT97+VKp/vbV+dfuh9Tj
0bKpUdIAw7gi8/V8Ez8epy2PizkjMBUaRqNu58fYWo+cyNvKD4k+uTymfPWT6pNFjgtsh9BFa2H7
mIpVh/RgpZWhSzBLGBCh0JOSuMZ1sEK9xXG9z0xI1hcTzkG9NsYaipoXj3u7FxPLhopeA0z9so7Q
rbwdGjj67ICopS4XkG71vPuF2cDDr5HmnTsv0u0rKXx/rOZ2Hz1mQxHfhIyFyhNAOS/Mdzn1/WD4
Xjbj9sVM321ZL84L9+SX38llD0XumSrZEeSnc44QDgXnbbT1UQs7UQ9BoaJWSoYBj6VsaVftWVAS
+B2XYOjEfYvVxavxCKemsQMx8Cj9Cy60B68BO/KSTY7E/mmjgBJEhthGk+GupASAGbzzU4as18N5
g9fhaMUY07nRrYWJ91Z20mRRL0JXa+uBTBdZVyORZWHhH0FVNni9zS6Z4atEy10+WkLgZj7+yPsd
Qffyp3cKnBUJjUqSyvNSKk963ucCtMAAyqbZgW8kc4GnAwXg/fJbFbvnyaxzKT47sh1/Q5xxo+MB
+B+PGHMeQTAhdm/v1QIO5YQDt5a33EoojiI8MIHYJcgDByXU7NlJ5rF3udY0Xji8lfwnd0ZLJTdC
9LLWj64QXkaumQOjxPDz5v+D3u9BTQn/7o7qEq2ZEpM+mTgAgxoqcDL868XVphHekz71YKvt1Erq
ZupPe5p75YsXz+FuBPViHC6x4vKuMy0q2MSIAqQmOrzljcjPkskCQwAQ1v2RluHSR+l5LHOZk8jR
7KEITzRn6a6482WApPjSS2Vj8PRXB7LtFRNgCGEbgNH2h8+l3uZd66Rwu5GdwoQzYkNudpEsGdyK
udMet+gS/gibneo6t0kD+Wr29QlE1u1I5WkrGOcNUF+xirpXMnIuhpdKW+v5z4bnq3zcRm6DqZ+5
ascWXsfvXMPKgV9XIx6eScYfCZ1k3DOOzNUmhGetbXlRCeNaC7qx8rEbfGoABObmuRBwVQee5LoM
PblQYPjhPrslHVq9D0020rGcg4UP7MeKSUzApzPrukZksUdsfNOb+6aH3RdREJGBb7y675VGYnbU
URhp7iBUbWov/SP7+Ku1kSgLE9W/MNwyggVPmdzKsqCy+uQGrbG9cw+z9l2bMKLDlsL0Ycu1CwW8
yRBOOo1db0RNqpzRZhWvKsxA2a+S1OhvRpqb4UgoDsE2x16032nHZDZWB+4xuXme+1ul6idLEYmT
vWOXMvTKkqM1eSmFFVVSI5V6ZSmENbX+PX5P7WXcm50JwtG7BrbyaSqYKzfZ78bubxVnE3hfvyp0
KxzExCQkb21yUCR4ZELQ/jiJH7gfmcp0Q+iUd+P5+wG7MH3Y6GNgGLiDHzPBX+IWrazBRWu4jPmg
YH/d6YKGVDBjBwRxzklhcvvmD9Z5f/EWfYAQBZEaYmToC14q4SnnYdxGBFpU4RiW8Rs7ecaeZO9j
cJ+1JGoByNATtHxJ3N9BeXxov4XQUzoM7ERBn82eo7ASebnMswLc0B53GSIyFs5TG3ptviXHS3CN
47vPciz3myHdiEDE6AbWX1XTON8gdcpEj2uExB8Rk4j679cm8NaTiKaXpyzWa3F2y28JMLzpNEWj
JApoi7QcmFSdxtxIfWOfzKqP+RceYbAM0v0zhcUiEOppIf0hv16/sewhUO29mGujv/bspHcOnx5f
PNC8QyHjWtvbusJOvxjhpZnfYuKQRdmklDxoJGT2N+FfWTxfd3hi60gwyoeV8Qif77O9Jv2idiBy
AzmLL1N69xKplpZrwOCUxyhJIc/jV/IIKZ2bsHw+9awjQpsKUadqwe6MiTB5ZbizCc54HvDVjAI4
jHrG3ZMwgPl9zS/6TOoc4zBvvUflLWprr9zta3I4djFwLCL5YLzLwIQNS+g8MsTsVAemaNDRB6Db
w39cBtJirVlVkkzNeYcNz2cwlppb0H3Mbmn25iU1NByL9Nc0ej5xYbmKUuGMv5PLtLHzGXk8kfBF
x7eUrDDMZjGLtpUGUFeW0P9lqAfvjM8bymSSMO1rH4hRBgCZBML5Rw/5vIrG03yJ+5+xHp2AkWXD
XC1kaSJBKShgjYF0xbm1Zf7LP8GlnsbH9qYCZkZ0wAq2MDu737cYdVPNHjbNgoZrhtTvkyqvxEfs
RtS3BVBoYDgsIxUJYa4ANQil6weW4pdwz9sgd7Ftt1uxsZ7yigkL2f0MpZj9rxe1E9D+anAZnvml
9J3UnW4rbKhtwoPdDFU6p4jTy9EdUJoM7vpXPh/DDDW3541Y4gZkMTwJG7VMmUDxsohlCM277+ub
2pLeRkFLkHZa/+PXl7xcoO8rH5XEnmOgtsOj/39H8Js4YoxdYx1jbgL5VzvVttXsnllrUAUnSSmO
zIbzSOHtLoJTET6/D9igma2vJbK6Jr3angq8KqUANbcadqM9pDGNd78lkmLqEJnJaeAbRQDECXFe
olYKyavZQmb8ShCtN0cOmnauv9jOpNaHbkQDV9wNgb8hy9VMvJywsGWI6pIdS9uFR1GhA+NarWEB
XNYCA/MOGJqn6+IQEBPDi8J4TQAOY5eB0BALTbhdJK91Bg6SXwVmtug48YNP02aVa9ych6H/NAtc
V34OAlCEbNOksus9nhmPTmo7SoW8qskUhtvnLiBo9dldJdJEDCW/eozslFUqNBIzwUJuuln8q5mV
6UgVkrg5MEjIvlhNFhjtN4LWoaXLf0HdeT6RoF1klEA1MszbnxCO/iavxylz9Cz75YzG7UpneZ8E
OhF4UNvkeOGxhnyc7ILGWBQVIzxptM/XlArIqleOgz3gdJKU9qBpGHhvHw8q/sjTOTHlGthguC/O
Q5ZAHsRa6fXNAdzgx8W6UHbnLn+lRbGwG+7q4u0GaRr0AUh831EMoEjPZNsicLZPsxltEooEgZp+
k/ujeqsVBV/wZlFPcQ94RAmR5O/urJC6gFaB5E52TACd5gwoROtXk+1jYXPEAcSPkjrDn+HqHp+B
B8v5zELHwx5lbyJZSHTqhiVimkCoNJZNEz5n+rIctAGmEDrXDMyWsLoCdpPrEBETVTCSs7xfuRPx
WgBSqhXd8VDqDluFVEzs+D/crKuERxrbNd02tqBPyxBSJCi4FaXs82PElGPueGnPZErCZFSJGWj+
y3bWECsRdLSlJZ2mLElZWxhubaR3hLGSLMuH6FHZT0AVTKUXMqsBcmu1gKcGJiln6QbFuOEYdw2j
f884PLnLj9RYJ9UZX+MIqdPWlX39e6CgEf5b4+iWDn1ezs23p9s6u+X5ucDbBfJFYSxaq+sdpjzg
k2N/0TBP4E/77BGbQaHKyQsrisToAxglziRNW6hPMxXqAdbyBLYiI+EQ38O/bCYTU4NNoqYfwSaM
zXDlt/lQvPrbVjgl6WhBKPiN1T84NwqDAwxe0S1yG6lXeVVHnmp7rhsu9kdqerafpEPfo0zsuJdl
aFFDNu2779WuEH1opKsStUZkNIGvoGyWzUMvr1FkUfW7oDu0iUEJ4j+5XIi3uSNIMzZmu+TE8rg7
35Ire20luDuJQyXEQiSZHK1ta4/d/TeDbjagrwsS6IGHkblpgm8Zk/Mk9aD9TVQysNr/bf/jQYI9
DLwJVOWwjMMiGByTF8Lfq9rme5CQ/fsooSBnduDQi6r0Hpn9d4cv/uxgtkOfsSMXbmggagySF/x6
H3bCPDJrfnVVCabBdnw5OiwQvozJkanh0achcQsuTaA7Gn1n2q/upRC3d7oIo1hzF8loER55kq6H
jxgGMB8pfX0VCnUxvWrV5RY345urFkzvLwwjGz/MtNAxp1ZPJqC9n8ogXFeIIA+/q56i2ZjJ/2PS
Sp0dvIhfnLZP7W3U5cw4OrxFP93eloWSUhPBqmMb2UY6FVi8Xy86bL5diygLrDANgHjlWsZVqMu/
nQyXdXAg8TswTxZlwbt+oSJwBpnfnLwhraLuBlJbpaqft3gSe9imDNAWG11U/KNkXqvX13CudO2w
f8kYMsDhWGE87lSRsOwI5SQyD9b0SGSReH+W50QPRkUV+lyTYqXY7NzD27oINNpuToFowMthw2LA
BsHykEXVHmRfHvT8XHovCXDPjqh/SU1gqTPB1HB39xsX84Uv3OaXInbAJpTrKk0S25iETXdUfd8K
M4/xzJAnrIkiK06PpsCdEED7ByBmNK/lMyKysg/mdqhZk/dqQtKKrq/ZacT4oYrM78SIJqraL0Kq
f5H0HwZsLLJvJNIYWHxzJPRV5xNvz+uK1vg2Mk+OZKPS4PYYNG3YIegCUNyMhzlGlSVUMEPmYZAm
aK7DAW5HWbQt6UlhT31VcOQRj2MlSO1yCmQiJSYwrQm/mR9ay10oAwh+plf0PjDgEd6YufnLW847
agYiUCWOTqsnlgKDg/fAxgssrEijGr2CByH7SnRGJrl6drCPsFr4lmMZQQVRRXkqKHCyelBxsO3J
N8zbuIig6bY9utKugmnxyuONg7Sz0lE70TSVlDZJe4+ItnN2IraFE1UH6Dp6MBf2asqHfWZ3ody2
IoJ4jicFkXbcH+LDmihRJcVvbk6P2cMMSlIbtHLxkPKZvQaC6Kc9bICdVDXl6AS/ITR9vA9RAdPu
aRnICLjGKHfiLLBzjma0x1FpOlBW/s6/Pvy9/zM41Inz1E12vPfevnyt/zLpHFT4srx9+UXbOKGj
pvBlzKW383istW9I4r/4wwoccNzI11oOcZB9k16HbGaNL4TJcdzCPOyUzJbTskWRFQ8DPNSBs6hJ
deHXG8TAbz7OduxdSddDhQ6rRM4kCKwLqOJKRGi0OGxcS+0ZpF1nKuMqdoybBf8qqdfahipZQ8+k
qBS5UBGuAXYK1rmqL3MKhKznXLAVop8HV1m3VvvIzIt48fuNgk+7TdLzODsiwSSsTG1N6eZS6YJ/
j/BtU3dQ0pVN3wMSb49HbBOULtaPqmYl1W2+fSXnK+IS8EXVAIPcufARya8pTN/zcSjj5G1bgCXT
4x6hcRGSht3ulUaXhEmNdcuM1yru52n90UUueqAemwR/7sdZY/hvPNUlrfOkdnCNx37WV6dxgSYK
XsZXBFhj16/OoV/UtVS2A1I0Irevpq1qFJXNCI/2eAHY4/LQ14krKJ5YrU8rTNymaKjDjcSrgEqN
HVobPLqkX86ppffkGaUJu4igeW7/USblM7/zi/6HWwvOBLq5juRg8Phzf2y2Xk6PlSeOb01ACAGh
WMKMjY9iHoI1CiTjcOcyMDQ0+cZMy5B6hRlXhrnH1Fn9iJiXqu7cQB1MXg/Zj2XN3BQY4WmgAqUp
E47t+GcmUan8Dpp5TnSN3Y5W8HTAOb6ctISXi0Iht6+/Q2Uh9rTu1ZwmUwOMq/DyU6GBKfnruAMa
CQnDfbJQqvglrePP/cnTrwZBTNSte7XxtyUNtnkQQ8aFJ1sHXPRgmHc6g9V/Qrljrh5ZrLfGDwcR
/5CmqWnuIMP52hN2okHr4TFRMFnu3OOLj1DQY/RWV3a9xkG0++QyY8zYqRC0yoGBaogmahN0cnIH
V5mnjzS16FfOSWkFyTexhuy2lYpera+HExDwww+AqFo4BArRvC7jWHzvysok76eXnm4ItgT7WbRL
j3RhyTfWnSeR3xKeqWHQWQjjPphtoEKQx/4W2SabXPax29xIr8ATyT7Ve/+zw9IpWFjAP0FS+AbZ
/tx8XOZoaPAAt5WLrKFFWjv26c2iB3SIboywOGYiv6Fl7DogQUg+ffPRMDQX2Z0GpFKW+/xaBxSV
DfyBnKhwunX0RLhxprMXGRCdAKONG9h5sp8Fu6N2m7wpr9i4CrgDK6PjZ536e+ALC+Q9uK94r3Q5
1b8kCo4Rm2KolE2UhA2wtNX36vLSQ3apNKatFluwd525+nxWz3mIHyP7DqrNwMoPlm8/1RR+ukhr
wnhIKIsCuhHG1+cutJ93rAInmpcxSMp1nWVsZKiSHK23C9coNQ2BsDc8M7cTk8Dxr/hDwQXcUi2T
R3NZ6m3ehxa/H22iNGPcMnjN0VQY9zserfGbG2bAi7zQW6h2nLlXep47NFFRIUxsRjE6/XwMMHj8
4zhTuRCKiTf5eUgnc3qrQuGxsDzer4ecxzVaVztovAaySIW+VLbHAWICoGf7liWo1xGo83XwpUwR
jTdeUdCfPlPy+1phdV2X3YxDZ+GSwjqUSR1UiNQFX0KIXplJXpA8azjcLfkb1UYb1fdcTolDFDok
N8SEMMx4o2qF22SGtLLI45ntXVeLJCbWntnrE44OWOpb0kbQyoBqIW3+VWvSxlTpl1YO58JYaanf
vrW9iRMEh67YqlTc4d3fY/KDk1lM7HjuPFsEB4BY5YwYW/r2cRhNKByroX5a1JhbnbKmhxvuD1ng
fzyI/vLRlYUL3SumSOF/L7SVdcy0PS07ib2icjTdBxvjlSJMtHraFaxVJLyEHLA2Cub7CM2xhaol
K9iQsZwwwN2p5zPLCKJdHGKjhLZJu7Ka0DvntqGMx+rDGe49cqq9b235DeUaHtcbfHWNQHuPiP62
X4UquK3SHDFUp/VGJ94b/ihDhJ2OqvTxTjlyDc7ApfPGnZY/tVmufbww/zyotBdCtCYaRFYstpSJ
8kZLV1xVUgKRFq7Mhm0aWlTvNw7IG3wAm/MAjO3Et5K0jcAbHWbwnFuH+gR4CNMKuvLa9UwRijuv
ltrxK58WIMR11gdkMGZ5xqChhXM+NH6w3r2fqnpUvR9dCxYRplELh+Xq74IeM3E2l87DNbVFfsfl
iYB/7qy7ROABxC8WYyxL/1IljvQ3pSDizd1d088F5AtOjy4Rh3fZmkUPBTME4vAdG4rpkbyLQ2sN
HXSYaw0fsrIsK/wJOHD9fDONp9MksxsQl8upUtmS3YMUEKJ6gir0xQ1CbuXUWgEwx1KpW50LDzef
orLL1A54zLG3IbenRBSPd371c+9nfSFvOXyRl6QqrZr8ZBf/QGnvBxxKXxTr5Ser/6Ja/lU/CANH
h6OGrzJ5kxW8Em1KwMoHAbnIUKa5MEAWzEd7tPtU2hB9kIyUFJ0d3WlhkrX0C5pLmTwUvxuUZYGH
ZhmYq/mSKJhTGpx+z7c+TNHmhQUWwfJXyo5WNieklFvXt7CkWsuvP+NyPS9x6FOZdGVxlLnHe1tg
aL5tuiFqTA1oJYmqoY9DZcQx3wIZ9qGBf3+UQonIvI22JmAUj5NDfdxkVnD+cMspQHab7I9bC4Ki
wwIGOsFVKB4xxnff4meFiL3ZMgZSIh2SlY5bBrDQZAZL10lIrgDBiOKKxyU+1a22gTa32RWtd0Zh
MSDu0D5PcrygwhHrY+LNpmskWui1cu61oK2nCs7X80gyqxvg/j+HPZmhU77yHBSl539L/EeQ4KDY
CimsBSKYdmYjK1IvFsivvtj2nVqfYVWH5rIkg0Qnra+BvuGDB2ZzHCqyLXi6fTBrJdyCmb7vVcgp
boyYQMoV3B7DK3O5SkquDM9k0g5oIOnRatIixTYIXWgofqaOXg4dxcYUCp/SpYZssxQOGeU5vfJE
V7fP7MsQzFiTrdt5ZeDy+OxARezreReTxj5dLyCd4q9phsHOZeO++2IyvMSFj+7xQcmTJ7swUw5U
dP5LGAs8eRuXX0agfXWdN4pfEGYFNPa+cYc2GP3C6ASL3WMvaNMxMtFFWCeAAaLXw+39BN5I09Zn
NecVLM8nYt2AYZQuua7jvhxzHKBVBJybhpynmeM4NpjYGNQR6moMZKZk/pSsDM8b+guH/YicA9ko
qkM8D4cBb6fuZ7E2lPf/A07HFfb9ePM7FQ2yaaxNAfnJkEvinw7/MkXXTck7TIKeYhbxkFDVFQO7
XArcg8LR8ZPxtLMPC8EZcZHj3SHN0ATK31db779q9h66OCA9naxYjlqyyjJx650Y/raGRr6vxCi0
RPV3wCndw1lWsvLnxPPZlZDmCvYhlKMZA2TS8fAN/QIn7OjmRj3mfeHbp7kduvlOLpZUHIcKrM6o
WMaejGf9SYPHGkkZBKHByKgvDRxmGndNgI6EeiAxtnLT6eHhI2Ss+Bgt8GNMbhTYDCcr5UJ8Q2M3
7HR1zhZqt+kR4tyIjYYWLMDIDwgheswqOYcWvvgJEscf2KBRhbZWTNnOTyto4W7H41QT0T9HVyLN
pX0CDD0X0Am8MMabaMcSSliHb2yEgYSWw5MYKfmFhbgTDvJh/GsS98bQF7pcU1MM2tRV+9n7vREC
zxJJdrRulyxEXcuK68ZFz5kaZ+ztGHmKDV3tClu9/pVPVPZTzZqDLZ6zVLKP3ynSd34mT6f5yai/
bXeIbx6R6z6dPDMMRmyU0zdF1nh+zyZvpXUuT41LSDnJh7NoOD60LzTqAjveuhFlVHjHuGPmjHg6
JimFyMPkf9J/yq6NXnRe4i8KmqNr23diF9KX2H6gMKHisDNpsYg7tXXWbtipPhgyn/eGsKQCY5N8
kRpr5JlRMvYAcEHlsNCm+RSMpxibZPRF93CTa9/pO9xZFFB0sD5qD+/mJl42BUoomIxiczRTf6C/
qgEUsZ8Bpmo7qvtvISd4w3ADYHA48hFV+bopjwgvfNyqK1ElM3BNZbqB+CdviDLgO4/eJoSnYzJD
mKlHYWiU3rPBJaUHW0JqbK0rZGf7HUuq4tzqedwnUIZ/QyuLBp/6BWf28ydySHQlrp7Q+1gkqXek
dmrSVr2F27ZsSh4gUHsU7yRXLpVx3S/g6pZuIPwU4sSJSAKiyo4mdL8B+fhvQUDeYKvJUe3n9t/l
1KnjeqAwvhR/vcaMV8dLpdaMFepZ8HddbR/ROyvpxO5yYuVfWy8h4bo23umniGyQDDeX/nr0oBFI
qCqFPWT59OK5d6ogyTmWd9hQ//ogTa3GFw4rzUYx4rRaRTNt6VVF7a1ZMeujt4sJIAYsSHH6MAPN
WuboqP1w3K/yPnlKWwn/cj7GUnL8ianoN7EdgbNSzsObZsngDj8pIvxeIJoMIR7yptGTKdLCHwQD
7p+DsfHXxJ0a9NDQJWR77oO5odAtcgqRycdLTUOdEBUh2sUhFImNQPXhP91GNVXm98z+yCR0Yj2l
6n663wnSos8uTynJD6U/af/LMkwV3So/RdP5RQvBuVFBAtu2e1Vq0f8/Nn8MEejQn3evZV79lfrJ
fK6udlni4oMmOXUPbdK98cOVo358MvoIwtlWxcYgZB2KTix4YFnKaUHxWrOhOka0bR8HkxLNEqGA
GHO7H49PP2csHy4Qsrc056I+WVnFmOCJuZp5coZ6ZEHEEZBcsN0h+kDEYKBxlx+SLcho4S6l7rgM
FVBgbSGGINFJblit35MgL3IAHZHgjueI8CvR+WcZ+dqKC/Y+hHFwPtK15ks8PDGsBJAgeZoz7ncM
RwO1rQwVWfrUim3laLc3ClUBEbpZVFAXECkLZT/pNSa2YS70Fyi29MoWbQDN7KmTqcXbbpF44l5k
53+CYtwT/p+HmIt6VACtE4xSEa9Ig0Wab/kQ2nTULJ+6IsEhMGfsFfb/xzGmhLcPLPReiR84PA8f
fhpo0vQH1ibr0NHJxVdvKKKhyeQfA4P3FcWOejA1qdSDiAgDlmOv7O6riOmzkV2PKc2FDjvYAZx7
jagsbeUWQ/fAFp5z5VXanwNdtMa2RKEArcrs5enMkMc3AHv+cYIWAYoRcgLv13Fc2n/FQnsJ4J/h
g/rm2Rpy+pW0dYRk7Oa1aVhdy7tHzaH5rvuiPGmz+45ZjQBj6dyGL7kRZs6rbdVRiTCORMBQWgQA
ynbTM7Hl9/EROwF49c25iCvA/tIoV5psdsCcJnIetQo9YITWQGHS4weq7pqWcZIMUQI001WgsHYB
/wWw1+Y7mWcWYfpuYRbHAz58gHbO6TDtHgw9+d7QOqiTLqiElYP6sHdB9EaHVJplhpHr89PyV9Ay
WqxT9xwE5aJBF0ouIpy0d1xGk5ZdBK8u8Um8IbvCoJCcNumWoUkuUhFak4vhYCf7Fqm26qDVXKPY
3ZHmt8fnGZx6LTgkHIve+3ROY4ewEPBAEmIVVcKcbwuIMpGZKImhb4AaT5STKiMoxsXE8PQxzxWi
0jNj/cApFZGKajdplQms2BYHGXqufsZm0IdXlIsQRpKw9KALz7gbNdfMwCDCBdCKy/y2Kisni2Wk
2AX3jRJNg34ml7NExG61NnTJ2x2fgAELqo/1Mti+4yf3u/yf+v9YBh9/oxephAR28v830pr7eAKs
82stCtCtoduah0q2pXrH4Sov1588/bY4qsz7WNjcjAtQnP4hyoavwEkn0+QFbbYzw8gcgHbtEO/Q
udYtVYtTm7eIaYizNUgZbFE0OjcEoF/cnejTcvpj3hocivpjR3ZMtnysSto8daW8EBXpcqISL0X1
Q0YL8Bfu28GjURLtvThg07zVVtbmy6iB+y6m7G6D28PzacUh2SC73sayzBH9duMjhv/iuug84R53
UZ/w+1exhAP0RIp17EertpRHE+l9gPPOZSiy2MfsnwXYJHy2n8GWn8fJPZ7MS/L7J2bTei6X9KSW
zlJUl0W8OIEGagw7MLdjBSUbyR5dQJzuDcX9s41rR/uL+j422DjRoBYLP/74Y4NSPTNY3H39UpXu
f7RhbQCnsqak7YXfD+wJtOGbbUynen5BC9iGfmw7PbP8CAGvDp9rL34L9tifU1NQfa4TgbXGh9YT
DsVYeP/5pexmQQgj7I5KyBI/egUPFIDwgAYojrcjH59c1ew6Mxhilg5LjHYKzuY6HM6T9toFEze5
i2FvtjvXURWTYIRChJBFuzqrlIYIfXMU4oLSNvj06VBpqeoe1ZQ7cinjGniDww0opzPlpwKMsD+d
cp8LxvkWarLpVODsAS6EhGuo3XDOBkyyGOUOKyklcSdRE2elwv4w5mYCvvqcBC/D1nqWN53k9YSH
YZeksnQIwYwcIyJIPmUx52j/7hQylCMkjDzKIiNZT7gxbS979OSANFl5cGdGoMOwGsDvezQ9zXeI
77jJNpz6bWne8Up5SjuYc0oZTtG80vekisAn9OJvbGDPNrAQrG+PZKeObEsh8u1j60y+oUUtpiPr
T1qDe5xponNGkivYxEPvCmU+yg2q3B2KkE9h87L547xZPKV93kMvEIsPEhWqaGV1yC6mjpFtgtt6
b1iVhtiLYRsU8weQSpBuHa+cuF0g8Smb2OG8xs1ta35z9XszveKPvkP0IsY22hifu3C+sMkNU+R4
n1kQIHtH4ZqnV7J6fdJnwbd1Q+OdHnAjTd7pahVOhBj9K+oNY941FKlYdyl2ieUFQVEx/Ylfy/lF
pM2JIiK/NeI09pZBGKJByxpwtTczbXKFtf974hBVx/R1ED7s4JHdzdaGePfHEvmklSD+sMQcjIIb
20rq+5mgc2euyDpcPSn1TaT6TsKZpzWi2OXRzCpS5S1VOMA7ExH6XgZCl7+qhAysbZEesPYkq/ko
X5NYZK0MISAAUEtCPZeVa9rAPnGnyOzk63t50+isrbxGui4UiPADLmRCjz1iDDT3V1beNxIMuZab
pxJE+dsgCmzVd89inks4J2yIXoGxmhkodtgPgcEY58skSY5YcfKCna3Si4i7bsGoF1PARUyfI1ov
YYfVBEcWxGax1IiFD9CCquHgLBXRkvlqu4lksGKfP/Uc9FvvCxbwHze2Ng1lxx0/j5kQuM2mUVRP
sNiT2xzeOB19OrA+n5zJd42n+wxEOK8NhFuCtnxjXLv5szEwZ7BeVvXHb6hxckhNLVrZk0+o6Ry/
amV150vhLs1Zu3ugdi+wC1CYjIw01r9ECzjAFz4n78J1cvknnA6d8nINIz2TPGCSAteNEpAlX6vB
xmLEzHyNBgyyWJG/yXAB7f+a1yDaRoL8PlJ2HZwHDg4hQKzy7OJ5VUGgm+TJ84BJyinTMoAGiNxX
gwz1yBUAbLcs24t7VFAUzj5xScAq0/iWqAibmAQNF/arN5XTt++iSLdDzl6cMRkxkbJRXB2M1KqL
TvTuFHWBdVm3L/VJBQcrT1TzhxolqdTWfocZfruZx93xbjvw2MGetJNLOAGDtOT0yxJhRIAr9N4r
eMpKEZh/qqLcXfoilfds5NW48dgv+zs3FEzhVdrIvE5eOb7O1/73CSYBzLRQwWGQ8fWtxtOvEKqC
A9XvdkwJeCCqxbIeswhfzmzzIcEUrwY3M5eiwG2aFVhbJ3dNB3sEbxdd+natEqpLxXGmImzTVwOH
GmqdQFnStnJH41X1kW7Bq5jbhHaV3iSgGS5A8rb9P5yi4/qST7Yg+4UVyGmPRp0WYR7Erb5xcARH
urXCJYuvJZfLIxNHNj0K+OW3jXBfhrb35QHY0f+ueDV04XG6OYkqaO/IrdNMcNj+0TAKCOhDuNKs
ZEIfUf7fDH4ZMEzWNal/qrTjn5yp+xaqD8Y3+Qxoo7lROz5zlzv7QT29jV1TwY3m17jKLkoffgXM
cljn0C+JVZqGcgczizNwWYqe846euKLknM454TQsJOkQkmrw1pJZJYrrS/w7OhkySCyu1OIQ+yEB
cgEyVLDxFU3/JxQwCc4I4HIqX6MDCMon43ZoiLW34H7urLe0gP6gxi2MCPbzNNUHdDrrXrE/uoF6
ZzWlHckuffWPF+RFRLp0RxaJR5Xw7aEUnpALg8aBBBMOWbekwWboyCviwvNMZlBYxdYrvhLm4Wdj
4SOBCCo/BgGFn6C/Y1lpsB32hT1RAPwEh8sG7NeFizn5AeeO6930aXeh4qPmBWUwp5fHhhIPB22+
1oHpd1JYXqg+VyMjUKjKzMDffiym7heMyUUYoed3Ig7340eERLtpv9BugOAPOvvW6BD6iFRtx4E7
i6PGbbVKq02Q9/Mgmu8k8mOxARkm39O0o/QEaeQbzoJfOpLyblMvROp5QsCTxaOmuFWPVqKnZDKY
8idoCgng5vAuDqaYiijtJ0FTdbgiWZYitA1jSJD6/EhEdU2R2AAsoatdC6+s7PqM5ZFovvJAoFW9
98YFeV1puLBmU1+JQHYP45arB22uE5ukhrSeQL2PmsZaiB/mmX3qiE2sDi7utvVBX6T10PtFaOT2
fJPuwWMsxIcGFdMx/SqJnymFwwddyx5ZKp+NNqw9WbYAHXfr72cIdM+9fk2Lj6ctEqkQJTyb+J0H
fge4XA1NPYAMt9rJvKiqF0nmJn4aEQ7zjDkteFDqPFbieizQU4LZ9ADD7b7DXaUQRq8p+4/Rkm7W
pR+Px9ophzqyXUHphDbn77Ioqd6h9cDaq5qFt2+l7sWKc4V5eqTJzraaxAmwOxxg/JUgh7CMWUD9
SEN9TJCKWyw+ueql3Slfggk/RarYa/QTjkKU+Wbw5d3peIegSWCjCjTyYQkP4OEfzJKGEOgRKsku
ZJd87ETVVa/6naEXzSnSjDxhzb8OC5fCRbtvHCX1qsiYtQos1m61DJXaspBbl1y84ReyTS8POhNM
S/o8hfgsdE0wCDlmdKG1Rx9eVVJl9OOPstte57dVmeHKoXGMuJhFjYznMU5MO0SGxl23+Wmmswxv
X8cGR0qCCIjQ7vLUjD16dRvuzxeyX0juAE0Q/uW9ewFxrmVA/Hx0Af4X7JtLfJZvsMWydxvu8SFk
2npLiw5PTaHF4LYG2o/4cZMd34YWMmj+LEQoSHj92Mr7Tf/XWVUVKVzg1HYhwxzG4eKnZ5YezpHw
j5JGPPZ7Xv+FN6DbKghmbS7gFQIKIE0ntrB6IYtSl7ybd7DsG9KfmZQMKMYGGpAJFW0cBQwH2EIj
W/wNfVfcw/v3MQx0FYsID/uWGrSBzfaAoK0fBHP1G5y7Lm32WuAi/HGGvPfIcOwWb9geHL25qtqW
4egfI9aWzFBclMRhAWWxGTwBOlq886NaZ3yhw2NkKrF1J2d13Va+C8s3Q1IBy8C33LdnyjLGjIyW
9I44VAv+D8qKtFVOnRkT8Eh6NJWs49n5t8/ICqj633v6QBaGmr2fK175cxbm8vPw14x77MvCg5kK
roRft9grT44hACcVE0cJTDs+5rcY9XNKqz02mGhBhHfV4agYHTI185FdoQPsNy9qyQ4kHUjPgRkS
lcFB6EquRVN5S9NvrPjAUykfZgT+6EC8hrbabaLqea60NFuuUMXRQuwopI0N6oO50t2kq/xdkL84
c6YOTI5pUgkPWQNq4Ag3d1rgDn264JcKJCeasmdjzX/NyXvIqStcJEdjXAb9VsQobt2hv5k0EPMb
cag7OasKbNyAj6S9JU186JBTyLFj9/b8O/QIcu5dCQ/AuKHBwF02Hp1S8cp7vVVauX2DmWguWor1
qkQ7BkPRD7E0428pGb+jQ0z09O9YDgPheogsQFjw+FBOOFemhFltUspUK8egAXXSczQ0PAZdabpK
SeX3+IT7InBhTf4kBfcSS7ei5agxnSiOw9VNu45f6mDTZJ12wVMNcpHA3XuPXkshBrjojtdg2/7W
pR0f66JF6t7JeHQXQihTqlNQO+qW4BeiKjKnuI0ePm+1ewxEX0wHor6SAxEvHY9X6KEezagXRpub
zB42VnstWNT3RTaAQfqx8ud+3/PKrsPYT8PiqowvvMlHTrnDwrvwwamjupXhtPtQm8Xky9ki4A5P
x5CGTz5Kf/FvkGN60q6H/Pu8gL+ItTVD3fy5vxScGgw5wzjEB8JmtDrvxv4pzbNYp9zxOw2pCqbz
PKPJkAPFxgFCGV+WiJRP6F69xLk3GhI4SHEHNj+bEeRvoI+AL2FCRWG4rfyMvPb9xySWrE6mVRSy
zOU0VR/2VvrTLgc/AR1x7TTajcrpyoq7tJEGJthc8aYFVAXuJkTq+nDuHI09IWWlWx3BPl7IHjGP
6h7nQY0bcdwcZblO/tim+4U5RzWs5DywrAzR2nxn4UFuZTv95ZTPq/RmaKPVy3FcamQCbrzs7cbP
upcH9Mi9elBzqFaEg7Qr3MTzgcDSjtKwCl6abc1Jao1T/0ytbSL/mAhTKu43m7LLyRBnsisQouuk
9dQXpcU8jRgrijxrobGCzcF5x30Yem0HL0phEgxAmEV4/iVZFYSBIzO6fZDEZ58D4zFWjLqc+2uC
FBrL9Oi5k1C1KokyWCIq0pxOflaTY0nL1chjKsdvv63W4IlWzp5QD6WAvShEQyJvdggHhYzFc7Vc
I5zX1zMGq/wRTAF1FmFtrjIaMpvia391943kWWkMI04fOxTOf4EzzypmLjhNRifrFXz8P5mwQpfi
M51l9sYfu+VHstTo36ZQjjaLvsTV/sucU2HqHEM43NupjcZ2XnZJtHsUhW4ROpzlQxwelkFBr0Fx
X1Gw5X/azO8OPTYYbejG7PoDPW6iK5h3HbzbGOyQnEIn3akAz6ZcnCuwPQ7OW/v97YViYMAaWoV5
dEIB4j48RHrsNl2iqWd1TCxiRhk5N5Y6r+Ym+J8XtQbe61Wsrnlhvn87dWy3tbLWEPUzPpTiwbvF
jp9BsCz79K7+W+bPhdjzcgu5RoCLP632NunL5obT1f12NPTa1YjrlACT1fHL77XqVj1LkeNz/eq6
PLLHdpkz+BFyogQb1KqeqY7Frq27wVWeIQTiqxnH/jFR02E4/5kOrxQU4Ndl3R2k/amjh/5TQVbA
12O+CH2aip5bs7nfzhWOF45EX/jcJNgA4haDm+aO0+Cndz57LjZzCzutp6UF0cRAMIvWSrLPOx6/
g6eLHtv6jLOD990B2YzDhgOyenQI/ASdLZg3yOEKSM2URATyY8BhYG2CBSkEghlC56iVUjCSjC2X
MKleP9ye62JEMGMoMKbbqg8giNtwDQ3xFDB33KGPCSraK+bvZaxS5SSJF7Rhvw1I2VFQNWhfX9Lu
9XzJyMMC9nm7cUPo+jYoZocMzRzPSU3xbIrEXP+p8oL2Wkqxo+2VSc1q/7FgAnuMG4S/cpRPNDdx
CiebFh5CSDa3mw0W3SGekq7yAwQLGjRRBsnM3g6OK75hCNteQxLFb2gdmt7WdMy2U59EgF0upaTO
cDCGqCY0JrXugzLLj8JqSDD5KHfWnh5N392zw6nmCryNLntSc1y5RwsrKQfsTnl1U0Xs7zVhKauq
Aw2CagIWf5NaKuHnBtlagBDCawqwLs9FYzcR06hp6Hbz5dvaeqZplm25gJgmkoVdGNywRe9pnsJJ
W85avL2wpajQn0bq//UyiNM2Bhha3BO1e5Y5vPNypIRtqTRSBuEVuyzMpx2ARncZ3z0EP2kWzGUV
R0nJzQYvEVRqcFFpe5G52oJjjbnm6ThtjR+Dfq8EXFAsLfWuVTdNL0YF9TrU2fMlKM8GY0e28bqg
mUJjeG6QJZDaz4TVCFJscK1vIRpOpyAnJCEkM0bgy1CKszXGvqlCGTylQvpvtpcAnb3DC9ueKZNH
Q9AFSk7ZGVBzyPuR0R4JpDgdoLa3dgapAtxEDb8lMoIaOvzoOOtKSJ/f2OWmAcREpAA2hvCpsEsS
E2Smy5Tmopx7g0p9mgxYfJh9sw2tUk+25pC6OMv5rbD7eLGUPyKG7Tde8+AtnGD1Xl2N/IHRV01C
CVqgDAsDs8IeSAUznsShG0Af0ueMZTFgsSMvMCnlebn2ylBqJ5vLK4VrC3m7S35S+J7lp+Qjmx+H
EF0SIdu2do1OEHzQLZVO6gKUTF/SAUHqrSkDorFpxuxj81nrkByMdg1kwuSoSRU7nS2FC5M0a7hj
HhXOZdqyAPrGHlcuZbj2rNAEFtC78ArzXTt7Q6SDeLME4ZH7b8HLJJ48nexJFyZZLZYkQRvZmGMB
5yCClmJU+zag/x3sZzrrkIuRwbHk3Fb3UXQcAuS4h1s/o/3z2lA0/uhcqUXtheSBCrCUsMpc6hwj
o4gUB/ObfbSBlf7Ca4iRs9mR763kDaTBV9zHjzORD8D290OKxxpsDmy0i9fi+OBwBF9Ie6/fYBki
DxQsbjwFEgBmMkGXhjxqePbFQyoszfXKJ/qon6rZ+oCo0+Go2s7hrfApvpWvLYIdYlYkklE3Y5sN
53lqueY8DIpoeZff/XzcaY4Pf4fSskDx7oeEI6jaCJuBaqNAWEpLK5gmuf6/NHvHAGtQZ5aZQtk5
EUKov57J6dsKiSqOP1vD7pOc4c4AQYDhGKwnYE4Ggbrf0mOx+ZCsrgaFt/jyNcTA+dc8q12NzBGN
fQbrenNyq4jRF5iTvLacR/nsKMjhtcQRkJaKFxBpCSS/RyYhjv1xhlgzoFzmJvqOk6x/KO05btLB
qWPN37y5tJm349DHlluEvuQ/6woBUIZvY7zu+vnO3qv7YXDulaMvfxYhczUop75jRtHC7AVXQK5m
fyJ1FhHEnTUypbFvRN/T2zfONSHjYRf8usvbgEzokl/muD/4HsvaIuJjj9ZNgSvGLp2mZDLGaP27
3DAtaGZkqkoOXB5ZVild8OlAnhrrLXKzRqzRpzbphkd2UIc/AJGunP217mE6Y4KjEe70kodkYG8K
31CPLlhscaU4ggAqOoaIY2XSzXxd8H1vS69u0UOHccohVbN0Qar7XwvJgyPC8zLVpNGSmuzWiGCA
ihJsI1SYwaF5Uv3/TiWthNDUmzj+9Hfrx1FZpDNhfjyUTRm0ZMTIf7KEfMpSboWNzMgH55vszQJo
nFDyXZWFuHQXvzpYQHfF6J4auuxw1CZWZz9S9rAow2W+cM17O60qjVXwzOCFzMZ4r+qEvOEHnAOi
nI0d+OCB3lUJMUYhId3UCcOOpSdK6lm1CWPIAgn09zsrlhCVLrhFZz3nP75ry4pOx993Wu3JxQVG
XE5EWunmjE3JKbnLOHqLWZgwvcFz6BGjhHJTxxypXqO/OshH4g+LFl7KA8T7rNUhrI6B1D3sEoKx
ine0mYEkZ8IoRJmQs9RrbXCXl7/Nx2wxCI9+4V2yYkYa68iSVjxCGNsRgA1JHID8Kl7nAb90Ae7H
u+W1llp5llAjM1T3Cv3OE1Doaj/5r9ViaiP69xz99224et41xh9LHc/yYE22TD847ZxYiw2VUzfG
+pJt5LBPPzx4UzGry9HPxJmowTUXzlApjINQ7UT5A6oNMjvHN1Eow9hPjTqxgJKd3Xp1rm5B+iHo
sJGj2Hvje8tGpujuQnVvgwCW6DlBTRIAfM/3gceb3Vvm2FyQ14EW1X5/QrfcvS7tFz78ll77vDMY
he2pRcOnZ9w1qmew7f+4pIT/Wmu/eU73Py4qNL1tpQ5VkHNsIq2eR2Fj+F879HyQVPKgGxibpQfH
fHjm6Whrnv4Eeki18mdqupfE8CiNW0dP9tXZDEaKtCY6TqFEIVt0zhEGH9N98AK5VhMkx6WTDQ37
jYA2xmH56B/X7OUU0OQeX8w9ydEUzLJZBnn7tswXJU5a+LwDWZPvwz24/qLhkWUTAFTZTYjFtPXs
SA8Cvq8CvlVwqRvJ9iHv1SWWJmJwyCRdf92Tq4pJOGvpIww+bEOxGzd2TDLDpDVWaY0c7MJ9nzQd
FRF6jiO6B5Gq7Nb/mxdzNUj2xFGrgSBQNFRr9aP60uViGwSeRmCHqVDHUSWcLcDMROFuZlEA0bEd
J/W/Oe4yNLQySj+yETuUf97MD/47xboMzPzXLXQw3zIjcSHq3sMzSfus52/6agWu1Nt7or4LUCFb
ZVOTZc7Y0bCOJtS08gBtL9uIvu0zN87RNGuFvyVhdYRhHT98nBxv0mCPBXPzNMgkFQZg6dwY/fL0
VornNITGJ+HS/PkTA2wPDj+DgCVk4shpgiRR3Tr1iTZikihpKWg8tU3sq8koAyXW+XWwf1v0R6UZ
SeCAid4JUMk7yznCdXt1k8Tbz9xaPMIe1aFAUZA6QWD/C51e9GnFkp/J7cUhbiGk2Cu+25IOfyCJ
UvGLXYBVDdYrrJBTCN5ITs85A11xF6ZJ+aH6HrW9gaY0fIENUnqLdL4jMrK3sIQmWwQUXMtOrxJU
Bf2u+S733C9n/DhKrhsfYkXKaDh1E2c5qLx3ot56kj5DEcAqsrAUuc9n6f7jvQYuE/JRmsTY/d8Y
/+MmKpeavS7YpSDjaL/unbLvUZjF/cZZKUWda60u6c8j35CrrWb4C0bxcynWq6DhbxV23DpM3eJt
y00J9aPc/vtn3qpw/2N6KrpU6SVhVxXKQVA6/BpRdapMtWSF4bnQPQBZ8ESOpYTOYe/xxrtMHax4
m7WPO1VbFRUofNtbk/np3Zzt/mmhQrXaIuVs5OKZvifmc1n9XOIVQ2RJdo3ug4CLN9mydIxYZIw8
nY+2hroIgRUFcuTH5P8Ed9YCj0uqolindRtUV1AGw+Bkb4at8vO2TZwilZFxLUQO8aTsp8bk57vP
+6eLa4GIBH3TT8FTzW+9s+mgC/tmeoBVj07uQdt7bql779B737SwF4vrFsn27oK9B0Vn2PJZBj0W
JlBD860bsGv87WUgVZsljYu2TZ4lHN/elxtzJSWdFp5K9nad/Dib/gXgXEFVyLUq79f2T6+yzfLI
HpwIBvc4vkR7AH7Zc0qyaAWpDyME+dWADHHmCNN5qZ5ZU9PZwSumKE4uneI5pqtHk0WJzxPx7iqp
zxm+Z7DNG2f2vUZJrR75OyZ0dK5g3EgtJO1xh+F7nkHHJULfsQ4wWkajSgvi8fMLwhIr4tt/xlQe
ZZBaKora3PRgmcQFhJeHV1KquZXqPc5gUGwien9P+L1oRuQQyqlTuNLePDTtgYcWCtyNrOKJXNtI
B5mlzapZ59M4b7OgNlltiy4GhwLXlOLX2MCrEqYYkzoZtQ5sHke8W9Qvd9GyQKADulaSi98/fiMT
XSnZJ/ZxwtVuBctTTQ8DWN9GDRtNuAN8dFXIVp7kCrMBNiwDUBNOD9mCRTWq2BYHEGHFqhIARwRv
UiZzrmZMDcFOPKof9e+HmYfwtaiAtX18E3b7Y5iEP3h0UvIB93RAdWLHA4HF2MTsyJ4QxIWNKCHa
J4uw4xxzkpMH4CLPlBfK9ol+hJppNMsKiNEefPReNZ5i6oa4tRcGsJoz+kS18Dfa0WfGBk3Fbkjs
vB2CNY7IS9o9+j/nZrrfuq389CggNYhpb9YSYWtl+hKGwKneEw6YrrkobTwhiD060nkvVxNP/wIO
QgQdLFIuXYwG//LwvHEU0Me+pMgOZRUslC9NT8M2MQm6lHdMgq4jlkZzcbXU6JtULcg4L3qNe7xf
k5cX3ofbdOYYwW4L+i3UlF0Hf4mDE59rLC40C0w0MFl8olm+LVtM4q1UBOeXYYZ5X6tkOKRNKzDU
/85wq4aKytfYesyTpivQm8rkJO3bvNGeNjGmjnb5kCFPAIvKVOaey/yOXzb7gpnhCF9ifDDyaAIH
9XRqx1eMVWHYzKbe4Mr2wcJrlT26fTXJJ5Iho29n70/xSTWOyyoXQjY5t6YZLqyLykIynhkLjluI
YJPO8wtKxQLgmDVFefvaI0s3fBeANaNvMitGXLAYPW1dMfUUdpPJq83KIHxEld6tfuSOfsBOyXe0
6mhqovoxxZioHqvyMSO83zerHFueDLiNnsk9t234OHHp4GLzygP7CBpRiFZbVXsPE4XIVKDCl+Xp
3jf9kZKTbCcPjVubkp4GrUK4kanyPIQ+nYSakqc95wnxoCNsF653aO+ACn9GNF/eIhU3PPXJWypx
SOoES5vb/q86/J4a1pt+Io4OqgAcEP0Y9iHSkpFXGS7AISo2KNGFb0k5J7vS6SMacT/nPpryfxSb
6ohqOMLA3CZM18cv4PSGN2AlAqqi0CnR/Se0l99yINb/6yzkm6THpabrS6MMXbE4T5wRRpf6DHR2
wwrPdARA7JjYXs800KeogbTbnUnfeZt8uk8X/lwFR6juGWBKtWwJujcu9+jcNpMPKgYPA7cvqdea
pU6osLGIe2QzJ0I7GGy15e1CFi49nXeFz3zls500HyhagYJJiI4iKSM9ZC3i0SgjobhYwQWcxX3w
vgFi5HuWl/aJ68HtlD9eWtWR4ZmG/nd9c9niiDV8tvVIGSYHD6c504a7LWYLKhaj5iHiFwSJvDv/
ge+2FM9DaJbH0R9eHCmYTsQXLOfu1uPEtY6d7R2Ye8pK3Im6lMa1fQ5LXNPELWzt1f7LI/epm5/Z
idG9bOnRfbH4vnXt8sUwIfNIXXJWU+R5D5eP91nfhg7oYdfHBlCV4MFOmwYXMK9hWvp88siSl+y0
WFEE0U8u7XUl86HZqHpFODm+RRP49I6qjWRfFOKQhcyfbnszJR9rCnsb/mr1LEjtyszX4CMuYyQM
M79P5q/0CrG+qZ0ApgtFsU3IzuydBu/hmVXiQCtlpGNSamGdAW1xcTwWcVNXSH+p23t6YU+fAijZ
7jgK8CoArhuy3Oymz8oJO/FxwsXyexiVbGl0KTBOAAYDMcKWX41crlA54hNyDqGIT6qE6O/qe0oQ
KCCBvvRcp5HBDTM3QYgm2imYqvNixK2DaV7aJYyCebxzHgQYacjYcpGBgLIZBIhO+QXsvtx3DK+8
rljitSFywlr8ry44Wz526AtJ5FfEpZCfPb9+z1urxA4PjDHpbl78Vz+pb5VYRRLk+p8ipVcyIqZR
7q2HQ7iej9RwDmf/ntEw7VsxQ652ho+HaMB0jje0FUxS0afzuxwMPYTxTjr+3lXjr3ZsF/o9Nr52
0tgyhqRqU7cJ5T4q2jjKSIEWAy/YVJE5pW6WCpLj0bxk2nGyjk0ewIL5bCwrRnvqFMqoD2gQCipl
ayChkLISwJRrkHAcqic6q5D3DS6TkZypkmTcWLZ592eC9dhswLAXFQXxhn95BYN9Gc9qv/H/adRH
dEbgVKOjRoKMmSvVgWJxh0lvDYUvpEB5kplhYru4O/6yUmtIImhPMUECoTZ80phe69/Xt8kNyG1m
0RrgOOwI93ZdvAybJB6kXg3pItMBS1V6WxR08iUGacLnbX+fXK6pJ/GYRE0SABJNgCcrMDBKGOJW
kZk6SJ24vHHQt3egrXad15oLq+yaNjb3LTiZ6ESC0kPYQe/nyMF4x8htdrGII/kI22PeHE1SziXL
bFkQnZSdVGfV7Hq3hEx9OG8pcAqVbllrPQZq3zFyneiBf6A0H1lbUCL+Xidu6D6SgxSTcXvTnHUA
6x3KP08X6UEm7dPG/JR3e5KzKqvJp0RHn3127+GnHjtayEbfrn107avZs6P2+nfi56S+6d3ZFD9w
93aOdpaCUP1oZr6KRdjnAr+OUlpSd9OrcU+xfBAiV+pO9hTSvSYClon5bK3UPLv2MGvt8RtI9CGQ
hGbuY5Zw0uPYJpiSAjfvbmAElTBdXikPBX29Etu35CqO7Wmh0c/hQiSySo+hMOfgQ8hdayaIGFMS
znQZSquCznNZ3iVIUdIpqpXNlE7zmdFPA/oQJWFGw7Xmn9XkOVh41Kyj4gvQuyceAErWa1KFfJLE
vkR1UzUJP2CSf3kImerUuUAj7umDBf4InnkgZskuxl9m3hZTkkLirgMqf3lW6e7TWHeiQXauuqGM
x/15oKLpg7F2kEsbssGffW6QCaDydLwUxUym15yEZjVcA0EZkNlXWlcKHGpZNCrCKj5qwW5FkP9m
daHuJC2Yt28aXhNFsamiASpL0UuRTg14UVLGtHqIa/AXLcxck4PveOSyoZwD/sMJB0FF1tmzzdzz
vgdK8dIguERLQNyqD+8aqRIyXCEfRyAnGL8tjIxLz6WO2EY65wD0SH5dvubRuweeUdQ1AF7yxPF0
RrL81Whb40XrlzundiEFbkUZ4CCbBa3UfFSPDCZRpAjULpZDPa21iaQfoR/cXNrY2s+cdiokK49e
yUmQA/ABVUjD1zib93BqdRrMU68Mf66mvqtqpvm2OcRNkX0uwWrfv/aOkk91SduNCbhm6EqXbYQd
jFLztHMR3pI1ME6yyxILvHWiCxMSoXCuz++RAvFlqcbBn/br9x15+lt3n2EcIxy9e1JDttiF80pI
sMk2XoLAJlX2IG09xJhgYWqv1jfqYv337QDV7ldo0PbrRbuh2w9OSeKfLRRzMD3EoQ00oSFueWhu
6dyCCNkZ2Bdbc+B0xvQaoMtV+Yvu3QH/8IgwveIaIH8oCZLd29x9Zx7vHOzez5kOvgqsyAWbqwWC
uYS4XCo0CoJ2SEvXYHEvmQ1ae5NZdDwrZcRz1oIHyV5CqzFJ8QV9M6Kt8hSq9uQAWPc2iZNHISYY
8J6aUQC4WOOeFBbAYg/xIOTbzjRWO9UdBQTNrd8rcJXDzBI5Fd+tBvfQGjBxSOAglm0RsHlXvIeu
KxArm1oQMp4myG1ph9Xia8sCAB/Ck6SwDLU3Eg+ylMixDxLqbfFHylPsSw8luA02GvPNueCSs0Ik
TL2TWAQYpfTBVnCiFO1OAp3TGieR9InkZ3sTvnvYQ0OM4S5gFfJKgkNWRLAK+/7foW4lRs7TUG03
HkDw4erss6N5PT/AN7ulQ8LBgn4cIV2XCKJF9xCeR1jwea5HkIM6Ui235d0dLEc4OFDR7R5RaMl7
Um4pZ+ivCN4sKuu0/KoIWmuZCkg9DXB1g6Jeg5cuRVWbkl/gC3mqr0bUvUJxwUT/Ods0QCwu7fnl
8U5MituLmzXZ/V5m4XqoupC1eur2XKmIQuY7gjuTCEbbwnSiO55MvDfqcKeO9jyJECYCK//mbY19
S20WL2WWHfYMBVyZfw9PHSsg1BV4Ths5AWnFAFCHa3tskrx0hDWgNNhT6ab9UCvdBKkI8jAy7mSG
iNANo52AQVad7SiDnSaKoboM6fXNEef5ByoTkYQgn3u+CDGjevCJlI0bUsGO5t2/aOoQo1+xpoaX
DRfbk3OAVUTx98sqGFsZd1TlP9mNCFhVmzC/pg19LcPBOm2l0VXN0GN7M0r0djAcaOVc84wAZThW
WOyDKlup2W44skLbFQqYbhFyG7dMGy7+mDn9E9F5wS4zTKqqAovyGUiQL177e7nX7qS2cE/B6x7m
W8YvN/imAclG15AJuZcJ8W3LVAnr0ucAzAZ26hx3J4FPtLuMulOcyiuv1P9UeZJ3LThDAmCp2a8T
lzFL0yIPFQcC8JCFzKsRWOushrwVWlMn1aCIVJoKwQqDtMPSyuGe7QVzfdeCIu7jexqMmf6YYoeu
uktvnzXzuSNA/BNKt4Eey6VLDnnYPOxxhbb7AiWlW+xov40w3+Lx42UdAxBw3iGvMJEowOqQIn1m
AeOS+uPVeEubVJ0RXwO8p5nhpFF79hrHZRgfz25ZMrr8/pt848423DqlVlnu4RhZ2NyC+4v9jMGi
6dzfIMDB4BU1IiYSuVcIkPca9Iqr5vaNuheV4UCeYSTlJz/Vx+ApvCcBW3H0iZpL6ESW8qFRJ8q6
AZ5WbR6LW5zFTFvWn8nr2AxaALpO5y6svdLhxRBQ7rfXtPG5sdLodQqb3JGKUoxMzNvuuKrSgwNX
MvajTMSdRuh29sEdZ5NgtNcYE5i83M5EVtH24kNiBFSa11skLXh2acDXaPNa93nlrABwyBon6L1G
flt7oJo5+1HnnIC7LLncYMZAJz84RQn839EFdDLu3Fp9ODYogAuyes7Yw30zv6DE7UPxO36XeD2w
miuggqYCl3AN3RkJ6NN0RC86dOWg9X1Qt6VpupfdZ/uGnFSXUP22j8RME0B5nFiw2naTnxMhFaML
L2zz3buQzFoR3tJRy2TBjBCx+hez7xQTGAjqfyJua6chkzR1U/GP+gdgYxiTzWsHkSUxsPEQaxmf
IO6y+UqSnyewb1hGFvZjs1fkiJn9t/8Z41o7OgaFwZFsDj3sV+pmYuyyGD77WWyFQlQSOeXXxlsL
VSMJYQVu3/OvT5EZL23JOjEnNoK8TNaEJbEGuUz4OzXjhRX2aAmrkmFsIkE8rYA4m0KoVzVI6jlM
IYgfiQRpdbORAhec+tQkDd/oy9vropwdfJoJs31ma4qRU56QQFi9gFzPhu0+58gZU/8NfdboqrKp
Goiu78EH9F1nmftVeNGlTRblQHHrAumLlrz2LezhFiN99gw8Gj9YrdruM+XNQXbaU12XsE4OB9iR
h/4BsmwjPdAO2clGMu9yAuoNzJhNscWxNS1jjOobqQDmFealRRkJoPLyvJk7VohemglFZ1pEk0Je
OvfFWiIsBue6dqLnahRGV2Z/dRlT1LJku+TbSF6OV+Xf4YIIxfMNa8ZmxHSwDDsNhPtGmX8ZZ3N7
pc5QxeTV+Po4kG0KLz2jI0IlLj49qe8iHGjmlZtlrZ/iaD+/+FiVI2D7wQW9JPxLfVRyQFBYwPIh
Z3rnSvVT4T6EzH3oOQdt5jXk8OaeBxsG1dT3ddjLWmNBBHySLSjNPyoYS83H81/kasv9/0TMvPSB
6WG2w0ZkTZt1CEQpFRQEKQ7HPhRySSIf+EoJElrvnlDVx5hOwMA3tGSoDfiEo2RMw3gJ2pHvwg0Y
rNK2DZEkSRaJQzxugBp//6KRvEr1pz0JBf2HxHAYZ5xBObczGFOTk+eonJvvtDE5hBsfkifrQ2QL
7Gu2SNtGygoO1o119cPJTRuYBzQN4M39RhuBW7zwAtesPphumNskxYuhbX6K68COd+aA0gCtj57M
K0HEzOQcooUW984nYX355Cvp/6kGFFvGw+qyvwvBerE61VfuLdwINIWN+4gqovcDRf1q0donEvnl
wNPhua2yub2l220ByVfBww9YfZIPyJvxdCZFsFUQxuhGujGaD0QWPIJCattWHzPVF2MezFgWTGNl
pK1Rby7M6Cfo1UvUwgiHXgH8vjfBGWypUHMZzKN7rMJ9ZjTIfkhWudQIA1sY1Flwiu8vx7xqhq6H
SC8HlHRoViP1+ScE2oU85/tW+gRSyi4hCjC48nrrmPWjcr18m61feEYL3d4e2VXY0ipfQTNXk9fb
/oWKqwr0Xj26i9eMwNwJeXVDRT1vz5x57qRxdRvvDmKkgJgQvwSeDbAuAl6eWumnZ4Xy+7NToZyK
UiJLN65kf+guk4Gsc5eNRhXN/4SJ2E15PmRx8pqIGVVZos5/LtUhsvTtTiqxwuZ/UZOkOGOPD+Ew
0vPJsiaJN97lOy/T16P6mRvwDAA4YzHuGU//ADRVjXjd0xIZAxmILuMY5/FheqaBG4oaI1Q5gFyL
2IWjWYLduuXqHLgTUcrSeFZllnoak8B61K8b/hMtIvYqI9nhHk3l+OJSU3lYLDjwOG0R9b1BKq3h
90UmvAeG/wGC3OwSuAffJrN4wk8yfK5S7PMHviztQ+pxhkzLNo3Jat2pgl+BthDtSG+i9dcPByZS
fnl9vLd5IpY23t+wkB+VjdyTvsjPuPyfaUozPxoLWyE1SB6IR78WG8TFKMhh2af2CVAZ5R4xuKkn
19tCnDUzsE076pM+SD/GziUT/G/f5ztJwJQ4sVm8grzVQydbClkVYl0fh6k9/egb8uPPPXlCXAd2
gHf3a0PktKHrJ9j3qN98s0DRefeNBy7AGYFY2CrxUXMGCzQFdE8HmY1u89d+yN4zrPEsfd+jHjLy
adrlCUTIv2/qJbhLkz/11YCvzvyaMH9e+O1Ap4wzJhwGUanR8w/fJuIWgM+1EBrCoUyqf+6xaz0+
zBanLDM4Np2Z+Qn84aBYmTaBxFtWrgsxQGTJoz4+AF8P1q/jeN96pZlZQ6bPxTrC3whL9AqHdF6c
XZrAFlro5TAPvnyGBNDv/XNlibclT1+V5Z05vJ1uwpOuwpJ2S25HCSWA5OdNDb3iRm780BCMPg8q
z+wbjOkK0bgiqRH9yieR0WN3cOOCezliuckFXAjrkW1K/f1aCr3mtk/qBAvxAH++nHdwkAgV6ROf
WEnSldKGsWY9lIiLezPIuf2dYQ9eAq151Q3C5ejSo1q854IdMiTyEOaA+i30g9huWSyZrQ4eoXfM
FOaIiL1ZOrSqp9EpKNNlNLtmcCIgX2Dwfx3Fz2EJ2UorFwZsLY311AvDgaeRSJDfGXpCE2IHpZzB
8jhC6eR1rJ2juLzTZXVyQa3YR3d4w4CoyLOirezuuy0yJ2Dt1RpdEB1UMw7PoOZLr3r8/Cvjp/mS
VigjgVPSET9aA/hNCUpSeISObHemCRa2DDxzfDwrOplqdgWo4w1PWeZjeXws7LClshy7Pn4M3OEb
zS1m2InDxz/8u+VlhTe9Ye/KtlP69+HmvsuinvL7zaDwQk3zn4U0ZkW20+JLJ9KkW/9ZxUi6fPWY
EdkdyzzJJRWzb8r6LAx0s2oxGB1H9t4msRLJ4Ge44yg25Zfipn+IZZ1m6Xcb/TWZS8kwEm6wJRYa
G2ZDcOURGJxrnErUcR+y+Ej71JL3EaJ5//T8dt8AH2WkmU9Q64eY0anz7Ee18a1bR4K6MX+zgneo
dQRiFNs/oE20n9Ym1K+9TgD8OJFCJaXd9fTaklvksy7aADSwV+9juHib3Yy8/DFspKEaAPeLMd9E
ncNsq6ljjEcWIr6jBCitK3B7975p6bb+Yo5MQV3JJjaOxrfo6g/jqQWMsKQlCvhKDJoLNEbpXT7K
BlslxEGllspcymxa79hGJ9J/caqkAlDlZxAZW87ph1e7u0JpMzcf5PCISir3v79BFFcxy7HX7H4D
TxADnqssX3uL8SxnFusg4d+OuqcBUXD+IC6JcYtdFoP6/uZAxTnEoip0H0ibUog9lDeDum9NZoP/
F8oQftfCrFlmD0hrMg8AY4UGCVj3T3+QTxYkObVRppB2N7CpO80NTqrQwHU3EcQB+Mhc/LSNxRBh
4PvPFTmacI0taPazXDpLDO/Rnoogxdk2EZHalPTul7XngQdyLW6CGPEFa3O3pr9FlCTTV+2zhAN3
4JL7sjfvpl/G3d6LgTOMjxUipCwI+U5sz8jQp0UsphONnTbICcpDFdOtJOlJP4abKBxc3xCUX9X+
peQDdsV0dva+/oU3CloYMoa+dwugpTM/vNwRXpRUSft3im8PacoRzjdCJRhHr2qWVGyA0EO5lntx
iSmyYGJwZYLUAMNLExWnARnmTcwk3krMo8brW9d0KWO4ev6z1XLOYQm8YETAjLw9p4RnS9LJE6fc
GeHCLAz4Ft/B0WGZwVG/ZQtq3waKBVyGOEwSZQx5m0hhIrTokZTOcUMf4eyF5t0m/CmBfPf7My7c
GNS1fyNsD8n46yR0/zzt06wZqNRG8sLUxP6xASuvrAGL9REx8RM1QO6ekr/dqjFCgSX/fxBa35vq
OBD/fiGbsjcvvicnDbRNa26i5150/EHBvt/kJPuArzs+jRcLa01tz2+/l3XeWA0QAdemKJs8S0Ii
DITTpRPP5yZ0o7uBtg5MDRSMhyShecBWM93Wsva4URpm+RfJ1eG4+E/h1SvswaKIPmBylEqALB2+
Ujd523yem943aVY+ZxVrUTy9WXs6KBGKWHme+xBgUlzsmPEaLwhW+V+R9yPru1IDrxt/GYMGwUWx
pb00VX0voAyJgyMLRkgVuRznuZJ+GFxNg3OxWjn4B94qsVBhHktqMTQsCLoZDmzzGzmbRVkLCmWR
LawuRf4Rsrpd0xYetXK5GboHoaRfICzds87WbVfFjO4DRJ4QM+H0o/YhLuK6rQiv7hKHzP9Z9FDJ
J0hz2B4Rw+c167Rh5sWGpm8L5Cy/9BML4r7JEQR6FJ18FOj9kXRbS4oNG0pz6eQe6WexVOOQZt6b
662UjsP0/HKL+A5Vb2FLJKSxhCcxdhgmpPYaLcD3EdKWT8uuqlSMxmN3XOC0K9z6FJi3Y7wAO163
Q6iSl6Ua+FKa5/oo7GL7L7E+46f1cSdZE9+2NFYOJYyDekncFLTyAms+w61bYYfvXkJ14VuyOgNJ
vBCMp1+mRQlvWg0njDEG3qpLnojEMGm6tQwIaqckZqjpt+oJcupn3pJZdmQoLPzMCfs0IWKGmGue
BrrPx4m1XjVWLh5zhASQiVfA6twIedfXh2CS9+IaQ47rM0eKUVO9821l8TfJELwGEuY3k2wIlw7m
yGdZCZ29dL3k/zVkJ0ZgmmOCbNG+FwKSvc+LiHVVuBI3N5x82W7YJosriOY/3v3IgsFidVYX9aAR
FpmpRWtuChjTVEOW2v5fRiksOg2MWOnBWBtP6kJ/Xa4L7+ZD4Dba9452NRtRnU6JM/JMKP5EAY+2
G3EScpSV1lWl5vaylgiUNZPKLf6HPO8BqIA4XuqmwR5m6yM3z19D7tJ2/S0H2kpc4PJ2Aq/XNI5w
LPg9JXjvKdHcCs0EppG5TiW0G8cRunrH74m/NnzwpzEDiCo21jW82y+q9fL7+UTF7N0ewphfSpzx
dIsi+ARfGO08CfNzZRD2NMWcu/jCPnRY/cluuhTlK9a43Yf8VY/Oz5DaZ+3mKRpR+ovS+1GIvAGP
OsKW2e3+W3FCI7sQob00nPCrHmASW/L7EVPTpaoDSy+6T2NL/Cxs/S/OCI76mWP3x+es+quwQ/+M
PgW016+wamoyoKtDOjU45ufg8LvXCCpqU4ulcT/GXG+0zA9MHY0lbNL/KsBWhQ4NCIw4BEY2XPUc
tgt/cLBRDk6Jg3hYPVEUXyZKkW5eehDHPezRuxvblJe1x1oi2ik1rvlUWDKEsA2vg1Es2VeiCns8
SBHOsuKQwvVpmE6DYey+21ijsAk3Rek2xWPrC9qLr5a19XInL+xX/vt9Foyeg98gbA9959elJT4b
HdXkbgJR64BxUT/Q0TlS+IssMS8ZKiOr6/+3OI209WPZQg+0X3AlmY9LNaJJpO7UdbRTNe3+U76E
yMDHnAokDPiAcKb+EkVvi/ArvosV8ETiUXqkv++6Bs7qX8BhEDgm106FEa4F1kxK95kzN0GHEVLT
AlTxe07zOn7o9yEou6LZpvXgpXUb+4dJ9C7StooP67LLQFD83kE0IZFVR//Y9/OQJvAiYULXD901
gLRw2DnFLwyWSmPxnc1J11/fBV4o9Pj20Xfbm6mlR0MC2RlW8VhLcv8ekkRFfutGtFyVVMaCt/mv
wDmyVvAX1D0bDcM22nKRgX7VtG0eg2RhXmk/MiSxDRHxhz0pFFaPumwkbKAfnGqYhW2I69OgUNdF
yvISjFoW/PS0ke1MLhmfQasUHQ0Jva1W346yovkUt0086pH8Ww5seN57866zs09D6kbq7XrNACR1
SJuMK+604ZmeIF2COStCFUNxpFCspexPV1dZyhpBkh+/k2Gr4C2Gzznd9FQpYX1RM1zaWmK2lkb9
qeFjEf6/54TDr3NIxzVX5oPHUeUfQ0Zsymr5VP8OoTuaKKZ/qGkJTIi9xbMci/dngEvEF+kmReic
yjm3ywX2PNyesVjcNcS97U0oJ+JmPUeH67/BFWGMgIHVBcQ9SIi1t1TJvtJ20u+fcTHJ5eiF6ZYX
MkJKv3+ac9q+nXKit9nfzL7Q63tO2Mc3FQjx4XJao+nci0+us1v9osN8RjeUFqBlrawUQ/jdbesb
gy8mJFYpc6xKc0LddW9Qt9lbodyr1MjdtRu+97nspTQse6LGrJka6NwokpY20WLuWGJs787E8ALu
Zkkt3nhgZtoQkW2zbmmtpHOR+4perkYU3Kzo/GRMWOXyf03vhwmf9t/6JUZkHjjVMDu5aHpQ9xhL
QK+Nlc0aDAj/YB46RqQKIdcrL4MBb/ffhjHHp9p9XJ2HPvUtD8ZMxiAsNMe51iWjYUA4pZ5HRZSe
bfY7q4m6+5IMpy/9IVsYAZam8yqVUIEyarby/mYi+IVA95gm5xFuMFEphdF/+SXfBWo2/NZz6JKy
wCYdOyBzhtVAqdz7G1fWtO6D4koAKpJg8DwctWXLjm4/IKlrfg0eungWlSHH4r1Q++TLLLbWRkXr
ScUncxPtetMLas6gf0giFrR+6JXex5M10RcfRt8WpCuFfIOwCS4wC94c9hDjyPDwXksclai5XJdN
/0C7HVROmSYWBMSHbPj9fz46cECJMRbZ+a29AvplZwl/JL5LLdmnu/3TZZ4pcEzaxap1A/bkpFuQ
/41YRcJr8gQ34spD2rny/sQa1IgWtZpSQK+nwqEq85ctayKI7M54PL6KBh3sr+FRw41xprbCz23y
5dfEEJ771bvM4JFfh/QF2VZUjHmwN1hMQ1Dl7fR1AbKG+p/Cfgf9zQhNMoJkR/iJIj2SuxxOLGTM
H1auTqcg4C7ZF8fTCHfMHjlwlm4lnA1TAmd7ulCphgb2/Pw9S/1NbQ/C2fo+JdLhiQOSiPobVT5r
Ud+ZYMC5EM/MAoaDCmxETm8RGtULALk3pvAj0CfS/9aTC5uA7Ht4aYfi/Lq50IcrZdzwcoaIeTWG
9q7s39Rj0+Pc1KyjGgPZmoypFN1ZyOiE4tVQ0aC6e55NbnACmLw7SQgz8DVj3jwQ6TMGHyFpkulr
pd1P+kFKiW8uMgpQgB23AjK8P3X0i7S99Fza4zrOR93Q4qDCW3Xy9fMOp8/YLtytJOHKtlurHzUF
5gjz4TsB5SrDcINjJ54IsU+rhxdVrl4oZvAZ4LTwLbVpQswFgN+Wx3KIWHhIBieX5EDA6ybnPNdJ
tcrJ3lGnsmctA3zsn0Ta9mGFNNDP04I30UKrSq+nTUnp0wGdO5DaSgOHuRxTudlGKMMHsOBudipk
xAps0SJT1izjBfX+OTwwbvDCovPCGwPEXS73MiAH86c1WkIh9cC7Lpf/86dyzF4Ky7yws0m1VPaG
FKNdRcdmUP0PFrI1iUo2t9xp48sXVq/xAEObBxg31y9vyYSVNz+Z39mTzYTeoURUs+MZCpAc1/Wi
yYgyRXI/IaA7Q7FjPC/MenShGBfvQx69r/ayt4xQTO7E6HuXG6eyAFbQ/gVksvsCbZJDAuRK0PQh
RtsuxuL6tea6M9OubW4N1s+k4hagUDD8noJYNqZj1kWyZTJ4q8RCDZMytCXAtmsWogci30wWGYrK
kmGYFyquEAc9MYvTfmaC6z9q6fPGlxUD+sHZBKRfbUIZ+a+q+HCYGqqorTGs02mwzyWSTd1/V0om
plRsZAZM96AdTmxmAzlq38QB8VnCVxlb+h2T4FZNVMgJpkXiXfUyK4xfLP7GirryWOf9p5Y22Fad
uIHqdrHZARWVKLJaUX4167LVV+4GUJKtvWBOkmkkNpKgSZ/v13r0A5jHIxiRkrE8VLZE6VbUQeJ+
NsVtXHxMRHyLdH2cVzEaRG5AS4ovCvam+BoKOidsN5XwmUg8widk8qbgXIOr4Ma2+CNjn5CSbj94
8QBGPHtmhDo1F9vLcQ12cacnjzHvtRa7vzyVZ29TNnFiAbFYf1ZOuhlOWNGMEC80KvTCofp0eHtE
+bT6UR3fOo72MqRYAMeP71opKf5B5bIfjipt4wwWR3hYM600lOClQFvG+oTt2uwcPFOTxyNv5/iK
8cCXrZcLnZvYeDwDsLRP2v9qLCNngfyRAJ4+2Yp8OMrfUJiwtSYIzpbfi+XopifdOEmIcim60L9j
LzGPhu71gYqV9CRHtBpnOIHwhkcuHqFE8DZ7UkhvDKXg8yBVtKDj8DthPPGx55hEkqgrbPHYVwz/
+TmjSnkneYZ2cHPaNP89ZAFqXUCYZGvVqF7wt0CkueAk4ER/Zmbow0dhB3a7PK5FZoLiRq4s1lOi
Gyfc8wiqmFA34B7VkQ44r6OxHg/Nkkn8vSEsrMd3/AZUhzbh20X1KowCpNvt8ldka55UA9WHwiT5
o9Hs40mpaxFzTeI1TI0NrwI5mOsBNqONEI9qX3ALjiLp5pyp75mO0b++1wAAomI8jv2am40arrlQ
fIeHED4MAE87PV2aYiGWixtIKP9jntKlwry9vCg0KlfqGTJr2UX55qAVDya9icZdlP80JM7+fJVe
s5CbvGJajliKGLh5HhcprHUVpRD9qw/QAr6tX6w6UAgtaGlv67nga6FPhwVqIFhHQlFqFyrTkdrc
H+34WEGw+lK4TZeKBJnR32bhexUj19Mql+zwQsyte4KK2Vijg23hJsZGoO54Wj7b9S3VL2AA/Txg
HHv4EHb733l5uqAHYSY+KCl2s/u9U1GOWHyIX3SZherIrIN5vwuuyyFSPv+EwL33ZWKKLRKJbiHT
+VX7uWPM8Z89dxz3oPJHuxFWEENWtgmJSLnZBQf3TrEP6j4UNtvWBV5vES/jfoQVmDnlKxasDgEK
IZrFCOz7dHd8cJxXmOHj+H6hTp6gf6qt+9j5qtNBdpVjI1+38RjL8q0gPCpVR1pb/sQF5Krzk9lL
CWnyWSPUhYFGXuSx65ON2s4TZKHFQWNOCH3xHVVDN0jZRMNKJ0f0o1uMp0VmMl43C5QKwshcPMBb
uxHTJFmwt5B0vvfweUIhndDQaAP4GOqTxtN3BeLX1u/Asjj6dzD1f4U1AaBmGm2xiXKVKr6DnB5q
9ZBAqnjD/rromgYEY8orM2MqcMl4tVuMgqYL5IO/okOxDj3TYDzJbOn4aGp7VHj/09kHHmvpmb3X
FkpOb4pOKLhs1DKbcBsGxVEph+5g56xCVIAHQuI7W1zz9FqrjwVR+6FwjxBFyhRaDVuEylIcjJ8v
L5/jOtNtsU+60sHccvdyEjY1cUU8Ro2jOACMyaHJ0VfjYs7lHd3iZL6IqjXoY5FjrApr2Ptfk6qs
2qYB+ZXcvCd+FwwDg2Tbe+90jPV8tm3AX2fCcepp8uuqKg9RO/zXAm805EfnekWwahd6k8kPIR10
oHQowroQJb/159KVz21F+GwINMMtQjehS0ATZo+fTvlWbGgelh9x7mqQSnL8ZZkYptn4t7bPT3Gn
qp96VdEEde61EqK5hXi6VERYNe2ySQJ2qh77eR/xQSujUlaPt7c9fRCUM/TWX5DAAFQGycofex+J
twarmAx813dm9gVY2rvXeraprglPCtuCTK+EMrAyT820stdR+SvZ5g5HgQ6Lk5HRbrLt127NsgkJ
Vnw15pCGTYPeVTP71jbLpuFCtmBQyeC9Ak4wgmmrwFpWw3yAaLoCfOucQZPM3L3e4gWTKvkdhUvx
ubHsc7DdNs3N1aw/kQU0LVjcr8Xnn3Oex+H7l430uuqjdbedLh693JzuwUmNPTTnBchg2++ePOrH
B6jvkg5ADkjUvvsKWpv1Y6FNDRrG7B5ESDvyyiwgCXwbZnh0X5ka9qBXUVFa/b4F0kIMX+UaZrfj
royQRKWIJkCWv4s2Ra8ZyyXnFMGAUE+EkFaiKMdIzEsYIjpsSWa1EREtYHzLJTdPZzLtQ4hk8DXe
VpGovJv1hpiv8eDQCrsUM5f6WrXKL1vK7VaMwR8DkOzkEJpx6fVqbdOuDy5dOBMY1BWQJofn43fX
4c70xjjkq3Z8qhPNFT2WlLJoqs4npbdh2VpILheovgAr1eo8wc6b+vWQE04IWnDUZfnsdeixHnBg
uuqWRLOVznGPkbKKIupUbnMvfRE63BYnytdvK+NAT3Zbi7fO6H4Lf8lvTToOwvUXRoT7aQAe/kiI
nOP3xsbksNU0vUs2Fo+cf1fiawzffUv+JMb6hvciDpjdM0NKthsMGBNJFPgLIYagKwvvCRHRDhw3
NUArpcP0SKKaO4ULWrDCB3BdJ6EnrKB7AjuMXkyq4CEZ3kA+2MyZjTCi2GTpAOwFYpErXK614bbc
koii5O6XI3/oLvUVV9KG4VFhKtT2LCqOkGW93y8Io+CXKJN/AfB6iaDHA40i/a6elbyBMFGCwXub
zm7b12CG3XYufXnExSpa4cu7qnD4qxg/pTmADJPS7p1T39dntjcJ7+frP/pitJkKl+mETw1d8wYA
U6Tbx6O69wTlt5NTaR8jyGpEcsbi01pKipsY91cw5MFsVhJPnt1/ia287hQc2lXtfbyq1dEkeG7m
PNbpsOGcCwY7mvMAJc5bVNtkjyLhdDGnLqHpfUO3IWl0U3yQaj4RCNtkR7TGinTUihjhrzM89COr
6cmqtJv8DTMYT9ZHlqRjRk9YS1U+wqkVFFDGpdMyEIYa/xrmEyfJPEw9WRIM1hVzwr/cSrNLxa+c
Ed0Pku3ltBCdw2JQvmFkit1ZL47Qlm7vjRtnXyHSWWL7xH50Vj2y6YAiXlfGuaF6ift3WTpr7bq/
crEiwuEeBH0hogwu1UF6MC+hw+1CYQCfw/fQjygmQiKsyw0omIXkX8OGfGYiDSCwJnc3qnjOh5bk
IBsJ+CVD6rLp32J1K671Rq892qHz0iDDDgf8TYM5PbrAgNe2/54/k3K4RRry1a9PrLeDryPJBHXm
T04U+2I4uKUZ/HDnKmAk90nwBRRY7y9P6njkxyYFC5MxohVYr639UwuCUh5zRg0JI6lLYrRBihK3
h1H25q+B1q8/ZrfhRpqwNs5MFb2lewJB2mEOjoUYp39UG8iQDiOp2vxKU7sS00fCW5/IOeFBCAmX
Uwi/p9vzPu//AIQpQ52+73zEkL2qplejgH5ArazMBTgZFROxu3IwPMnqWdvGZ4ZKYfctnzFo6pli
LNSIwU3jMdOEpnsBHNm1BW201y98DSGgDfzsHiYGT5N6CWwQuvOqOIrxfgO2XXw6aZfIu43UGqur
bbs50J38A6wxPYxUQGg6F2GUB/WPti8Fzp+Z31aqkZJAYTxJvlhiTfrlTvBYWkWpBfeL/sGj7qBK
axAXSTfhUZr9FWAVhz3IEWx4wLc1K4Y/mqi9/cX3+vAlSp2R/FYfFKw9W/XSNBrfMCvanB6X5NXp
eB8Z8rJFu7W7XkM1U5hMRlwlvuV3j/Us0Sn3Y09ZbdD+Rdfm7hkQ2VRWGh0bCOMmqkco6Hw3zoOP
54pJ1nIpMYrInODCwhJnoXYT009MCgBMk1VLppMC4o2rkgVNwF0Wl8whnQVAoRya3bRJNZDSjTGb
R/NNnbW+T7lgj1CiiPhoerliMOhcv6XrkEMxhFd74VtddumKrwOpD5ugJGNI/lNpoHIMr9O8pQ2A
haDFQcGcmgIJXwmSiohDOju1cLaDwfeYWqcx1hYG2Qk04gaFf1/9GE2IyO5RqEyMNjtkxEnF/cfu
NOZq1bhLWPphnoq2sN7lIAJ7xXewrThRMfLNMRqWTnOTEpLKvZ3XxcoqLKOfkSv7KAsngzDHJSWr
9iT0Fn34bQMoizjt9HSWUqx4zoQ0BbIQorlULg3L26HTvtQAtF8e5fcZEwL4Ls2yuGfmiSlp8I3n
WJBzAtrut90VT5FxFI0eAxFau6hn8ByA0+d5077s2HNZw3T5aRUxDbIP991g10UlxLN+OTC3nEEa
TpfyK8JHIl6aEw9oCuJ/cG/rMZxns6LmayFDmOLUL2iRnISfqtp9zBwFLr+mExtbdgrjtTbiPdad
/mEE+664+vK6+PnC3268v+HpuLv5wAopBk158qTMrKKY8oyTeQVUekllopD1rNIBZFlnETXtAVg8
Sf74qgdVyrjPZSDAUOHJaxDpqfLMxw7R/4nKaVsQStJuqs4SDr2wz3U/CI0G5rxdtdHtY0yfZBvP
js9hWn2om8umWCdmbkh6QFrEF0T6ZN88pcS8onTLqVAHKvoDwjMp3u9QEwC4b6guGK9hR6LnTxc7
6SQha9YIWRh4egpnl4UoPpoTEgTixJUPdd960IQ5aZWLhOuwk+O+T7wnKkdJ968xTy1Lkujb0FoP
+KMPtrZ6WbrFYEwAnpX0J9i1f1HvAp5vI7tPnHkI6jGtmDu0ibexaEHh0JlbWrQ/VqucrSQ+3y0g
yK8yM+AIgzhmDFlFaOOdlRTaljgyh7UETC0x8BIbnuQROxssIyM2nlrq4VbgTvjWOzf5Etnhl6T3
qa96d5UqDfAhaOK6DFwhWuOMIBjxmJM82h5whDpfhe/p2OCdd3rukk+NMVGNsJBm1doj8+5aI3fW
eCSfnclKHs4BJp0oG+ZDDoXZhk9N9ozTKhIPbIJkhVGV22104cu2+34D0KPpRCqycJI9rSzAGCCf
0DUWNv93BlnVa5YWmv/XXamUISBO8LbqsohIDHWViq9lWZh1jdtWWwU0xG1nragoD8v/u/UhMk2t
HVHjOk55F+l/nec838c7h/JBbxxAdPkLyEpAhfwB5lxlZ2W9MVTOzasA5G8QcZFJsfJSeI+eGoEZ
A6bYfuNRgXNeW4xoR1/YDezO35VPtCjp48hgS2Tcq/fS+2xBii1BTjiWxJnLKsSdxbpdGdq5sLRT
lZYR7BG6p/ZBKsRKJ8uepxih7b+iDKh6bczbaLZUCvL3Nes1L9vBnUQZgDOkdjjr86PijgvD3j65
KNVJBBe87G1/NjJHacH1VIMXhBK63VNmmsmb7V6qAw+ahKVk1mS3UsDNzlrmBi0xlCigjfGnJmYc
UVOUpXoSNvDpo+SFgmI/8pW9a4bnxExOHgarR7/qwaRwyvmaVY0J3xGaNO6JrQFBsovVvpnaYKe+
Ye6LbvFHkhumiUkIqSgUU/RqWMR+2VW17MTk4GlE8oBlD8Zu4bBne0Q3x9QoaPv9DIALWSYazuFW
9ZsYslYO14v0FBwMZsSKe58jxwfj4B5vNYEBg384yk0iK0t4C0+3qm4g0ctm1KAZxHRNcK9kXJnU
/mU//5c5AUnp18T0H8RyRrB08AzghVcm4Yk4bpSfznq2QHLzRy7GW9hXr9NE2Bpjln5mGlumTYNx
5AyprSNPr798O+GJxA5LGJrtnXw6COo2KFIu6ejL7J1jnffkEQ4kPIgt7pCBSzViVRp7aTpB/Z9T
pYaRkF26fg4PmwOPehNbPXyXkaNm/RgYtJ+ui8oVCQeLdWcchBbMIq/N9YNNRJdGUxE6xGcWpo7y
8WNRB2+LxjTTO0S+NWeN0O9QTqKCKoPwa6b+msL20DKKdEnZMCHrBa5rWWfEpTXRmqRig5pby+Oq
N+Ky1+M4LTwCIYM+TrSCMQRnVDuGw9/q9FHtb605YudhqhrBHGjJ80L4+0vE3myADoqFcuIvxbtK
3gL2A2pq/wXWlo8i4USCdEUpNaUDKlrl1Q7xmdBIZwBTZ0aZsZiDa+w8pm6DRilkSjrjrLCF22QX
Clh/XAgu9ZW9WaOQ8smWuw+Tb8wjmwPW31AHBdGfI4W/oBwqPPRr8CCKznLiK8Iv6TOZM4NEidb5
I5kuv5ww+KTxY1Ut+n2Fk6TT93l6PLOx1nM64zcTzUcfGG0emssIOnhogr4WnqqHR68ogv7NQ7xs
v6b/vfOTcTCB3NPHodtnOpLvyLNUCQipYEtsf1CvbNoB4TyeiolNr9Ju/2dVIHmBfkIQXFEa6PCB
I8mpZhla+F+wCKXRiKR+kiub4DJ74NeCi35NBO/Re+uFfhE9v5q8v4LSVpbCHrSNVcvLy1R6d1B0
xsU2PH/jHWZJNi0VY0UvFj+BUv2ewQvVjEkuclefG/wwM5L2F6NxSFzOhJIb1ZY77nSMobFX4tsj
gghXL1iJoO4HOt1RoiMS6/plv2HLR6AojXaHovUDyOhoqqklNfR4bHD3tZhqsRH/sVrOffdqJPNS
tbY9i8DM7PWRnrPNh6MGvylSZd2sjfx2ukVIkTIlMfgSYxrVS6F4fFiil8OoRMSdIo6zm7rR4pFG
ZmEW+CvsJWd943Uaral/hXnqhARlv1JLDI9QxpW3Cw6bRLIy/pzFH4/1qDC+BthUedBsx8k6eDEf
U+xXx7mviG3kaxrRBVCJnk5ES3sl9AHvPSjHYbF5Gplqcb+fmjUXl9wZY5QPrGjrKH59V1Ngp3sx
yKfRWBMz4SX5yhzXq1nKJNWvkPWDuULVI/oGlHn5AS5jHV4gIm27HvJlUmTOAxl60UHba/Px5AdI
lzO6i/HGpBNDRIzxpzoMwpIVpNKAQZRAgM+/qj6rPAKz/jm0/CQk1x2oi16KW554E227dKEktKh+
oXHw/iswPiw2C8chO5lU/mXgQoBESxaC2fxaa0iPB7JR5rkPqJcHpMUF2zUzE7atsQC3VZ2+otZj
QS98W35yQTb3gLWwD7YUrCFWznykkt6Vy+S6sVo+tusl4lKZT/moH+3B4cn+WI8d3Vkjp9lqov+j
T0oRs43SLMgdsZFTva0hH6xFXy2Mpjeo7oYRvjgBoihBBv9TkagJVdA6Ug+HwdlOWkkhnfFnZJXn
j42U5b/CJ2nzgCVLSgPc8Pl0QDf7SoBydM2F7L9prRa81KHMpUSmnNxiACwWa9oVZC9jsGGGr01d
bVwsWr7UkszrK7CEn0Gopq1nvJoHwF4MkPG+q1wf4h82RdkFuK3/L/RlztQ3mIAX11iVvGjJ2H0W
sGzJFRuQF3e4Cj7Bm5GkasMlQkNsMgC137kY3aYFKaGVkaq6QhTYo6GPka1CXbNJeSvWwMo1GgAE
Mv9AESfT3kG+qugrYKYA+eIII49fQRhr6xZl32/G8mMtEtp7FwWatFIUQHNbHzL+YLcrvPCuh89b
cMB82d5ikvlUMwld1LPwxqa20x82DobMqyrNf0GVWrZEEzkJHVGxnTcjWpf6PBJV4kP23KV0AgVI
rcn3rZeM43xq0K4TUx0h5XhzrCFNsMdnuXVmxybp4jv2ovelXXxZ2Zte7GKBYUIsG9t76s4NTdyk
ezj/u6rxKMeZyZqcGXgdhh7cVm/FNlMVlcsn+fFeI5G3ZBHT0rchP+HIhUB90nVIDiOXgJfQvyUc
f1P6PSOpGSKMjYFfPFOwY3AFU7jZZcrf4UVg58Ju3Z+a5oiQlCcQdizzAAgOVGbC1GGEaVYHm+mX
mQ6/rckP7Bfc/zCwwaaV2ut26g3tzIEDy1e1gBHhtHmrJ8YsvPpsLrCMTO7Odcs580zZ6P6Gip1N
HGBhQeqOdag6kq3fHIId+ML7iMQPn/zgnIwTV2JU/Qn4jBWqP4eAJjO/K0bmqdWI12F5yQkA+rij
Jw0ezHvqKGxu5cIwTGrY0FDuG58MXmB4hUd2wEEco6K9Fjd4bw8kDmEpjvktK0lpyGAufkTDswU2
JwapRYfOMmyf1a/LTz+q/rUnkuBQEzkkQSEn0x4ewT4qGa01A+HMhySjSsDwZB6fjY63EaceyvC3
SbE18IebuaUdO48r/71plwY3toJuaQtjeGF7v5G9sAEadKKVwAtp5lf+pMJHaoMrOc4hGhgD4yoI
8piodAW5eNaGxfhBpfUvPukubGUgubc9rTgCBhWNKXhkB7ULUpznNK8ELfIbUXTkEBzwkwGDNGG6
yXzmy7JD2AYtM5zEluI2PtXVz4/0y0TlIuiMzRSv/FBVz03/wZy9CpMTD3GnXXsdXV3bZ8da7Iai
wlkq3sEta1oZMAPBdI+hQ7sP+LXcP52lIKDe5Lnsk3tSFOQyLOcMXnCnbRyFGqPPATUGR52nC4aj
eWG48HJAgbpzgrB8n2lH33W3GeJLduodyKv8fIy1o4GITecoBNO0NCMBd/H86+ZBS+RQ/xeZMupF
bSqOVK4M1RTXawD3PeOOOd5C5KzEcoV8S6vu0dytSgQQBBrb2IzLy9z8FFW5F2XT0al2imZG7w/A
gl2cke1SuoNbU0qRrg4/l5eUCzbwtyGVwcxKiMppoRp9NdGGO7P5/CmAF7ysiYMp2MpXlI7kyFYu
pwJIUsweET3bySEndysHroxv73OYtWXx1hNt+rog99VcvEv8hxkZvkdFKuZ8XOGwX2cO/HF0HA/H
3Sd1Y234DAnhZaIP2JJQefHUK9vsB7MoX2hTZI8fa+O/4JzxiWwWFX0g4oz9gUf7HVEFZhODNrZ+
wsJNI4zroo4XrZKxvDoVFa4xN7OyTzHGRPznHn1DJg40v4c7hlrDbnYPiwAmrpNGLkqOAiYyeE0z
8RmI9/OQ+4p5Ka2aGXKZf4ThYISJzlSznrDN/xkW/qeer7OeVGj+PUlUCYFrsoyrMppbUIkMP4OH
yFI8N0CTX8U3iP7resSt6v310nsC7o2c34xCjuRb3AQxlqLqK1W8KS6OdT2y/v3pKVNPZYGfxg3O
lLmz4qvFvO2QW9Cdq8PgynBHbSDjs5vprInVJSLJvjP6jAuJh8fgpHg1q6QWuowKMjQ+cjbaCwNb
N9wjvlew1WiSqZZi374jM/wmxFOHzzSTSry215sKYxvzC2aHftwpwI3LNe+qklU7vYX1qDFE21ZP
31yK3FYnb7TFzjxhCa211O42Xv0hrmv3BVrx3jah3NkOIXKd3U1IFlf7f1GAeq6CWDeBdrmNGCvD
VrDOAzg8oBxsgdEt+rgyV5MqNDxavmFuYipgZQcbBHLYbvRuw3W3eRXkjff9OkYZLtfoeJR+B13I
QAx6466jgggYVEndPifKZnL9CCnpYaaK+3OXhOwCeg17HaxIyiPNFMErYpuwZjn5wRDEvvse1A8W
dhxdr4xVAUf+Crmms03hveSaExllR3G7kE4MQ/9Y0Q2O3miQ8Da9htfwN1g+ECT5vkSeHG4KEj0/
oUFSHtcN6YWLhJO/Ma8IvMpmT3N+9vvU2KgFBlyhGZXiSkQNceHjGxJoGLqrCwHG5Oj7N5L1kwq7
rEPPCqS7YFD68aVZezZ0JCSwpf2PlNqRdRt7FYnfBd+Ix2ewenjrgH14Plv/fAEi9H/DaCN8Mq9t
/gQAZotH638pQKrxjyvDqfCkK2Pa+0bqr5SKFczyPnrTLSkCFhd98AZ+XvORvhA+jM9DwOkUN3OL
Mjik8LfypHLcx6WK6OhL2KTZw4z4LcdcNartZiTcCx/sKAKTAxnGEtz13Gd8MRXK4STtgAIlsNcc
E0N1k2xXGTULSolgZgqLkhSsDBNTODiG+2AC9lDT17Ma6YfJ/H3G1mvaPUgpVgPJRejc5Gy/+e5u
2P9TPaTs0KMQgBdfnr3l1HK7OoqGDCJ0IhjhvdpIb98fdwxZHwTFPGwaTWQsjo9OoneAN+F4d3o+
uU4+TGyXmGJWO/91PxXr1Qw3N09gX8rA88JgvSMC2KfYUcWpdyric78B/oIiOsdODDVlfP7SdO6F
PKxN7Ezr2aWH29T0WUPj3crhrpaZe327gR60LgblWIWCDJMDMPdaBpZj5EvECLHEdbxCg6x7VXFh
etL6XUPB6ZoDPKJ4IlACL9pL35AYUItwo24qfMRhnCfKEDCxlVNzIopMkNuIkugrPV1lXWqNBP/2
f6Y7HwiCUrApOGkk0HPBBYDQEEUv5zO0ApWP2WKzJGQcNPXdDN0CuE6TANcpsA07qtYoCz9KMwHd
YSR2On12Dwsr7OaVKpGlbdsC6p5NkQbxnjb9nPHqu8LdHwjAO5CDezML5G5yetwtmXdAN6q/7B1E
OBRtkLfdG6aB1+hevVWfRLW7CKMavPruSTeTXP7qBMtzpWpfZzGP7RxMTLjYyh+8Ilv8HLRd4FzX
LBGWp37YKqgOpORJV6/yivYZuBAWrHfsRF+7mcIvwxI906fjRgppCQrkcGG9UZ76d2thxHJ7BD/E
rpa2BmSo3SY2UFB7PAUfH8doWjQbdQ+DL816k07fryFC3Grj/w0Rks/B7bA+8CsGs0MwzMX0+v6D
B7wl2KS2HkQZw/W10ykfVtaX54sTMfyki+RtWGRWCMaR64JCmG5Kk8GoheYKwh6Hb3q4tH+f4tY/
i4/Qq6Kq39GyaICs5F4gXxPvGXNE95H6lVNfn4FbVq/4CXY8rkbubgnLwAOhqiTQfMbLqd3WM69I
GL0c/jxDhP7DwQdbw1rVg6onjIeT116FuINsQ5rpJECSHQPWDaaZhwtJ1MMxzPIthZuWV0My+QFT
O8XPg8RuZYCJZdaVSlvfdWo+K5tOMDM3Ce37Sl+VCtl4tBwbVbOmYpLyvjFZbQDZxawN6lrCpjAX
OYb7kv57pLUU7Kr5le3dToyjfQUlCeeOJnfstgkW6Iyj3R/maT3M/FZbke05xnzeizn4bwMuImn2
MuzYYMEya9PRr3by5MZrlKPsxYdH/TMMhY5KN+UsW/HZFzMJQevlOs1/mPLlZaMl+pbH24aE+wsW
ExD15Ci42QrUYO0FHN6qpVZYmFeiZDsC9uRXfz0uk4+gzmFdBE1WyNxpLnip1/EjRZzyi3trWUUi
IxFnQMR0EIkfSRf1vPjhFkBLcqH260rZBrDu20aqDBrpcSS1ybakHVHlCs8X0y8GOEscVRg9uWyE
lHIE2pTO11wn+4B1wS/orBzmWeef+bGKtyUMI1OViAa37QmIPb5OEdXpojnyjYV4P5v36pOXnL8V
+SU9rCGKVBZZ3heMfchlVm+UDQbmcHdQjXvHPHXsqD9ifnUpSETjI7TAkiX8gQi39GOedfQNuG2s
NkY56XZqYNZA9yTngBzBB38JAihPXNSgrbWtUoNwpy6EpbShfULgiso+OUIVcv+EQaIwhNGaYAvL
9Xv5oEWJpWo9O2DxJyEx84KwaLUy7ahA1sdKLfhAZZfRVQj54J36GY/3mdeNsEYh6GEiVhuquKYj
3Hxe7kU2XXbLPCE+rkaIv6AdH5H/iaKRy9sP0lV/67hs3LLi4wnhexAFK03mzP24/OMkIhNo52DP
FplSGPyUsljfF0bIi478KL56pouvG6kzRaXepKGeRNaM1KXPaETBV5UB/u03wk0x+16zmz03oA0o
acZi8PeqPFsFcLw8eV+g2pE1EhFqOSUdJ8StDG26UMuqRXui4VzamBMnZfCXPOJr7x12a94b9DGc
RaOtKI4Q0872IXEFi4flIPwu/ieM2dWPYl/s0PWWj0m8uBzcGYgZYs2Tfqf/gS37bJNt4LmD4LCx
njFeoqxEcW6YJFsYE2S5LG65QIykwfPyuP51zHlDYL3stVeSPmDIei+ODnSfjP7PbGkfJXU2zQ/y
NgVG86KTd/f0YyudImXAlpdtVm9ZPlI4ZCJ3VeZk5JMtDearB/433vm1hng3zNgbSALqs3f1WNCs
nxijrgxqb07dtTGBu79aURzY6feQvZGgjWn+Vhw+z1rw79LFUb1oq2XL+y0G8u6fgf7MR1cf7U6b
U6ndT143UGepnOA5swPFdqS2bxuzbWg/pgrCT8D7p6Z4wCEy4CDjaiGFSD57oRf3DwcQAELVR3mC
j0uJkQS2L0brG2evnuXXqjBCqBZ8Jkv8TWmx37v1q/hqnhf0m/6GKwWoFG5rh/DTNzAnOzXgV7i9
VD2JZwlh/QvAboGntxgWOb7omdNvGeIHHmF98uyZ0BtAnwIsJAScWbBdOUaZ04l1Eew8oK7a7Ukf
o0dR5aVmO+vMHI5IxZ+kdF0BWUGWbmk2rgHImSpeudsrTiDBiZ1wzJ9VwxdsYg8ekNmrTW7oQdA5
K544jZOBDv+pBGafbNgzgIWcbPai/nu8epmFG3IRa3j3yb2sFPCTv4YwxBAvJySEcPYTuVNpPQfo
CJ+WoIVglEMj5TP6meZEL1go2aIjNXa3yqLhu7bq0LW80G5QbCgDCSb5EIWRpFkpk8fnxXr0MlOI
djGfyeD2GpUti4tjiSXOaCe7hp+VehkWqWEHTfXcJYsGXFqrT7UMS93XfPln8otq1BjM0k2u2Ho7
zoWI2HLGHLKp9NJsl7tog+xZ7xy8gPnP27jmerUFyodIbJgU+AUQUDXGCnQsFPoa0sDdPVi6QMOH
12Vc2roeIKI4jwl4+/65deiW8gbs+rvlHmzlbFYp1KpyAxhdWpwsr+uJerdGijIhShQuOLxjjjxP
3Dfr4jA+eMCJqD4Z2Z+1Wyi96Q/OxX7LYIY7GMULbYBhMOcW2e2S4ZOBNq1Ig5824CfBYX+J0NN4
igZ0vf/U3MWEut0h9TJD+p4F0HinkycmzzAGURGDB/mU2DCYY1YKZd2Mb1RZaNETGBFMHKt6X5N3
e+i+LWlFdH8+lESOCAcRhcXhM8L2cjwHQr7sBDwHfpvvfHa5bsLjd2pKzjL0qyHo1f+7Vw8a2wn0
KeKRugE0Ptft7XQ/4nAtUDlgjBpxYa15+U4htk//vsbAiM1xZpGnVvuT6Arz4N3Zm3H0p/9Tg83N
1PJU7uYHi8Cx2wW3XUP8KdOwlJufUbVKs1jphuoGv8lDcVClO4gWhxzmTtYHpJV0O7K0RBUVnbzD
dlY0yKRvV/1upJ1md0cJgBuLsLd/nEF190klVGQeXRRPExGoSmw7TNg0dpe/gL2XbQI6Mo934RFh
6maELwU4XGGc/GYxdYTdFwkrLi7SkwOfVVmkWggrC6KY0+x96bn7pB5Oss5SHeHMcAXSODoSNRyE
bfp45folgx6FfgAnjfPm2DN16Cwop4TuRiyAt+6D2Nd2XJhzV7WC2flr0im/dgMYA6yZXlwpFsgc
27Paiy+8XTI817ypUv/6rvwoDonY78tSMdCiUXPL8IgEzy0/tpe9lOHppQ3mbghrPaF9XXGQ1f4+
K86s+/2Dh59FNDPPmqYtGLSd8rys5f5cnuKm9NOT2ARxYsgSYBI0aZVT/g6Y7ueSP1UkDYARb+gi
rC9FDkqFNbO7bTqGSKf6Z9HMmEN9qV5x0pwDJcOX5ltUjOlOrzgiOigEhqRw1n6Z6D9YZAZk8JpO
riMxnOX5Fdh9WC1skz8d7T9AwjtI/r5znPWn4T2MWrQPcbZAniDy79EgN2+LoMDoyAeiIMNeG9g4
Jrqh3tmVLS82IYGezTB8Cu4d68upTUnjyo0yTLDYm5ozuZv4PP3farIUNEL+KXDLdXlRuagQFxbQ
RfRKmM/Gz0Dsweyo7/SW6obO1oHpHQBYjv4n5I19XIJeoOU/q/ba6iSTkLJDOGfdV6DrrsNUk/ci
YRz1OWmGjhqA69im6+/rxWrOBYw2OohYFBtHjD0sBrKWZNP/6jIWTKKf9tsClUEkB3xyhxHviuLv
/QppdlhlgXQQ/NNi3nRRRVqjab1aoQDQjjtpTRHisrebAIjJVJUROvka+qajlxrcPewbVMAeAWha
/EoEyS7KS2Mk39ZDidJ/RRde5QLYaTyqSg44bV4By/U0PFKC1GgymiAeC+qhKZb/W+Rjg/kIje07
c7wC8iYeq+IJ/CVAbF/z4RjOBxoQYSM5LFOB2HvF2V1VC+2VL0cQ1aNxdWc3DhM0zhj/NeTYqw/B
F71woiCOhCMUjlXd8kHW+E1Lt6B7l4qGTF8K2Qz+10m4wxH5CWYiKdatbLhcoZetJnB1Mi0SnI7B
IqoOBm6f32WuTKLPe3VgG9WG9lah+s1Apt7VodXuIjtlQAeINK/RbLtIEh/hom39xoZO4KLfrr5g
UsikEuvD0/JEZmFO4Q4afKsIpEJ4LNRhbZ+x002juqnjBJSZ7Qwe72ZnFGvA3fWcD3QHdnJiOe9C
MRVaTWal4BNV/1DFgnYGMjNU5Mb9UuDJt45fHShDOSoOKs711Y4aux63rVPo91Zl6PD6Fp+iqA1E
7mI/9EJnWTluk+NyiGQHDuNcChJiTibvdfwELo8ZYmlW8B60Vl7mozXc/oEmm5amm3CUosJ8wsy+
KLyVDJG/YecUA12w/Y8LpejvMWaYk6IuIY7DtI+m7a4MTLWkClX/Pg2yUHmzQ3lDm2hxUEvKZzZ8
Gkpx+zfkkvKzi8G1LSGDGsaSmeqLy4gKwGFXqiUoiF+TPzDHyNj62Ly0qwjcTroxyjrKzE1RROJ7
xeR/dpprcM/jb19VRf+AcbH5d/r3TEJvZxy7hatqylSW0lHEcvjyxHJEoFCqGeznmPIZtZXkRwSX
ZEVO5eGqpIrJLxY4FHHwOyDqrk9ySWBiZdTIPqVONQq1TIdq2E/FUL9dExQsKSBoXTtMKtGbtSJ4
mRria6yTgR/nV661TFxorhtwq/TmBJ9fmLyFF8sEs0U72FGdcxnuYLwKphzTZul6KKyT/FD+vM+H
HsinmrzQq+AkX6aqYuybBD4okPWMe4sX5HhlMV40UcSCOwmQJqLxPPw26aUypDDPt1mniyazQIYg
vDxOZnm6DUSTHNzrFsezLxTERifkw6kNFbb2g+3ECTzPNF/6zjp8yTuybQn4yqfoQYinEGOuTKRM
rJk4pbnNSwg4e6PbUh8yd5f7a2EM5gpe37utTSISMKNn7KeWuT3NgE6p1kAWSSoGTe1LoS2mA8Dz
q12c4ODqAunHlFgrw70sH2UOu2m45k5J8aolSQUwAwnqHbXSztVZBGUCqzOcElzHSK1R64p5YrCy
tzbifjKEe7sVovX+thNhYsGE2c1fCyAU7HwA3axDnE4wlQ7kTaJvOiltu+wr3ZyP4jo9eEBx/lv0
eig8JUzCLnsFFhmfQn9hK3PcSVi/KvnOtjUo25r+2s7VC4OBe77K8ACota7DGu0hrze2XWRohsz6
YN2Lb8Uzd7uN8LnLgN+TzXldr3QeaSebX5NRYNHEAyhjdRgbZq9DWtrhY47/MVTswHEPOjt6mEwR
kpQCZ8fyl6O5KI3jxy7T3n4C+OqxEcD4k7ke8bS7EC51u/vPTQm3CqBaLFnqHxlckWzUanvY/P1M
xxJDTYiRJ7pTJZF2IxVHY1KNTjlHYBFZAzDrHqptkhadOtXc7NbSw0EQ7ady0naqfCfJIf8CRRW4
7gFjzisGXdB3g5/pp3cA1C9S5O1jfVV9PDh8wArQXsZ9pc391/Qq+JJg1fbfmZt7GeAXaLt1MewB
kYzb9R9V/HpTtJGNneYq75+YmrCo0NVcoKgFbyGlaI9XUeSeXpuSVbhrJOUPA/bsVFWyrNC4y/72
mvAOoAAau0q98YgoL7D66pyRowLHKrj+Pkkw3Su0yrilizhg5KrWjJ7Urs061wvvyXa6Q47KsBDy
VwFAK6ZrH2lvpwkdlMSf8kg9oENAtn5yUUTBOWXiEDW4E/SSELYA5iSW8/n/Fq44Rcm0gTGwKDPx
rbVvyFELs/BXlE1KH9dHdal6Fl7QGM/MLCFU839I3k/d3BELg0bpb3EEFp3L8XDVO4QdG0gIBLXq
lzhqTMAiocozhukK4biDAugvcfCBTjUdmcfzi9MBuTLKa6uQyC/0m/Wh6+Uw6c6wJpljM18lSn2/
pwhtYlDsYiKD91MDBVMl9u7QqlfB5oU7KoNLpiO+Iwte4qe6akxmF58xK+lrJuvPOT5jpspslEof
SZ9ejMwOfk5jwOZZjoX2gol4nKY9SmzSViiW9X2SSGrEmdGDfFX2aPf/G5NCDVsqpTSR1MzhKvNi
BaHuj3Comko6nmwqqOZZE43nws5fxUQ/v5ml7VJWrLFup7mdjBUBrqoosqw4sLstDLA+gC+yyjeT
ixR2ApsOpWXP3et/PhbdlugMf8QVI24Hbr1Uc+yd6cPFGBm+cKc+scXy5PcS589KS9Oi0e3F4bxh
bNxZ4fZtYBZqtL2rFZsF4HSk76Q1lTJR5ybdjKCz/wI7i5Hwxd+aZgLPEOkUyuXWhwUrptNOxqwH
15oeP3p+CfMBpazPamIiYdAIZmVpyCiQNcf40aZ5I/gYvMZXZdIMhmQaeuM3z+U5QqPf4UFncyFG
aH8FpkovL6Vf/gp4YpC+UD/Pq3j8J25IqYBY/yxxzGSY5nDI0P3YjJrmIyBDY0c30YyuMbC31YF7
wrczSwXTrdADQjKADd6Yox358ARqTgwKIyYLo5dgjL80BcM49XOI3C+jp+3B+xhTnAZAMdUgMYDT
xu6Hl9oJqrOMi6rNyb4fJdis3igzui0kKAW4jqQrLsR77f4PCgm7mp3nEP8C4qDip5UiNfGWPy4D
p8xuyiMKze2erwlfjPWlcBxIUcO3vzRAYDbZuEDBX+05p4SoXdb9/yFbeUHvkr8vw90naaQ5b4g1
kYIDM/pdS+UNWRAv4llbrz4D/nSzjkDfbP8AQi2z7JCkH/HGjZEJZST9umUxIgLvuBcqXjog3SUL
tkKuYMNHyU8dGN1aTaG8J5GFyP3ejUgfCZ73Z45cAXDYrII2Vz+SwH/lVPVvDFLwFcDHLR3uwZxf
d8Q+AQT66xap0KtXkolSpH6oRPjvPU/qiQ9/71xztMpCHuUanr7pAS1UIhvhOerLSTWD2rzSDk3Z
fXVtYC58J4vV12jIBPSb7Mm+KC/3MTBsN64qfY3U+uvAWJtU+yTIy7yvGxcLMfkiM5tQabprR4G3
do7G+Uprtwb+5rCZb6cWCiQGRs4GtyyGgotLikCHZKbN5I1zg2ItuUGGX3HBVWYTucEvMvBwYxFT
mqhywGhTIbQqxbMc6xLsyLK0bCXI63JW0mgoPV5GwchE8Yqvl63zy6oQxlwRcCcGPLBtI2Y8SUEp
0QsBG7914VNN7IrTawmE+deu5CouuPKInyh0xzplwZtc71mrruTLwb7PN9Z8VJqIJv+Cobt0dWoB
aI1n7E8ut3gt2L7Y1AljsunVYEeDV5Dto9Azd3XM+GF+WNO9NLyTQEuUhkXzcjnp+JydqdMSHNUe
u5Xl56LYFqTH1j6xXpNSAkvfLon6jwSFgoU/sbKIvvVH6bMXdoUBbZv2r2o6/iARvkFdPQGGggLT
xxIJnStg1EglynQyYg+bN37m4td2VY+piX29bWATwPIpw3nMCUZB+CJWKfbIgJH0NFV58pz91wh6
BTRzdJADgR8AAt7dxH+MQk19FrWwbWtPpeauj6xVHYftl3rD2/K0R3Qw+Oo1/iZ7g8HvAqoFjqcx
NxWMp4IDR12BRiLcjtZKCqrg+UqN9WK+JExmPeHdYvsEx2WxAj2PF4t4L+EnzY2vo2eUpCmDywKj
7iE5iiMhBAFPdazVOBgZGNqFLehEMCTRIJgsMlXpKPKBvZFPFofRRCzEZNu4Pe6uNjxSCeEhybQn
QHTbOFCaY5Yy3bgETTxvsNnJ1p4ijauM0yputBqBfs4baBCeP2E/QfkOF/IDDpcka20Ms8G6siJ6
BaiEOVqnz3EELP0nChTvJxXYBGZPKArv1Eomr9jh1PkIL2Hx9n46t4Ss2IHB16pIItleOfqzQ13q
SWCekxm6rXOd0x3kmLUxJ8f/8adV8iwPu0aMRpbHdBlWXa+ykGSHFirZvBPkbbPnCILpOgaZbpPa
VH8Zik3vLqOYiVpC1TbtV/tAuvElnIdrbJj9H77hLemFgSISyUUkkuTt24+5vJz9+INH453BapgQ
4bR6UqVqWH/NevCXfB/jHmZUF3jRJTbsdpGMhAjvD3qFTF0/QvJKi4kHrce/TEsHtIxmKvhgtASN
TOG300iSWO0GbJGxHcv82xEpzEqLPuPRHcXAncayx8SKDjcuwIC2fFMmERkuA1liCOfQKFgPuG9J
dJRkbckrIr44NwhbQtGIxD7fN7Wxytw0EuHzBUzorwK6MBOitjHIFKUFT52P25gOLdkK632WB7q3
QRr2w1ZN2J92aG0pbI2em3DPrICiG0mdW1edJXRsxoa983nuOMZZF59fIl3QimaCLM6wiqVTJNjz
aZsOH39bG9Xkd2PocSxnnqKK+OdxHf7MaCXFty6eK5+VMzJWRF/8EAeNQe3pvNChDvDZGAF8V8FH
uPkAcVVoQqU337xAMsmM/LCRBldjsM+vHKXEglVd1LwcwB/qMIqqMqa+Rz9VxbzKKDRUY0v4dF45
a04h3S96LpEIQPd+wyhbnRaRf+gagHUcdcoZh7AnqEOwm5tYuXDyTytv6Tb2fNOicmmBWqo58KRu
eKOcxe+1hbW7A7ji0Gblsy8GKxwRIr7Ab8AcCYbVycvW+qccQQXrI2jeql0VJzMOU81MSj7VELPW
wDJZpZ49lrMhOsRa2CDEvDc2ZwNXl8R3Q04k727MDHgiA+ZSzpQAQrKVpv7thILHIumfmmjnV2Oz
YeFZunln+ABZIfDrdXchMBHVVm0G13eEtV5vhRIc3hqyd2DFhVv/p42Z6SS7mQokPP4fOkAvG0L3
ZQ1v0tbbNGdSuK2cNP+YNaE/MAzf97osLq3nXYLZFcQxjwuBwDRzR3O9T2FD2KqPp+4SMbbPjxp7
BZUqQD0caHFSt3qHpoa6gy1/GXX/MwyFJiPYiHPxqxTziygaMumMQJtre8heYLqldTpe6HMZelem
jsGtFMS0KiVVfTbbm33ggy4cywrAeaR4pdNoUvsbnZcqPAbB4gG2d4kfQbTS/Iow9UNEmr8UYAgO
lfU6d9U9wQ6HND1j0k7+kyF5eavygIKZxlkx52y5/2VNvwXPTo1MBLeGdDVaAdHuUsYQ8DG63MmW
TmT9cZo0m68KDkNUP/lyR8jN/5MfITyZ7H0ABR8WcvScu8fhwS8T3k/7lMOEpIiP86Uz7fOywOui
GVkSRvzOQWShe7BJrnwaFpy0E7ENwFad85mYqZtYgj7ee6BI87gv/qDzifpnYOsCOlG4gbJMerrH
zpSFJJNh83QPoZ4f+FhIX1kShxekm+pbMKM8kckFtILvrY9Jb5qTG50PUj3YyU8r3/tIByfGNtLP
72FB9MNexn1S9ajhbVMiR/ImlEBB6MzN8ZcU05aPbhwt37ykUDs/sBdwXCgnBfwq6+4P5YN/pFBX
vcUpO/WgeqyjMpsot06MVLHEkhv41u7c1kGvWG2PJXWRaA373S+hBknlKNeAhSH5uWOi8R38fkeA
FjLYk06vUj9z0Q0pnl16x5k5glmuOqxfaD2NVBiwXGXL8cw3BOjDw45ZpmtGCCaOMRMh9VowBjfU
n+GH4wl6a7nwQ6F/SqA+iJ39vq92fdoGUc5aY2aO4NV0/SzQ01kUtUiWvev1xQ+M/t3izvCdwHr7
+/fCXvzqUxvnvG6yTgWiBnRzda8mvqVh+lPLfO9HEqZIZhTo3TC2IckB6QXKNxU0DavKHTqKIzMK
8nCsIgLhFS9+AhhlpGs8iFeQ6JKWajPIGkpqH+f951+Xc/aV3V/gzM7UwXj/cN/E5FfdRZKUtk+U
Ri6p/a8PnwWlVip9Kxi15qj0VloQztKhOk0DxG0lqiQaa5qXjwLXmvg4sTYTgTrE4kJUtQRpdbcr
ActzmUb8MAMvfQMK0pNvu7knzYvfjdTTnPywbpP9k3bpwHe+lg99OKuP4Ao/kfrKifTQXk7O+Ztg
g4tfqFDwNRGhZvnPs8axsxInwy3JiEuqKTZqlgQ6NZIjJIFJRd3UPAzvUKYmxJyppzF+IJd8AbCO
d0qkHlOSqzd3fb6dQfgbF7hy5/HeQ4t//v3YA1BlySeceNj9/Rd23AX7osKEGXWtpXWlMD6iCP54
0q7lRLpZPz5p8sOfmaq1PdnRnbwr32HG7265xzfcAKIav3o2jT1DfeWjCQbz5iYaEl1jDp5wlmjy
AUjTHTDG8pULbTRy8n3Z/+GHp0d3dNnRhRgFev6l8z42n86ozUMRn0p3/e5+ALvVDd0h4ZMUDSSE
PhcfdTnOmy3q97u706RowcNcv83jfxLA8osd61sERxTazYAVXPMh+TJX33FMTVz66fnt6W9b3JuD
HrPv1W4Sv+DlYAX6ZTmHiU1hvMYbVsYyE8sTEL6Sgo6V4PiSkda/Z6zi9cj8vPJ0r28ubif3J2Zi
aQuM3GMoXZq8jzSq5hps568pf2La6UgUqYAe/399i0g5C0pLsWphNsib5BqtOL0cyR/Pqafl4ruG
Fxu0GFXv5tKbLTTQqJOFHNnJJ6/eftdsNYtJnfIzGmhyqD9qb4+JydbGskLGFyOXN9v2YIoOIBiD
SPyM4JtUJ5tAQSDVjBNGRg0rhuKejVulbo/3SGqsOx2vNjr+KjCCE1ck23qrFan1LujZ94aDqPjd
ZIct80OhMNAcIglPURgVqxIe/aN7DJeT4YmxvGwg9noncSXsfeaNNz8kiYZ8m01vMHpsiKEb4Ykr
l14zc7eJlULxjEHEc9lwaCvLq3nodOc9XWpRlqZ/fm3PH20Lyq0T9XloWxmypqRsvkE3ftg4ZC5g
UmEODCDw44K4etN59LDxJsfHD2tHdxQdEp50YvZRp8n51H9QrVNt6qL8pGxxjjmOo4OgBW3rdyok
ik6nVef7j7wPeU1zoscDL5qHCiN315gf2DP9FaRgUwGiF2F1NLzk1h8P1PRm1x4jhBGrjsXLTp9X
3ICuJqOggJ1D/N2c3VPPmdf7htGDlJWCf4FhHtsss1A5Pks1FTUvk+l8Q7CzSLK/j6sLYX7WC6u0
E1AIO2zFfUCVS98EdjNpmKzw7otsYX51i/T6AHuMUSh3Sdu/qHrgiqN/Lraz6bqDcy3XUXnlfp0R
ebnB/4Eb7NM+UrnHtTBa4GsCamSXRxJXOdMS7tapqXEOnhqBUcFwvHYdpimgjfbYA0WiZZZOs+bU
imR5brAw3LYIY9qpLiYk0wiwX1MJTnSz+U7Z1kH4S2DA02+gJcFxU6JslCdziBdFg8Qj7ei1Oary
XuejxvCioHV757XCi9UmnD+bEzwTIhDzu1l2Ll441fp21AJbsDF/3EPA+roGeIzcb5USNe2Fwc09
Kv5JIetN6pf3PINaZUqJ8ZvcWdemaF3y02s8HiVn/k4rvwQCLskJnfU8lSM30QbwgRObdV6zcVR/
/ujV7A6UL+qO95MQoGuZMj0qYA2mYmZruRt72KYVXijqWLQlGNrS8JoHaPUHLCY+qb7ed5Yt5eeg
e7KrcFBpdqLdhqSsfl2iRRnV1jrIPuJpTsYj12WGhCYfH8YGtsoTj30vkGt8u0zJGoD4joT008oG
oDP3Ke0qXUwssx5epjtGYhBH3TZkKZ4uEtM5I7ZO57iw6VvANoKTJAE2WaDONYbqzilyCBXIpeIK
QfhLn/e0NI+5L9VXd2KMSsdSpgHnrwi+O6TmzmLSiw1raS4zVrgpGsTtm6UbM6iI1cnzI71WAM/h
PS7SlH0JLwt1OA8ZIHXoTUv42mhfxzght6AYAH4HJLjRbqxHCykaFKsX3kbR8DifeziiP71qiJEj
9Dk/V+z3urUHU+7XwtELO4eX4f3xah/ii7DaglTsK2lTy0ZSrDmclg8jnSzC91ccAEAAuity9Rfd
IEuAypPhA6Wlrq7TkR4xIw8159sKsXTSLV4BD9kCPUQQ4UtPcHx7AEWvNASuXmC9lEvVA7xSK3jh
X+XyQuf1wwXYpm6S8iLLOEibOVWShYCvsL+vb0lEYmcXbVU1XXzTAgcrLcwDZmKrkjmpb4inWJkA
vIUzn7e0rlA+NVIBSLxRefjsAjGYxC5fSwe2rCZeo4dNetG+XlpOuMl7/w3dDRM07vg6GtGjVkRI
abcpXT2KTguGZl2h0ms1B4BN4B1HbcCeSS8Fj7Zbdqwu0TQv4eCsOGcHIITTnMInLg34DyQeyMUJ
tIKCqBefvtv4wh3Jjvf56uPVyQHzGTMdIB88JviIt0wH2ARapv+FlR1SEgqxVxtdGjQiLCWtdKIF
mkqos+68h8GbxpJ/HRqTRNBss1r7AF7ohxUbZPCia8fHdNdL6kM5EZSBWiYG2axhMN40+PfSxZw6
+MnYNc0a8ByNpF9QcxBSecLIdM9rsv+PcpCzoZDBLwiiAsA/iQ9YKyhXqZqRA3H8EO/zNdqS6HL4
ynBqJ8WtjV4BFO0iMZQAR7a/XshO3FTlchii5RbZtCoLRw0bp6sngjNdX89NnIUEl+p8I5PB87+k
4FdbKqvzPMfNU3bfbIWz1I4KL4vGwkoUGbgcBU3ulf4joaL9xIjay7BTXo6PQ9sptdP3hwq/gITs
Cg5kCCH5qCOTFlJ8JKfueDcJoSkavLB2IwgH/GlprtekazaB1qXe3QC2z+tiXOKXhoTmFYHPI9I7
MIpQfslTcY0GujFcnuPrmgcDHsf6TU059oORz8dZEyYXjx2Ifobge6j+XpfU79Mo0MWHsHj3oW4G
4XY9+lHCmKV+BOncGy/N3C6RlF0IXsNVq3tkR2BL3jo1fSlCBoXMK7wdCkhl/239HTFHuEf6msjQ
+umFnd5FiCaxFjOXIn0UbHli+zKiEFqn6Mxt2dAzKb4qYbD25yXFCMdQ8ec+hg7QggR5X6tg/eW/
bS8GwEBf46zr+oB/q+9qZF6ggdHpIxw/t+mW7/zYDl/HdAPayEshxzOb65ZLmNCIwXg9juJORWfB
4/Oj2QT2kdC4n3z3V1aVj9jJXwAYgUfHRyYil/epZ4IIzifhd0JcRnPQSNdWH9uQzdwnsWymr8ne
lqfOdtHkpSj1VvKzhCA9TATDnJPcpwWw249GlxX4gFc08XfEzUshHpMGNZBL+k3BT414DclZGzaA
AEzpfwpnsyyXt6A4AGR1px6eBoz03dh5aOmnsWF8VEOtOpHyCdIgOuNNaodJECLaaLx8XJUkg7tS
VRS6+m6inQbbVpJpOTZpsfaNhePd1iojhd2C1HWqf+ygeL7XPbPcLKdEYtlpo+4bm7L5WYOotU8M
pqwMsyqL6rrVIa1MelQmV8K4RwLytOR/757fWvxM35qTWMGqFq6Q2DOc0yCQGFaZqMS2ZXH9EX9Z
jqOy8mYy56bn3daOCDMaZL1uY1wFNIOfI1fuyp0fJcZCA3KzQJQI7npJjEAWTW4oH2pxxfEeSzAG
srjMmxxhASXAesVbIShNojk9wS26pGbTTTDf2PKSQKX/9DUh/O8/SswXyhfK2/LFkMsy85hs/abF
Ai3UHT3xKydSD1p8uU0XBVBHifXBG4kRZE1MIgjlL9G3dC+PPgSKCfUW4qn5XEExfR+XN2GVtXV3
cnZ5/iclfx9Z19DiPJ5Ia0SzxZt3uxMLYuwpZoxWMimNfmoBc9XzTMy6ELTQQuPEh1oKoTEShm37
sjoRPnO/PFICdC7UPH5dT9nzILDYvz3BN491WMDZJYR5YAaDKgpCFLzADeaSXl4fZMgxfDOvXIy6
He/d2TMGUS8ZvvzLdJr3W9Btk8NtgN0pdSJVdi0JDOGPrPD5izDRJJlW5xuiag7YeS26Ex4clVvf
pZckCAJPPhAzbvCt/EFnmlc5xd5WX9/eFwSXV3g/iYn+i1AjU4HXD43ue7Ar30DPYencpIIexZFk
R8EwmttVtCqJnKroeGqP8kpdzv/8SB3M3fby5hRDlG2qsPOmQy7dvFiTUM5384SmT1dPMDboohqd
wZNLyvSw/YRDltddYEU3Oloz/yScvOWszjsZUNuNlhpCEnDATFUmkKGTyEqoyDRiZKDsQQkCFF7I
hk6yNsPWbpMqnwBFx10lTrLXfczYE7bOsF38KYqpMPrzNq+g6urfn65btuI7e+DkAwcuBj3Bb9AS
q8Budsk359hhWo1XxkAVDu5T8yLUKeQFYwCv3s9ZHIiSOjFUZXEB03DjhntUP5AKgWeHP99XeRuv
uYaesdB/dXonaoPkATqS3Cnks4BhkJ57VAeckm/MHqATXeV+ZuBz4QVV3mclCjBV0gKOcRdgKpGV
lEUNgC91lCu76wJ0jLi2V83Wc+ZqOTIwuggq62RgYPdjfSLJOp3Nm0nVQFgkBm18h7lSNHEgCBHH
QdeM4dYENXfBsdkTchXCBn6uTxoFgudiXMVejL3ghT/Y3k0Xhs4Hn1nEkhhTJ7bkfQH788D+J8eI
3nsLwZhDdDPZnAU+JTcFQaIBwaOjB2799iuK/+CP8SP99YNenSIJG7mo7tIT7GrpZSWSK/LD7jSI
EHPM4X3g7qjuxYRRsy7gopH5I4dRb6q655A4V9EuGDRkfSw0RV03IWfZ5M3yDdI9bZdfHHCNIVE0
LRDS/n16j+s/UYcmG0kbMzBE7vdNyagGFwpFEAovNfu4UH/Q9X2dtLjSIXDr3SH+Q15wgILG9kKs
/X3mb7ZG52r0TXakB6cESDexx6AwzsPjRto9O13ljS6SZQ7LJ282hzkPdB6dQPaZAD9OmCbBVZLq
zDyOH+1eV6AeRLY8TklxiM29cEVu/roLGWYvU0TMvUl63QyCoHCxVFISFG9NTgyxef63lalNEmnP
ed9pe1tzwfzDwe3j6+GolidO0A6zHxrnrBXTzdTB8DEICtTCaPJPzfcgQFlN4ucTrnyzzYU75q/2
eNTvFuYyKPCr5/DEgfYHPKXbrf+t+MeeJXxLDk+Rp2zjJZ7ucrXLDTHmHCq1VhlYOfXpRjwQcH8H
vHwJDqV/FolagaMK900FY1/eLi6JLu+tYgHNkX0TDHzBVb6oCVRTOx+xdV6T3fpWrgxB3pRyhb+s
zCmgEja2NUVhBFLJrDWKvsKz/9KGnGO5MU9kvDbr8zT6zxOrgAiJBBve0DONeBc4/OxnKlUkbcog
VOUTeWpkjsjE8av3ALeHyVWaBcW8BevuxezD4/ulqUc+2t9l8W+eDQVcNILm12DUwHASSdZB7p5D
bWpjcqJYttVSTYijqUPlH+BZJgPQglE/0ZC1telbuoBB8nQ3oLSvI/8fkKMUivFEoRd4f/W0iuCN
Iml1u6D0DoiEwSlnULEANUOmfHykPXGxMIhNZK1+5X4XgUm7p/TXcFTtkwE8sIDGxYyDbo0X8Odl
+MNuHT4MHEcBg2+a/Pbyw3Qv9OZJ8F/R2Gu+9wujOYt158FNYgsGgQHSQgNlEZYh6bkDzHEyNj9M
gV2O8rvF/E9YUEeH3kSi4JekFm7xUTJRzB7ZWcRo5Gwx0HtuNhKT6g+zLq7oAk3/asOFsV/7YlQK
JrUUo/a4V65nijScewtZQDCz5gE20RmK16q/kjni0rR+/QSSWiCaGIftUnARVT/O7JJzYCMbBAxj
kYiZ7/GSXxYktG04wLBhVIsWoTjDm9bnbZFYeyFlshoM7lUR/PPzaiATD0m8d+JMMiN4Wne+fwb8
tz9RLN1JCD0gMaaPA0CbIp1TDUxumfy14CmSaLalBsLmCYcvAuDrzLILCYOjZp8qAdyjZw5yBoM3
XYQ4vRrON6t4liZv/ZvJEyagTR3fIGrDGF5+TakSK1uCnOptYR+K1k5zGhA5uBhaVj2B3zvBixeK
FF2RxQ11CCe5TkYuMOKIMJhtfAbLBoDrRrvrK8V5c4Nnz522xhsGgw1yaxvHpziwVydaBMxo1UKy
eBkWdbHwwiVzYCye+OGaXq7FS0VVyF9w/lgEZJDKVp4yRqBiBPrysBgENCCRqx7kGJpbYP43v3p4
hLzPn26ONUplGdQsGnKU55sV8dPFCY/tfnfqiN8Vsop1WoSbHh0Glu5Rb4M5lbthedhwirjj1Dd8
o1j5rct0zXcA6Oi7NvbbG3GluSo+R9fEoX8ams5P64AVPq/VeP+CXkeJUqEiW57/NfU/DO6G04CQ
4sdNMRNKQWt48E7+pt2LP9F8hT6oYNFd2hxpxVStL1A7uDw3paivaO+iqD465mwYC8o6aFiF2Opw
FBDXWYlRYEZELIvKDCEC5r3mjBBGw+/l/mN+NMtPzjiy3loviUwnkLGDzzLA4+WbydqxVVz3mwJB
34sZ2WrT1YF5196Q4kjfRuTVJ2ejoZeq28se7SDadDC7jrfYY/dOIBynp9JPFYIZxi3IXq1M0D5I
4MdpZdJF2ryuIUHHNaebNIVxhYC55e9yiA2o5Vs3b3rkuwXSa7G1WaU3V8Ng3RsPO+FT5nomrlVN
c9JWgsdU5pUV5LgCL3hroLvYCEz6p7n/4rdVwRo3T90EHTu67fhj0eskQNwwjgpvVqepEs6YAu8q
G6Hewja/9fHfZhqnpgwbT06Jh5nhcZ722qCvZne7yMxT+w57ehEw/UPsCwIJouhw21IKmjwlp8w8
he19UQUrQHSBLwUi0nHekxOvpDqkhKrkBCET8nm1i2C3JMToj7OiHMtwKVrkJeDIOfYnXbKUUIbw
s44G6oPYGewMMZLcBY9rLt0Sih5WPE44/cv5j9KojErhrIlhokuqCfeS1koBJOvA+uYIHq4rGYMO
BkNMDelFLi6TJ91vFLXc7LyVvg2ACRwxsE8dBPfLZvD9zAsGV5pBbxvDE5+7OyYvDgDoBzql2HF8
idrXeejUjqqEULW9XVv5BMzC9fM0tDRy5b4gNICnZ0uh4a3yJdjUmo1105GGa+fifp2ajDt64lGB
tVPMv5YgmcI8oqLgFBYUmr2F8YRbVbAaIeemGeQx3D4uqBURGpZOzHg/3k0woDWuxns3fP92yr5I
pXdrFU0BUt0kPzhdkP43bH3lRwHZRtb2i7joMZxut6WreVpxnZm8SvVD2yLzEtjnnJXryn4iRXgc
oqtkrNMUDBrtVgdUcQjfVc0SuMSGziyX2vu11Ipj+ehA9e/gI/gJGcfANTGJyQqlp4BE+C8JAmkr
7icM212gqdkcfm30H2BGqHpjpK/fOY+LTrfy3OfJpEXNsdd94cTtQc3CMh1NNaM/HSjKAACwOGla
cw8YcDk8rffnp7v7ZJnsVLtA5PbUi3oRIszsCtmBFgyINSjS8YzO8jOMlUWUIiWIYVIiFz85pCRP
ma/9PG4nVNj/aOcmLz81Q0j6AUEh7BAGp2QEU1rV4DsOwJfrbDrcH1zXgmUbC5i+V9P1Qhw8kTi3
OiTpz8QmN8u0gF9gy2oeg/5+Hsjg5cauxXvV2PigEo7gor1N92MDeCiOGMux10ljEvsUt6LQADw3
4of9zQpAOm604g1GbkkZgi6P+zP0Nm7/cYpAUpa2a3LqElUMYp/rXXI9XOAab5KUxR6gq0FT6A3f
p4JzZO0FgdcNV6lbVjTMgLqcx8NWYAbKtE5sHFj1tXSYKEGARZ8t0hAiGZkluIJCJrN3lEnfNIoj
rhNQIRrLxUsdg0uurMdBvBH6FHWYarhmNpne3kNWrWAXM5ipy/bkxu5l/uxAG+zxt8rlSbCNaSUJ
coTf2MrHhtBeWLCW9+OC4b8Yj9Ue7Vm9swMFCxCwutbbjiaUF1dRMcIHOkgyeZXPcJJZ9WA6gDQC
BCSM9FSc9BXne9Atyhiez3oj4ZhlaktcYahxqu1G8EWH34i5UlpnAjfgUupD+rI3G9XDtH5idVdE
AwlTd4D6HewAJkgq33jqVJsoDt4S++MOaq7MuWt/Gt74QzmE3VsiRuU7m9O5qoy4qNbkUuR4hcHR
pTltM+vyPZ3s0K3z84uixzSQ+sFn24gEO8reZi3HauA7bNWtQVRXEAA/snwX0Pdc/H+Fte9Oz4D+
VbNwl8WjKSNN7aM4nDNSnyD3N8J2u7X+gZWUfPC7ev6eGJJGaV4vz5c8jsxn//+eirfKzDGJdW2U
MOHVmLnosxjIbRBP2O/iy3RTzHfl/XTOudAi8oPx93brSdVpMNK4vQ==
`pragma protect end_protected
