`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
ZZICQMsXw+5Xkeq7zVzUSW/PWDSV5fByr9BZ6tGIPY0zC9F2ZKivwt7dS5u+V0moFOUFUAZLg9OD
ktcuuwhwTYcwgX7b2Mzpf7u1PVuDe1U4D0g4UOceIw8gpMbcfN2aDJ+fNCKUVECmEq+tUVOMXwtI
alZml1VusGX0Ih0fvbu2dbDgyHUBOhuVUUaZVvUOeIAE5GvCZSUsIqTLH5cIEBX7bdwR9rECBLKQ
JEYsqttzZ8iLMPL/FggtV/qoS6Hne3w201PRRnz1Cbu0m8etJyetbU1Sp2oMSUAV47JltqN3O5ek
DbEST+7HF/JFehAiPUhQ6pX4Fi526phjnw6Jsg==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
IzRErwiDENDw5uQjaYO0V+ki+jOpDsca21Wknp4F47vZ9q9boW9PTuE5X91f8EPnjzv+OoCjEwV0
oCSvJqedicap/PpzWL2ER/qEsxrCPRi7PKyklZzv/e1IlgiHIMpFBxAmRYHJo3M8nqaB5B0sqnlq
K8BlmNUAJThqAqpG/ac=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
Sd82EFyuRSPrpxaffmd36qiganOgkNx5/Zdw1cyMeYdQQ9aJItuYRokwHrOho7KRJgbQSh54N2tu
Y6TQwBh0eYqPDOwStW3fOTjfcCyL+zlb0+Tvjv53DuN7anwuiIqBjyaiVzim9EHJJ/QpezLiRf/7
fKKlhiKtQTPEImKegRU=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 37184)
`pragma protect data_block
8uCu8Nv6sJSgmfv5qjfgA4XPuEnGEwl9GpR9S3phZz/mVMPtStkU9Q/K8TqNES9RqSLN/vu7z3ZJ
/K7oZvhEKhkhTNVAqueaIvfO0mlKy0ezv9Y3yvVL5XouMvIpSeC+AloATwIVjP80ttYlJSHOTLOL
QRnZ/kMoBQ8AFd3iCN7C3iuOM9uBRoAHMjUdKCe9XPRh36FnI+9yB8sPEUDJJZvQl8j674jS77eY
mvuXV/kGQdM4XCX2kHADoi+Tt8UZq2Y0u1aQ5/FgZhjiGksysj8mxj71LAskLb0n/VwVo+YtZIa+
f1BPFv63UZQkctUgPlpyrMvP/cGXwKZX6BmwlfUsVoNm4eOGODUU1AFDSX7cu+edlKTFghSiJacA
ZFnMgveOFZhKUO0sNW2KtA4XhxODq5MKz7IUThEWDMUnDM5un58TbbFaPGa+wgqWjE4XQv3efaPu
NhNcGWEXenOUo+NgsNdVTdfe8yhkd2y0ZFgMTiH5oSDIAFiLrFp4VP6dtqBQtg7axHG070xQMoG6
Cnv8q7agYI29Lxz20yzJ+O//tYgTW7UX9ySYGBejM7p+/16Eq98jJgd/7VlWu5UuFwPX8QdHAQ8w
Q87VVqrYTmE+/v5m8Zw+l2z5zkV2dNnA0az7gIR4/JCWSQf/Vpca1WN+SIwaTaqVrwh8GjeFO9q/
lgvnWbnCU4F0enXNkTT3Y0/0DOScMK0E/NP0aan3o/i3p2PpBpBYwopgBpB4YQF733YYYmDxOwOA
dIxY5+fMGWb7+w50Pk0WKzOFvK1+mnUaDWGGPtv5LrruDtXN2fqlbQADz92raH2T7vXe9wRdHg/e
bOf4Ol1Y4cOhj2RTisxqR962QbWO6hgBU5Q1BBJFbBVmu0AMqCuX+nRddyaFA6KjVUXT/mTqGhDS
xg5jICsjE0trDTVliEfYW2/ZP08wCYlofuuJ45j+ZYDnnexPk8TZ7L57bbJUaDItcYvrI6zjvWzm
4nQJjS/jmZN5VWCFgQGN3gVzNnt22C5hS3e6E2HMtRGFrpxVRiBLg6mSo7gFLJ+DT7/HHAn0NloI
l8LXhX1mpyI7zGgZS518qK5XMcIK4LhR8xyGsntdSJ9tej1QFiYM+uLsxwlD5UWcxP4AaALT7dHG
BItwuXXLwQ5AMY3DkaVTOr62MpDpxkFsvd/E2V0gpepPs/rXoYdAx6yL4v7eVvCACrTO/RcS3jNe
VZjDDvzIGiY0+vB4Bk9c+GXqpT82Nx3vkYCJntc36dove8DTRJ96cZnNzgVHXv0AH+zqSoQOE1NB
tqAwq0PRIvqLdHObG5NhC4xEMZIvuLs5gN9k5IcF8wlQImQ3DdP9UJL+AR2Kyt9IDf5WSyC7DgqC
3yBtSN+gTEGgtI5iIwtwlf8l0Q3SJwLHsn3zH25ExoJKcewQhZ6jhcwld7YdUEeWZKwBtxoE+7P3
GN33GZTYGo+KRk5raD/Ztvky4LTejEuhW6Gi9D57XHbL0H+EUHZXNNBGS8MBtW6VMVCdyQkFtARJ
pMHJXidgEsxfAjobMoj1nKnDN3ArXCShrLd4tG5ZwVOruZ0UAdzl5ma5eCm/F1WAiwfrSZ/V8KWo
OpOAOiJAaryl0tV5Vm5NQMWdwk4HinRFUebTSSTSOsja/tpzM11bZ4F1DZasHMHihqP9fa0Ugd3b
KKBibSJUI94ssyY+E7zlhHPvPlX+vdcvXfNzKFvB5LQzIf1gREt41g6juafZkKk9h5xhV+GIENQE
0LEofuCL9Urk+2lq95RFfKloWpHpiLh19sTvLRlqOMtDpKh42aGjpufu7tQiBNIfi2vxOTjqc/6v
qvvNiUiiMylQC4+1bFigRCZF83wiM23Top9PbPe541l1CujygoB2iUOamFr4vcCRyTOK8QV4zdPG
YauSgkqLcVawGvTaNSzi/hj2HWdiUlT8Nr6E2PryiHsv2xEXzew9LsLg+3XpaYC4g2Jh97kewTB2
8wYE2YXKxIuUn/Qeor0S72rIl+cPepQwHfg/307OMgKLVvkVpuEd28XbRCKiJd4XQBr3ws6RIF7M
8eeWZaO06LTmxP13saKSL7bjWk1DwxEttlUzWm7ImqHI2rEKx6EZp0HwCJZCbbzGr/vTzU2Hr0tL
4dD/6VwmmuCUE09d4ig0P7kFOd442wj0Axuj5uXBh4Xctqd0GvGCJukva8ZhXJjNbKuz7MfkNNd+
J/VSkDVjmVUqEbXw1zVdGouiN5IKMiTIQHObyuiuWfIxYqMhXcE73awBNZ08yt+FZVntNA58e+Bn
PgTDZtw4X0NAF82DRBHnsUXp382toCN/kSwQS/mMSG6ZxfnK3vx5mTIuKYMQdfHiHtjZqsPgEeJs
A88jnATLRz4Rh8IeBa6DPCY+SrHbdngNe3SmwOqnL72M/vroFuPDTYABeLjU9cq2uE70wG0AtYon
cPu0P5vk/rMAA7pCDlU+UIKEaz6KQGF4XN2modjLQvY1BQkv8frsgHDdIcuoCiRDt8wGOh4EFIzy
l1zA7+6V2M3J2Bj2UpsQW2shwaJcfmHwQoovJOmt6P0kU3Lpin3V2QAGt2Kl+XrIpz6Hb0f8m66d
JEHM05v9KpUZz4yuijtTOZmFD6+dghCyg4vG7DCwrlbEf6ejAY8hlaMQdHloY84xhgKsXKmvi7Oi
eeBFeO2aTufcyjAHKTS5BUU12eT/cVyh2p6x1J+Es6CWujJmqCx+lC3fDp1Gm2Xl3VbHGWZ7OmYl
QJ3GQZyCOjE9yWQSkMbA0uD3pnATaX6olzvUO3JoFCUCACTg6IQZnmlsPZHoxZRprbC/FnWOZAI4
tcLSATyZcTIW4puujvkqA5Grs2wBS0e7z2Q69SdoamCiShH/o/NvRHks0BPwca7Nvr3BtWU39Isk
5fwIAISWxa40NsrylzoFpvXo344xMaO4pDxTX9x0We0ebPil7gsgpRuJFl6oEL7zRx95dAZ9tmhZ
GqnwStYBNk8mDMaSIfY780VcjDqXoCQ5praclcKTZCqdCogFqeICg18N5ooixGZz6XYS1OTN+gjK
x48/zoRFtUUmDKH9irCMmKTPLWllC29CQVIpy2AD/ag1k8bDnu/3LZflD109pMEZ3YTMxsP0RCeb
iYZJ5UaFF6DdBrd43FSsmcKJgi2aS/EG7COICcAbiNYx4CVfoIbZMWqGdjBobZu+JcPlxJyq+3vN
/aPuzgTV0jTDrk/jHSdBjF3E3luMWpIUi89NOMhD9L1sBneA0ksGwOHT8E3vukGMzwVRMz72bfl7
1d+z1y3Ieq4p1JS6D+eN7XlvelqFOucgzJQGV5Agba3jdqIE/IVwGU0+Bu3A0dGmY+xqGKlVK5Bj
QU1wZTovuIEXUS/mviRxAF+RboBq0SjEbQJ1X5mZISTdNmpVrcFWns3Wg080Wmqnttzteh9p5PPa
SNu32iOw1BKorCWK17m9kXb+dS9Q3+D+f8jrPS5cTWQdjsrP8VU2X1MWqFPm4wIlAfA2u0bHgMmf
YoF4sRWZdomZCrc3QSXMxHCOCdSXa5sD/2awkPhdRGzhSpNeDPN//UrLmpTgyUnj/zU2653MZ2V1
EEJQzcHMDrRXDBUKZdT6dGsxcrsrXiq7AmT6UQ91qhV3Hm8VmmamASTSfc5fFrBfk/yr5ekSRCO0
cHyKXun1qIcRxoVyGInGB9DOVvFos4AMXThj1jgiDE7c1DjM7RvlDpZ8XTpFf0e3BKV4q7k9as0e
xwRObMljvNi0aJRYCfBefUhQoswQXIIwa5/wmY0AO53CiBEb+gBokNH6zA5b4UtdmeS6NjOq6vkm
Fi/ktcql+i47H9xV2x+K8Xzj51Rz3S+cugZAaHetb40zKdlZ8GypV22HYx7jFa2QKOXye/41kS+B
itS1sd/0UhE54ic5QuEGGZ8bnreRrYKUble4H5FEaMrJnbMud9xAD1HYI2mahkF3roy9jhLiXT6U
Juv1K7pKCGRBLJZVsjVIrvR38FZzpFs/WSrGcShnlH+SPJuJPn6o3clZx1lkiBRXJ1CfduOl5Tmv
hlJrCZVog2s+NK633kfP4qvR0bxCgLhs5m2pqUlloaJipWAXn03nMrvPE6jKKqhl/mwNVCJPxG0c
vTdOVhKYTWCfNUM14rVZ3iejAuAleqcL+hYO8jC7MtGWT96/EUlFPji+hkE+D2n5GjDOhpBJjGoa
BHVwLDitbn9ZW/rhXQmL6fYWl1L+uAe3PZJtF682iCr6Px0XzV1UbVHKvaXRYeucXOdI9DIqKXd3
Jg1XDVDk48IlbcxF3HYCfmrJ9JMB0hdNMm+N/kRE58/n27KX6Hu0KK305o/bLmBqVRpwOIry/dmW
QQ0e6eClY3jeCu3LGX/n0QK3RekyPufnLrkvJ/tR4fBRQYtuzqUKUAp0CZbv4ddIaZ/7RA5h7oER
9+irqYpkU+zPmIwfXF9gDfSyvDrn1p6RMFEzxirP03fLu+U+l0cuuZesOCVO6v/qXtG8rFs7AAbl
+D3QdyD2XBnWSWaelDIRflDLrAIQwXl2PsR/53y6fKgqLnr20PwITuNw4VJKjnFhzLiPA3dhFmux
gpVuQMt2+V0eN8DlcZbtt9T/YNnI5GUu9F52eAb9RASifPo7LPLgbO056j+KG5l1CfvpAlHAYGT6
TqutjHmwmmj65STkBni0ntg/V/WsSMeHUWhKkbCoMfVig7HK9b/Vr7+E+306pEW56mwliOaTnf5P
qR+T5opYRg8vrlHCrEKM8jHWX0UEyfp48OTLy+Ylh1HQYGawMa+sOM/GAdKJch7LQy3Z9FPkWjYT
sU7HSDohFuk+VZxGt03d2BZwdHUhRJCtwFjq+g0egRRt2UlaJFwoLypqjies/me4qdmJzn1SsH+z
aAljcS41j2maizRACqEQ8qCldrqCn6yKh/B9BduVQLgiDj9af4Msh6ntDtuT6qqPJMRld0uJdlwg
L08Zug8VIsu8EhGBqs6vU0cBqT2PjtNfWiHd0neYUDtSHNfX4/Mlz+OA2I7TCr/alp3aYiuVGQES
qNj3E62PjyF+Ias3RnMFtsjhFm6y8g+A0rMnVJPKAI1ff5WXGVnlFCXqVyxY3k13LeoFb3d9HvZZ
iXF78VCWBdLZx2p+3Q4TZBI72KZ9T3Rx92pNcafKrqRmn9UXCgQfIjyDZSfCb+bfMKzzdpR5TO/1
Uqom5IgtlOnCmLJCdbj9d48iLT4mPKoJ4s7j1GAvdaCboaAcc96iw8IrrRU/dkTNbnElHv/TBsOt
e3iHzPGopCrfEsP8H6glaD3+ABSoHTGcXmkvzKN2AIvjRZQoF3FZ8p1pxFsXRZmKrYBnx8fo65e7
UrxQtdaZJf6T0I4D7U02nfqThN6yN3/Pk0IToKcgmaUQVim4eIAXt/SHW0Qhc1TVrlmzQ0kg6jSf
Wp6tqrPUFexSkLufGEIp1yP/r7TtbncIoI2lXxKw/MF4lFkSUiVzouLSmRINHhCWw2X7UV7hTDqb
PErX1N6N1XeoSJzv+EQmCdSw/A9f57VjCuubyOroXCsJsZSJZAoCm7wsQuptwG9i1wqxqGkc004t
tC+IsVxBN6ulCOccKiuzEQMpGgAs6IARGjedIRYStpSbWDQkGXbn9vG2n/G0K2bM27D8JsZ17CEC
S4i4qSSLCfJthPRZOnfXEp1M007MqWPM9yA74dRw7wOw9TsrMyZ45g5ULl7vUAXvAD6hYjYaVFMf
4/225J6cTRBWb+rtORgSbEjQH26/4DJkns7Wr4NHJrpngYin+q/ZkvLkJEE27aEYmbjzPA4i0YGo
/P+i+I6FMvxKRmovbgPcaLSpmt+TtFTZtOL4Doy7Hm4eg6SJJk5yg42Y58uDJpikezXrAHw9MXuS
dAzvZgPu9eCufdsL3B+CbemgAr5UKyPAyvanu33oxY/re7c7PNGOZfMDNqWxv9Vm1G7E0xGjiO5q
HYbotsKHvzNmal2pvpwyzPZfVk+hVlnGLbRrzT00+6F17yOzrvx6dNcqGtmbIv2PZ0CXP/nVAP+T
hcxM/lsBo5SaTY6FSSx3qPouLFfmBR4e/tmJH3Njq+697DSb74o7i/Z7btjZCRWUoJ49HmjNjTBl
S2MwP25ZsGeieSA1MXZCP4zdLHQKZ5yG//Y9xBtICqIa+rVU/bCCpXdaVpXJJg/6DT3PEDURODn5
Nf03cwX5+167IfCJYvdO4W2RBuc6mspq62k5TDsg+tdVNoPydH3ZVRLkdQL5wt4At5PfTYSW1HeG
JeUGrSYO0Gb2ipFmNXaPeX4QcOT3DzwPp2ZcGUUX1WvAGX9pa5xR7ag9hDXFLNZkBSktN1t86Cbf
/X6pR1jUMt/kJILBHs8x9+oJJwVrPWntDwT3kvUDei4zx22aohBUbJivM89EwyJqnnBYyulPnRv1
vmUo2rvercYuG0MRxft3uaRfB1Uk2lr70/nJ3gzI7BDBfOrj58J1hMxF9M+nUWzmlRjj+DRwnwti
WnwAVmD+6qvmZ2oWD/smRFL9gTREFAPwzsnRQS3b05sZxrPFFK5ejpoEepcn3LrtWuTDCPLXwVzm
2JgMxLWgSC/LsFPd7nXHNQ79wil39+1Qsv67hi/70qgAtTqDo2MzVaMi30hqTaWpOVQuU5LWh3C6
fNn9z5mjU7rFSdoA945dYVSI35+36MI3pPKgts/FXDPFHmRt8EXY+CHHoOEPOjdOMr0S5pZJPqpr
CXCKBiCImG6/cXAiBSmmTiBnBoQjPAzNJbkaYVQxlsIUWZy8ABKNcD+hNpKHQjfMFyMWDznmJpoA
U/gXlccnBvfLXXd9htczbbO/8Xv22YoumKpvYVNLeTGSyFZoLgLhrC+fklTy3+COPk7E3o+y3Ctq
643nXKxboBAvIPSYOTxF7m6xq+3qvl0MJ9j8n3ADtgFsszRnOonVASH9xhyADm2GyhbMwA3FbUb3
Foh8I0qplly+qgUDQcD8Eqo+fgUNyOjbpGBeqO0fJdyoL1tfsaZ79WfNC5UBFZKgK2ThNAWtOBPl
jLQ0I5dMl7REpmJctIRZhX8TSMXpFJpczCyXkQu7n6oNPtX/n2xOmzC92aBCtOni6gmSHytoYFty
baIKnMFIyV8MOlTokQSNo/IgGzURyPrslBxdDgM0bi1L18yQONdoNfZXpzszOyh/O2/BrKUp6CNK
MWmSlOInjbXTOEqLuQJiW3tcw6YExPLZ8ZhC8dZsuJUP0SNiKyuLGrGFeRId1QLQ6mB3iS8+Obu9
xvlcINLy//cGc3p7UknuQl6VHJR9/qyfX2enatGeH4c8yY7NDgZ5t77RRGsuk8ColWN3yussh0lI
FtsN5rYbyw6qpxqCDRDsRJa73SzOVUAruO/Svdcbj9zdmG3hlbidMOxd/9SnQi8IEktQM+4lU03W
Uf/EjPRe7CtIfomw4dvRrfNYdO10XQD0kHOBPOZT5ph4+otyXMiFtvr/M38Z+HqUkfixDeJ6i8h3
khCh8nRTWJMz7u2iL7u1VAToUETi9XstOGSRC+Fjg9U2+MHkmXb75DSmL12MGv/c8gdXFBn5Ky4Y
vhByosMKAHz2BIFwWjIz91LpylbppSTfOM9T64v+s+3mSgBuLbSPvM2wIl82IQ/hyyhj3iWCJWrI
TBbPqJwBTFHkWkwbN/0j1pWCddjUMKrz2ldFXkTeQR3jb6qweQGHlzvsB2CQYUFlXeUy7H/nvzMQ
/kB8NyRKuVIuL3hNIoTXp6DwrYA4raAWc3TDFFjE6TRSWjMmQbhaOgH+/gbSc5orea93/syedyPw
TbECgLUxwlV0cHtoRAem3fBYiTBzZQmWcGQOCiB3K2sR9j4CSFpdw/5dZQo5BawDhAc9ccj6a43I
oLaI/2GTd6bIlzZMNM2YsAWd0mX+6exv4iwdyPZfUUc2NpI+Qq1LaUPNKzyeX8apWu730ji9E+AM
US8qf90pTmjmIA4d5qvp9h3y5VHjhX2f03f2/zkT5qYqj5NrnZY9bAC9cfI7e/BcSN68Ti6T/mgI
oA+bC12SsD+SL0amL0W18yNhUNij0jXVcv2rDW5p8iNkNuLe2rPWUJiPaDsslZLwUkaN819MkBJv
QCp5QQxh42dU7aQ5CTvm2P0BsMfVy4WqRkjwOFVZ8BCysebdM2COFs459Kpdo8VcrcuKqJoqCavV
9RVHWXJGbLFy6V3fnAFlKokPpVbcm63IExcUu3quQIT6ozXROQY5wmQ9s8SCQY+7EUNvlin2aDez
hFFTqnuU0icjezS2HmLhOhZ8K62M+S2SW7ctcUT7R28jF7vfBUSsHHHmeZUQ6LJK+qbSK56kDzKE
4IERfMq4Z6FAhwoBIPSlEQaL84JXBZMd3LaoSiquAxQswKWyeJaTdAY9LFkAYb8LtHgltxseB96q
RGFyU/f0iYVDGqVIhv5LzoHwdcTcfmDP7ypn8chr6xCIFjNdML0StCkxsTQLxRvZJVt74nK6QXJu
pB5VVI6nY8ffxsr/ekZIvubDJPYmTEXKCdrTkjGiKV5Pi8tEDnaYkT+gyoRtwH+6NzJSqHRpWs/H
FQvl4sbt5J/GFfa2VYT6khn8YekArYbelpx4FyVEf4wNMv29MaCCWs7X7ws7ww0GZwRXj65U58Ku
ya6ZOp1r6AT8pwfaKPZ796Xh8FjucHQS/uM+CotrWKc4ZOfmiXItYkZi2ocRq+q6qlaWB3wDWRkW
xVCYh3dav+JNyBxAz8Xt4+gIeQFnzV/tCMgYKHk9fuhtKAOmtZtE9f4NyyDF054kWuPsIDosjmtc
Z297dZ9lptPa2umM8TKhKyeN9++qhE9BwyQeR/Dee9bC6S6dW3s/eL9f8EeUt0He9mqYphE0VAMj
2bbK6liPSaiOcI7ui4P2NoyRVoqNRXUBclPXnVK2V0ttz/TY8THU8uVI6YXKD7sBfxQDKvy7bnWa
P+jL9sZ/rpAE+iIYCnpH78aHUgupM2i9M9eXDMS1zvMAdedB6Vyikz/30becQNwmKi1lNVfeYp9E
PuC0mNNChziuQRyISX9iyJme5q85fjhhB3ewmeq0EaSzJgivHrEisnXk9TAqIN5iY+2nR5b1CRUv
K+DA+CEtPjuzwXXwvvUby2kxLVuyvEf+TndkWLZhwqMsriEnNDH4gvotozapZ9caou20jURWoNaq
fbU0CI5Idz/W5km18jxukU/UkmaDtRDlLJMzzHBMz+yvREwqLXlxq4lpaqWddL5jWrF75xzLyGyo
kHhxLnKgDEuX+gXwtcbpu6OhuxqcENaQdOxGz5P93Q3SNkMnebId4ashAwwLi+xl3rRy6Ln9rvdv
tEDUDOjQ+Xz3Z4eISB/+hjKIrivHyRuib7pI1+BbhKPCxnl9tHxiA7KBZhUhcj+U67OZwyID+gso
f+AXJA0KP2KNcy+SOylBDxtMCDyMWzgyOxOV35e56GUaoHiSUjn292LhcVzbYo4qqUZ9MEYGj+XU
WJbiHrAesUN6T1TqYm8YVBuMaYcyqQcX4SzrqvAvKUog1QSOpLv4yLKSC16wqobFMPeWPputYHpY
1yWlSgHrhGxDq4vr+tZwb2bft2V6NTqGwS4r+8FDCz8ViO0I7aDHzXoAzJrqgSFhUL5WgcB0XbXs
jicrHKfE+OymsvtBIxRrawPWW6ZEZ1KEUUlho3ScNPxp8CF8J2+LUQesCxGT9bsqD3F2ZBtV9Sni
SW26q+MJFAEJeMUxAycOTki4vSMVqk3nHKyzH9cPh2EdPhEYpFXUF0rbFLMGm6iEz9H8XsdRYqtl
l9hNMbBtBHo2rYPS8oyyeOMqamEVdykbgrZ+fePD/raMSciVNKD8wfubsgxxo8nQ8ysKzEnIOPR1
kBVzlHSiaJrzXJLIFVIcv+qqEyW+DazkCbYIKo85htBAok65wnTuo0lF8rYpO5E40lkbKMMZeBeZ
cXcdW6W/L1e3zX+YuzaKT0uBDME0mdoGcgM8+59//gn3/CKc6RV1XEtHfygaBBVYGRWpL6X1moVc
T0WMsLVotTvd5Lq8OOSYMfet4os25BHAvTL/txDeWn+DIY/oJqk7TaTaNCjtENXg9EGM3XVzysd8
Yo4L0R/VPOLLnOXTcFElqzsQxtVWlbcNNEyqdKntpkUhxj4+abXIV4M1kVPGkJXMB0wO89KuCVvE
l/fVC4kDCH+pRmFM3vNKY/a2a9Uub/A5Irk2YRC9CO1VSo0O0pYeNgMcl8PQAuY4950arbyw02R8
/eKwZetb/8smVFptxlZFhaZfjt4YEe/wOKyuZK6YD4G0MPY8DX89jus1iYJojg4qiDUNUoKP8oSq
lXvao9aucVlEIFZSEs1pHncrOYrf+30P6txgZUF24u+TfAMIzKONNPTHHJ+smxwGE2LBPPIHQNZP
4A0i6fi5ZDEiMvm8D5kUZruoikAV+WoYgEe+tRfU5XbBjyJSgYdQBOD3X6GPOOK8rcBiZSsSTLFZ
29ufkEoDC9WsNWkoBHBTjiomrx1nRUrXcTQK01k1i8scnwqXYm6NRar48kIYdQflEeORjHFDLk09
uCgcsDYlNfU3Nf2rYDdt3XAB4zWOPe4/ASyh9W7b3FZYu6oRs6qJIrzJ6Hai6NONvCNKOB7SoVGX
Q7BeC/POLU4KJAPgota4gYJQ7Dgqm2sEcyLHXhd1ZGrm0HM+OhwAUckN3imd+IctliuNm1zVXw53
b8W906e92bfJWIoPDI8K1Kcd+QEbCYvAsb4bfndJ7LbZwWuqMhtjeXQowZkqazpoYvamAgJ3vQu7
nAFqL3Wnhwos6DVy+HTlv14dyYxxI3XDIokOoOASRP4bQY0bUVycmrY8cAyyrKKwMPdrkCxZkcxv
tdWLkKg92HnqVn9ZlES7cdS/t4LSRfqeMSbwY+ssKYKpjNOt3WAbEKQGdOsuA4sbrKZIzC9zVdKb
XqRZ4MozYbQj317mEQUeBKvm2LXIDhvS+nlCsNxQ3DmKDXtM+gZElz7HOhN3NvhegneBdDJpKepT
UOSMdrR79Sze9KgSGe7OSAFehK1QJcAPNliHa68yutXTBYbJuaiguTZjaMw4ia69XAEBPi4Q9VNV
o7eOwcdZirKk51rkxr0nuHT4oWDNT7VYejWbF7SMpL6q/sUER/qRwl7wVP9ovzHSKF0nPDJuUBhG
TP6iVFPb2qHzp1mLVjZHWb0yQIJ6BBeRWYvaP8nYXTqYxsHnX5Ew78ddlsDoCYdKC5CNz6lSx8by
esW6jHcfbz/ueTtBI5Pksnfhvwae97tgaT2cSyuoOwtS5fgrG3n8bYjb1E8hjjmXBGX2ovn+3bMz
J6XZXln+AxGFKXadLIE15CpADW9sjU2UFvMOnFFeoM5FCORdFb/2KwZxjEM5ng2inI4ES5N73iXT
oI6xLI1DMDmXNrxmi5T/2SX3go+Ry+JpAeb6BaTWdaGHnympFjsUzjJLSiPK2tgCC4qJk/PChEyA
iPRuEc5Q/lDwdt0HYtZ0v8HsmYP2pbbXC7P0bC44XY1oaQFCdhuPgL9pvGzE4gkQwYT57DJ+wnmp
3uVapzNWbReFraPy9iPK9QKg0lEWaxJSZAM23vl/sZB7DuVYun09GwYJz5SVhPshRxXaZ0KPgbZ8
ouvfEmVK51pCyb3a/F//qpdT9dEA/oWU3FrkM74r+lDSEA13W9k/sSl6MwmrLPc2xYnPsR8pkDc2
hgkFj1Fh8N75qwFgA61bfgv4ZTNf8oCbfbKqu7eobkA49j7B5UMYuZb+ElEvtPYP9BMsYdgGLtkA
TXzJqGdntbrns1rh23jfx9ZOBPsdFlfypWYKfM09w+ZJ+N33fQghQTuN+4Vmr4rgERb8YLgkkc9+
VJWH08hIel+nD8VdGQ8sO4wqmOqeu83WdkHPOGyuW0k4gm2fl3K8HxjJd4wUY6phAAdnIxwwntm5
QaGcyFU1/P62LE8TGBkwZC8TygqV9prwhXsNmT1wuqFT9G9IpUfiHkDcoQXf/RNgu/LuRcEHprJ/
9UmUe+seXLAMIUf3QBvs1nAsmePlrcdrMyRoijB0lUMSD+e/2bbkR4G1KL5UlK0qt8P9lAlS3XU1
hk4ogVy77KnTwSzqKOunsupBb9R4IiY7KWwFaq2AYKZweuRHk4QxVC8ZuPHbxP6RqcMSvumHEUc7
GA+lati2ig9qyMK3ifu9ABt+Wl+mL19xXLcwPahXCBLhwLiENAOdnhOAZqp4OXZh4vh9yC0vtETn
2pZlG3sETvefr9nsu+uhV6LojPW6gMEKQcaWArIJStlW+uOy78YOTJUts84Js4kPCIn54FOX54jv
BK6YQOggLMeBlg1goq6hDymshS/XhccaQ0d6ThPnHIwV0kHj8JYtONRWkWpjlkejnAXLTRj19kVv
xWO7koRFQHKUi+yK//GH9RyN9ZyUCNjtvr1Ljgyw+jLn+uEDHJB5090wCSFf6C78H3nFw4kqQ9EE
bDiSP9lp0JwryE+vdtU+JjZc9DNmD6JdQ+/pH1dfQIGTA+pGrGuhlMXyT1i3Xm0349j37WP44kk/
SU5wN+pUZfpwC06Gbas+kedNgDgzg6l1poKW4NzV6YHQWGNGMW8+o6DdiKtIAtXxNUSDPPuWSisk
rKYFaM3mS0rBSgMc0L5M66c3GSfCbVmKChUNnhhinZ9mpg64NuWDxAgMckJYGBPW7k1Dlw3X8Gnq
eedpaIhBLwljexHBTcKF0Q0bLHUvOUjOKBL4tKkG+WChxzYnoPchSjiYcX+Z3cI0LdaslI8r67ox
mC85xTmfacEyEFsLEftHHfx0Jy6WhAUpLjZ9H4vc/Z2iOBuxCt0OknjgFSnp6hC2ePYEd6nOSVBN
62U6nJDf+lnQi8SoxKFDeaPtdyBTeZJ4qzldBjg6oXxdMsi5aLwXp58XpyyV/Td7yZlBKOYyHZd1
Lu8hsH0CMTvz438KM4zrTY0+rstBHvIoYAC4Z/nLdOl47SH/oF1G3oXIIZrxhyBJA815eSPtD5x6
+RVaVWLFHlMAmYXPHtGfHuZIGgiMjL3OzG8PJGIc0NfK9kH27hKirYxsd74JsT0YoTkVUUu1EqnK
suBY/NhYWuyEDGDW4foLKx1kPtmxfsq/hzI8r8vErqnpNWDte5svKzTQn9k9j+w3l3U5eOFM7UTl
fZi1+e73UyntwwyBSKXwGTJ/9j7wI89AoLw6MreEi4C2/zQobKbm/HQtoIiRd7Lm8AypajR1cWlm
Z18O8sWNUuvK+Pu2NREWN9rH9Mg/I1at4cwNiC/DQ+TRPCuac+co9Xcm91rqvOZusEb4z5VkaoK+
mFtkfc+jSzXy/6RGiqmZbDw5nxQ8wotyt4qKcjsijmZbieHpzyx1wSEv5z6kpy24O1s4XLvRFPXr
FED+wwVrt8vYv6nVRILdPTg0Y10HCo8HCSGwIOUeQTueWbvh1PxBeZCZK+nfLxHRdRbP4fVPR6i5
0uJetMIeiGiL1DnJu7QgduT3kaD0J6QBBpl7f+sktRKy2iyPyPv+ClO6mepMAGZLwKWJpOoGdMgX
aUrnTpwMVQtEDenrNfFA9qLLOUlNfZkwSC1J3gn2ZXyDSjA4zB67CGHrgAYuXUBLu6ly+qtcRuFf
mROPYSgY80oyCDm3wufeUGq5HBsAcrMxJbEYQQquuAg/v2lY0LUgM6PFqwyaHlxCgvkhpsUGFX2u
znAj5sLWNrNyczvd8VKGQADw0dgGt6UbhCBjdKUYbnkfio2mJkbqdf4D/P4HZgsRJ1sAD0EFAY/T
g6zbxvmdWSIR/xJrD/LadZGYXW1AQv7HVUORhkAE+jVI4ukOpomsbERaDgbyEbZP7rCo+jPFnwZp
nMTi7iSNj+7zEp+Ut5L1AVlyJZ5une6erdZeb3sKLLKDjFaZ/F6UhB/L/5eNsC8L11y8QMI1tpA8
K+4lrfn/dk3rOOdYPWnLA4ghR1Y6hjaaHZQkZPsAAwc0AW4WfIuhwasPb3xU4XqcBWIFTRZXzvCN
fCRoarjW00tTLz5J8Npc7PiKwMbeUrk/mSdmRtxqciH1E7V/F2zlIusF6RKCyn1SKVmfXITxsB45
jVI//CIrkjz//vzz34dM0LufeboaOtwuL3H8meVJeKTGIw7AzEpDt9cWhv6hPBV5RVEvCwBkTx3v
UkTtraekGhfrHjlQVYSfS8jfFqA9ldOy134UL1gqbdyv5z666NSdxL4qj36OuDqQ6kUql3G5MdKf
ZcQkV6CQ5JJ3hLEfy1hwJQklNT2qHveO52EXRRRhwo+zLKRCD4brMREt5NLSB1kCs3t93oD6gAlg
7dbStvYfCrN6Y+nfZwurrvbXY5HGoB3+Yw1G93Pl+l3KxG+spe+MoDGPabVXjDh+CI2iu5CiWAC0
VJMmEreP55cYOSVbqTedcbYHKy0zQ0Sd+MCiZDuZ1KQC1YMsKvm87QW3C41aPU3kLdF2YQfUYEPO
xBGY++qsdCc3M01FGMAAMhiTOhyNSJL2ds61BddWbB25Sz+aCVXufdd5I8IOHL532irJLCLJErHw
tkbfTfSqj1/gMjlET+uNsxLj0ueof5Ici2U51syBTEedulv9cNeTnsC7fN+wFf809JuDmsupvcII
t9Gj9j31+OZ8kV0pYgeDIjfbmXYJzNqbfL0vLFhLGpyH6TiXdNqBAb1iVPvjVm1P7vB+9Z35hXnU
SGHxNqn892lmX1oqaMDUCB9qQEw38CRJjatWcs3DHn46vp340ryWm0ceSCnRpcycQJ6Ss/6b5EOW
hYaEC621llLiYtwQRLPN/wtyy3CQZe2pzJmKAFPe8MJ3S8T0T0nhzyz4FUWCKjxvuzSXQqDFIAan
NXPBGuc1O0tTNRnCMU2+IZjpb5F74aZP8lDuPHsAuCHOmFJEX4o9rVPu9PbPD+hLjoamTkRNKIU6
lGpuW0ILSHPJuGNq9KT8cbem2z0rBtAt4Kt/0Y/Q+YwEceOvJfJ3DOCcnMrYLtQjxHEDxe5DTQxL
sDCIhiMQDcPwvMR3jYtQV5ZotZ5KJoJYTus3a6lTsbvivpvxKfdoqUAFDvT/7P0Uy7E51Dt4tZXv
I0n25KpO91N82cVKq/3IJA7qppxv+AO0yO8SrpB5jrChMSUJ3R/U5UJhBofB1YL2epQiayboDwMz
ySiOT2EJyqu5Tzjt3FHBKhPPH/DyHPi3sWDcDXt5OD4GHzBQHJNcqtTtPnd0N8KkVjyYF28n/3Wd
llYF07H8/GsQ2nFtSajzuH6Lh95zjE4bk+WDXpqcdRL1hn8z8KvKrBPffSp/xfV2o8AmaBlAsF3s
k398kpAfkxkMECcul+bzFdv6Stpyt33Z+YRDJA14fB/6HlDMDd7DPSolGQP/YTi3euTPW7yGHjmg
rNVwi4JpKky5cEEV6/N9ygj0fEzsYICQfE80jatD756WWtj2663OKdgKeiLsnYrjgvSULZyXiCtu
WvkL5nWRIL+kJ5KqAEWWKEG7iMqhFDgL8c5cPF2PuPlu7B8AkhtavqUwR5Xea0j+udAavFUuVkKU
8243BpL1MNgdBLeEshcdGilCRnHQU3MN7Om7Md2QYT5UOIKkku7qRY5L+u6PHNf0GDpFldQW7KNO
iM9ujA2cZ9iHYti2edCVP6Wn5o+0b18fS8NNX4t9ett62XAk/IrPpUgjg57kRhRPuIIt+7dYOwD2
wZtyULc3hg9X9JU9G7FquXtnkxasNag6qNvJ3hFVwCrvfEzfRcu3ulnlsrMB9K5NduXvZlGDCfWE
ISPrxWn8ZU+H2lO+G9XpURYYLOBRoluV/AOO6C699xAZszAJ3Zk5dKU3VEw8O68YnKA3EgQmR2c0
1zjGR7ycLlgUgDFyzkJrtTmYAf91u5OC6xTq1CSmECrbeg7JXDCHv5e7cSBVyFqFw+FUXQVOAuLT
CrwJ/6az+7KMJMl6Ue84x2s6j7bsATy0a/jMymNfquGaN6uLLTxqtcZ8gi1DvEFBOzI/GiB1LfT6
x+pWj2x9AaZ23MWF9jD0KsBMoiQZ1+HYE27uI9TEqwoCmJ5zqkQb0FV7lA0BTi+O15VqK23Hejtu
eXiCyiqTs4mRCeTC6lkW94ydpH3rpV8JFpOUZGEmsWlVUQJEt7LtZdPttAYoQjiuXvgfb5yfFSMA
qIaM5hXeY4k1IKlJmDidQeWl6xve05tXSFTDJBlyqSD42OlLmSC7OhaFdOsrVag2GJp1K+oCbw2z
KHKdTj6F0xwXmz0ZotbE30ewuoXOFTM2kObnF8oo1/OwO3+oEXyXIZ7w334OzD5t/sb2CkHBa3uR
qddcMXHeUiYe6vnx/sYN5M+kHsnYHZITFGjt7LNcCiNV1JMCKNbTc2mcOmJ0KkZ3bLM/vUauiLdT
NXzFWzeeC7o+S4pBhlCpuAqDPIFpgmQjltaYAI/+yNa4Iik6SRDRgLpSWpBmGbrWNGvoDjqk8ezv
rFMdKDbX23OBQpWVRzN6tbvckxTSV+cGR4D6aeivybjrVOe3TKg5t4H42ThgmqbpAFwczUlORU02
Yf3nDwqLxY4gYd2sweOrNmPtRZaMrgUPDphYf+8jBRFOS0cmgy42E8eeK1AKVQ1RVJP/RUrqAXZT
B+donOWme4TEquD/vUZOVtLikfcAfgrpY5zQanZatAF9VFdHIwLKzD0wfswpJknVywJlNNA/Y5Uo
n8pDD/GzLAUBXlFOUWNB2vUpc7r7dTd5pJdvZc/wdzSMjGnpY7U8Bl0rXvVyZqUVaqBq7G0b2758
HYxTsndI+13xxQehXo6TMZcGWXifPWO2ppabN2bVCS5JUMWP7zAO4eXMCktdWzq8vjhtnluV2ksr
qHGaKEte6sivmdkPwGSKfXbKXH0Dorzre+bnHHh4ylQ/OM4xqGIas/idA+Nw4S6zS2iIWmMEVm0Q
jX7fgSLcCYxFKCfEw02rMqdxYni6hnu0x1oBzCT63OWtQlpfEhtMTv6F4KykuriJIT+Hnp5MfC5T
6t6UfXKPYXVll6RmP40T3WNRp2UltQF1BL1gwbGy78gySz5++wqYeiNsPW4Ebhouem5LauDP6eA9
HqLbPudVGJFMgQCGplnrd6yQSwiWC8nYEqPAuAXgUu5FprbeDzFIXzGP6vsQdXygRMQo38g+ifMR
RDkOuEfKrtEyXZwHwhnGm2a733eoEoMkxcZAkcnfU6JcaR0UWN7WyIykqFsc0P2vkJbSWMYTjXyN
i7aGBwRZ/kRAaQpg6bUgim6g4VAxMQkdqlOZXYC9Xd6zJDwY2htO0bDVw6iV/0La4DpLilNnoL9Y
vM+AtPySGDep5bz9HwY1caqvDFGHYjAF36pkZahOoGdcBNF7odvZxdaannEo4z/tUeHzf3OI20S3
YHReG1iQOKp3M9Jt2VT+HNvwEYAPOBfka+2VA/YjrJFWwmEZZFFGOufL6E18g3tzVOLd7b2bzBqf
XhpQW4ThJ8p73zOrNzY7WGU9g2LYPzZf4cBnvx3x9eEfCVjiL4V9gkVxeqfNVR0yX9RAIjqp2nvN
zSMF0h2n6MLD2jvXsokQR+jmUcaGe/2f+fOwlSrWRpr/9s316TBgBTSJZa8zGGPCFT1QVlz8AcUm
G8/TTx0XjVHa4gl6VkSxnx89Df/BrsMmPG4j6nLupxpOHZKsFYEi8Nr7trhHj92QiFi7LineQ8rk
+KvvCyWyD280Cm4eoyN0qfmFGfEC2ANdLlnf4DHLJ8VDUj0uTuv9k6O58C2LhGPkmJ0/7NqWoxYA
iqBKQk/bNT/6nJ2lticd3OrWI6YGWOInQIoVj3h1jcQdP6rbwCImNLOeIX6+IyFb4a77RlPVKpEc
aQgCqUZy1Cr2nswTyklfK7+//7WTqEFtgleMsvdE0U9CCzIPvSFAZGsVYOt8Ckyux8bB56LSU5S/
JlE3Mkk74X/9I2BAYAEqIw+h0ciU+fvrgIztE9txfIQPxRN85FoB6pBEx9GKuMSXdclPMv8ANg3k
D8j1lxiOhSu33FKNdAgo56XHiNAcHZqu8WCgaYyixx5F6hVBIn7IBt9Qw8IOac3fZHwai8WNfMHx
pSNtxj37SVwh6NZpW4pfZcRR9lC5+6LcVQKjtzRypCrFABqi54/3VRBRS3corDvNDYhzI3RbMOwF
pZy3R6Y+SAwEZBkUehRyYsG07dn4hFwP+3VQJ1gSNsmMlLLOkhCHSteCl0puYDW0g4qA5jIgt0Ju
8ljhHfbSL2tdSeXouPSSeGIc/FJpTQKrree3Jx1KpCkUHUDhBtvKZHVLCutTJJka7emjyFnHtYuT
EpM1cZZenpyasWpMYdk0Jq+OTi2MmRIKpeZWQzjsD1liRU4U6ZItri2mkSn1msl3m0cVKSOvHk54
P6Ew//wgyuJS2ak+099ZGe/ll2TWFrrtGm9sOYgZ+S8+8oq4X6a/fYAamdqXR4egFORRRy/DcXzR
/DTgNXI2GRn/HUI2PGIZnZJyqNYPJ08oztC/uBq8tGmyx8Ohai0hHvQFNcMEdPP9lriaTK34N0yE
tZThyrb9pc3vgCU6XoMVj0gt6Zxqqp1iAOz1lOtYfXsi9nN5kR4cqKIXwhFBzNgDtvij6fp0hCvo
zE+z1cuG3CRf3yxNqabk7zyRSjG74RtrMP8/6vUSVPnq9s7MqXRHB91U8S/++28rpCnN3q0HdeSY
k0yR0I/v+YJVz5uQCbmhlm4U8SSDvnz9AeHg7ZBgOj1ibe+otRADwQz/v4LztLFmDAyD5B8JxKf1
OtlTbQiG1n0hd/i7aYU8GtHxfBE1wKEXiUn4/YRqHwteE8c1N9oF+q3h2+7emkwC0ZJuCG3Ma2CS
5IOYi4aAQOjNfHYxKJsI7owon/5XSxvj7RMXrpKq69BeX/hHa3E0T2YpAO4arw8VNf3YFbKCEzel
jR2NINHq2y9nVfdGTmpmpWBtrBbUWX3qp4tdOOHt0XJ7uNaMHrSFhi0LlpzyHsX4QVflX0m9MeHm
Wg0+1bRSJJR8DQfHuCesPI5098+wIG0+38qUkdKgMqJm+zsXj8mHuI5clDp9V3a2bUB+QWBuvtVr
I9wqZsVRVV+eMgXd52axxjmXgqesmJrEe8efRaK0OnN5nRdmWIrVkyrkft3/b1YM7lsYoaWAqT1H
OwHTtX6xlzzZNqiGS9C+toV85wa+icXakEcTFxLnJLIfcEIviHA70pt+FHaITdwg6ad7Z9UWnVW/
y3di5mdyR/lpiepsAVNlhzLxQNYXLkmFq4XH8hbTwYp4UKydnP/qv12rUJanVFyZsvLrjxiCUeKC
x5vB15+d4AEx6UKoNPZVgqrw0mc2Tyz1vFqrUU42KDsxfaQSjhfvSLBgGPAD6gXOAgvw9QFBvrsi
3oqi65cygr6JT8RlMZaeK3Ym8eVLUl1OHXVg0H3pq3mhVWs+Zki9EznqlFO+995s8rq9AfNQMHJB
9aHPI7hISCyzkKt5aVqrsVNgKxr7yo7jsKSLZaYnHZLBViFoiFJdrL4mP5hP1T0pd/Yg9Be8e4g5
sBDjJ6eUrE24F7I9XkDFIgfqQIivLUxm0/zgBTWEgBzlFywWDWzHNGY9oe+6DpsCoI0wpVjUfLCm
Up8MhHYdRioJ9R3pWQwVYEhzqCrg7BF3LGMT0O9Llrt6BRJEII1ZvT9kQVRXYrWgfSMaObmoRgb1
ctxN5TrleQI8xcMD1yKSUAeb+KFFLhL/2DdLWcopjkEKWbv33qgnpRQhZ6GTy02BYy+N/CASfuRI
ezmePqoawVnhdvXbSY4g7dL/4NiEZN1oLeLBTWTkR/vSQXrDEYGO0x0tBlSa9u62UDtVEQuvanmd
scM+NtVmhdycDtt2oOFw98u+16i686Ml5dlTHZ2n+kchLCDH8yp14Ra4v6ntBosg/mVfEeSrcsJ/
oZohD+oph+cNYEnyWDhAUKL7X7x5oVtY2XKz/oGGN2kpYFVZmUO5dMNh4vBnEw/m7dWfDHWAiubO
+bItFlNVhcd5RsmXYTg/uANkc0weHpLpEbIhqB6awRIglyR9sMUqTyMRncMhaFCYbrlqCuHThRAj
IWnKwgj4Axt7knticyHKVGMSSKejsqVben9eP02ISv99TvMYpWsQZe8kuTHBaWzsRGxLYYjG0upc
wNIpmgpI9kUsUcHe3e5TMu3eRs7nsAINXv8YK2myF/xPdroS0KRU7knDe7f/tFgMXxUYlVvXBLTY
Upstlwc2WuMtHZ1ogDFbZv3jTk6FPZTNt7PUELlcprXldubddCJgGhWc6rRZhe0+1o8nY7iilVLf
nWJubDWYBbg0SbKfQSU0n2KTlaCyDaFKXvNz2NEeedhDvNTBgxuKe2dyn/noNdJoQ/Y89MxGqbNw
QVKl7m7ebX+4p2AZODcYOtNccRDpv850e7Xyo8A2c8jF2JKMVjS1cQqRXQwj0EmLG1O60UzkwFdr
5WF486nfhn/Yk86+euAjkwDmACR1M3/H17B2Z7aGX3zaR+OoRYvRD0puJWrpb+9J0UbjmfIn+hu8
JuNoWizN/wweuYMDJQxm3cPOFb6zrPpq76VTAPoVtJrNri7bgsFPmX3GyCG+SAyV3OFDBvZBjB7u
u3EiKWH+ym0XqfyOB20UFtw1rJg6UNJ1CQpAVKmMdOUgY6RZi6pvXZ+ieLl4xU4uANEWYz03YIHc
33M9yrXnJOGiiZv6uizRPlN/v4DDYytTllk3QydIiNbB7T0QMWE0vUtYrVJvbag+hRvyWm7MjIid
qfw38C8k0zYexbMzryNuqTAbTUFDb5UV6XtpQWfazNGymIns4+Ef2WDsYD3TNd4CPezBJMzZdEy2
RMkTqOhPsHDd0fFjn2va9Ags9vNoBRnTcRnJkMcn50Co5QEJQKgFk/NcbIGIk+QnkF2lIYxidDJb
h+4MMZfLuYcOyQP/e+46OpLvw0LWRx50nU9/1OrgpEAwaGrwHy9GxVJbiaWv0kXeJsHTaCdsGU6k
tJoKTPBAimbYp+Y2DDF+YgdVQbGCkRohZvlFA/60fA0ue2HJNp5ZquoKo2zDOorKwPLO4cnRoevP
2MQ31T3g3Mrmc9UF1exW9WyJzjMkbMNj6xm73PjA4CD62zs3ETBVCfsCbTQiJldRr/c6PieJKZTb
lASRcUpbt5MbwTDuFpWn+Vm8hNYZKwkhvroJ3i7xIsnQbLe+Js/QfqK9ky/1W05F7SVW8dElo5uV
UOl+LRECotPM+H0EzxmSg8nzoU4x9cKUSPglPQeWWqkNGmGsfx5lCAmZ/twte5mikpcaF/ZGgZ38
7hpsXlzk/nKNiRMF8NrCrJNuVzNzxgHXyURCduSR+ifmZJkrbZlufulcHAiel26tf8RsILK1vUYU
ooUnemScGrfOt+9kvH75i6IepIf6mdRigCyTuBiNUE9BupUSXSCexZTZPWU0zB0fznXERbtam3gT
+pp3+vNidq3US0v5rpan4gmvfZesnqw8gQEK9tEN8DtXWhagv65XzI0v3V4cLpR6twZrQfP6vmOm
m7ZrPsktebijJ6eQmH+S5qxN19zCCR9VyyP9Gzf+J2pYS1/RNNDDMUuGLgmYiAj8mX5/ZLa3gCT1
obf3+hIyP+iczeUyynEEqMa2PbOb/eEJ7tLAkeNRCmgdo7w/xlPC0Z/fydA3m8LQpyKL0X+LvhBL
UPgRnyjkKQRJ70qL6hO3clETXTCBg5dl07Zs1owlGa6hSsbpBYvHxPg//0cVC4ub4F4+QIfw7ST3
65qyz72jdah6eDP6M91aA4Vxrcu9MYGQGE47SqAHxn7MUkLLFjyVkkvAyrxBc+f4Nt3O0U3o8uKC
SqHZFAN7gwMGbJtULjP8bDS/VEpknwF3Swo8lXNmkseSXhRv3IDkJXPauN6Hb4PCAYGVKPz310Ct
8VUsGHAgFRevrUefKgOfo1xRcBsnHvDnQ2b7lyfvVpksRDvIwTNleID49JInFr4Ddn7hXqAGaQdj
1rmMmjHCBDgrjbd4KVv/0mSZ2/PTelY09WeR8ntQ5G7hEblFLcvw6d7kuzKFnV0JnDu4HCRwf+ee
9o2XN3cbAnH3H8svbcsMqcSdFgWifzo7rrt3zCEJLNq78e1+lDldmMjYzLeLxM3rOgjvaAu3zTD1
6MY4VpLZJVGsttETzE7lAK0iKyiEsjTatDiJF9s2aH3Ld69ksz8OxxGn9iuvW9oPsyDbCxtfSWGs
wmbB+1HDpb0BzX6eHFDoM7fR3gqpaxxcJGuAaKihTNQikR8M2eqs883vOzASLhmiKEGNAdlfw11f
/l8kVxiSeoUO1G4+gl+aQqH2PKRe7iU3mNTYwk3gSv/C8B5HquqTvNn7ugePJDw8bQ+mrEeIpbkF
D3Xa/Zm3Nsdi7dhuyMY3zetLaJsC35dX8fGWvjLE9v+rk95KoIIlYYWzXAgq2OccguSHHUGFcytr
jeAwxPiW4NmoBJEgS/zwRwQbim8VXr9DzE54HNGZ9PcMGf6kqMuqxHQv0VsPKlA1YEep8W4m3t4j
LimS3UZCmVwiJHcXF6cN0EF5Tn15VXW3vNBchG9PGZ2MA1FEx438EKaxRmVBNRwTByhsoUSW9D2J
wXqt5rNKs/oRkVm9rPSCCkwtY1aT/QMTpMw0lvwfs7DCIr950X/8aGt5S3MseJ+UHpIHgcOLnnJB
t+86/gFkTtxPcKRYlfPM4cHDaob9Cx1YHOYB9fnB4ISCKmpeTBa3djS+PnGgRXUXOnEPj7TveGbm
s6psoEWMCFgGZSWD6W5yJJiSB733jUz2Rb5iVMKOOtPkrEAzf4AHTA1LdBGVJTJFP9EMGKTiDIZZ
kCdi3vtOJ75P3qShjU+8UJtHg9nDldKd4WI2I2KP1xyGOL+XfgP028qpimDCkaqcqRDYQdki+rLj
0cn2atEslEI9Ea7lghIQ3IO7s7YK/j9pk/tuz/NmocZt0o5OOMV8NwUNGla2kJRiQ364BdWcisUN
7GVT9rK/dT8+3EWdXtFi7hIXuC6hspmiyf3w9rh7zekH6Jj+h0Qo7yO+/3O+WyMpua6Op2mFwgA7
9gVSfaSoRer+99B9OqDcn5Zi2hn4OVcNlKVSaW+B57kWXdr5G1JsvNg3/2zz54rH4AivfRdB3VkK
wzOcOOOwqybl3umU0N3ypSTrWEdSdS7SrN06dcL+oloDosJcHrxzf+RqgFIDVA/hPFxcTTd/ZsHj
r3BG1mxwvZUxzdBktjy3UW5ritiCSrxmooTPGwRxVab6MCzapuqKYmDWT3ENB+h61bDiPD9xCOqJ
mIiTePWZdBfk3PssrqiwcmzZeVvjPnHxbBVoBznlHnqYlY457dPZvrYa0kuqsq1jm6CvUv/Py6x3
2FeSfjhzXaA+4HQ4KfFAGYCKIlYFG0GL2VDfdf5o3gKCqtqsXR3uEVPiTxFdV5dzFN37BVofYN6H
krPAUSypnDr25qCxhXPxsem89zxq7RvkQ6xMS+bxJChjPG/9hZZbYRAs8zauxxuWNBJlfU8mndXX
mkmweefJRvt/mJiS2f2GD8Wst+yYL/31ynrB5vl9RSLGKD9BFQ6ZkUOwC2FcCA14ieMhuXkArkAd
gbR4A2adBp0+14yZZPC3nfgIXWJI8fd7bv09JjeYHNkOphlXHtAWXwS4dvPnTzZaVoLsdYXNt3Kc
F3QIEJJcoklKYF2t64X63uDsL6iUa8D8baECM/ZWcBILHL9q7X3+zW5oibA3ga7FiUzUMUVTaUyZ
S+zgHobAYddUJXTaEBtlXshugKe2uL6fBSEG8GHjII8W2mtZc+Je47TY70HSI8biaopT4PFHBNNn
lHGEQqJc5gfnFr+9eZB5/iXUQ2vJI5KD0GAJXB0OYyNknQkFwryFH/4LP3hIA/E32PDXsQzpuN5T
uT6sWviqMDFApmM8G0Zhr45si8XVh16LI+LuTh5gVGh5hXqFjXalehZrd8DAMU7L5qgW0rPiThJl
puvQ/q7AwqW2Lu+PGF9XO3OwegyT5NL4rlpACD5MgNlUCfKcuLDHax1HXiEV0zoaHZxkyuqjCkMs
L2xaMjkzsglt94QZdrkN5zB8pPRQomCXewzU/xqqU50maRRKZAvzHBDhkP3AA/+8zw9SaWSnx9Fv
r3hkR+0MXWgl02+WsUtjpgMt/nN4rBJyMMVDEvPl/Er1OoHyKjIPqoaCFPw8zqfrc8SSbVIZOuC2
PMrDTN1gRFGVqbpD7gYuPW7cTPSaCzqVRpQZTEpJYZwJslF/n356a+V2DW1fvoV53X0yTuJnpFYP
OuEEkQeaT+qbJnpGjLU4JO1Da0nIWgvYqtnhA8+9v6YhlTUlwe9fQeoiUumEBvQzyHpl6n5ESAXP
qh/RKMDz1x18/EX/BAlrpP9lmdsKN8207rzToK1nFN/X7eCuezFVQzJAU7lUb1C8XOhTkdnv7Qq0
KSyyfvJ5AOMNq2kkTRxbC1Awn2qJw3tOYzYPfQRIq5PqNZNPvlBsly3hhVisReJ/jpWEKRLhD6aA
xPhGck7I8aQDfJmQUICxqVodAWEJttFquYjEoNp9kv59f5b0EhgoNsyli4qaoYly7qu0Hr5Mtfgj
EMuGY34/eLiBt2BsLCselGZpVmhUWdYJZUzRmywBoy+QAaSxKfgQsyedwmpVAvfDo5zxIsLNbZVx
7fFdpaqA59zOff5AvpnwTFUC79SBuVwq33e2S10UFZw3BJtFwdNIIMGhgoY54Kx7UIZY4v9J2N5W
60qtkabKAFnARabLTw8zimrFAnL1joty5Z5Ublgos3DzkBC5dfxzC8uBlo7oEOWD8NW1Tluq9Gl4
nldbYyr4wwKgydQ4NhS2Z2lnZsTJPqwllr7J8+GmzXdjpb8mjI6l2CD8WK8tvmohT3Y0hRp6NMwq
N0awqsFr7KLRSTnzx5rk0zyZX4S1pff4CWmaHTKDU2P0WsHRXo8WD+Tu2j4seLt7urzudQUQwezs
Bg87BwOnwuXpno4hsjkczQkI1awH7tvuieSxLEstLG7Yy/3Chj3YUzGohu12ma3htUFt2K8XOpPM
+OfZiOR0QsemQlpQcTj7+SSlwixxskrW6mODjo0HjMC2HM2H8cB3riyOMyE6mPYOOEdQtv155Jz0
8f/2NFuGuRZWhoFz8DLXU1OLc5or/yvFrZ1g5MZL6T7rujDdJtJPJAx9TxUHDuvhaPesmLZCH/8G
AvseZRosIAH4ERbgh9hpYYA5FmA0E6Qet4aFMVFTTtuPyhvlzt5Ql8Of65wqifr0DEpFJoRYB4PT
ybL3FSR2vwebXuF+KU1848xiV5Y660IZpFOYlZ80iC3/fh0wkxpsUPUQ8bztRqBQdaGE3uOnSv0N
PDnc2M7RH8uqOsBLAMBXd4SnPoSfp3L+FPhhx/srknM8VjwfuG1ub4vqdwlM9zVwdPOTmYqM/8ZC
g47Xc/6gDyCafkyvCBUjx0Tv+SJvnD8i/AwSO4/R2fftGu8O7b1EMzE6VYKm6bqIn4AlD7YGEmn8
/zVyDdgFZ/o7UltID2/8fRyxbLDhzwg7tD8WHdikm8co0UUhHaMwv4NcWRZnhvdan+sNyS+5oSGP
hmPIeUQ0IrLsjHDg53x2oeqD+RN8WwUJZdnCJqLgQGqBUbfFeaLJiVcVWqQ/M8Z22jwzZLKlvKMs
Z7iE3wjyW2dnQsfp8ZNLhiBxioXh9/aAY8wScuDpbFgifCUffQFlWXw5+RyxRUHfVgxtOF/12OtB
m3Nl043HCxNR17sl28FJh+jkYmLz8nwLfch30kkWTiODAnM7vn/LsCNPpXbJmOZ4ZyJfo5grQ8uf
FkJz/rCebsGJn+VEgxs06vwXrYJ1EHo6aspwHepueS++46W6jIv3tPcCOF4ZpRcE//NQnZcUGsbO
lWjhnqkTyA+oC69+w1trQtE4UK2BHqhlhQBRCFy1gcRn91voWviEP5CmELA+l2lS9qmI+IStV1P7
oqw0DUxdiAeNv+gEXX55mk8kLx0dGGtNVezR4vqHCM8BQlTsVQDwFx/ZlKE4+9B/tSg7dgUof9+x
lYJSBW6BvkWKyJSLituwuTIMUbPvjHdkM+Kf/0vXDqHPIzYh109VCEA1ZF+LfgYa4nGzdlEhR7mL
F41q7ljK3XrtZLuubNgK9xuvGs14eK+XrJceo0NE7s5YbxHQYNVCvmB6CxOE8SF0xvUU99wyt6aE
jJCPItYNmWz/9O6HcOKDXgQ0hBe88TEiNOjBpxrIT6FpLxvAxwJ4mI2aOBpbQeHQpQa9qrfkQxFY
37oYoedbB1ZDl7rTyw05G/G4QdSdHTHqdoMMP/KNoXTM9bgd50bjZsUdrTD1gvdIUHLO4zjYmtH9
L7HTQVxDGnE4AasVvkFuVahemI3/ToTrhw4PL6guYxHupBQfgzvV4wxP5RlrYbFEmRtrchXXKiQN
O3C29nupSwCMP10a+Qil+0kjn6D9QmrJqtdYakbCWkzI2v6rcvfhxeLpNkqYoUeBFGPrG4G6MzG0
2GmRwdbyVPbjCqFlO+O4FJuJuu7xRZjwrBD/XQXxZWMpEhHmMTnGXvi5fzWEJXdUpr2OBedbkgAp
wwWWLKtbrsT6OtMhSw58UmkIz/wUz4I+UjcyGKXhWngswNodTgcJfTbsPlyOpO7HUJ4ho9/pV5wG
AesNCgWjBqC+r/rO3cGLtEiVKVnRiKd/Eg6m7VG2Tbd/N4Q8ba2FddLpYwNVUH/FDRyfVcTDbRqZ
5bz5fpy3EZCTkHy9TrYdViAQen+Qlzv4Y3tPq4N37aYzHrxnlgAXLty096BXvPzrvHTn3TQE1jg0
Y0kOQtxSDaoLxTGx/U+fEpGroDEiE97Xrgx70T8CKLfCNDViaqJsbc5u98uVhfNKotecht38QSsx
M2AXN0hKMJMZgCrrz6QiBf37A9gedVumi6YiZd6G/YUHBskIfgaOxntHT4tW50PwkHbJSWazRpKY
2fKLqSRMbWEF9UvVrSE3fLvLI3dCuwuDaoeIOuiPTe9JfydjG3cwIzsWXcCJL7zmxgZQJOJYRBDI
jncLPpRAKbVF6UIUIFl4AlM0uo7u2Ge9HsK7VpI9gFGHNktGxOjd5IFIf9oD/gCADgSGvnk6wClL
uFoSpOt2NHAGkrqazzfewZimYQI9JL6LL6D510C/H5rQhd4PiDLi1moDJr6STXh5Aco5bjKI/52V
NFx/6XacXlls0vpgbi8rzgSeL3NTLl5sxL9RJled8OxRMkSxMTp4wsotk9KTbRcCCeJtiL6ioWZJ
RmiQfgULaPIfqogCE5+5atwCzJuoeLOR9rL/UuxjOJ1jDztwNxXkEOz3ZvFnbpJQR7irLoj9gPGF
F5QqU3iq7Ds9C45sVT3kbQSUTJ1CLjZIZaAURigB7PfFHGStkQd6POFIDz8B/Uq2yZ9CJ3uMdk5s
8/X3oWAnilJFiL0oSNOXtD1VB8iafSclrBKGtWDDy9UKomBPYBxG+a1xAsiCBSvrp7l5AIadCFch
PdtLaaYhrmX2Z9RYATZhOGjAd6tjbuLRKYwrZOtaKyIPtO+vSJs4qXSU8ingzb9o130uPWnc/1lH
xNjn2JHZgzdcTo8VpXe8TY6Uz9yLca7OA5pqmwr3G7+Snk4bg6AJLcLZT7zS+/IlTz3PaayiF/6F
OJkGBAx5IyU4ykfhjpINMD0Q1Pab0tu/AgE5CHWqvhNjM9+PysoQXFQold9uKIQpzxeScSg3Ri6R
bGHTqk8SdfQ+b51TCZKR9Zz/s//94RGNfSA4bZoODCl9QhGcE/ZC7pVYX8psugvpZirAbM1ozNhk
6W72Q4Umddc9UXGwbQ0/itl2KXbjUqmdFL9ojaMa67wr+108WLE31d03bPf0nURUt9hmgKG2QMEW
LeeVa9miZ50xHNAm+4ih8e5BuTadFaryfoNSTpEl2Ly4dQ53cFvtyiPMSQgjJAD5Suij64CgtxQQ
QzKJxl/h9XHb24+QE9TSrTRt8iJlcAp+w2X6yIInE5wuGcYp8q+Pv0LUjfDN5oV4elQEWSGNp9dx
pNz5FP0bGs/DkU/z1b5C5CQlmp1y/eHIM6lQIsJMU5d5ZIs3iKjRuA9Py89dM+o2/LPHllivAnVI
BesMGuabu1TxZ2iB75AOlN4hn0pybwU4gqj/vPgMT5ca1fLy6R1wBibMGkckVVWDNej+2CY9icF2
uS6GcvNSajkDKAMQdum6RygyKy/crm92fHabp6VFjhJS5TDTIxvdBEfTRbY/LBprT04NHa1Ey0Mw
Uj20YIsoU89hbo84a/FnR3VNnudDqZ+zzYhZw8WXPKYBiEXrSEx8yElKA1aEdEuQrOR08YTnsixQ
aaFnuFp7U13YiQ5NSekgVG5tujBUqZFZWWmDVx7l88+Qyx0QhtkCk135TEcPhxDugi1dEI13/lJh
tzDqiGi1HAHA4D0DNmLv0RY9BniW+N3xgqq27jvg21ZVt7dAFJcP736iPT/87VoImpt4pWeR7i+Z
Rjc5Bv0wRbp74QBd3M1W6xUdgljQX1OSkUSwwmEoi6OcjEVSLIecJMXtfu+2mTXu5rskDs/DRisN
2ysKR8psc9Hpa1s68MMALLg3ALJHu7PLoOed6rkGPQmo1vvDPpGRhuvpw1k2mnFkWwATe1aPRH6N
iOSUVUY1h7YYXXzIfOODTBqX2KkQr096kTrZGcilc1aSgfWUny3mLrWgCOgTYrDx2Lk6fhcdTH/2
0kKpAtbP/urNEAGO7hfLUaI9fIYBtEP4qpnDF3HUoMITTRKqiYMmiui0R36HaaE3QIx0erAU133V
VgOWagz741+njvLshfvZYdP+NMT6PEUrjJ4Fp1F96sqCW/TEpDGZF70IFmkmKaFAXoiAtKpIpD2m
SgCwXCinGHz0swVovRLBAo64FDpL+FYk+BuAqZDXHcwAR/XHgUswOYtlXwW8bbSIcZOxu/SZQdDm
5HVlmicWU0DX+XSjDxV0lnLwfpdknvbp5tbucYycTeiB9BC8LmR4A5hhnX3gpl2cnkeSS7goAu4j
16m4LV6luO3hLLPgW+oPTVsGawTgMWMyveo3AU6NWVqqwhn84W1IDNEzAare7rECYqkDjw6TO1w5
YkqqKgup1JV8j1PGpt0yL9iFbp3IwyTIZuYll9Qa0ysCXSKAQD471VkRo2onM6BIv8wDveYLgpXm
jnFzxMpHWfoIDCeeVYgpkw1mkcybxcp7YS8g3FeRmedCWul7YyMhiBCWOAjw4UD1m6I92RplwjLH
JKUjVmzQRzWVLN8aFoAR7vrWrDOHpDIcvLi9fZ5xcs351hnmbDCuXEF2oDTw4GuvylBSjVFoycxw
DtR2+RRmQTgjCAzTIYbMMtlvlV7txq3jS8ULLj2HTzSUn5Ypdr/rr8qa6GI3m0H9LfjpdsfqV1Dx
Qtmikjz/AxSH4F9bZK5cD+MuAR1NDnCBQjxayPyuySE779NIz9AfbCOYmvaWLOwER2Pd/8VMX/oa
96sRcITPLKSZXCC1sfyMdgl+j0CSOFCOGjZW8K7ga8dCE9TIC6R25A5ClQyp1GqSmV6KUVqL5N89
hkq9+xNn7KWW4G9xf7BfAT+GWoWREmN0fJ63BuIKUhR9wNJggL6hB+o1+ZOG9ICzocMK6VjAequn
c6GLPG9q5UQQ6pijuKcSOaiamWwD37LdjDNAxZo9e3U/kVvx68gN+7ZWQlTxi46VGne51DMe3l7N
j9Dce3NhbT8oW4RlKnEJvi2/Pa/PAAn1EANz8h0AsFHCxLyxYlHC6Jv3hQ9QSzCcINOeYqm3Tf54
CoalxhtxrrzlT0nXrYaraCUkg3ELsx0AIS1LG6eTIYUpkrCDB0flRvWhH+NNAZUXO+C4TFeolmmR
T6Tgs8+jrlBHWb1rGQ7ed6f83a39Lpp6GzW1dkYkhfCVx0ssVcooHWsdWf8KJ+avX1/yoIJioLN6
i6MJZo8kdBTcLtz5r3bSdw605pecCi88DMw6TVPH2ub69CXQ50lXo7JOkxbCLej2S6fjMfP2DpOW
aG1Hm6a/xWOdslZ8wdi9f+OEEgZEUdRs5HF5MK4FHj9CTdS/dS2fJclKFjed33SfBxgBBeqBHNFb
fQAly39EIGKju0LbuTXwuI+t23rh+FTFvU+M9NQngDu4G0loEkYM9AbpuO2Ezb6AelLGVQSFnJwe
slRr3Ux5+Fv1TyotPg3vsBZXGpZC+s4HmHqa48VFjyyHc2zNhknvbOxeTJw8v/QKWSmsEwMS8yXQ
oULQwQy0L+RQRb+AiQTD/w24q2jlQzdvTwsJXwp62B3lGHdFApP66tHwKYhIiIy7zU+dAFUPMpZK
ksDGOmeUMnl8gqPa22TDbRrIFSFPeb1O9FeEr0i8wIPPfHX+rM07FJYPmQmw0COwWn2+hr5Fgq47
WPS9/nABtMkuE3COjW6ohUKpulgsmxc0l7DyNllimLe+NaWB12RITHs8hkhoORFMQ9XsEMpZ3BqA
2Cil5p+bH/95zqJLjqTztT2nbG1Eyw4LBIzFynjGCchxizMq5RZWOmj+IbxDKYEgC8cnD51x9rl/
dlw6/IMNjDktx+TsG6muQ0u+rt4ld8OjVsFPf6EtcRgCcNF71l6cjTLMyDnuX4LvMo7GP2ThJBxN
bJR/CatgPnz3YOwXBclkunhibglxSJkt+ygC8MqOHp04Ori64CVKNV+xkX0ugZi7rGOe/gSmMjm5
+4qgv23VOENKEOcNmKL/NnAaB24F8+w4V2ra4eK65ufcuLAZNoAB3SpROu+z07Nm7I++cx1F+yZa
I/+pLVQ+lDvzSpgSyJvXvwqGfEX+mV7071XL/eF3iHD8HXBjB8DcwjqjWnJBmDFy/OtELFVx11pv
NgHTNF1rh7JFS0w+TvpGEw76VTAjniCZPea/Eje9TwXbcR8L4qGcEnsyXOlUILjmoMqVluMnNVWK
ZLHEATKIkvUvqY8kYCTO1h5uZB7mKavjIOLW85n/UITWtimKF8DZeQutztRptU5fEH3ct3CLx7MW
yVa0zyBG+oNw2gDNn5RphX7pQU0yQjiUKfI1V6aaQhkFl+Tudvp7p1d81QpLAHAvof954angdTAL
q4NFZ1adLWeAdgMpST9L5hH+QcGSjhMgif/FcxK6nGn+IqdbkXeGJcZZ62j0dLixMora+5FHv+l/
op5iV6DAExd0AueALFJiMx24upPvZbFeXotYTEYJ3GPzLOgwzz81w4JdKwnKAmW8L9wSXL+4rXSl
RrHNh3GJzXrWsmirG0lc79Nj59oOVkRmrRoLOTb32dxtmT9Ct+po4/OMSj3rP/66UUpTjhMTuZJZ
1/CaLFi4C6SMsVii6Um3cl4NCUAnYU8QoQefskBik1DMc9pSxqrtm00QcUxOkb584FmFtvFDLVZN
ypqFY9icKDnkWWf5Exzx4wh8cLcpIRMpdi/Q7s8ZwuunIpCNFVGaZG3jwu7Qni0icmx5OLE227A0
F99NVbTpAoG6o+ZEk+7SQ342XwJjUg+UMXAD1jHhz2Ar/CGP40j/3lVspFhk+bAPMIRG3o831Xh1
1Hl3tdZ/jqk52kIKgRSFHqyvMZhS/mYsxWjv4oscVR6kD6osIyP0V3gfc+Ww1M2plAagRCe+WfJe
RtekZOZkvgludP3r1W6WTbdNyhkzgf5K5npWBzUS5z51yrXupPTKPj+InB5a/YLiKKsdZAaoYxet
ICeclqcqXCEtChXS8z9MKb78NFy35EKYm+bZ48ljxuQp6xwUvVGDDIvjOyE1NyFTcHIAv2NwhqFr
9jCjVOw8mWSxDveNBscnx++1YYQRRchWtyzksvWlupX5yGdeHR452M0/jMn75NSJ4VhEMt/29TBs
mqWmsEmDtFXybvHlYgXOJ91nY6BFlreIao+JuJ9kguQ7SoYWhyI44yPdnSIYy8ParE1d1MrL0vbr
7XgSK90vop2Aj1wjTSGy+/FVepD5LkXZ6nnorvkH9d5d+fvWulEfqmVJfm6aB4eRmoitG/bGYbLS
e/ygqjpy3wo5tV0CBq4Lg0sbfyXZmMeFXzQpWI/4GWieibGi5pBoPkJYqSVT1OW4CeBXCzTK2/TV
cPrl/X/+bwfWUykKuwi/5gYW/v0PyiZN6HqxiGetuvoB/iY4E+wh873gPgt/ixTyfsqjnIppjvXI
nucnLmtmMllhNZ7zSWXB7PF+B7pS8fyJx3ZfdgB7PyyvG0oN9+pis9aFuX4vq8Ric8q/3UTwk5bO
LlWr+2vRJC8oq1bfiwMlfw4beTwn4pCI42FtkhdFpFKirHcUu7bxlsQ57d7nmhQEEpflApGZeoHW
Pzjr7fnUIQ3rex+XEgGoTtYSKneba5SnnbFSG4dS+A1ITJE/tBDgBb31G/c/ZqDI4+gN5HMky4q4
OYbhzr8pn+HmHot8HBnMYVUkcfj4GXPNfKCfytAlZNKrp7KjhMUhYnWBmH8q6KsyxMmmaKe0kh3y
nJbSRVvakVmWWvycX/FoqwkYwFv6X12hmY9i5eGAfO0nwYt9LcuSf3WU0jTzcKujD0qx8nra7c2n
RGW0KWM4tf7PhVwm0C/s04AdPo0VSe3/RNk/Tx9SOFxg6k/PFHT68t991OcjqAcO30sjpGlZac60
vuVuDhPd0y69/QT0QfUB7v/SNN0vjmnDoR777LZ1PW/Sa7Ix9edQ0evbhpcoXNXZhNVW6Ink50gx
3JqiOP1xas8cEwqTrU3WQli2zAMYHjZ3DXoG+qwdPsjDCayetikG38cewcVNtX26fdGb5pSaB5Dv
VzLAMd46YK2Y30+ylPPGYt7mzMXvYJRNJgLHxrAi035Yl6Hro1HMlpTzXBPrDu+NEoM4lhtd7Rfj
5uiBz9RYceorEHKB95SGZbFXwSdKxQWNJ9jzns7c4Ylf8HS6QVgm57MmsiPl66waR1kmhQqNv721
Z2MLeznQdvKaZ5MvsAjgtUT+fE1uz1lGr5oog3/VSPbavZlddJ8D7ZQhmh9arKePwpi4n5H+RttF
Xy9vGhx1zigdYQ0hBlo45bOA2eR7Yy5qphUz7CHvHbzEuEigSbiEY7qK+3xltgzh8M+Z/w9TX9DL
2EJjCZprxtOveJ6Di/hXy6VDllOJqEqVQjve5kCTIIrfPQ69BhyDPQrSyH3/0iXPKrYDcHWjvBHo
SiIEJhgHhNHCUpiefRL1C/OCTciAWdNTpYRTXs3TYF+35gF+C8YLZbXPjUfDSLsHpPIoYZC9KVao
BEq1PSpCydSn+Zo97UOyTv204znKQmVKREqTFID4qCG3Z5AHihd84ol39zTtBt+JaiKcnlaVTjBJ
kSKzMwCpwUl0TUF3vmCluioLRRp7EIAyi4qjGBgOla/I8Aa0d81vHUiNb1FUsiHNbhutjoktE6tc
jheJNesbNr/k7PkU17yKtmQJJwHWdINWFmwYGn57NfYrcUvrqgsSWcxkoUdo4yL8PPV0eoxokcUn
BOOQ90dpITlAk/cHmBYCQ0eFdc+nLNLONEJqUkWDpIeoJ/VvG3SdIW/EO1kcUbt+VFxna/e85Tdp
eLWX1tcjGwaUYPXZUo+Yk8+PqJC69iFzc+MBZXieijbwhVzR5Nw+hG6PuK9pHv3HwKV4R937ZYQv
HMJ99TlKwBe/nLwQ280UXsflX920SLUUjjsL2D1jT48tExWmKqQtJjj/GJ6WuMrwasFmT51AaV7p
+uYVgUawC4OIzI42EVs/RKU6msZtokDVC3uG/8SpiqR7A4Jb5TYRejVjzL73J6/QWM06oP6SceQG
DPfe7jQ0bWCq7gDfUldz2UfbdbCg0svnlsfmUa7UbghSUqF8OH6FM8lwitX+pOF4hJSkBAQ9GOe5
H4HUJAuH7yyobhdewZwsRquDSXH0S7Hk50q+LY6/FY4L22zGbCWxy3Zj2FJUepuXFkJJsyd+KADL
KYD9TtL73AH0aOCoV5tCx/RXZDnWD7sAzStvyfuIeUe1Uzce/zpdkDa9YuOtyPzpWFgUlWk5sr+4
CgjD28cbBf3oLjZBJF0LcWtw7LBkAMtB+2+SbK7M3Wuc+Sbk6roXDZAk2pOX8vUo4eoRVxgKftZM
UyQ/AyqkHfkW4xOfbQ+lW3XTfytE8ThOhweCIuF+ahb5VMOOzcAptIj9Dqtfop7odEaZyyDUF7L6
8ARsYlEF13vrbRZhuz18mzHDLFmPZq4IbOtXQTqoD3zLEfx+SPCG2a8tCzDyXrUdWB16oSVIa+5a
2zyUh52htM0ywFGReRMxZphE0pt2difSa1n8C9n/HKIwodXb/uKoSc2UtLK/4A/9Mm+JUXr+IdDC
mvErVqtM2YRnvG4CbrejgjTwG5gMcrhtUVWay12NLQIAiQkkV3VsUzrcaTUwPt34o+yWvPp7IutS
RHiv3PyIR2u8kwMG4YHyc05ynTqWPE/6WW0qFYZ8304CuhmV3qt94MIgGjQWsyHxn5FZmqvmAnOs
ouVAHJSzqASVC3htAgUdNVsfF0eqBYXPQsBLvrIbOxLtfiON/5rG1M9Z4+jLX2avpfKQEOwT7ysF
qtOEhE/hluckVcu/sC+T4bNFCX8hCAK1kDdbWX7ORytdocrkrhiNdkQ2YnZ32eLVyx+MxsYcxqAq
OW8RaF7WqSC34toLUdcivXLlPvEHipObZzzFf9LEvZAx751IP9y64iqRLYAEMxTL5ioHZYzRLIFJ
2sy4mgwvzDE2xIcNJROQv9D1e/8EzN4KSAFYxc1MPg8WKWsr567eCWxKgHKE0yt2oGYXAdC2lh1F
Uuxl2rdmZWiMrdg8y+oV9+sx1rE8/l1TMIY47eWo5yxzQ2Ftk37l91MB6dsQEHLt/g1nU0Yh0wmO
9a/CxljB4pRI90ZLx3xtd88THoWSn3iriWJkPgfqC0mo8KmdTox515mSwX+dZ8e6ikF0wETstDrR
96B5PfpyD7KrR/lTAekKgl6WGLznflPrFZXuXl0BHlRIDKtGpeAj92aj6Hk7CDm/fda4e8f1qu58
278rDq2Ct3RMPpo5nQ2a7wvrVqA5f9T7orNA/QmzgkMOVmd/WJBgLMejYQqZ+9ObJoVcqmFRcad7
kovBrzZbhcCInnBrYNmDDFMNwpXTezyVrG3Z5wiaEDq1GPTS0m2ADaYcMPka8YX1qDryHLfRaF4m
vTeMn4KIUBRhNy1fk1UHH1WuAQ0WMXJP1oS5n4T7qT9hFqku/MzponnkWePX5wKspqqCa7kZvuQ5
W8wyhDvhBU++XieX2eSnetNB50CD61sLhGuPjiBe2A21eRq44L5tcKpEJVbuNstO+F3Em1h2e7Fw
68491QZMi1OTYmGXUE4d9T5aAliz2ofdHmvW9Np0we9nZ92HU/Ob/0Ry5sqpQx7CfnlOS2yk/WkJ
qN9oyfHh54HNCRTAkFLmc9AUSgIxG8un6WVKLczNogS+Rb/w3skKBv3vGd/NTxZfQL65PkGrwYBM
E+VO0ORgqbOMFYlfrK4LvSIQonIYQJqPcZcE9xOREKZg3w8m88xg+OChBZ3rbiYSVuxix/v7HkST
Hy1dmddktnzwlSfapy2VNmlUQsIGQi7/FqH2YvA1p2cO7gyxO1KrcEDDu8MWGknNDv/O7GBwyne6
HkAjfx/RcPEIDThP2DlQ/GBDPPwLX2medefw7b2NqKSusLjyj+opvGLcphrsoGo5U9yDcVAWcAFG
kAbJtAbUzsRyPSi4gJ3IEbGETtEj5VuDcpJJZujFWHaWbfN7v61ExcdkVFDAhs7uDcP0IYWMGuV5
EDNevu92b9jvF+6bmXjDQGj6WLg6vxw5wbG4d7M1IQCYlND3fcm7vsQR0aRPbn1W0DXDkpFijiA3
f/oEw3G6c0FX/ldeyMqkR/64EGaYvt0UTt08gVtyQ2FriGJwmuQ82vnixlfygs61CqFY60A2qB9n
FehNyXKBpROqWLRW2+F8oRc6vCpRXld7Ch9Jg7ePZGvO1Y7teFQ4X1Gl5fn2xhP6rwP6KSVXda2s
dFsCC/vMQMvBgTRJNnC5nU35FURcMmlwsWRD+RrGygo8dTeDA0iSe571NLfc29m3KxvUqn4C8NuW
AZtc2Njag8GLhlo0pyVlbMS2JF10p4t7GSv//jA9LZU5uxv0gVjSIbt8bSs2sERRwMhVC04se84K
QDXKWvd3pK4BvNGrq1fNtZ43hTz4o/TYbivnEaLdE7UhN4xo6W0tc5CiWVzO8vsuL+7O07eH9rfg
kD7l9SsoAdFSXqlql6Cg0L1ujFIiAXsU94Yxc1DbVaYb4ViuJpW0qiBg+njzUeNpd4f16mRjPH4A
9CAwZV63ed1FeLebKuh6nRGMQSkOVYh5fnDVPl3cqje3pzu0Xzsv9n3AB31CLvhpST39mpHCSp9U
8jKZot9KZX+C/RFMZOB4+2AwsDDg2ru5E+jC6irtiOCMISCgksczz7kAOOE4Hh8fHtObdSwkWuQq
SmVBhdoHbQFJSanhifuegdkCBTHA99c8fAZ6O41vNVrPW20HCTAwp5snzCdogoNz9A2n2I7OYq4R
qx+9oILkMgwhogVL25lXVwKciH0JoE6DlkP4Al3PAXt7pLMCX/ervXnoRJ0R1JPqfFPc2VS5rGjO
w11K7+Yao0bZxToA0yuc5b86DJNOg1LNrGjVICt+2YWOCHPsdpa1dbS5iF6ZcI5O+PVn8yRLL2jN
CxLSZrQGeFwhu2Jg3TyyOjeZHDJNDcF/wOdhG438ZTPtzyGZA5CBCgonQCTZO0BYsu7LrHJNcDyy
E8w+HttzCKObO0W34Bs4jMMcsgJSm1wXjzZti57Kj5nRxntb1JAgXijUs3cm3AKRZKTVe98jhCCa
EBA82kZr8ZkjOQntm3r8ubMJ4ONRd6nSJE39IZ+01RutetkXOg3B7WECoRvPBSaqtRq5LrVtB4fG
mHRa61vzKcEV8yrCOBCkorCo7qlVP1rtZcmST9KrlmzOpE+DD7zAoFvdGNLihYlon6p6PWMSNxl/
BAfCVwVUWXgxj2wioDmpQa5+4E2IDLe9WTPr6x7tYyDEFVvu55BNg3HQGewvgP0JZJXi07g3m/6R
HpzSPaxNlNMAT9dRkPvppy3CoNQaOZJMOvVpkQHAz4gLiWohJ1J9VAO7MIIKPm6gJyynl4eNIx7E
CxJm60Xv9uASbJfLYVvPMU67qQjRWD6bHGbmy8sLVAZSR0r6K1wLtgHQq5LpptItvFu2CTQrZsl4
p3K9RNO38InwxL9VD97sAyNC57+kRuz0ykMooI7X6RV2SmZRIoiwIevVfe9+AfQy6eh6J7XwRnk3
Th7aF5w6dh3y3P7ryQZJwe9h+8pa+U6E55EyXBA4eSXB2EGzxjEmI1o4WuzwmR+TL15+XE43JSY8
H8GENjWXBCT223CgRfiMHx3m+tbHRukYMu98waktYdyE+NcIs9fk5ApYi50J5T+qgFbJMkJgHeFj
y9GPOIUwFV939F68ifqjS40R8H0Bd35XWj4zM4qMSjHXNJhGR2Zyh1V46Tp4SvClz6FAmuq4zNHb
9h4LNt1kIznog7koQmhxqZs+ePm6i/0z/IxrsN1HmfTpI1sK8bv8pS0lWWugmqNf/PA9SlRoeLuS
g5dimXmz+zyXdbQc729EMxatgEAad/13vYzGC6mN/0pdjX3ocK+Yv0nTpogjL6OdNXVH4la6GHCZ
zg7Kg03GPvRECEhuvWnptxtAmY/R/NTR0wju2W7u129o+Q3M73/rHMaXoLkfPAxTL/HfLyiXMlvv
Cdzj7vzNCoNGRDBt2jYjQoyqky0CM+qQEvpmWpf1XRn7eizUbK32sXL1A80rL5KejpJ1Mee+Ey87
NuQCx15/9eHuP+TSm33tvsD1wk+gjjJxQwbo4yEFyIlwwqX+DSyQJN2BrIQBfGm3p5Zql+iZSlvC
wcNAHBnXP3pmjfMYlTjSxUYkAob5vxe++I18Qpg9Uj1xJpN5rfB+eHTVbRLz5gqRk8i1SpMSaMQH
amADnzz9uv84bWEPo6ANCXxd1EvApEcqR86wQFRzaoJP8DqprBz6ntoWg2n974bPcwyLpSN3E6xk
oU/bBYy+gA7KuY1Gb0o0Tp4uatPBPgaByV6d3Gol+nxBGASjuncEOeHrcfPYWhFJH9Y6IUyI1/tx
2AdX1pq8NihnnBrBcIrnS3tNRZZ+nr7BN22BKDy4N3g2WsmcmVdwf6QfVmaMuh44x1bMbuaSVYxP
QmYJM4mm+ijUe6uFqYGnMsXSwVSZa6rxxsJ83F/t9ymr7pYJrzQBnvEVzIrvl5ksEEhoEL4lzJwa
GndjdSyKA+sqcxWP+fUrXmE1mVGMUYlkM/GqC3HCLNRQNXMc6xM+LfGi6WWmu7Uig+rnfo7IJnfE
33+RicUcBuK+meqdylBx2wxr0GxilOwx/JfBvJd1T+4Qc+ktF9AXCkeQdzQC6ON7iovp9tvgpVq/
16cAG77yxcEeauGU8HgQNhL16a3FN+A591GheH1LBTow7S+ndL19vwk+MgieY2xvYQ7r9rQ0R40j
6xfBjbBoY6qRDi0Cp7u078s8p+Gp2ZtxcZaQQxUVFtwQ5eapCxcNyD5rTT36d6U5zHtSBWcMaLSu
YbprO9MExwZ9iCdFV8+28jd3ZVNNbaJXEcgJFGdZHkf4bk79y9DsBH4uOUbyZRDSCU2xN3AF/5Su
tY+8fE8VVwqp17w2cHSNycviZJ3mhf/E+l/gdQJtRKVuef/KEbx93csqp3ep0MHSHPAfQidsCoga
Zlcup440mbCP6L5TNSJ63HdXPQK4oAL5neFUy5+54oLhlK7cPliidq4yHoNdDTeKoeC6tXxkPpS+
YMVGLMiqyMYKl/+BtqoiD9TR0MFWD2ijJkR8CpH7ORGAErgqoCm4qoh6eBz/xMnwOAOV2REOCtOi
qK6SzTF74MBaBnmsqOu13pzcRq/T+ftHgQbumHTXJKsoVxooVPunqJxo47cffFDtPz+IeRxOD/5J
VJJxK64KLb9nTjabFQmjP9lSHvke8ctOHAeOVRAhZ75Eoj5LjMyNHXu8NaUQuVUrRHqfjk3sDV6g
DPs7IxiDpp5VGpI50PS8+ItwplIFN10IVJYXXXdfkuHJz6Dq1qVTu4aZj5/omU/3ZqcityX79o33
NyUSB3HsoaCjujcd3S1EdmGlWG5zaGNRDMrEsbCE/PUdEHl6Z+553MiHSZEMjtsxaU5rX6F0FMx+
1qY6r1K8WE4w7JJazS/qDRM+11MUzEvlGuiATjLP4GjKzN/pCuvCDsEQh3NocJ1Z2NKNRaEkjNS3
0SY7SHm1JFUIg8QD607wEu0ZKFeLDa9RWSc+h6YRUFbHk7GJtzB0iSVo6FzDFr1uah/M592Zfdah
8R+l3VSzmd5NAlIsp6bTiCabMgXLhv79MbBJTSZhv7KOmsyDFIBFiSoFGzrPGLSaazBu9eNOPcEI
mVAuqY4ocR/vOt8uh0F6iYyqeEwtxPITuUHptJk0pzD6L+7CLxaxMYqQT3J9noQ4fviBkzxQ7ufF
rqhH0SKPEvD+nmYdWdg6ZPflFoX5OCtrO1EP5Pf31vI5bxPp6IQ1uS65oqpijH8OqkaHYebAgt3+
9uc4Uqpk2eTbfUuCaVuCXO4iYvbXCrHwDCrCaHSIfD80k9InA6XMNwj577L7Dhsn36tICuum/jgy
kAxyQg5AV5prhRhzIVPetvRGoK7V+nsNzOafpQ9JP75/KiMRbvR0K92+KPwubDgrLMoTMxL15ITb
mayXkXooJ/XojsNyZuqwBxEs3V/BZ+eyQKWmgEhDLv2mpPDOmYKw54hBR9QNGIt+GKmo3s8fitQo
t5xAqDp9cKVp+4YMDydndq5Ll3RNSYnbdxWZqm3jN9gcaaHAs3L+dXKvGOQpgj5TzJtNwE84OuXN
nZzC/VJqHT3Qgm9d6v91+PM1qODQRS0pd1J0m2RlLD6fAL9wb8k68aY/b95BZf3KdR231VIqsJrH
5GiPnIw3B19chvY97zrq6j6jAy7ScR9W1ZdiTIFUQaXKLiuvkpzh+Mu09+Mx8p6Q6jSBqZgzJcsy
6UrAiF7fMFCXlLoaPsosdK/MhdZ+isDbjyUf6J3L8Ut4QU99gcE50TCvsNvuvFoiCLVJIfxIOa1v
7sKdC0SkBbiVgiHYzjWb6bmKPdA2KlQ+sjcOU421LGrh2vTFsey6AtG5eMK/UNo7TANbV+k7A+X4
dtUxNXc6q4KLO4vts+BRVO3o+d6wWsmnjCX7azcfnSMlMcFcZPyTuNUxS2LFblOtY2aDFRUXjIYP
YPNZPr+9YYNGLeVsj/Ri/4qyIhQsiqrXvGpjWIEgyBtwbTVyE+eNyPf6Rx8RwYwdMJM4VMbVWHU7
H5lDZEE938h1CLHrLEHQIxUXYEajFEplGUaMGfAAPxDth/8F+O3gPxDiRSMs3IwPIdw1fsVjp5yU
FBGRjjAr63TDrn+l4ce97IiS110EdBKHXlyK9HpVDuXP+u6Bxua3P1G+UXw2kB50pclg5AXV81XO
eGVhz4G5/CJwAjUw3PCnC3W2jyJkyx55aHRRHLZO5Fy1sYBg7PkjXkq7PH1EEYwEaNXy+kyy6aKG
ZoTvag+ZNAPcoB+N3d8twiv25xstPu4gHDgJPStO7cg8jz8Ywuexned8cF6vCAk78ffoLXZlCNHq
yhSLeVrqR4p4/xaZsXKRdiYDBxxJyHbEwDpS7xVpDThSny4O8BHYfWFVAan8niCJSHFhtrd0PISc
a6u4NR/u0MGb2i0+OzPRdA42Y/2qBO/IPKdY1z8ZzIbcraNVDf1yEyTYifezFR9dX1aQf6skq6+u
sIQ/PCMi+kuwwlMcyLwCFcdAL9YHB8G7N7ChxAfv0+0BzcMzGYJ85BHe0xsYmZUQfHfJ3pWm2jig
chDUDkfIFeTwhtcXv/L0LeRKUQbvhUg8TGCo4PXllMYTz7LZvQXKJOL43ZE9dgkr+z/1/WSMQICs
ed8BrdsvP5s5mdaxpldQHPj4lyFzx0Uc4RpcFts4BpaPWC1MZQHo0VhxJhZUkWeV6LBQ3Tab13e8
IWH25MrDUoZRivLHHR/Lz4CSqXRdBf9GP9zI+ge2DLoaEthUCkWeYD79fPIKU6mzhgWniBOgO/q7
Oh79iSHlcOR1V5pjnnafTGsKLTDuLfKkxAAf2QiGVU/7JYaDzis4hFKmg5QuuY8UJbtFxv5PBb23
jCgGUQog0vIs1an7zD6dHjg/e62oRQCiTGQl/Z7s/hNhZwRR7Lve7sUgdF2qOPnFXQovJpX/vjxp
pUl8JYIKeW+1r9FIP5GwfI73c3lLNQ9vVoNig/xa9I9ABDYrbFc6IXwRqqoWX+Hs4M/gO3OawECP
VN6wflqq0KOeV4kWIRXoGQO8xiq5IbMYb3teyXg9c8ej08VowhPTRp8XyM7a0OHBEc7X/F0ig+l9
uz9JlHYMB540a/YkOYbzZDJbKJiTbJjd7+J29rtOBx047Jr+xQIFr3iF6smAcgE1qFZwI6QMg6ad
OPpEFtmacUD4N7tw0RqZ7odUzf9k+vTjgqTJHUitoyHOP31sW+IKepV5T8KrIh0L8jZOCAeFlEpv
55QF4NVRXoF8nSiGyoqO/awS/Z5GE9GvkhHqFYftX64X6OWJX0Gt9doiBLYYLYykxAeWAU2ElaBf
CWxd7LVV3D5yrxBcCqZp7ElEiI7WB1eZoKXkCayKl2iH1hZwJWvQ0bE751dSsxiKhR7A3br1NCpA
TQh6uGhdS21wCyPPl+gDsEeL36Z0WbYZdMSJ+YqgIqugmCAwNWgMybNbzoLY7dSKZbT36OSpKlf4
cDh31NOz0tW9S+ybcPpwqm8pIN4HOfLETmhQy9ROJl/FuGzXnZfWsQMcLpOcvtun3JX8Q08BDgkd
CvuV9AgJcnKzxkX1yRtFtEnwNP1q+EplqNxnykveWK7JxdRpm/K/Pq/elELwp6nJ0F4oBW1F4QtL
SJHxMOMtv+qqlOlNJ5B9BlMy9B+HtW+b1j1FSlShvw8/zRzb7aCzXY7ThHOYoij5TT1ng89C8J+U
TZ/CaEYGGknM8v7sFCLFeHJnt3zOTYyFUJfdLjE7ObH8xg8+EL9msuMXvlfiMWm3JLoUHIlgFt5f
/zVuSDGVKPdgdBLIx9y9TbBwOfiR/G/oVo36kZzLDcT2tVdeDWBnRVBO2bzVTGLpOL7d+mNdYP/g
5d8fcJbS6Ka/1a0SXGbuVV/9qZT7a4jfksDdXL1fapJj5K6pfEpwmr+wsvOkR6xGpdtYaC3URoH6
mnwPX1vqTpd64aHyW3CU52BKNkJMWyVKHU3PVu6JXgM3g7Tj29BXOICfX/Vj5U3Exj4hiDK4Ygwm
RuOoro/63CkzWUszKES6WkQU5RGkAbB0Qo9bHjayV7HQA+Q/x5mwFdpohs4A9gQVx331bvHEsM61
c9peTSe+VIgGyKRsCJneH9H6hVI7JlES5wvVSQk9JGJOiO3tMGLfwKpf+9ta/Bxcm74GAxdAoZU1
Y94jQ5OisrhEwkjJlrPi4MZQvklESjoUU8UwS0MOunbOfHoDeGDI0b/m0KH40tD2Dq9v9vaxw505
qW2IO1uprBQ4nx8Vo3q5e1YV2xH0KSTmqMggFWYWeBiO4PetLcx7J6L3amj/VDROR2Sp3htafoKH
UUIJem0Vpjuze0lPT8pU17TQ2SJkMMIwX7ChLXwi7/5h627W2bznjwkREa7D0qWI0igmG0Nx2x0w
7cAIeHHcurSRsNVa+ptpjiTX+2XClgAOdZUa2nxBtffPH9DNIq55MyfG7ii7jtts4+on5l8LBjMH
BxPR0CzAeuC4HYBUFvDzADibBZelTfw3ELz9lhDmkkSvdsqiBe4lFI2dZBdxFXgbrcjeg5rBS6um
NmLOW/inqj4OEZhQw4Z9GpvtLIdN2uN1diBsAiaBLCZi1/Jl7L0fYzEd5K0/tuVBdv3cYjuqitKC
2IV134JJoBXV4kZEasSdFBeafjuFLuLZO0uJywYBymBuQ5IQS09CZhkX2o5Py2sYZD9PhOG/mf7z
CYvGiAFXdkb9qElLGDjLMTTJazUu/wsKE2TGLOp2p58dll7gCLcTNjXRzBVvryDdvLAMHRjM42ob
3NE2XdPDWQsSbMgPK5Fy7WIfQk9yIKjNsDeAaIerpmrVlXW/FoXk7swA6RPRXyK9L0rfJtUoKenz
mhV7Wn9CWIrCuWpLhyaGXOmVnatTsNsH4MC7HvQIp8CsKarzwFpoBN6XkzI8J7exjDZ2UYgqmbD4
RQfAZP99cpL756wuR0Y6f7Zn6kT+i4nzXg+wTIHoGwPQBRA5uy+kQpIS4L2U5X/PHJB6v9B5ONV5
C1zOHswfI/4G7chpiS+cnhN46EXO5rq8uhFKicqy1TH2q4q9yuLe4n8fcNJ8CGY48P2uz44Drk+Z
WgBAA6KRZFG5+lDhL+ctxR1sx6qMzJ6wQjTfWHeT1t0j0P0C8+sA1cglSkJI/+z6LoLh87jSMbCZ
NXzUVoEvi2Qokkr5CpCzsULu18UkIaHvigucF2G4w6jfReT+OnzmdCU/ziPuwcA0zmlpNoUVn0+H
HKz99JOGgoZBo1TTEZ7+2fsK7M63nZxzMv/8qTzXFERoZVd07KJJMfr77sfo97A97io7cXkwZJl1
287gVs1bsisQ34bKcWAxHGnU8Jz9sufxEbMHBYHhAYSp8JBJWpzP0tpC+zbCLqcxFBqRscOiJqPe
DjUKJKyxE2k3GJBytm4l9JnIelO/dX17uQSX8yJTBryo3I+L168wZAK+AiamnmDQs8ZCUs0WB1h2
kirNvu9mmofWDu5DMXcLUElWhZiuK0SKjuaZ3JHcnQU8EgrSP+4LQKZWAnoLkPqKK7g/qb0mH9bQ
GJ4LxIPLfEQWT3gO3qKF0Lkhh+CknwlGgoklrcqgAdf2MyoUV8pDu7Cm18lx5he1S47NQwn1f41V
PujZdxRI08cN9pqG8T2fcsJOd49cqWmO8xgZnWjDbqLf5ksvLgc5jsiVFlAg6kAdvnHwOg7dTivN
zbvumE3EwW/1C+rOXCDHP18aYlDEvoF3iz7O2ZOCU6mXH6lY7m4kHrrEcv3+p+4dqLfHqXoThpKt
+kPM7279Km6Z8t7mETwvWcRw0OdVtAiQCdHecqsaEhzXGi6xX1az7qlaVlZT4oxJokuDtwo2yWd+
hWO+bRxtLaZDeODCpB+QlZQaKyGzSi6THwFMrIuKcnt148rqS58+JBHVF2M7cDOKPn3y5kQsQ98C
cbg9wOv21esctSOCPEhB619Skjk/VqXouIHiGryOrAlJmxEVZSKbygClj+ESLjxnmWMnwJJfpM2K
yc+4lXPGY+2pFviUJ0/BxpeofDqUYjOf3WgwZDAwqP9Zws3u/hFr/5F9oQ/jzvTid/Dca/sAR1Lx
vhQKYJ2ETIlC4nVDtonNgYJZbvTSZPMp5eZQgFCBk8D3iAw5Xuh+IansTMVvQ2COLKGFGNN8HVcu
8XJViaIVRC3HWctEaTsB9mM5ZVZes/ECrVVtwlr7mhqmOW0XLtHWVMPb4ocrXX3oMShb53xB3JKy
IudDAsLvMvreMw2TxDjH4XXAXieAnwrHAPXyg03SWDCLvBATzp4j2Ow2m9cPN61rTW1vBTKIFgbo
1MLvMrPWcpjxpYCy0M1HlPyVuLK6WTgI+otpRiBHsHK0WS1zTf9z2FwZ/m24Qk8jPjnd46OBKzs8
sVvUHWvtwwZ/wupzXzEt7s6nDRF0FHMVlHcvDElJtwwIzR/093e+ZCC/3/jAoNqrlXfLkieqCVDx
nCdoQU+9hHQ132kDYi5nFSeOPRwzQH6lxkI4arPUbLx/0dciv4E7OevI+jpXMNyzbKrzxsdBIo+t
pcdxlbEj8wU6T/+JTr8jXd1d3rysunmXvmo/C+lAZG+Z4Gq4/ITL76WnBoh0Rd7C/IccuyRi1HQI
5w0AgiOoZncQBxVhINt5m74zPLn05qehr3FxCqQMwA3+E2Z+vad5BnShsdXwqDTD8sA+vFJrJpAL
tQq0TiU9XeDsj/jc2BSsIaPrNl26LsC8V9zqypib+UBjsNL5Q0GLgyB03oHXKev9tbN627d/p6oT
xBzL8FQ9NE9qXu7xBOKDy+P9Unh6lNeKi2P/161Fsc8NbcCe7kRD1EztpOo6H8q/Hd7F43lb+3u+
HNb6wDz0xL30y++Qw175SNEaitjA17uK4YEPQIrBstEM0OrNs7ESEewCKlrIEmrEkdSWFxVZySTX
kCbQibYJDu1bkadDB+MVQGYhNUPG46tVNnDBKK8Z/Qe1qmDFI4zS6U13cgeCQL69yN+8JO6JzRNe
SxK6JGsd6N8FLcJQomHjrFlgI3HoA8/4kwv1v4d+C4Gzmi2/59o/wrD7Fm/DNTlsanUUT08SZl1P
Gy5Nhl+Y++TSnC4OAEQZMoUHncG3WrrPIMDVLJIekY5reLIU/u4tKBcGUXo+McFrgQxNa6828c+W
U2gBMF6S1HTHKAmLo2ndGYCvF7uBn2kuqvOoAB5CjUo8HBNKI+MbqppskYyEdr4rpN94ZbXb+Mkb
XHQHwBHfgunl+t7nk2DlR2Tp1WkP8GuwhyQUPLHMhq4Yt8P6EVUXcJNf215Wsgbm4kp+L46C+Eb7
+5I/Hawod8811HaRnjWieIEYoyOGevWXwnQiWYTscV9vR4rSERvZAn7rrzJ666Zw6bfvzZW/j/b3
qvc60DQepoJ1GRMxQYrHmVj3KVLbXkoyE78B+EainDZE4EBPjWLnpYBu63LAbUt81G77tC8KA9gJ
TNiAK7g89xhJ1CkUlTb+7sAwOq/JfhDUzZUdXJ9BGgxe44A47p6umc3mpujiaP9G2iBtvbXKC+r/
9vRrRfIPf6hkuZNsRpS432/WGEwicKLDsYI5UZUzeXfjVU9gHEY68xVJL/iDxHnPBuxeH7ZPZimB
8H2ERnYnuj8n3XNamIgTZD44CnmyHo9R61UgLz5MBbwrLcVHkf4eAPnOKizNbW2UJV191siUf36B
XMUvc6xswjhDOWSfiuJ5suXgEOkES3oTPsxatmcKYCFNsmXCkfclJcEqmLjvRlbFIvwKl5VOxUYW
wgBxrUcIq37OrJi09WVm0QU2GbsMkNriBxbyinOskuc11kaT9Ka6gHpopIPcTzfEhG5NytuJKonp
36ULxA3tsDgKdY9q4/9mSnNRLg/4FMDaSJqabFTpugmd7leWijmIxvaYa1l+QsrFkKJWLB2qNJRO
3I7KyBJXnHoPQNFnQTGo2q9Cj/HC4CROiZrs5trkrjfkadDxTJSBcvLMs7D30KVVF8vrP1fbuGYO
84pfJzqw5jTxtjt1i4COCmKbFzfqMkjup3VyXo3OAXvrSMtM/gYUXNTDfBAAvBy86ssIjWelPsre
sbGMEYG+q5RlnGlj+PSHi+2BoRYbUQWn/dOvSviApJXYvd85Od2MWtc7apT3De+9RnQEPn1mwVCj
V174rVSXZNzNoMP6dju7gv9F40BMqEnFvrTVyGwkgBkef7fwRX+y3wz7/gxzrhxugrY1rqJtaWU7
qw7SOHisv9m1UHYHDx4deu8dbJxUnoWH6R3jpC+gNgf6HUaLYNnzWFFIz25c4ZGZ+wcLwOyPsLf0
yLrswohrNOwu5oIAsbs2Ew89llny+J6iyQZUAkBvK0CiMXdjIRTh34HnX80xke6IcYp9IM7RlziS
V2VB0ABtB+dfECYc2NPRCYCsRSQvjAxx1G425vetnXILvyzQCi2dNU6GTw/KSgSrTmHdFxOOgshG
Ti7QluPppfdCQcLDCDMGperZF3gfg3L9Wlm8ao305cPNBJw76TptEi4h/rF55Pd4adaJ6EQnGilt
SO0ksAmYBx2UMvfOFyNIh4xTUbeiAzcFnSGQTlNZSd1o9zhheX/rB7V9LTMC43JjKLeQLvQhTSlz
6MMepGyIpJll+4+UPkYl8SWALA/kYnKCjAne+dQj6mZqd3/3kk020berxPV4xQmEbYFr+KsKP35v
3eqbqzBLBLJK16LuNsrYCEuqls2vOYBHwMT4XR3/++LDu1FtZBrkDZkP/OeY5aBNmUYw7hSnY/3C
poWAPod+ufwDZBwQf3Wpl86+aTGaGN5DYvtFdKkHrEvbiIIv3QMbYT+9UQo3weSVN3WkLqnzMrlU
9AnHxDlkBeu/ZnHg3TyYyOHpiRHD24+SKcd+LktM/9aUTkGxG0aX/qAHicVzYvcV/OxxwAMbZXgW
AM59mZI4+og27B4eHFLSIky1llJRUPAndvKLugIRjbEdTXfn42vs/PchJrvYdAGEdKgkElbAnLVS
CPy7v7NRcswBIx0mE4H9anavxNHksqOZPY5GMuglJ+PLZlQkTJdn3q2JGt3B6uTWxwX+hJ2z3pyo
M8uQ/NulADYVk0RnAaxIf4LbcnYYRSwwi6MojftWPdrF/56wQvtWBbEMyqZwk0oLDuo+s/OmkQfK
6NZS3Cf2e0dx0bGjpQP/wzYcXNRhzjld3KZYR7hgYn2aiXRK32ATa0w3XKusyZREg+y74/2OL5r4
7vZbk0rCVBukpuzDQENfa+UJNGnkMmbLEHhNVOkAA0R2HHdm1zdYc5IHU2GCfmJOKqYJZ4h1pL34
dldTxW2g+H+T+ku5vUii4Mxw6Xf07sPlmpU42PfO+bxx+5wx8Yazs1Hp+8vt2VKNxJFjWXV1i2Nl
B2MGlZ06UKAjVY0UZAyJtX615u4Y6XlrndQj+YhphvSA1U2NtJsoDWf+QZQBHo+ISE0qhstzCXbl
b2C2H1IjVHLw5vqESlxDBkBJKlB2V9wNfrKKllnGaa9FJWBSmQ5+EPK6lwQnEAm9CMod2hljBovK
f+ryHAT6up5i2mZ29a8Wadthi1nAH9rEPh0oOrsxI3W6Ot8uipNwo46022kjjfWKU9uOBXYX9s35
m4Hko+adAoUczfepXft8GWjuRlqEh9n2iIKbT4rjDa8AbaRArUc4bpOfVaZC2AwcnqgdL/jJyDHa
2cUpCqowjIYhVF9DFHfdiXlXS1Qqc1DecM7ZWisO/IOIT0U5jJO5yv/98snfpwTs16MKSLE4MF92
Uo9+TLNb7L7CIAblv2D06hSVUWZ39ALgXYw7YGiyzlCF9nEXTywzcFBwD5LJWQLEf0NCPaztc8Lf
xu1FfRJ3/zcrNaL6Gf0IaExUajA8hgGuhpc50Yhth0Jeap97O6ro+7lNP5jiFiSWyi6ArMfOAJad
k0xV20sdKsjjb6r2loCav5NAYyzgTUos8TyE6fQwVdq77rCl66iKisSjqrVpBsYHsRKutX3aKpPr
BO4ih1r2bd14/SA8xRDPPxY4ibfNmyHDM948BnRrOGWwEpFJ3fVm9g5HijkV436R1X1/+RsNHF5N
aXtGFsm3A7i99a5T9a1S2UWd8w7kMA/pHMkCKNvvvrsJC3VL+efAO+qefaY7+nzCU/OHNyyLI5Gb
1JB1tA4i7a1MibzviGgPcarrSHALOkyfCLFsrabAmb1wNwmCCSOXeTghyDKQwRJp+sL1bkmil/sA
tqhgMJ045hWLlutU8f6TKOu7C/8kYyAjuWA1qx3IcrI0Zqj3nGiP0CnBC0M73wisTDjL00YuXyKH
TzhNJLJKPg8cX9Ags/U40ajRwmCJU+9azKmGDYyBV789ahhiFVKIkbjLMUlLFIeMaCJIYaWANFnA
yzTglIuqIrR3XpMkAr91+i7SxlO0MSFaZSe2ZubgoweLsKJEHGGhqw1F0qVBGMvfZP3M/Fe/gGYU
m3JYWHriDkda3Av72uBnXj3crposCZsFEL6nCZZK3fZ0qReEMy5dt0juHsRCI+BZYfzI4dIrvOQJ
vVPrUIyzcdEpEh9lJDh5ftGUIM2m+3gLrxgZKItA9F78Aqzt1cCHwUfZ3vARDgVBIAOBt4YG6qL/
P3Y18XGqYttFd6qC6v+HN5Ydx/PHJFyCaS0Rrth926YlT9cQeqP0PQ0aEIKYnJ0ZIFqyhUAgsEHy
Zsdnzqkk5UdO+325QTeEdCVtf07vRlT2esYiC3pLR0SNspPJW2AEjwE+nqYxk0rd1L8CeFgRDTa8
fPwFKiA3M0M1kn3Qg3sU7z1FfhUCo1gAr58c2eAoJBjBsnwjfeqVxZTXhw9bXlKMFG+21TOw/OId
P+6pDa5acvdziC0d9rbjLk0PkAECkP0gUuRYmbKpj7I7v2tEclNeSe4wTuW5Lp/dd/HG7qq2a1Oz
NEXwo/7FxGKq55cuwoqDs30LzngGT0qOWf6SnzS1DPTE7QUHcvWEU2ofYsQurBG9IkEzlMxpC8CK
RwfPV/WUCAneqViyOwFM8IBY5M1Si5cVqnA81SceXRbHrz+xBydNzIwL9vNC5v1ZMqViH/OjI2Tv
ZT75d951QhdXAqc3Czbwv5XwLhFpQyInbGjfbXrC47z6czrD9KX/zh0rZSgGfEGaZIdaxPL1EF99
1j8vMndls/goGWmZAD0jH5e6Sv+8T9OOpV0kkgt4Vu119A1CcMBqM5E11Jii1BlzUHfbHZntykpB
PFWVYgIKDghnsoo8XzhfsaGJpNcNnTAWm6zEbRUaYlbo04hIHkkoicIeskSpuGswY94EXQmwHFKb
HcvIkQycHZZCkMcGgiZEqMh07HwWlmFUmdkJSEu9+iMCtG8rttAxk5KToBIWr56ziimu8qGkhcUS
TvPoOJFK1rkrrEd0e/f2aw/JkFRBsb2PAByGguZk7j50I61rUG0z6ggBClbX3v6n/O8/vnEQmP59
hpWKWQ8py2fJ8Xr3Uuqq5LZ9+on5yCY+IKjJVwVu1oVNqOLkBHjiG/bGFXnULWO+Ag42RRmUP0ib
F5U/ztjmIoIwdKDmfZO+8NmQrGVleMiv83x5k5X4agFOt17hEX4QwqEBTbGfXNVnPADukLv+KctJ
eiTPEzJ35JWW+Yewl+td9vOap2o=
`pragma protect end_protected
