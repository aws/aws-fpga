// SHA: f463fc25b8464dd6c1672ff28a603eec67bfcb40
// =============================================================================
// Copyright 2016 Amazon.com, Inc. or its affiliates.
// All Rights Reserved Worldwide.
// Amazon Confidential information
// Restricted NDA Material
// =============================================================================

module sh_ddr #( parameter DDR_A_PRESENT = 1,
                 parameter DDR_B_PRESENT = 1,
                 parameter DDR_D_PRESENT = 1)
   (

   //---------------------------
   // Main clock/reset
   //---------------------------
   input clk,
   input rst_n,

   input stat_clk,                           //Stats interface clock
   input stat_rst_n,

   //--------------------------
   // DDR Physical Interface
   //--------------------------

// ------------------- DDR4 x72 RDIMM 2100 Interface A ----------------------------------
    input                CLK_300M_DIMM0_DP,
    input                CLK_300M_DIMM0_DN,
    output logic         M_A_ACT_N,
    output logic[16:0]   M_A_MA,
    output logic[1:0]    M_A_BA,
    output logic[1:0]    M_A_BG,
    output logic[0:0]    M_A_CKE,
    output logic[0:0]    M_A_ODT,
    output logic[0:0]    M_A_CS_N,
    output logic[0:0]    M_A_CLK_DN,
    output logic[0:0]    M_A_CLK_DP,
    output logic         M_A_PAR,
    inout  [63:0]        M_A_DQ,
    inout  [7:0]         M_A_ECC,
    inout  [17:0]        M_A_DQS_DP,
    inout  [17:0]        M_A_DQS_DN,
    output logic cl_RST_DIMM_A_N,

// ------------------- DDR4 x72 RDIMM 2100 Interface B ----------------------------------
    input                CLK_300M_DIMM1_DP,
    input                CLK_300M_DIMM1_DN,
    output logic         M_B_ACT_N,
    output logic[16:0]   M_B_MA,
    output logic[1:0]    M_B_BA,
    output logic[1:0]    M_B_BG,
    output logic[0:0]    M_B_CKE,
    output logic[0:0]    M_B_ODT,
    output logic[0:0]    M_B_CS_N,
    output logic[0:0]    M_B_CLK_DN,
    output logic[0:0]    M_B_CLK_DP,
    output logic         M_B_PAR,
    inout  [63:0]        M_B_DQ,
    inout  [7:0]         M_B_ECC,
    inout  [17:0]        M_B_DQS_DP,
    inout  [17:0]        M_B_DQS_DN,
    output logic cl_RST_DIMM_B_N,

// ------------------- DDR4 x72 RDIMM 2100 Interface D ----------------------------------
    input                CLK_300M_DIMM3_DP,
    input                CLK_300M_DIMM3_DN,
    output logic         M_D_ACT_N,
    output logic[16:0]   M_D_MA,
    output logic[1:0]    M_D_BA,
    output logic[1:0]    M_D_BG,
    output logic[0:0]    M_D_CKE,
    output logic[0:0]    M_D_ODT,
    output logic[0:0]    M_D_CS_N,
    output logic[0:0]    M_D_CLK_DN,
    output logic[0:0]    M_D_CLK_DP,
    output logic         M_D_PAR,
    inout  [63:0]        M_D_DQ,
    inout  [7:0]         M_D_ECC,
    inout  [17:0]        M_D_DQS_DP,
    inout  [17:0]        M_D_DQS_DN,
    output logic cl_RST_DIMM_D_N,


   //------------------------------------------------------
   // DDR-4 Interface from CL (AXI-4)
   //------------------------------------------------------
   input[15:0] cl_sh_ddr_awid[2:0],
   input[63:0] cl_sh_ddr_awaddr[2:0],
   input[7:0] cl_sh_ddr_awlen[2:0],
   input[2:0] cl_sh_ddr_awsize[2:0],
   //input[10:0] cl_sh_ddr_awuser[2:0],
   input cl_sh_ddr_awvalid[2:0],
   output logic[2:0] sh_cl_ddr_awready,

   input[15:0] cl_sh_ddr_wid[2:0],
   input[511:0] cl_sh_ddr_wdata[2:0],
   input[63:0] cl_sh_ddr_wstrb[2:0],
   input[2:0] cl_sh_ddr_wlast,
   input[2:0] cl_sh_ddr_wvalid,
   output logic[2:0] sh_cl_ddr_wready,

   output logic[15:0] sh_cl_ddr_bid[2:0],
   output logic[1:0] sh_cl_ddr_bresp[2:0],
   output logic[2:0] sh_cl_ddr_bvalid,
   input[2:0] cl_sh_ddr_bready,

   input[15:0] cl_sh_ddr_arid[2:0],
   input[63:0] cl_sh_ddr_araddr[2:0],
   input[7:0] cl_sh_ddr_arlen[2:0],
   input[2:0] cl_sh_ddr_arsize[2:0],
   //input[10:0] cl_sh_ddr_aruser[2:0],
   input[2:0] cl_sh_ddr_arvalid,
   output logic[2:0] sh_cl_ddr_arready,

   output logic[15:0] sh_cl_ddr_rid[2:0],
   output logic[511:0] sh_cl_ddr_rdata[2:0],
   output logic[1:0] sh_cl_ddr_rresp[2:0],
   output logic[2:0] sh_cl_ddr_rlast,
   output logic[2:0] sh_cl_ddr_rvalid,
   input[2:0] cl_sh_ddr_rready,

   output logic[2:0] sh_cl_ddr_is_ready,

   input[7:0] sh_ddr_stat_addr0,
   input sh_ddr_stat_wr0,
   input sh_ddr_stat_rd0,
   input[31:0] sh_ddr_stat_wdata0,

   output logic ddr_sh_stat_ack0,
   output logic[31:0] ddr_sh_stat_rdata0,
   output logic[7:0] ddr_sh_stat_int0,

   input[7:0] sh_ddr_stat_addr1,
   input sh_ddr_stat_wr1,
   input sh_ddr_stat_rd1,
   input[31:0] sh_ddr_stat_wdata1,

   output logic ddr_sh_stat_ack1,
   output logic[31:0] ddr_sh_stat_rdata1,
   output logic[7:0] ddr_sh_stat_int1,

   input[7:0] sh_ddr_stat_addr2,
   input sh_ddr_stat_wr2,
   input sh_ddr_stat_rd2,
   input[31:0] sh_ddr_stat_wdata2,

   output logic ddr_sh_stat_ack2,
   output logic[31:0] ddr_sh_stat_rdata2,
   output logic[7:0] ddr_sh_stat_int2



   );

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2016_05", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
PscrApznik8KIAQcXmWmRGZs995twkxENAWiaxDUhF7Rvm4WBKTODc10DdbXBXwIYAxGReEs6e2n
SnduHQFx+dG7okC5Faodwc9ZoS2vm8oN9+hs24zq8c+VwAkbsRAX6t4y1BonYElbNfTyJ3AVtSCo
wf1mdra6sOdZPpD8RIw9iFSebexLfFiaqYiwE74u1C13ZsVo4lmpPmXvnKd7Jk01ZORaW597EBk/
KC9N2vvIPtjx3z2FYpfav3E4E7HkRXZE567+QbU3puEVeNfQElWSvOcpF5ZIJe8oA9y/36kL2qQ2
QYrNe1ZlQDweHxQDKOKY4WwCR3te3iopEdWzJQ==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
cP5G5ft3MOV3DBwKiwQ8PrgOj0BFYNRFifFucF6syid9V+XHjxrDvDgekKBdB90SMTlb94AQO30s
eyDQILuZkBnCOHNYw5b9+S5MmMZC3ZMTHYJQHLt0y2Uf5DAVvLTuT13kRgia017QDOxInNeHW9DA
yz6pz+IR4G4UPQ2vemE=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
AEW1v7yXx4tRSijCfEVM+QAUlMFB+Cc4t85SfQy6m8jvbVUpStLaBxPIajBia1zRzxDX/eWOKEOD
rvY9jJkZceoIyzxkfKim9IIjqCaENOMRuhfCZuN24/32wOZM0fFkXv9x06j+dcWfN1TSGRTTdqTw
YNeyxl4HcKC6f0acb7M=

`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
ocXE5tapOYRBKrrAlwmaFZ8jJZ8frTMnH9lYqyfqbA3Mu5WtQGKgKSsHD9BrUZhXifYubpvlkKxc
jeip9wmPFg==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 71232)
`pragma protect data_block
ax82JA5Yz/G39jpKniMvZ0fReXBJ/5U1xT8wZSTITNelxQ6KNHt8Vplj+WUiaPQa0T3Jumx9u2CD
fGxOV6wEYhfnMIb8UIhKUN1GAcl8Cm3c1e0RzzydqE2z8iKJngU+OcqxDDQH32RLUxbmjitn4ysk
Lh0BnGwO9EF1q97tjDtEmt38HEcKuLmlYRuzt6+vp/dEz+EHuE5AxB4cZ/iYa+exw+nWYmS4Wl1Q
tUpxLhDAG7r9Wjg/lJown5tmT6Z1nbJlLRbiQlLH5diF/jIPwR77QqTe8SFWiSonHsHu9w27n3Ck
qOCwsSp43XB5gpJbDXgFKkm2A7R9pqxaRcf5+8U9R0VzjGQslk9bINsvGpRulzoZP7Fc4lKmLB1A
QqFjZ/fWBvwa7kPTeUNysjwEFWl92SsVNXpEZrS7wnsT/CuA35qoYAvhtCMz/HkdPl97ummXhn60
SM6Ag+7QJor5V2t5qYSEjNfi48v9y9RjXckSbLL77LE3Q7vT86TAM/lQ9Qt29afOYjAngsybXEVe
xnYxdH2zrIMv3gvsi7Zp3QkMg3tsYCMPTfItDGchaGLiU4stUlE0TIpHG+zzYlTrVzh9+zUVkfUU
6P/eIRN567Ua4td17f2mdlucZAugBIC7K7nhb+OwqSk/imVmld7BKoLvfuxYzIBanagT6NKE8L8c
Oub3I3HKF2adUbBgFIqyFB1JlClWPE5yLZSm3BOOK6z8/xgixCdQ2vUnpW1ZtoQHe4yLquEI/py0
+wFw6/5hP38Bj4sml3XQ9ocwqDpTSVvbVhFcZ3xyyrtLTKA9tom3OWneaCujS6s0/cny5ExFAJ1q
kUixiU4QZnIA5BpNjL0Ji1f1/RpSMhrDby2SHhhWOXzzH6CnjVln6f/NXQbfYtJK3IttwmILgaJg
M4+0DLkVs4ufRIcjPweT7QmYU9YKOa4lrmhaIunWNH3O/5x450bJbIdnYJPPw996rxzSdMOsbdZK
SMau72Jj9aTuv2AXjk/rvMaRqaAzOeeyBJuULP9vALgQ0xAtHdPUrFewmFtyMtGxHZmV3O44fUv5
1VHcrukWLIzfGvfXBitsrDDWi9jr4nL97r1W4OMt6fjhcb0GvPJ2ksfkyUEdZm/gIbVU4UWswJCo
gzDxgTPhSlh4vuZjrHHlovXSeHIw1Q3n3XG4tTTpslF8OEAyRsmz2CjX0fFpUaSD5tPXBeP9GEAf
f7x40iDqp2rhxh/axkfJskjXkFO5WMA+gHqfldusmRkjrGJkQ2cDGQZb/Q+OpMCCyI13b83NPkq2
siR/71iAxG5XY56HEDiDZxeS5aVfSWahN1ANbv8KgZ3j8j/j67wvhOMgXN+jT2w8HvPQgVCuA4xL
o1BSqZ0ejltpJX5iUScYb4yX3g3drnt5+2nv9CwT2yyyzXkFsp8dkPzB76xTXoQYCrBAaHjen44o
HbBaxclvUIcPvvtXm90b8f7DbW6n8gN1zicVdmRFmmwPjlqHIRoJCmIYulIcCfbVL/xhgcaYx2Iu
ZXFjfobtHLCsjfVxVTzbwQe6cLkwnVWGNjo4FpKG9hfwMpvYNmKlZ1Ju2pH2sP/OIpzrhdRI11E8
h/tsMM0xXOBwxgYzd6mEyvt0Ssxh1oicLkqvZMM+/U26XFb8MwgNRnlBczajWviokT/f87nKcLlX
CiuUa5fXZTo/I6ez6760TAYrROtF7uPt+nSIu90MJv8t+IwQ1qoI8S2AE63vN1hzrAq7y0zqwKZa
U6Q7GNmcTnXSEq1uJNHlBLPu5AsbcGE4G8iBExRtIe3/ik7auYVlwU4GO7OIvO//0j1D8ccM0R1b
sSKm7E35ZAlzHudAyY2QugRr/lvGa4Yg99xdg4K4hUBbNsW733rS4SPvVKy3oPzVW2T/N/BgF9Bz
Fk79o72PW4tFJrlrDEFaMZ1Vstua69Qu8hx7YGmYhjh+3W78e1h3rT+k7+CmhyRtx4v2qWZRNHuv
XPlVEtfdveHRqcrnGH6ypGRPXklyNSX6OHY/yuURJ6YVhj/mOxCJww5Ykdp8puX73eNCDA7bOzx7
s525YEWnsyLZEAj8cj/HYG4igJbBXIgdypKi2+0ErvrR05w5uFXTBnBmRNZO2ghvZV24SpOq/6G9
gYbK1tfnu+Eg8lgh2la9hZ4Sarwdy+6x+VmrPmiILb6wDXr7TsNHnoJYNwrADSwLRJr3RfHyKNYl
59CzrB5FXKUGUkTP9JtEmmCbnKM6+f0X6QHz1HY14ebwl9xLg458G86cTS7cYEpZQ0F28g0i0Xty
7FkOSTEglcu0GmR6h1FHMaeEEH6wkZnPOQvhUbS3m/JsnJtHnURqBr+5SKznWF4wx4LxiUJKaXrc
0iV0K1QdOuq+VZtiHHUCPtGWKRWDfLyaOdIlIE5f6zFm7JTIw8LHcw5lBbpnwsuQP1ZQhNEKMqdG
GNqjqeXxDAwrHJAfrPznIZAB8Q59aA2xyaTF8SkhM/cQs6dJpPh2Z4a15lDv9Vs0/RhE3/peTrLf
CMspDJE3pRUZxp2bM6QXq/h1iEZqyw7Pq6TQrCrqf3RdOyFdSEKGbz0yfG2WF5ryySKA5cDl5B7o
u1Y0IH4eecCQ747+HHzz6NczvYK2zvF3QDQHQDzErNnAoYLIKl24uvuf3QU9Lxu9t2mkJ/eAnPjc
kAdPVQeq0zjkEmjS/w41sI2mQ872Wll/7qeb7r9JpRYZCNV+zZLUAZLctnDbdHxZGb+QAL5WoDyp
Hu9nPR9Bvu/kvM8sKFScTOaeZh9LU9InT/jPFx9E6pyU+tSvrfrBuT+vko3iCFsutXKtxAq90Qhh
ltXg4gkNJa2TbuhrcLtarBw1XFAp5jOjnemJoYtKhSXyiTpijVsJgh08VxB9RG57PWuip80gCxY3
z9S7uiJRJ/jf0hf59j1mfdae84KISY5IKO+hXbFmUTal4hVW/8nGSngO4oDGk5y87aZBPAK+hXWb
jWDW50ICYImYGLo9W2jBVkEQOi5nC7vS2CwOvxQh6oC05PXGpLVybb2oIfUNNk1Bc20dG4fGv4mG
yqkLxFCcPbvNOTFLGhQg25/EA36hK5j4G9nayd9lN/NZ8ZvAMjGaxDRvRmVHJ0wwAA6ElIJrVwm1
tzpqFt936Hm6wBSc78J6lbfM/lbOFeLcUEIy8mSyn2KTUwJXEDqWBX0PAXRy5AoOaoCWGN5V+t61
Vtlefu2OWgDeNVXKs2pXf7dX1uZoQK3PtvByIoG2DzNACYyEc4P/yJomIvU8jwPjUGsNApXadWp2
0xOctG9BfRiz1yUuZn1r89SmYDULle7Sr5qgdFvnHGRPyt2+FRseP2ZifvAH1cuyYP4j4Gwg/8Uw
hwaRiVYEvU78v26HNrCAe/XH207acC4jXJYl4/I1LlTVizYfZLV43PG39+x9z3VHL56emhIsCetT
gPdJ8nmhlzG6K4qvTsYQacZt4ichO7F0p5jeM8fvYPggHuxwEKvwmP4iQTKilP35YSiAu1r0UmB6
KMmzmB95ZwIESdUWoS2rzdN4ALjkt52GQ/Y5otwnBgcEO22gm9WHA4ukgaFu23rkQmgxdQSzuVnb
lwnSj5YWcwKX4xZu++OZAXiwMvNPsbGF4Amcd9+qqysEQMoMWuBVhVg44k+aERb18bzyTgbEOyy9
Cwv6LtYsXgkti7YNuwPaZQ+QL5shfSufwFlR13cB6CxyEjvgIAOHQYg6aWu9ZSoi+pEirEbX2ZBk
NhD3VrC9gFBWsBbGzRWcR1GBGnRQLv/RV2Gfc5cV+1X4TX/CTMvkM9laAzT9puZ12ZwuIUtamLqx
h+ye59xtLLv5gn0Em0VLa0LKsuDgLNud8ang0UNIw4cn6gOEjVd8ya1H4RDEO+xrVWekjDDS4sGy
merSBCFSy0c2nkgEOxJW3iX6C/xm0RddfGZririFCDrqp8d/BChdD67v4Cp5+5AGgBhIVL0XvYKs
xqjLXc3jAiXMDtjhTubi4+MRYdkAYXd0HJgzW7tuKhkf3gTz2yTbZrjQQzioE1syDuAGMvXid9ZV
1flmFUL/cS6478piJ/OP3U4Qylq8ehi7edUO1DuAzeOdESiDQnwkLAXYTFuAS7ABdAy/IJyIbY7y
LkKdsMT81YoMb0hAYdgZP0uHEysanyHId2KEAy86SuI8vhRIeCU5j6BCNXR0o2mQSpnLSY2Ek3bF
K2xkWYDQwQ5ZcyeDrEx6jfkPcZeDih7iTxUU88Wkr2zqKwfTw/t/EveQuDcU50PiF3I4thsKzJjP
KZSdDho7p/gwjx99aWZPViPh1eCKxz7VPaBzlD12Wt8OwOfouJ4459JSYRWOLGA++7cp9dkWfQRs
9SN2c8GeCIMGNwPQM8vAMBcxq1qNbLwdUFup5Qda1viJh+0bZswirXhNoViTOsc1Goa/Avd6FbZE
l512N+5URp1gR/CPcA9+M2rET7nfwCJ4XZ+7kxnnaaypJTVTw0YOtk4huhCJoLw3dCuhTLr5VKAo
alGpqCxrHMnFK7CFLheuOlH5wT5MYLOsemHb5SIuAo4uPxEz8Fu13TNTzM6AksB8Kf5FlwBRf7b+
NqVYw0VsqgflzGO3HtmHGs20qrt4bGThF4ERNiH4uwxhdOh1tQh8F5QN7sQk5xndiPoKheg6c0dk
ANFokcvTnQY6dhcrBhC74L/FSJCGkpqd9p9VOUpeksmc9KtEXhuPiFa16IlKhbjFN0JXAEsPwASh
+QZcAIwkvw6vYeumVVetH3q5QsQ+I0QuFHgDqsX5WFyrXwBW1w1fsEr5JfUh4iA2hQseZ776dCpb
f0P5hQvTqhRCfX8DEoJh2rMsirlSdyJFz2cWU08Q0S/HCWw+UaH3yM3oZ5yXrl0Zba4sEYkX0Gr6
tbwbkX0973MZiRNRiZhT2XhoIkH+1syVafh2aPUTJ0dayLSCWZnDtsuQc3tSq6MHtZDmvn1OjKQ9
E6qr0raFLcF9ufHzOT//T/NzYXWFntT02i4lTAm1eY3TnpueWhvKxv+CQL9/kMeamV9EtQppxcrW
VJdK41ctunM73wilzaGDPjupk11+luwmj5K6XT/PG9Fk97t2LqTjH5fKfNF5ZmbzPgbOem9/YiUv
3d2WcHpfxAU+eqMuU/PDCs+DsX62Vghniod6+nXPdsZwrZfV0BfO3DiMqYbYQ9NEH58qbTLbJEkA
lBIYWDlyyvo+5iwVZ78a7VSHyUSs7SiNBpO0AZJuUiwkGhtSjV5WMMB5/9YV8GPaxQBVfOMWYydI
lzb2MT9jdrtvYJb47PBST8or6HgloZRZYVlPd66tZdIEFzOhw4wIBR1K8czc0rT8IJ5PScz77OEL
UOCDnPFxZWTFKvr267GROGnYUiGD2l/VHW+pWNoRlaqj9Q6it1OM0VnnRoKMoEd4w0W8hhbn58VP
9AFbn3iuIE+JL35AYs9kqhNmE3hbLv/NEywoqv28CVM83sVPCHQuvqZZrnCwhc5cRDSH6Wf9Y8lE
wnOqjMQouYnxqfU9EQHKwXBbUEnb4l2L4hZ5k+p/qDSo5+kGaH5oege7UVMmdN6crobw6qvZAJ84
9a0zk7XClYJ+2wqlt21oNxHem1dIet5e/rOtItiJoHdMG3Vr7AkNlczAjaPDkYCFhUmLV7wPjDfj
bV6AxfK5+13eqzH7NQUwNuhU4We1QIMZ5fUvKkFo6Dx5+1S6yPReTRbBoI5CdVnsacBEMlUm4uGE
IxCjqT6EXhvv+hI8nDw5I70S0de3Z5DrKxeHuESdfTZvWjQl+3DQoX/aZ7tGIr6vzL8hc9BSTMaA
PpJh+iqm/g96r5fmcd2XgFHFqgNtwvmI9se3/rLlAaTwV5aR28eqWRCpA21gCzCqzYC8yJnwk/I3
uJuwh2RKVuLU8ekDGY2xydKDU92VTYmhoSjzS4UiA8lKB0IaGxbYqy7GGP2TKKmRwHEjVQjVfcKG
UYJ2Qc25l8+o4YmUul485esYDS9r0RI7N8ughGNWmK6kqYand/PT0mRvqtTLzBMpbLYx+ycK6+8n
f/SSubLU7nxeUkM8OjDO4W3JRuGDda3Ssv59Enm3bGT4PCdvZV3Ig1Z2M13oHlQnZLlfAj5/JaID
ged7kJbvAmkD2alsRIrIryVi3FYrQk8Rpv/Q8XWeqPmdEYYtmFSUTFAwpuITJXhKTF8JQtPEnGPd
TF0d3GlsUIt3nVWfuS2D4I4/Ekay0xI0qQUEZftVFg2L1ChpVvtoxExUgvGm9fh15xU4zvU4ztzs
n95uS+aRed5n/W2YaAMjJJLPCq9Ecq2luAUbdwzn0zwTYU4LEltIprl7noyLRj6QfVV9CuM2N8QP
S9QY8cW3Ha1X1y23zigPsQE+MWg+wxwAG+lMbwHzCQUCqYCzicKLlNw5xP4mfDBJypsK+UvGG9X+
jr5xi95bZYmT1oBahp2jkVaIXQn25xbRR1tuoIuwjJdWicYQzjP8OatsgGmdIcG58Dx2xouCBy/q
4ndvp0puBYANeGRNMnrfwAN4VmU3kCvZ4dCDhe8hNAKavUMj4N4FNNDpvm+d+92ATiY1fwwZEtuI
3yUF2MFWF9H2/r+IEaT3/GXofUr6EMLYEeqtK6aFRugkZp42P9aUxNppHFHkqMWjS/+YQrF2qvTa
H2xVxGzDgMJvisNYeXiFhVn9ZcDSoI8kcTMFuTZcth9LfRm8gI+X5RUfCgRGx986gc3rAD6V8Z6+
Od/vvUG+wh4l4neo2SP9cs95ewxdtU1/L/Q2x+gBXPZXNHcjsXcrgM3R+hgTsZ27YZSWvYO2iYkc
RFc//Cbpj4cjiuH0XZwXvRm2fMMN4bdDlPpaY1YYCa8KD+9vRAoxGCjsjQwgahlkW1EZgjB8zXH6
jrmzGCDVE8llwwjIw5hXI436ig1y1dbwf8VqDrXz6+IlE6qU8Keh3cDh9r2v2jIGKfAK4lmhr8zW
rp6Kk50g9Bejvw65kZO/KSA1DqQaL2jmOnO6E0ovsotRtAB8sI2ci8OYowI3ZSfQqWnwSL/0YQz2
1Taqn0OIFF4NZ14fhyDJFl0z+ZoKEGa0BX4RTqXP/tY/sJTShJuWCtPe3e3NOPFqJyMaqFghBCI8
TUKEOUjkxP8irwmFJpeD2bR0OgEHCqEYjYUx9rUc6C9Bc8VWZLtajuA7GQZBv9E1n4DonL2dN+RK
Q004Vrk5Ff/FITRM4hoP9ATLv3rl/mTX1fIdbs/C0/W3i3/kFg++dGnNGyLH74UH4vB3uLNNS+zm
dukMW8KWjpPs7Lb4QR6QufSK6evd277GYezqpaEqhRLHhOUWF/0/dcLQh03ceUHEBEawuYO76SC+
48tL37oTR+F4Cv14DruD3up2i1u17h8JqbGLllHNOlFgJx3ql3J2KnbS/VyJCKrjXCzn1ysRuAmq
HPXw1JyQE31MsE7JNNENr3ywFLKGQqOf3Fq1EPoZniaLh1qOwlg7mwzjarsYAkQsI6jNxTFRzi38
ZVRkY9r9WsKpFxWdtSDjyEbwDe78+CfjLs5eJ0fDU62ir7FeIBveMtlkYaLxmhkpkbPLa/S5ZKnq
OQAdvbmVjvf+5ElR+QaeeRtI7blau4KBwssf8TEB+6ezrLU3tPkYNW/T2BTnsaKjgjRApixk9ik/
Xej/fxpvrMNkrSn6dmBLWDbIfyCE1z+KL/kDkeXQlNkEKxNrmLez5mZoXJmFGNBmjt+vIGiyOIUV
9AUOnks2xoON8nhfPi4XbMGxHWqqsYjzj0cYFj7BlV0iEI3//50eiaPGgKji2+M+uzg9XVcZvbDI
41W5FOIso4mkZZwtVgeV3YhTfKdD+COADUvC14hF2WaRUJoMIZuPbyFKn3rAWVPF4F3CDRKEqMe7
yOkH5oQQ4uDXQj0DMaMpDFmQYXHyMxq1s9h34ufI9HMFnDbn4i8DQBw3Npn9XF1aI63Bpy7atfOh
53iBVl4goyCZhqMaiTOve6mcPhEPozFkyEQTGOojNxjLvitPfY4I1c4JHreWNXNu+g3WyH88N3Yl
T7N6B/VIoOy+qBwV2ugpSFPlykr0ktn3eOpReAuamc0hKvi/PaMni1T2fIOrq8Ifwker7Ae/PGhP
cI3FhP3PKxzJ8zqR0bhK1SZSnCDb7Axpvb6HVsqM3JTHQ+Njd4mEoXcnJzjUuPwHCo68pdFI73WE
Oea8uVVrDoRIFzXmJcHmhyfyoOIil1kNxGHMhbrce6kgKw44rmeURQ9M7NZYnkh+/8yXHTaGIQeL
Q0D0ghoScmG0qsKJSQZB7rbSzOijU8HQ3j6w7kZ4QgJwhtv0T0MfUIil1ZKy3f5CjxvsOCB/Qr/R
hgPF8TyiaWRVEp6fPD1zMf7OXPHI/BYEYEN/smWT+Aju5e73d38yOfrWYoY/0snAa0slBvr1Rswv
0ouvut63gOuhTzdyjgAuYtYHlOFdJ4yhBajIYZCJGhs6p26rvtnwaVyzUJfE+9mGzrlzhlhqRTVq
shBX23tkQBd8q/PjqBvzctf/DTgr7soUmuOhGDk5yo3ARJ7fnJaY77lt1clN0KGnNTYO1XZd9Hre
my383ptVxw61nccI6cxhr5gy7KrBFLicemY/WKaigPZpm5OW4mboKGgI3QxwvPW5o/fctUdsUKvX
b1eBF+xcRYKSp0ZoNYfMbxCfLF7ivZCepa/dRX9wYuvM1Wl1hGJ2S3+PxRQ1NNV+avdQ02pFiuqW
YhPeEF97JNeY+9XvCEVhWLWjxHa4o5kk9TUytS2xwDo0Ul4eqam0KRm4Q0zWMxmNLzqPG4vGzBZ0
PUcBK9thBoE18IJKo+z+FlRG/3VLFkSWm0dNmOqKacvDvZLWRP9hm0LwViSZpQIqB4b5arHPFrFL
bMk6TGNRaGxGl/GrJq8FgzHNL5TKIlkHddmkLleJN4zGEYHM1UoyXkWk1tbCc/UTZyyI7nf6YEH1
cr6VtToDkkktqhFcX3XeXC6ltnAHL80E2avV2/+tF8Jcq6pU3+RWrS2NNuC88BSYVPWP4IiBq/7F
nGWGDRTHiYj1jPVh1m1Uk5oHJET8zkeqpRklNK9d47BeX3DdgoR9ylVqnz51/znk2pXuuPiIviox
3yEfW/le6WAcgZB/uVCwiYlnrxqERRmurF4JEYRsMXUnuURObjNABVUjlhA3wczVMT9SC/OuPL51
hBywycUFIm6Hivy6DtOugQdt5f2dGIQzPLdlQSzeT6Dp/uYyNnUXdU5UA3nxOH57s9fZadeqEymZ
3NA17r/pfWJoGIUR8GUuhl1HXP2Xscs9zai+wbvLLoPuF5kfcjUAvNiz/ncMHolaAF4Dh4eg9gCi
s501feNG/dBhT68K19ENxhii5sxu+0o9XxwEM3ci3otWXvNlKu8wJ3bONyp/HwkOwxFDwUlxGLIF
pLAUbhqqXoFgQjwzxwC/AuAGI0ysFHC/Ce5bWJZjOnvVAz86uCe72PzUDYkz1JE6zub/BPMHjjhZ
QmQsp1v/qeH1mB1gpFxdcZ7l3h32KHEHoD0iXJzS4i3mcaQhHGvQAIMQj+TKPnS6uVE61hFsLNlQ
AOcRRTsPuUCy/MXqIE2xYusNV8FFrtmW0oaMCpwwg97hlqgIcgl65NNnNTwYSm07vO3m7vI+w3O8
9G8r+NX//629kR//OPQBVJg+SdoWWQHOKysoy4IGA/XdkQRvZqemQ35woRu34VR4Jk9aLJC4zxWI
MAZVpSPLm7LBvSvAeHLNLHaSMySoZ3dVfyImgbjNgciRHpTuE75CwrMuRWJhd/z6B+DxfVQGv56I
3Czk8S7vGxQTIDNWVH3GH3CxV+2RDG1TNzA13o3ScEf9qVX4KHj6kRqYRBuwvpD0EnpPdE8D8XX5
kUtP98uPBE2zOy2Las/cP5jypFFFA6m1dcC195hhJGg1Qs7TGAN7swa+732EjP26sFN63sICZPPG
E+p94y0G6e45Q7VOsbZoZL0KA6RLowcDUVNrjkTEJ6jUKbe0GcY3hsKk00cul8FTenN8ijZWiDIu
0Vuuyed0oy/OIjkNVcQ56Y9E2rqBR8NURz4aWrWSG7pogBo2v9SmTqrlw0anc2BeQsFGdCkdyjp5
eGkCx9S8F9yZ2jkarGSktCN+ydxE8UBsLUu8XEZWjzbivDuOZp2tKJ+xv6LijRuQs2/3HK9ovSKo
RShGGcDCTEEU50nVg9waMIXUD8elIDlU+lj63pd7polpcAEq5I7qoYsLI1LJSS4fgPuexgTDbH3e
8Seu+Wh/bHbMT3yAYdE7wZpK2VQMpJ3FfSk0SkLuNfyjQpRu4CoYaFlbaJclluYD9YovbP04N3zZ
Cbph6+96NQbgpZhuFeLLcu5m+IF2bAIpUiQIM6ab9WVV744ixjm9rKDBPDgWGlShw+L0BeggdMJq
4656O4NYwa+hmk6yKO+YYAM96oByx1jQdyNTe1r1hea3GyM8f6S4DOlOnF/eO52SK7NvUM7SEQ9u
IX33Wpu7upzPY9oppYxpnTeJ3Erbh3rwX+r+oVqWmdjujdNbaAlIZRh1WVRbIdgNZEa5u9/Y311s
G0/wonKg2vtIQ6NbcvnD64ocsMaPYRFtYi7EgeHt1m576HnSxBLPsh9rlGvm/zbmo1aMoItwm7U/
97+xtDmOisr3T0jRSkNklS7D0Rz0VAIr7NLyhJnczDiyE28zhfP6eav1FxBPk2VDNIcuKA7zpo+q
G6WrboYzIo+kFyvJ7X+VX9OMddLtJZGuQzhyUdFg+YpgM3JsPkc5924GsOjMUOSvqDhHAK5kubOf
2uA2wX6FSKyNCUt0KBq24IutWoZlhZzZLwgEO1Mxm+Ln4hdX2PaKMwF1N/nH/Trsx81fFAuSSvGy
01uyACcAWtgko6jpqcjg+kqK7AKPM/BQvvA/gCjqvKwUSRKWbuxpflzm+BM2f/5b9+UGRfwSV8Fl
g5BqO1td/Ts03aN14BppYk3wUCoPlGZSGnAoveHYxrmhyH0XIdtefRJvLB8Vh5Kinj6ji/k03SA2
Q6DNQ6c/C7Ph2lHlYajPmUEP5eMouP2apzePNSt70/KtRair2a2yjgtovuENeK43cr84PYynxRFh
zzK2zMEVgx5FSAJiMWC7lnxboEhCugCwrXadwtUDbpFkUNVhE5+NenWsgMk2tHGfvfAmPmo1iCad
HnvoJsXSCRYTUQSf3aZRgCXf57E8dRCzxhN+zM8JHsIARA9OOPxLEQso4E9nugEPcpPSzob0Z3k5
LlI+p5SkpFyL7M7PA14muKvOYtKNzXuuoQJYE4dMqZ88hbmJY/qQuN7kQeL4aAOOmI71vtEeMbaY
eYHdUJt2cn+TFwsVpf9AJfpMquuZHX/InZWmiIx/3RgxkiNIXxNWOXTBnCSEFWZuKIX7aaoKk0ZZ
q5/rQKJp+1iRLwSZg57Hhcf4uMDBoZ74GChVX9lIbb9NmgoCeqjoRgAer7hApTmNuG+sZpu0/cS7
f6wgj+ueQZK6Wzise9eX2XAEguKxPkHVS2HaO9eRWBM7vLL66eFqcSOLWKabDxIGhH2kMwq0xMhe
zebljR9PRiH0MkiCqdUaTPTHojrKhmcG9K2phxEMkA8q3CSegXZ3b9NvcLmkeCAR8LvpKGEOskSX
dUhyKPgwV8izcKaG8vClwekSfQ7Uh1eSi3TgiDIXpju1Chd9BthWFK4vcrXPKccYQ+CkmbT0l2QP
AuSm1T0+tjMWR/SuJXjuo6N9Xj6ZkUKZUYttX9joJe9vuo/jegGM5KKLylZuzCwyMJxko5/X1rkp
rD8SiAOG9hy2sqTuUv5XAcaKjEExiLpU2xjPHvFuIyBnHUZU11tRqCEW36/kvzEW/5WjQ3IMjQE2
1Bx1UeqUxamReuZIIuq8yZJ4y/j9MTic3WxC4GUUOWwM/kBPF5qnfRBMuRLrSIChMJEEZ1EOoR1b
KikAdJ8ms4+tqrVNBaZskzzUI4lRmFTW2GlhXfg+AHEthbFztHaoQh0xL2MUN7LQzz9+IpzxCUJJ
tU4qqJrbv1ZPK/XigXHJmO7rNcSlEPAyHZ3G7EfNviXDUP7molYo7kkp6kApgNbPupypKcgDcDlM
cIGMUhyd3ipTUFXMyxVVLvGR/H3s21xmGQzw7a9ti/JgwsPbdPA1q5qTVxnf05jf9msDbhTu+pgU
Ly5GsF0E7AC+ItFEd+X//4k8afmGYKoXR3giRfC12CD+SM2ameE2CEcLOQCF+w/0aTkPLOQmVnEU
0pufMaQeW8TlSuWdtUBw5E0tdP4ybhET/PsjeX/2VWnOEb7T/TDjmdi6FDbkAYuTKf3tls/84WFe
dRKGLrb30C1Sa7hzddip5DFZ2jVHb+v8mqJcq/48/8Z4Se8PhCSrMuuXuhjkKExg4f25QEpoAIXr
nzRseAa4rtTVBulU6sxEwbWtwhQEMju6lli4MFnuWATSNPxgKdZ3/nxHSvT8x99mvYJpv1HECMa8
5jSt4pDAP4H3SItJKSjqapfP+jyR30vp/eolYCzg2umu+8AXWhIYYH+l//HcDqRQBpp/6OwY36CE
cLv9z34NGJME6rD8yDO2KT37JHSUJdLlBaYU2JShTFXxQsTqVGMpvoyspsZSyyjRwjgbGh4kQZqh
/xPZY+K2+FMitKCfQkKerNYDq6uWIkMuwt5PB5fGjfCxnqtHghXS/oG+jdEoSdORVrL7KyNNrZMM
GGXcUU0A4yt7Ma0Zu7ICOkQ3SDRI5R+Ax3FOaH5/pa1FfHc79hF76+240L3NxgTQINds351Q2Lig
BKlCOD2I7XK9jUepcFJcUnT43Ti2KHfOxGODi0oX4QW0HW0ZOmC8hd/RAzD6A5qydKqs35F+au3k
qSdEC7/quJb59yfdSNf7jWlb60AROTdKdBPkXIiiVyfPRUwviXRmCyvrYHMxIxxcwdPFFw3YgOQl
dkGHIBRP9x+C+UC5wXhZlmEgtujs2Stp0FkecxqZZ9irs+2UmQKaRnEirbHfRYs4+YXqPI37lEMO
j5J/XYs2S080q8lZLDs4cQPGT4mACKC8Y90zVhviFd5DB+6/Kcw/tGe0TrfXSc77yom0Xo3s0gla
PfFJJ1Bq4bKw+YvcLO99wR2k8OSIhPfZHIUrVpuZRN8xDzBdy+Vv0W1HZ5NTh37p+V19s3PMPXKs
cQrRe6ujLPw1VZBELhUDzPuDu9GjE27GnevnZI84+oO1xlhMrKMCcwW9Zok5a15jsGokXScdXejI
zjzye9Cw+t+kZJ6UBoLTfspbZsbCF8/U3Ku2ww5yCttv6nWtBREnGnDe1cqTYv6GuYHQr4u158Xa
n2IcQyMabnJ9UifeiwKWel7c1qPdJZulBCy8fqDc4jHWsQyad/nJdYm3vLF0sYa4fv2Lqx4itx+r
JEoff9RN5RkfyZlmnR/WlYfCEzO4o+ifsUU9mJJx79AxzsyPH98qWHdpvqVR6ERWZBW7kqZZCVZJ
/8EYaOZ8OVuoBl0rQpEuIDXwFiNC85xpP2dl8WbjyCdzB+Tx1Z/IuPVYYgWSfDcuQKx+INZ74cvg
bByT0JU88tfVfyil2uznFlNBOyT37u1BpCTv4s6NQaWKLW0DY6fhgn1eXko9N0P/HRXWm9QqEWhb
qbo+XLvxEHYkTJe1MlDabVq6/h+A7aI84m4jkXjQSELLfjh2XcIeLQucxGClFY0CG0kZOeK79DB4
PSpAQ+0VmXFeUCEcnf+MHlBfYfW6SlOyRkmATh4UvI7g5pWcKQ5x+2r+bMZgCSj+GqlkbVsm8+GN
Yh83kOjOD1jHvp1vuitoVUr6v1sg9buJd7e3Av+/4X2tscfzNO7YJtRKe1LAwV00IgYoHIQn3wYx
BiYrBPnPD3WNXAufng47qM3Hfn15KUSNw1OywuPhxhe9Z95/zKdWMNU9ZTmnTcR/PQ67OhbVOCva
NOdeTaZqUs/MKCq//hDHI3IaxiCBTzQf4K/4jUA8mO7cFNkF20ZxaBgT4trcpRPQBOWGKvNNQ0Z2
r9CdOsACHukCHjwTTrpcPNMim8n1xOmuWXTtFmoM2gbj4GE43b6KxWkCElZ4djR2SbzNJ60EYXxM
ThLUn4Z/NDKHM4GkRWG1mJWje3OqVdu2+SRi7xxohgPB8KvHdN6FXgpWKH8De22SN+zKsnn+RtPp
gMP0krPaEZg4Dp2RJFx4OUhNd4Q4vsM6x/zStl0D77/BpDgVZXWB9aGCENfSzHZWJTtHn8pZshOT
SU3EJl2OUqlyWqVyeT5HP9kJUU4oNkAVhpE6aTQtobsmWMdvu1WVqlAx5upWxjtXILDgFBUodqbQ
/k+4ICwbLMoEF1OHRnJNGWTlYhFRYhqMX8YTUtnFEsqUey4eBytpTIIanJHISvCMANBDFI3A4aOG
C4vJAfER726ys5mnQJJjWQK9T1hnZTQZAJdX+6jMwUZJZXjnSnH2GJzV5Ze/5UMWRFIRrUm3ykcZ
NJ++bE+bmWp0N0NggX4+ZFH68MZ0G0ChNCqK6LMHvUBJOr3UmHpCW1ZM9w5Cn9bRs/bW770JHOse
v198zeq47PqGEv3s+NHev5vWaT3sUFtI3k0fDWf42ywX3YCmO+LbQnhy9PVGarAuc496SIjLNScL
pCmjzqrHUP61XT5j0tbdnXQDzEUZ8bDZuoObpTmaqfOWoLjQhhZIj1450prwPWcY3ezEpe4Iaf5I
+zyPStIYSFyl7y2/WN86e2/zXtRf5JZXypJ8QUSV2wcqBy0R+wKGu6AuBNdUBUHvmZN4I9wSwZF4
WOsHR8QEmk+UM0DO2uLuFenTPn8QmkBoBWcROJJPxcPpi9n4k/cfSpmHFCnZ1Ntu7YPFKZAmArhW
2NzSBUMolvAZ8rf9Sgp1Bam/bNhCh3R2quS0bhM1rgbNc0XGnRxnUHh0ZxhWqXyIZjOH0qNifcDU
IKgwRXmSxcdUTLdX34WKv43M4OB7bv4Ib6PJLkJblYpCTESaP53N98Cbjh2CR1dIjZohR9iwQRbw
IgYxO7mGAedPBWtVMkG9zF2R6eiDgO8Uj5WD6EBe8C4sKu7uGDySkVb/Vmnkj556OIZ6DL5GBAuG
ujwQY2bc97nCsW75VaOFN8RgURdPbOp7V9OkRmWQDs/kmbud8wNzA8pHHr05QBdCiJWvb69itUSx
6klTRL6icoRBhaCwp63W+WKkcp+7xwu/pAesphHUCw7npVOP8O05T+5aY5aOHQpCjtOdFE0s8fDj
/fEpg8xp9Of3mlP7we6mDhZmrwNji74cNflPdRxTUyQrNuiZYhSDIfIIu6yzBSM8+1CI5zkV9Qo/
3xU4nvk77RJkjMpdBkaEvX8oyCePCm1gg8BcZFveE2mzlojOCKy4AFKzE0RMEzMppBDFW6mxzFOr
qukKnAHDJfR0Hh+kFwvYZt2NJG94gvdSxPrBisugx2zo3Crn5f9fuDw0eaUmsoQEM6+mHJWaa/yj
jw2aDRxsiJOHp0VDWMfGcvUBykHu/DHNTv8fW2ApvpferYQj0JdqGRvH2O038EyxinOdLPf5AfLS
oVlRsIZRJGDUeRo9+iW2sEoYgTxKy8MKq/lAN5bjuNkEfwBG0/UdgIDKZlJm11JKobF2ohp+gwgo
flu9d++sZgy2Iqtbd+MYgeIIXRf4Ql2ewdAa6AgV11ZerOW7g6IDNzv7rwtJdUXfxlPCLjJcGmKR
UtCnhQezocapcj7cnaxRN6QB7pd/d4dl4W3Jqb2gF8Jv48eKiYyseghRewzTI3WbDIs7nLHpaOlJ
BzsW34DmIq8RcYQduQ7PPoz0y53v7NTyuSbNuBZzCgf8EwytH8XUL7DZ/3Q+l8g2A0aEMSNM4ouh
aQdWGsMsRjPgc18FCfOfzHK3HYw0RPo1pt3RFMCbM6TtQIVu23X7FCtxHW8+/erXieWUyoZyaRc1
Jcx9yHeAmO6T+bKmhUIqArhAxfjlArfCVMda/drpGKazH64dA+YbGKkk/IGdLNkiS39RDNlehuBZ
4x/juJoKkwkj5zGgefMgCud8O06Nkrzq52/v258z0ad/unVJDZeP/V9yoCawFK528wVe6vZRoCQf
wWRr+9UmSySFthqHLGlgh34edvScCX4QYX/1z2lpFwH6HeMiSY9FycwGok/dbZ6lsYtWR9BDj9Ud
iI2e9mEYooGiUaDite1W6lOVjpkg00KQ5MjGmkTqdJDWeyRKU6+8+IuCRAaB4xb3ut0XIFypLP+d
vohXvuTEm2fBrDgwqxZDewZ0KXasd0ZJW9TmNxf0Va4oLSPsJxoLh4jobn0aOgoIt/Sj/W0sqDO7
Vx3JIxcscUcEYELN8emKS3YNfrhZHe2NfCCCo5ofe+GfJie8EmK5zvmBlES3rJ6MGt6RldhuSn3J
5HGRlS0U4TOIYn3v7b9rsyqocFMP0Ghraj8Z2wR0IgxIkjlE4nh4/+O/xcXZESJGTIR0sTrxE6bF
u+PeQ4izjU4usmIZ1G3v8bIhBv4uDEhieN/3oH75PwXeO0uuUZPSD+a8PgmW6b0+404kvGb7jmdd
Lvta1U5yyk1MLRaVyurw4bAwPUXB9npTTAyD81m7nHEVo4HV1JmbUrgxD2CIbdDV5En2CkAW/MxC
yoW2/L9jfg/Tqr+ZMGrLfPJeitI1crY4BbbeeGmLq4FjfvtbQJ026+r1yIPFvRJS3fjhNnDFL2+z
FOCrO1j41ynJjouugrGFAM2BxpCk/CjPbeyysP9IDIPT3a4tAQLP//wnSbhfFoHz2HnHvHejU3Sr
2zhsOFg8cJMntKMvI3DClxaWPqB4hQeRZoXYhJ1Iq/+jBiFXAWesIjoSYsUrVAqQAZ383YepC70m
gMmqE7T5cx6K9BPn5OlGk4EIiz3vrXGOfYdrBwCbgYCjilXmVkHuBXmmx3h9wvb+6Rtb3Hv5nrxJ
GV190+pRiIq3PEs6Af/9GiigG2mrH4ju/luZtBbbMrEVriUXLWZVhILe+AT44nlQn+z1IGjaHeAA
Hi0r32k4VV5r4KpgfQ1AfMEV/A9tuHndfcdD3gMWHdq9H5EYgsxcm/TMG2VFwIdG43IFCyncOX3r
MDSc+JuTX6bdMx5Q6hIv3jynrfqikjpQ29Vz2TkT+h1vfF4CEKu1YnIzairfvA4AbjLjS8r9aUDV
N3GV6U9R0hH144lSeAtU1s5LBKml8JqrRNpg+bQkbnv/OK2QvrYak1/xpv6COX78XLFOYU170Jtz
LlsFnZOZzPwMahoDV57D1KoN80YUfts1tVC9kxRzkZgcuEennWOxiAOGWZAZhOnVVifUexupLlNi
+1Qxs1XoOeiQ7rLLG9Lx+QFLvrk3UcAmT49qYi+oKhaKQu0e09V8HqvHPoCj9Wtgk60BTXPdbV6y
mVT1j0E+qbVWY6BJjqVQTpUo3ze3ibOfoh+4lrGocmQgOcWNLv9FLX16dV45qjl9tGN2swLBH5Dp
j1ImM/AXqtdEcRFu3CFojwh3eEOuAcjim5vlomvfuPMO/8U9c90/pyfbYRjIxQy9DpEzb4l5QoHr
VquoDduHzKRvqqaCGx0SrwM6kD6E7eHUwq033S+4ue/S9jwsxnnr/QiBVRror79RwVvcyw9SS2x6
PjJC4VZuQrEnAnxPzgAaWe9GMImb9f9j8eTTvUW1mTkm2cIzj19bz++lSpEz9CUM4Ibtxu4uF1gY
mt8Ne8XAMaqNfEsdxmpWI8rS1iDqNxzLXY3bXx0DbX0KrMpamzoz0EffcXBFFjTmtxQ8addFMktB
9DuARtFSnmaLr/ry1ct+W2iaFf5hcaT+HHKVtORz7LxZG1EWURVXnIlNW5x76kOLRpd1fJ6knLRR
JhrFKTOv6UfO7eD/B4Xn3vUHEVB3sp75/HCYpilgsP3U3Dbf5IuWaPKRxrqJCJYWa0JSzWwhXNA4
m73tSRK+RF7Z3BO+nfTwaZHXfgSDu+0TRUindfH141cI9aw88kxy2zoMbaTu0EpZPeSYQnlbnkS2
kDGvCMI9uYoOj+zUYYAQ7OplKZynrNo9xJGbmVJquI6kKlEzLTL0GsJ/ritwUCgWhDxjS4sZtA5J
TXWWDak06jdRoyacHd+mkTOROF0XDbrAODTiNtkx7Qgs5CerEmuJNeHNZ5j4o0om1KNUckMUcMM2
tNHWa3JWYOVUqdGTiXcJqWj8PmrF1NT0TbCIaPX6O7qAiHMSOx39aSYhQ5O2OqX6I7LHSO3VCpGg
FGgEFiPsgNNBLyklqnHgZ7MgpQg8gIrQiN7tXmnXgmZyE72tjtiUogVyjrshfQ03suudN+sTyzZQ
+ByqqUEkSemaz+kmsRioxaYK/BzuURhav3lHpa5cPQ1HGpr5iiF7U/5zXo7YMxhMD/XTah8VRioR
nTwbmlm8na/3miju3TACFHFertnKDP8eh1ohXxijuF7tnLwSOjfAkMKnbp9dFPl9Bvr8MjkGVX0/
+8h1QefDgOcTjtPV4KLjc0mR0PEz81VZ/sS8t79KI16NJGhWEh1ffq4XVajHg3IrBsE7epBSn+Nu
lPc89PkGe3ZhKd1evBBlWIqKYIK7+NlM69kMk7/MjV3tax4aQyQQLpv5MnJFJ3FBL8qBmLKzPJlh
0Pi1X+4ptjgod6GmjpHrpKXRl/xGCbrdh6gqBKgjApx+Z2HNP1768F6SItS0WaOC3kSlEYE4Lr81
NQieAv85s7oAH+KR+4z26ON8JsV72dXPv2uOqQ+mPu6GOospJuYfSmZAhQLXJvelQ3ZVPu7A0vu0
wBIxMMZDrKvuO49clFWRs6JX552Bw5WCiiJT3hVlMxdZwo1JsRiBcEf37fqkV7EP5qecadNcPknp
xy/2kCFTbyp6pS7C9gi/64vNp0G4+ZT3YrAOGqfJXt67do02otPn+RuCKIaAumy62yPQW4lx+GNi
aZHAohgMV6J0dlSz5Sv2KuVAv1+ZUQVGAXRBuYH4JEgScpe3IxZmVh30NDqB9jJTQ3DQYmj8pShD
23dRha/Me42lFtlUvNTZoBJxU/xVwf7/WGAIJyo6x1GRyxkS+AM8vSyB/zzgLde/y5p5NTsA909c
X5TKh/GZVtSmvNExdTqQj6ERO7duUZpYzW/Ybx+ng51Wh/UHb286py2AvJ+BfC2rlr2u6t/AN3GV
wmgWNw7Xi9lj87HRxRFMkjl7TIsGIZOyhv0FHeYj4uC/6ZenSQVGiTMamzUkKRPiscgELbuxEyzT
lWi7l8u9NdqzymQmpYalE/VcDq5eYmqqgCctuoIUN4dBAYe2XGgJWyHUz/1R0eR8EeBNt6O2AhKN
qffY9HsbD/FaLtGkVTDVsrZl2JmhF+KGRhhgPFldcmo4vh+2ZPgqNgPNLqTY53eUu2Oxap+W4JdU
9kf6hico42P4EcFYUXjm56YgKK2GWkVLWoUJxRWrXTb4Zc5tYG1kRMHqmTbl2W7kdne8v9RnV6+R
y1gXHwXX1kDHTDqMtANILbNXcI7Sov5znSeH8BUSfaeXrrh8xG8JtXmtYWBUUyU7ALgWqzzpbRHF
2l+bncWj8WbTzZ7P1JetUiKTRss4rMas8PqYvBusCfRR/ETiJEndrk/TNC6i9vgbIK+FdRFEqZGc
d0EZqX4UG/VYBGi3mAG+RUqX9FJPwE4kSGdJ9udVN2OD8LP7EhtyK57kKxBXRxiSQtxcsS3F6MIh
i+cByH8HXS83HNNdAXgPqKnveJXWe1/EB4UalAeaBaRmRvdXeNUYftH70pMTrS5DvpNNyqoY+3PT
BMSMhmtI+7I3SWNsPABJCk+3RD8UrS7ETSSaq60S0lO9T5V03uYJeLWa/snd33ORmyLEWhAjtfcO
v8gQW1ju+iQ52RV6a8xirc31wt2QXyhBXBTVYzzmiDxda/1ZwnBpsxmZ+OIe2vu31RA9gWHY3GNh
a1Ose56t6bHv3wQxVwMnMCS7Oiy4R2hi9ryquiUU6ISBscA2t8LegUVVKFqOfB9xJMCVni4Jywtq
cWXW+CAok24W+rdsuYGpU8RcMtVffUg6azDFvDMUvqW/poU9nyLv1yDQf5binNpyO2WMXYUJU7Nu
vsHtQvImSUUdsic6ZmdQREq9XoXJNDskK5v06bp+Xru2v2oZaOeqMsOBDBr28Rd+fA4/HcB/xOB3
xV2zyp1J/u8Cko7ER5th9OO8TM7D5/JWS/f/mmGb94mRsg7jat5WKnTJS9wKlfP3eoLy8BQ3hVUF
rEG5lzZiE+QUgBYJ0ynRLpCVISmWe4Q2By2qmNskpzCMDdla0w5c0c162dOF4NlxANF6H2jBFa9Q
pqaXW7JaVrFaM4w5gaWp/jMHmhdH11QswaEIMI9rf8y25NtCcHgEgoX0UlGKWDKLP7v49yMBXOCO
tSgsIw0IuFuwCHsx3OQr+pWEamifcG00BOqoAZaxrYLOj/MJyq6ggJWvv5wwSwIxlP1Y0sSQ/rri
xNWBkCcYdBhxXXP1isMTzh4QcZyMLbwwFm0H1JRkbf/0Baud58bTD8wN9ObptjK27wblP3bWCV3/
Wse7WCMzwtCN85Yuj04l/+tFys6IyoS6KNb94UgWw1hw7HkubEp67pA52iJcT2zil7/eKbQHaZcx
xtTEzEF9XDRKbSy1CypUHolsnM/b4vWUUf058Rr00harZ68cIwv9MBwuoV8Gxc2yvbz7Q0mQUc1j
AGFXrJHeN/dUINBswIpeFj9vIglL3S5YCzViH7gLw4NJEbh7BKIiQBFoD83j164O8DNQNmMXdM8N
msDwzgv+w++DVZIllRA9rBJfzQR1WGw2HSMF+cHbkkwTaMQT0L3+mi0BzowsaqWahCoIRhVMA+fg
6WdukTNsLAS3JypSvFqA9i1fLfabhvey9E2GZVerlyWRDirntrbKU25UYKvXEeDTOmadNWFvrRaN
vkz2ShklsKXeuDUyQqgUfO4j3rB92Y12//kThdy1+dlb4U0ihMhSdAmUEzvBaGYTDdf5X8dGVZIE
RLn3qft8oh4FbLwu2ks782wVh5l+u90NNnbRcjMxv91zixTPQ5uq1AbR7eGhrFSpu9J26I9TrtFi
KITUE9ir7sPTCoKOTjhBfFpGKwi9Q1lOGPUFT/sMOw1yzb6sUc1AQHbkU3GfyVCAUJI0pO3yswvw
XFV7cOB3frTcY3Ie3cnrSHPhOz2yfOot7NmGdy/JgAvDsYjrijmMqw2f1w82CIl3FqXyDRV/zqEq
7RzhEDj1rZVFZM6qPr3Z7B8CUz+cC0QayWfTe3LeyQyerMWT8TG8nyxxtQdWmVwfZXIqCMszuAWU
igSFGdDXibHEBBerlLA9CFL4cp1HX2W1EfsbGQfsitaCyIGvREgTu1+8/AuiYF24J2+pPfbVdb2A
w8E3EbZU9TU+gMf3CP/fev7hJvFuHQlY6pyDuKceUX2n83FzL/MobUJr10DG86ARKF3NyG1ZdhQd
YaTVHD97e2/BMqBwCj1VVkuz4fLwTjAtyhG3IFjfT8hSx9EJx1DieC8e6n/fYtkfkSx1ZxQu2Mta
GR2EaV1VzPo5rNYmMnDgDbeiD9mzbZT4wNBr/Nchi7+oeWKDrULi02qNb7zC4rtE+Rf1hUvMVGJS
4O8Q+WaDh2toNZnrxMGQUvBjN6mMa3fZIdgFLjfcr2kxBHTStiJhmeMemdXz4AfEiun2puDkAr1k
/SicHKcy81Ihhee8Qm54aDLW4yxdtGdFfrQJQKAa+mYetQmZg6IH5i6FXdpL7KT/l7fTVYLvfmcR
qiR9oxdHZ+UtAyN0bgkWBhZATgfmsGsnzgnFcgqVgtAQYSuDl8rBg3jT4x1IJ9Zrj4mzzBRm1izM
IVn1XU2V9spVd7qOIBodhu3HR8d3SIa1IXYFO14qDSdx8qMt14PUpZI1lXdjOdte4BG58iMblxR3
Zyh/fini/eQD9S3Mgv2+c6B0+d/8pgrEEwkEeW5rL4JqP2P8w+q28J18Y1SV0VewkF/duWaQfIsv
XVj5BS72lxaLpc6RDjJo8VJKNOOHfUAcmfxhJDhTTKKatzbwYUg1Sk2D6/aYUb8QR78ygtnHhX2d
xtMdqRuOmS6T8yUmcVliVoN160ay5cjxZpbnm9gnUiHSqI/QfHIfzkejywK9bLJEBxABuT8sIpwP
18TJstpvOczWiEJBtd4z3vNkDwgkPMULXZJkPK9Y3/EK3wpXRPTS3UyRtS2YP6JydXQIkMJZO3BM
1g8TwWB4ALlde7gIy030nTkgyLzTnt87Fhqv32A4lwpwbZSAOysrnwMvC70OkfxGKBjnQ0hjMJlq
C4udOL3opHBE5uYybQ9hGr8bsbH3VUjA7+M/nLe0T8/zXAyrCvlCyWvW3Hh3gYgKi4EUDIjS2xlY
3UCtrnGkfaAZOvHIj4RkAOAD5Snnq27fjoQ1RHWAjg9SJ3zz3uh2UOIMOEe105lZ2uWhICmuXeXK
qn5ANisPaVyAZV5hNFGpKmn9flhHvUjobItVygDYfloV2/stPjwctplNSNbwBZBKQQWBuLdhJVzC
LjAtzPtAfCQJkH3yN7Rwk9LXq9TJ1NWzoytRqHvTwZIyfI5mOIBKNdVUvaAg9hOUFa67vZ9psGtp
l5/aX/IFBVEHpx1tZIvPZPHVnkkvk8kCSf4xsibZ6+BdA+Nivun9tzgxxL+uh3YZE1HWq5vfoyso
y8AwtRNMAvC7eBivOk3Afis70yCHauYwYP8tC8l3JknGSr9grk7kUfrcpRdzWHOtAwt4OgpY6FTI
/ZEfSO9AD5t+W/eWwhVUrHGyuWa09thYmfJ/dN2gLdGEDzdgrK/J52OkFLvIUprsN254mJztSoi9
SnEl32jax43i2QAPDKM+oAHLS9tAH6YpGNTTl3CgjFLQSLsdD5YdSXX2Rubvprhlf7O42lXi91aK
7mSuuNyvKc2B76p1KJgo0DItqWW87X2xfKmaS6hntRyKY1CPmC/fkn/T2RuJUxYAxxFH/NzA7eY7
z3W6Q2y3G8mbGwRHmafzxtMFUegY4Ysw5cFL6s1zZt7sECTN6RY5wyxlS45GonzPfGEp3b24lqpB
iTkKcqtPKtTg373BLnjwFhbv61wvjnvpdHhNeMvqQHjC38wXjJT2QHqxfDUYp1houI+LEP71faFJ
V6PTn1AVTvktycrPKh4xFyWftJoOJZfsAmzGfXcLot9nTEcvg/pw7dy0ZUnNLCro+Jt7skALtqcj
h/x0AGU4Xcvy7Sbpfb40pF9aWyH0lZrouOpJXZtrKT+VW2htqkJo/4Ajl+wSdxYgDDB2kj7blh3Y
5ZaOEOKkmnVNjKvdRzjoz+m2By9QmlB2JPdNKQNt2n0ySFAc1mdFOxGvB8Hmdy4WkeC7LfcUQlVt
7NaHcRUYN7CKLu8Mt9qqFVHh3n6Ub8f3IFLPNFIYvq9xdQKzhyarVMvbWfwh4E3JFviSyvbTi3BK
fmcd5fBkSYxHfdeVr+ZjG9cDYcN3Gw+v2UKS1lUX+DHkMS6pJ/f3dJa/OAV0s9uhgRtkYNTMiI4y
2CNHt9SmFuAwlKLY9y+wLMN+v9vwWN8Q/gSjesNx8Jnjb5wo2ovjxHQqYa+IbBsRLKrvzq3N6g64
3/L+oe92f7dBXt/85EpHBii1TNaf1a+Ha0PbLhDdc62w0kaQ3YtAecvItK227R9o9AfEQ6dHexTa
dF9bRQP/pP6MZHxeSvMLbWllMeMuE4+NspzRty8UUSOJcXD+FMsXFqLZj4RutRA0lofPEDtA6fwJ
bi8BHusn/FqZwRfxDuzOXGaOVtrN2vn+uWhcqy6EWNp5of4naF0zQHpJyaR9rRpYYmLjuRS9Q9ti
roA33XGsA2/Eay0UHU32rbiWTZtCFTxpiQZXMDJbUhzQ7gjz2N1VbT/AOu+bLYjB2AhlTomXxSv0
QFDUqJYPZSn7jdZg+jfe4j3m/aLFbJLKeZoY7I47/pwZ2XMW2IYR6YsTfKxlR2PQzEyV5Gqu+OIq
NjzUAjwd/6LprBkADRLqas41YB8lZ+HOusAiSxnCPd8J30fkhjPxTcjQEw2efrwSZFSbIOGURF3P
F3v5rzTPWT7QEeQDwwrVwDwj5OrPS8/V1E4Xg4B4rC9X7EASO+c/g0qxJZtavFOEZ6vyoUas6fnM
NmDT+hUUODNh226hk+yjMM4eyfFTPX1wG/sod4VfzQJidHiYeC3LtRKBkImtHCg/vZF10sBI+PR9
l53Qyg6dz7MOSqti/lgtsuTNy/ORYka8y4pq+hWrNnLSMCvdQh/qGowG9OsVjmUO0nDcGBNNoE2h
Y5Eaarqxcf/lQ+VElKasSqbBRzKWpbQa08+ExkUKvCak66Ji+C2s8hzoUkLg4fxZUpQK/feewrSr
d8kgipIPWjCYNZ5qnWL56XZVAk78tCSWqyVL4px5OLS7XwUI9VzdNgyheshLgaTlrR65AK74A67y
e/GaG33XOK5ndjwnUSJTZhxf73dkNwMkzwX70/ysUEJQ2Pp0K1t4pd6aO7lSdsJz4kV+FFDhFHi0
NDW2mr9gQ/cGkMPpRYKEOEgjBkdY1tjsEj4rU1xuf7vTKb0qesfS4+gulKY28ulkXMz/dv6DqGOp
3i8AUOJnxbWqYpVj3nR3X2OyiCaEKBTwGfv2Zo4+Cxz+nNXutBfTTV3IZ+HYgU/7XA1TXIBgcZqb
ksznhjZ55r0y2BbHOAVMMZYECu5vAguxp353DN1QH8VoLX+/00W5mbwpwGD7YpIWvVnMtLpjnQFJ
5wDjhjOC9BgVd5aqSX9epJ48b/q16ZVRRHoXRO7pYMhXPry6TrZ0VoHolMAv5RfXbeug8EQvH456
H1SPt6Lb0cw7rsCdg51k//CUgBHHs+tfyG8LNFJaWW7MovWozsUdIUxRHxpnClO5tCXNKW8Omeum
VVQzJR81HnM2gXTUCgtBpeJAI+SbSYR8FDdiszuIYDcLcZwDNh12qjQDOOYKIFDU5S/Jiwyv4xDg
LNV7/86pflHj+31XKdZFNj/av4VrVDDatL2KedTSsN9mYPdOLa3hubzTzy2rUesfVSUMTfK1Xhuo
GKhOG08zp05/t1BCYKrKone+7H0IJbfQd6/nHkQkZJdLyAE2y6KHnYOhI8YWveONcmVtZp+FpAjC
DaScSYAtNSIVQLoK9CiVo/DfPwb/RsT/4nDHCQ7/jdrjaYfC6ZRD/5GmJLIjUnDi2/LfsDzkjchD
BmtRG8z1YYmv5HFrr4Erxq50qQN6iMSi7WAv0MFUioDZaAYSQyMf/KruRljuBXOdl1qZJSEeaI0X
ilaN3RYo9k1vXrji+VrJ2S78EKEDeru3U/nXvSGPoqqpBHNAS7RaniNNq+4SyxWXXf6A1TL2EQBQ
ocrwcTDx5jIW/gf1Ejz9DQpKYsdZpvwmu/lCiDoPLw31qYME9X0bR3qdTht+yMYCPVbk6ok4j6mK
d67oMw5WgjyWwZ4yYw1GvCwUca0R3Av52GvPOg122d1q+I6J9Nx+x6rX5Yp3vfIP275G0PNL1UEw
2zRMbdHGqHz20hu8E166o112ooq6HPgsERlwVfeY5sNUWkg7epjyxl0HnWdXHaMAoBasl6vzvOdc
IGGO5/P8Qyp8Evlug32B57RBlRqy/c3c+tj85/ZHNSDHF1EZtWUOk9CjDX9lLZGoKgyrxeQxkRKt
Ahx50tb8mDC+pbHXi3UH4S7LifFPTtmlVi1tQr9C89XDKQLYgGRivi2G2p8Uw6NY7kqO5STj08N6
RlwR1cRzPYCRZyBUv4RqGx32HuK8P2zLeedC3lp5gqEUM6Z/bSmOia6MMnteO1Aml4DABivBudWY
qd6izgt6kDZoNefrR03L/8go6lmcXRtmEWsU4P8eEJ9OLTr72u8Q/jfor2TKgkOjbaGhnQsYJU8V
7QSrbideJQM0prO3o1cTLw5zLjuy7+aYzgreBhmHLURwsv+8qw4eGzrNNNUYwn6Yhlv2ZaCPjkUd
x0lquTJRVGdzhTELXCNEFjM59jDUHbVKhwmYAR3YRbDoHZZt+t8xoUw48nW4ys2U89c1xhuPmUvL
QAaW+5u7727llHdNjEj3rP92m5A/v6ZAa8N8xgXXAn6EwlfVzD3ITzM1BwJgTTPa25az0tHP3SVT
qezqT2QgEjJr0zKefztUjDLOAY6rEWy2LmHWuBl6qhNVlY/pjlR0WkDovr7C//uUDxyt11z+udN+
5/Ej0dUPyqfcmwLllm97t6oXaVMcjUpTsEScYBi5sFcFLULAzlv+0OgshVbYSHOybttBPqYjKP6t
DfSGfaiHMqf5rkitCO7QATu2l+f+2CW6zP7Ulkj1B6Oe6ZayYFfmC5gnAlQJhI/KQLjIHBvUJ32Q
TX4w1Y/EVDjXiOT5XRu5PDs+ygHQYwu1FUIjbti1dd9ZSv81e7c+lNbh9OHqLYPAf56cJR2mU6Fq
EvBwys9TQY5ylrt9a1kAfgU5BmvqppgBBGZxAN67wn8Ur0f3hF5ZzV7WSxYFxqA85q5Mdt28lQ0L
slY154FuhzjiaizA0MEL1MDTNrCKWywesbalJW6xAH8VfwhMZ2sVETwua3S3pYZTTGLwFvjcVauQ
gTj5Fw4Hyr/NOPJd2aISW/QViELjqrBieqPRH4TUbn5j+pMbTtpAff8h+E7qy+fNpiOfPzJU9G1t
CJpJRgw5jDU7YocNIWybcrnZ0Bezf6XSKsm5tDPtv5IyqFkWWW/jgNNNLzg5M7ZoDh9mMCEznbc0
9I8dThMe4xVB6VfVRhjgOwSqEIHp/z/RrdDis2BlPqcLypNavFyz8FhsDdrtzbJylj4xKcXnhXr3
l6wrzroTFmII8t0f/JBzVeAAwUYPioYWFzO6skQwAinpiifoNHzeTRKQ7qiIpQZyDALYSFIkYEUk
nxwHgSyUXzozVQpDeNjsIwFJB9xQ1lWJ3ruLdyIyhvkAIs0G/L0MM9SUz4uH8U+F3mTZDpL39Neu
Dh4y22CR9upnIwAHWbmpxR19jNb91AWhS9x5E55VwIzH7FWdsv7NhOFzy1RD5PvZ4nBk/HwKMPip
D3EoXt/KJdqawjGJtyLQI7JSO6smnVNOJfrf10FxEPnETWelPyso1QuDYE/PKNYm1txuPpDng8uf
yXctHQk5lazpAflTV2BA7t26jR8oQw4xPkIYN/GWPHbnEHZ5egnTK08f/2CpoNGvt6D0m7NjeL4h
ylWsyiTEkIknjlJvvS+bions+iDCxKFzJ3jEgul7AYuTYsrnNIVvEOxbw6/rtUdTfhoYSouu91k3
8J4HgKaqxQFJLIAIkdTxZMZ4LRfhEOJ8TD4ickCTe/2iAv90tvIegF7ewlfnCh6ZQiORTwYwdII3
RtjfaT6cNayFMRUdWtk7jwcTDIVuzUdyFkdTH+pcrC1uhErofwAJyDni6HOossD8BoCHDmxuAZ+5
fljVzkn7DxIzSVcOeg43Q+r4tC6q9qvcfMQmKHli0XMuk5KXqZwYYyVMDeEZ96pqdm/TdUZriUcq
O6HmmNfFini2tIQ4mv2cAcQqedpwVfeK0PQoY8Bm8cHQFel2WTJXqn6z41Y/BfOahgp8EnFO9jpj
LaT5REp3g6l5yc8ssN/hnCsPhnd6G8Ff8OK5oV1LFvBZtptKIWMtuuDgQUoSJ9jg3bDzopd44uki
svKM2GrW7122XyKFlOfQDepuK9WO7K072Rbvzi1AemjyRrFVdV3wRMsJJoYG2tCAf2h8HXwnaYtk
0LVQlu7UwKpY7ZY3KUlyTRaEF+AfIYRlBEAPeD6R/aACb8xVJyjzkz4zfoKeOdMfkkFnMq4em2yr
zPXLrS6tVCmJGx3FlLdcpxmypQdDWhWOTwTRe7DZ6OppL0bzlDsFq8eRfYXWVQhrHy2qve5k8TIe
Xd7Hblqx0rSj1DZpnqjDOmESbN3OtSraKMjC1abX7cim1uARgiXGflTCHlQ59qXzdFKG5STBEgdu
99hTU5C+bn0sM/3XvKkaA0HjYbwtZOiiGK6LT3cehoeYbPITIJZmZXounCeMm7lgfpLyIHM3TUXb
hTl/ix9Qfxzv1D3jEDmHRDvjbGrNkmZou05stvM34YrDzrux1Vo3CbT/UpecIxtUyCo5MDDDXbQa
WeAUiSvfHKVPCqctw63+yb2LsQ+Z+75nPnsNAQFNYJUFaISzIvzedgkjdyMP/8Dbty77+iQR1D/A
VO1Cle7wCDVmQ1LJrhaPIuqsj/dhIwrbs4f2XYXJ1e/Pj9cpK6Hcr2/EKiFyerMje43UYjYeoLq2
jIal+NHwrZk0X0cqtdJlM8WPfGc7jDroZ1iotGweO0NUbKjmn1mog+6KJ6YexHjT0OVgtR52IEld
XjMqqYNvsdwkkaZx+7Z3U5Z9Rw9g41/neyN0rJ87ZAw9Jodx0p88V23nzKPbBDUGaKl9o3b+Zx3n
eP6vYfV4Rp2yJxfaK36cvjvTp5dQmT8nzVdI1jDuHKoi2Kt/Szl+NlT4frRkN0N1N3a+3SRwucty
HbepyeOL9w0iHfRdtwAwbbyx4huOvVTMWKCL7vgu+6kkYeupZShj16wh3JWQpzuxoF3KSRWwSycB
PXi8/C0bDK23kVHUOMRTzwTM6BSa/Fa6yC3WeIEE0lAzKXuxGplZgc9dFcZwHMu1UxNGcvodh/od
1yJ01KWV9iu4Tv9q//P7oQlUYVcnmbbRnkM7c1H+lshG+sWqkP1GUyah0ZZfyrSFznqu60nUOkT0
stjNzjk/P4kN8iTDE0+jUYL+xNGFNopo1Fa8lsDTyA14KYKW1Nv5Y5jWtJ+1lYViLbYREpmwKpkW
1n/qIwwgXPuxASJpcx8pUJekmIjUxgM+Czoj1UcMlNEkk9JobgbfvqyEPwGUbwWWjID9znNUqy3s
rDulYfSxxn3mYh97hx/b7quS6r5Sfezh3+cYekLV8dfwRd/6bHy9kHx/m7gJMBRtvdIR9X+PHJ+y
MRHGJ6f71ToYPqBwzwX/i4YatoFaQGDk11oleBSQYbgZhEePQNiID+Ev4zH5Ov7hEWZlulfrRDJB
8L3wjTYp7jAFJue3j9r7K3IL7eIvGuFA7dbMtJzJTLq9cJ7RjvKAv2lcnniy0UaajZ0E3hWoEroK
rnU52XVYqHHaz73iK3KssuGeLwyvOsHpy98bNwFHUjMNtKFKwuuP9n1EP8hXicjM8dvNv3AGZv7b
olVA7w0FUo3PGVJR/JMveRNx2snwNR0hsLnylSplptJ6kJzsWBCatLuH/Yc4Y1pvD07hokHT/DDz
B+gIN8WSPajGZndNbShl9S2q1W1PkFR1eu/pHdOektsblBVODzJPHHZXB62cTJS5tjXg1wv4I3un
tUhX4+Edmw3cDa0RJX2PQuuZo3x9I3HHs1HepV2ZRxBMsPdB07RAbBDUl/zJUzNbaJbAiGTre0QB
McCZQSj+m43IJIuhoLZySbI+tz/10dSJ1EedYhtSZqt262l/0cjmDHwUs7xOmEElRIoxkvjKsK9u
zuOxBQ2cF8C284yhRmlGuuv0YXExfIvnpjaU26zB9Ud+J6JB+Xus4jcf9xEMc31y0h6qbbnpxJ0u
MQnT0LkkDCBFMyoVeXqyROff91odPXq8+TxTJmqSqiZAdkTJmTrz9WwBRPrh1EkU17l1l1ApMrW0
IKXtmyWWQ6vJIO/ENF4ddHfR6GTj6r/sAJe9aGWyNRK9k+yUO9i+1augfXyJWc0DUv2LSsHG/0Ld
2LxcGU8RH5tXat8sS+6KsfKiQRp0TFYtGTqeM3cLRwy+zURI51uU7dDzlrSevpE/473NB/SCSMGd
TONBStzanSAhDGUkskCBIT3bIlrNlBMR/F8xRjzkMsfczrJHatnzaTG2wFOdTnZv3FdqIFYXhPc3
g5hJtYnuwG0VFBZyFMjDhiiaCzhrvKyIlhaH5fExf9WxDsmAGi0Yqdb9SsI2nwdLZNdDDoky3D7i
ULcAfaSYJW9jjmdRMUog6Lbh7u0rTCLts8/qb8dBcy021kxZ/Wo+jQ9u9QgWfhB0kr8PtlXJY6kD
1G0g4yl6nLmEhxLORPhQQewOf0IXQ2UHda7cwET7cmWMhlPF+cTjTe6kpUgK4hkfBMFzNut0Uj5T
+qlnoU8ZR3lSlWj3fUjMX1CeGCAVSi2Ii1uPggyAQV5GWmAe0Q3vUoFN+j3WvEf0X2CNsb9Z24VI
wiLjdIrXz3LYSg5VWO66a9pupv8ije2aoJyUzvq3HBriq/eKmcpJ6xgnObXH2sJ2RQWd4mU1XTWY
cNrvDQjy6s9aRiF3J3V/FCevE+F2IYMkiv4nMCI9UEYeJss7/dCBDzBA+27esQp7T2KPwwMIUA0Q
QBwRsN6kauGeJuC0yTvhLEeGO8+jBlxfKD/f6+EgAT+bGRccSAfvHwK2fMU+xJlD2Efua9vle1QL
J+RJmCUXVB5hM/L7vmxNHcI5LFXVIWh79xSutzoRl4GcuVnNED530zofs6TnTl7KNjC/An01t5cs
T75kY8MLt6zcM8oZWNye6NuXymwGiixUZAWbH8UzlfQbRFb8yeXBXlM01mpyXP+g4WyYnaTAC9TM
BR4TZl5vnbWzL6kJY0Q7yK/uVW1H7QW96lh7lP2PRg+XU2P5RxxnZwY6UzlrNrFDUtNjzwUIa+4r
vzjrEsGm+Y9kF6LI+PIOMevQwLDA1+kPpnIUa26a7WOTxljYdk/R3ljtkZ5aF3sYn3TNEFJ3k4up
vVm0wtdGDQJMK+heYrFWMO6ktQnCvHcCW5qDBSbaveZTrHurxBZmhfGKzomaeklRwK/+uEj8wY/4
DvTDsMRyguMlvclHYDoSWeknQq8MRgiYEHdEBqrPg/0FlKxXNCXL2wreA95lweLsoDE9LL8+QrQl
RSc+yccjl6iEIx2A+7P3Gx58FqHYkj45Y4NcO2KRjh8XcWKr3x7r4jCT5RwUJ1sG02qbPgdeShaB
0QT7vJmuqzq2tyJ4vCarjWJa24npl/rR/tXT193zohdb1Tm8GMnlnlK2Q+ky7X2ZZwsnSQzSkt+B
dZbOTYyLfq4aBGoRcc5w4Rld89DPjBuudX+kfAnnxolcBg3p+QX6yTUauT3hXRuess2fUpdH+jow
83tREym7oSoQLvJwwZVZGweKzy9w5nZN4r3Y0bn/Hdr2l/KSzBNNFL6latLqXEqf5c8OlEPPsgTi
iIQpdvt3/gjHZGvvTkXm4M+bYxr11pwoP2FhKRP9L+6qC/byVlN8iH/r6yDz4g+vpDl1Y45sWSHi
BsVWnwGdBPMSbptntmxDzlP9qcSuvv37IdsspUykYEC6BVSL797AqkmKha0ZpnA2ntAYNcOT4gYn
Iez1ELjXZparAw9WB2wA028ovxToLDZsI7X03e9t89RdL2sYhHXoMAkLMnn7Xankazv5qgbn7zFa
vulkOBEt1noTyo4dblBEeRNWMDehDA46Gj5U18D4kmSiWLR3K29KjLlgS1vzNJxpWddLSgRNT4YV
v1Ne4ffVpx78R9WUZ+djHfNjTgqF3tYGgVM9hTtagOIz02RpR7Y4441CP9lGwHlurBxIYWfGgBpB
Zr/t50tVoacHW3z1r97CGtz24G4qPPlq0OofF6t1PefdPriY3kni8IZElqalfzjunCrd59+r87o+
KcuKErkbV1lkXYUNQcMHP8rZjSmtx2E8ega1FEpT2ORit37Jwqh8Bu4zEdVEn16sxWwJxxplmMtI
G0Hr0I+na1+s6coodEdY2LX5Ld3HWpfGDmAxWnNTP8O8FC0dUlQocCmv7I9IPqQGlUPRrkypPXxm
9ywY+eZuvDGsW97iYgT9UxB5uQ96LByeV6qe/1p2jvSItaFpPYJ7rE2kZwsBmiPVR8+fzylQ24dw
RxTnuJZtbHP+2aJGpYvg8nN4Xxr25oBIg4j+3XaB3j/ZGnt+Q3t0IDzgBRsZOXZRimWdt5th8fuv
XYhQUX42VjUa1zAY7BRs4a6Tu6Nuh1J56Sp6K5qj3D6+0Xhs7kcL5Yb9nKLnEfCjLH2+IPLfnuHA
7DyVDkL5tTKghrje90oIWPXSH05rMK8p6l0fajtFvE1n/eLntX/rZJeUQt2g8JRSh7kz3zshLka1
JQ9ooc4S9jQrkEYed+pkz+RgdZvSX7E6aQL+j6xurTuhtHz2517PPbbv2RSAguljjaqrDBIq5+Ow
2tBhKGg85bv68c5WzWxQ21+K2D1jfQ6Co+3mzLwTgPH8PeElZQrmN+ziJIhAOAolhNOWJN+O7S+s
IxW+b6Cw8OWZEsjS6a7QkZorCI4VZrVw2P2h+Z9xSjkOx90GHzyf3SJnhmGWKT6LxTZA8oWl2KiU
Tnc9rauTp7nJtFyWmfMX+ENjRbaUbHpnNCECnG9J9DCEL9f7tRscYpDiiFDcc9a+PbueTGM0u4SN
1myjd6t9zXKFRkPL6X79wHKOkommIGzSYHG+nq74AilqW887tbVe3BbVmJMnFfn3yjimPjjQQY+n
BX+TJyLZmbHHM+v/+I4mFQekc7Bsn1m/lg3YcZ4Kg5W/tBzMos9V6z9zeorDLzaSjb1NpfHnGJdG
ayy90Twt1iEx40xXcHd1azcQ2AMzUQX/ae6n9bleonIIsD9TcWw8tSNgT9dCZzH4TiU9EUNgIHDQ
BIfkZY8xx53mQRczz1LJrWGH8Hi1/Vi1pci4sjtZ4H9lAW4yAVaxeqD5Vb26bgVor3N/TSGmZ42J
KO/78EAHo21YEg+ZvYTtPEQw/iSToJUHWdI3h+Y69UoTFMHOXcFiRa0cqIRULqq7MJiGzSa7avy2
Ak5a0eBkFu2QveRs//R+p9o5V7p9Jxbx6xcNo8aefO0y9yugPkjFZKWoPIGirBGEhcjiv+gtLSvz
Aws/AerlhWsddp3kHpqzIBfVsSjuY+HfTzVhFZ5OnywUSoibwSqvLvSr8YiLjEj3iUEf5wx69y1p
s9tzjb86Q9VdEWjrueZgLxuKYdvwCRTyawlcs4EkcHK8eez7eYYeNT3zqnPHUrZe53cNj7aWvLbR
4aiJyDPkIbxz/mEVM9+A3eKhmQloNNhhXU8YUYp4RCU0Ja0979GCYwdVxbQfEqYy877KjbWYCPNA
DIXck9j1M0euozlBWatwMgRs6wodIFjbmw3gPm6BBpLQn+e/t+daxuDhUOW5Wpq6/KQlDGwkAm+z
BXHv6g95OFU+FRVlldacCYsAJeMg2CtUvbUyLSgWc6zSymk6T1GIHRkp2Y/6tJFBXR+ZjlDJoA6g
5a2LVyPoVBupI89Uz2apqkAcW8l9uwaJqklSWvcnWl1hHeolvpXQjrdUUxXEmeptKzxuUPmBfIe3
GANMSFTbTwbbejuwWEBWcfF1oiWMpiiVeIe+YQPWjFkkT3ZjNzjYqn7Yur9ojgGRQkvWEYEMHqmb
aChf+n7Sh/GJRqczUAU18Gqd/q4HJZDmZoHxciDwXnwMXW98bTf/j7uy9yD8AZ3aGckXTKupUjaX
xKaHRXfRM9c3jOKURTjaLBvXIpZu8cUNQnE35sHlPxNVNZt5ApMOv04UeOOZL3eAA5WXVRQrUdXH
YGSroZf+R0JESIVM3fj2NjoSAN7jGVdAgKXnlY68g4vUQ+ZZAHRFs7HXbEZMjQNrVybx16bKbfWI
1uDEx7HxPO7c84AkJ3LAoGixctqArsq5tSbIXV0RJUU36UiIusMz45+su2DjhwISHHuVh60pgpQ/
2xRjQtwPq4O2VLF2nz+XlPYhmaVi7Mt/pGEoQEA2nhtDhzgGpkUdayMCMXZRZ18QE23TjAIM0ekz
zDLH4nELegTkEAqEcUa+c+90GdJG2X3ica5Rc46ooIr1tpMEtw4N0oWbgJgtl4NKYuQYZRNdIf4x
AJQGhDaD9+LxGTlsJQ0XuNYbrK9S1aVR1NFWPIozsWjCN7PSyEU6JQN8cURjJiOlJR53Y7OSuaaj
3e8YufD+4NCKLVJaO37As35bIQNIUQ6MtAVxDc+cXxa/KJQAqKPtIq7MbtHGU0eyQDPS4TA5NYEL
vyXnAKiGSzvg9Z3cUSnsVL5nSWCkcWDZFxQTxs47w7Rtl6on7xI0LG3Lhl4zliXq41uCcpIBJX6Y
BEsSHqUgm/QXnT+n39wmg2hgybxDPByAo2clDd7H3+3DcnjKNRsGmD+HCFp2EPDhbZp6y/9KwesQ
A7QITk25V8SJHUXPmmCwYRiulLUIPG4bWZBmbgk7B+UDODFgQltOGFiS/0QxL7qDpMZPp4XlBL+F
uzocbbQqfNww+uMcJN5vb8j1Lo4333K+1EhRPr5S4qz+Uz73zeGGXENsGRzd+1xQVEloYKLkdYuF
bBOV3axXB4p9Aa4Cjg3VOSoF7abc+ILdm7whXodRyw4NySTcxYH3yeSrIHiyLSvD6RSkHpdMPVUm
3uOEMYCtzvpNBf7DN0Q2Zqcs7ddavL1CvVqBA+eKx+oHEOyD+M0UZ56YK5GqBp4ybbIhR2g4VdHO
vXsiLW5E7ZCgeFgTgRyOhGRgd0SonCqF5wg0LLHBVCQFZD489HuLxs9zsCvGmc8egjUu0uavlUCn
uFPAAdIcJfcexIr8P6XnSzEop/QDA6+aQdS/DozhWn8rZVAmrM57XHc5LTRvojaF5T4PXpjQ9QiL
83TAh2d78Dev2Ewfb6gO7x7qaCJaVmBrXg9V2Klaq1GO4XwacTn7HU6ZGnHu3KFtOaAqTBGqOsvb
Hv6xw26eiOBYMa+FBsdCng6tdllTyAcbA2iqAZJBchtW8CPeoOPb3jjdmyNZ97dOlSDvu3/r2UCK
w3u9JLi8cyP0VP8F6EIWpUpN0zPbu7l0FqiKudSqAWiGuFvcLhv5Koc5D59kudOG4HkaInR4m6TY
Zfd+9UvGmn/36Pq/lFOGWMGxUqQ9nUBGaIj+zZSqc51zOMlpkq+HsBISBbrpNI3ePU9mIQliO6zw
7MAL6Rs5aKDbLz/a6l4jo7A4KRK+Z7o0zN4zufUOqFC4c1vvqqxpjODDUyRzHUW3P9TZcj3QEH9Z
KaKJbbRPzrEtMSwUCIQmcn653Yxp4qs1Z5IzVLdNMak+NZzzslbn0nYzrC+7oaBit2bnPqdccfsK
9lQYNSZs08fPECWG1hj5jHIbFS6GwpDIWy67TxZuXU7uMzW+5iuhSTBPEvm5dE7U6OI9z5hlbb2C
X4hO84VxCgKeUDoi1znZq7GbTCxpy1d+P/OWoZSu0JSNTBhcXRHmhpmRkL6LnoBkAoHuXet2plRZ
kt4bPDF2a2l9aPTOpcjILqZV7zf9aL2lasXlYhaC0rHOk4vTAnwoG5p6oBuL8BoUVrbz0lX6oEzA
mM/aZLyzswdwcTpa6GPsYxQoZmJ2cCFLdMNbSkOX8UIu+e65eUoWsQMekt5Z0egnNl6C3DIAt0Cu
3pRPQS+H6wZbxhdMXYy5RL4lLnCp86TO4wTR6YvrOqRB8rxY0ozsC0VOkb3rYH7wIJMryJHAlIkK
Cb2xgZEtPv8YPxlgQ34Ti0npgZEu/XogpICdSrSDxAy5A9Qj9YuKN7HP+kUVlfLBoDgS5ebGiNT1
iK4BsEJf7IuK3OKbzNJyUU0mwcTanuDKZR/V99Up4wKU1DLaNXHDo6isvjuYsr2Zb7Ubo3XK6dNX
louHBLcUaAa6mEiba0sdIJhYUuDCLUL0WNQ9dhciUPCi8SZ8GZ4sjfW69vRRIt6S7o3bUWHig2rJ
gr+f040mDDkx0Fij/m9wNMsgV2uTEqknXyBXd+uzwvculEUs1y+z3y3WL/HD9akvPF6seqDshqAo
IFWH7P07FBSN4+QXW+tlyIFlJkwyN8DF8YmaB6o3waf1p9EKEjXas5GanviptKq0AbitLKXbql2d
dCpjr2KDkBa4xJQtErk3WaquLMufF+TPmK0XrFSvhcYAjbMl1cw9AnbCyl82RMNJddTcoGPhekoz
OLxo7NKwiMLlhTk948ux/wCh/WsPZfl8H9Hxux0vbnwIt+DnWSWU/gDfkzhJPpHq1YityX8Qignu
MB4EJY3G8Z5L7XYri15JeYopl2SG4fCCMTZ+FYb2CjxpdF7Wyas39T7fyOi7KN2Hkbgxd2zl+DVT
3Eyy2Lc39Fq99LZX9dvxpoXMy53mB8umwnIgh40eHE13xQ0t8te3hw5DS5dqINi5yjjl5ws79yQB
labKj5NjEeDOJnh25/Kfw1DVljYlROGNmev210Ax2lJUKARi9uHvqcg766LqKV9ZOTy03m0BLMU9
KO+4KA66Risu/qMcYU9jo1PTt74EQIVBg11ocDNw+SGQmW03nOy6BHctuIW3F4gvwGF4FJq+nGFL
bIvNG9VGINb/J46R92Gg8fCdPw3feaPLx6bwFdqJvPc96uSJzNPNLsuEKK+i+5cKQEhuaiDrNzzf
pUIc8OrxMA3Rs5KTPT8zjlb8oRe3zbmysRioKX059LGQF0jPzsKa3MLuj9+hUzCFZOTuGyxEoVc7
ZuJQuSdYua1VxRbYhR9AMCcQwMua3mbWv7iRsn3V4Rl5RAQLYNgwtpAUGmWYhA0CcibTkuUjzP42
xRHIDbwfysPp1q2Bk9czr37XC883OBuCWPpK5qtiE4LRF8iA0vMHIjmz7lF2fmE1xLBt+NR/2bjo
Lkw/4ybUbv140lS2EWYdifQMkf089XwelbaDdijBIBSxSfUmxsJj9sxbhLuN9AdnP6Ul7dOqZ/fa
UhU+XGOFtrNrtJF+QuDGgAn3umIll7VzQEK80/SvCK6suJvVWgQz6tA9a4A0Xbw8b+TTWP6LyhNi
RgfvYKxEfGcKz/bNvpZ5XGGBKbKe46dOIr1M7KCEIRF4j7y9Ep45LEeL5dRt2qw6XMBw6d8bwRoA
yo2N/cTYx99Fm+g/ONy41Bqr+jxsw5tmI8utNrLXd+R62He0WTUbwxnGLUIuROo/v8WCjcSoV09m
fe/vVbkY0IGV/uNeJLR+1oC6pVqzU4p6TOZMzhAlLNbBSIOqm4XS55Q3t2JSz1LPzrdvN0+ML3cl
IQrfflQ+hKlFfJgeBWdGmpC1SCdXU77pcVd7vtPrdtgdm55TxL8KaIEgs+iMvq69Cpx5NNKdGRtk
zJ375oVC0/UWwLqTmf7wMyItccvcVbmxu3gKIOegc+A+MvgWwBKlX4nR365idt9BrSEAQSVfqnuO
XEqbWHeA8av6lptSEAJ0Gf/3Nw/MD389r0+mc/YZ0b19CcJX7qf3AjSo0i6U1PwoGiXX+WztiNRS
+3Fu55KUSpJxswZ0lW+phkVaX9DeLBoCLTnElOKnZV6GYoeYDpbMGT6nfplm/JVVoqRf/WIyoJzr
Mhti+veV3F3dSGMWgfcdfTSYkR+LzV4FPT5e1yrF850tEVxcUapkDMVNo/g5O0pNVsbGgxb6c1Cx
P6S3RoDkCJg7kdP9C25PLIoDnhg9tw7sz4FqrMsR0KeqoO++BpyCzcc9wAo/TrRVbAykPQzKj0+F
fib9V+3qzrOLhpRdj2DDEBduhvcGmxZNeFDIKha/Wd63wJsM334l22Dd/3YGpCrNTPuHBU4OUkx3
7HyzovAAPM7uyEVc2w2k6z0vBAlHgel+daVnykEgaZpCa+VrUbTQkjFPdbO8ih//V7WXJuix2Bxk
YDDej8aPr3dj56jEDJGodtwMdMLVYCPeeHH3x/JKi5BOjjZAeKJ0F94S67BeNGxKTjDFjIxUOzIL
zp4F6nKWkUtgcUreL6+oogkpSVq6td3bkPK4TFK2umkSr7Mo6IV1KJVVOHrflydsA9edN30qCa6T
RkbZKgbsRTD857yIopD87JwXK5H+4AJjesRyqWA505BUBVQVxu6qY0B1Snh3y22qkmC7e4iYeRml
JFua8TFqCNZtBMqg0zlE8ca2f04lJnOpKN5/41a8J89J09SDvuA7+5D7aSpl9iQnvsNHjPUTxhOv
MSLVrSAA7rpYsJokXjQbMVV8Z1QduLtULbxCOQLCOkfOrYj/rasEta3FuiG/bx5ENnVXQCLzsiUx
BDU8JusNZT6eQdX/nOsOVv4jPBRTPk0mhpEI8SQPxkKvEGamkN4GBmgEFP9R7g2qAhAEcb+cskQW
1m13KiQcWSgzwiLAnP541u2HseuH5dZO/moYaWAd+746dYCSqSPyKuIg052B73QuQBEwHSz4szvH
rbMNAw96Ef97EA5dDv6eY1EmUeiuS4OIjK8JTQhrrqcOc79qUUlZGSyc7p98PzI3Dwv3fqhC/QNh
UpvIn0TIwAIiUSADcJWxsUKpPomO2y/q/FCk9vxWgHIJzI/zhwZhPqza+e7Hozud+vKe1vRr+FDM
J7dqm0LIhlqKqMDr+4mUK32JlO/iNqooppAgaUGkmyFdPTuk2IvGWycVSWCQ9XKXtASyo9jjRAT7
tgJTfTN06CpU+xV1Wf44CNJW8aUKCvIEY0R1cvuX55s3NocmgZo4cITYN/D2StNgMBYa0qcykzRQ
iTbvGuKUlfSoGYoHnz8yHr/4+o48PIWcv1EDBEIgfV7ZU4rrrxN+922XWtC/m2hY6PawsKsVWq5M
oBgE07nj7lU0C/bjiDjHTNACQv8NygrLL630foBtxfrx7sAkOoSquq/ihW9Wb+2sVXUG1aiMZCxK
3mMJIuuYDaCdbRG9RghDy4Zy/Ub87CIUcSKQiYLoWovvbGwCRihnze2/t1dohpsS0QtBKcia9UeV
EYhJ8HMHH+qY/69H0oklrggcmYkj+shVLfpXwSJec5UaYbvmMZvNrS07HwfXo4RX/yH3R4SCiSvI
rP+nU6iQdmv/xA1mn4eCHfU4d0KZW9yURCUJRRPNfEBnh8+GWhLuAaJaGI/UCRTAp2fbg8yiR+yS
livsh99GrxaLlkCaW8m24SqDiMkajGkqgbEDceY7cS26bomLDNT0x95zx1lRPTD7NYFwUZzQHcap
4BDAytULxxQuYrEL1MkK3L2VESHzXd63yCtsD5dgCPv66RQqsyBwmCG1kfj3AadoVUHoyfr3A0Sk
tn+5vC8JUBmWovHqpaaB7tRBPiCgqEWedqFyJF9itA22LajsiR5yiWhMSBkJqkPsJexkt9cqjg64
NCPIgGJWKb/8e5Zp83j11APO0+fKR5hUiB53gMbD9Js9e9YDFy0cGKdbnmJ5btgyXCJtFPVGLftK
/srlU4PQu3qcV2o4EipFLIaXg/mcvyavlbzisX2IQD1SmORnWZVoad55rj+LpCIv6aIdo9DHfvTU
a7PWRpI0O7qIPuegn0mWMpA1hhPVBIdEOwLdpsGk9PAsmgar0m3+ljHiepMHumoqfJ8BbdIuuFBG
UU8vwb52Mn8NzdtWJSgb5Cn1ikbFa1SpPKiG1AvoyWNEOR4NjX/tG9Twnky0WhFpSLcNVxHmULtv
/wv55pzDITE+Nq95GbrGVAHVRXTMtsWt7uh2J/OU6CQBxBUhEUC0nbiCmu9BPHU7mOJjxfRb2yPc
miqy9rtSLDBTMlVo8K53z5lLBB1UkUenx2vgz9h4gxDbplgFZeFDGt83GS/QVPafKNoLQXjpL9Kh
AJ7oiCdsW3Ie0fyfQcippqk8sI2d+CvOI55JM2/1WIJWoX8+WXiOYdqvyutTDSUXzEpH72F8TDss
WSvA61D2iZgqL/0nSdQaSdQvkVCgMBdyRqijQL6xoqSkISBC3gprJKsETNZUwshIjP1nxOMfXv/z
yaKpyVQ/pZFzu8GwwwCpZLGLAPCGP167c+bWj4Ab8majVBsL/U636WVJZOCZsaQO5ULKLi+zFv9t
7s0QQXnxpe4zv4nqO+WYhc9mm1Ml71Pd51BmR/h1yN6fw1L7vdmcmADQnwt+sBS6/Ds4xjN6GE/d
j2n1n24K6TADT1iU2ubrcKRU5AddUteCK9Jpcg2+a2Q74yV5ntJ4flPXhSQGYH8lyr5WhvXZperZ
YcGyNLT4JLZ2as4vN3XUkYMJKVlW8N5dwSvi3YxlSLc6n1p0ObS/xA5+Ay1zYhXtXr0nwxb87mDG
nF0Fx0p0IYT1UP/ly0KVXzLJpk4lCDizy3EmpGgu5FIHIISMncZxUR6HKkdbWNhHDHxLdO7oM6bW
YiUnu2cqSyndLiZhFvDlJpBkTle9wjqIBfT/GocbEe3ML6Dn2TgCwOn/4MUmvyLx4G2UUw8GWW2e
fwF35E4RouvizRE6VYsX/bsZw41UYCgXpaZJEkkK8s7AiDnWKV6iGEi3QY4jas3SfEiUEkK2oiX7
iOegGkijCdYC+yxnoTpbSsPTBsVA8u88M8IcWZONNArgrvaYuRqcYXNu10ZyQL+u4EHGY8XEqVl3
FPVpG/wYXRaZRMSRXpRIiVH7TLZn0GEV84aHf29g81sxrX1IW4V1p9/O6hQynEU8xOAKRCXBAjUr
lE3LsIO0UDqPqosnuvVepL4yQ1MmTFjoZgxsHdl05UnpkDyOm+iJ/NsNp7+ZfOon2+KFZMeW2X72
zcdNK1QJP/MicaMVORz6koMM/gaEyuxt7AMENfw8pzqYjRMyyk8T04yIjoNW+pxx7fKNrRqwFJzx
bLR+XSa6ta/HX8LXLQ6t95hNJg59Mua8hpwU70Y0zFhfDUQxnCaLFLp0mq1b29Q92dB7QWfNFywn
Rf0TBxvxtyWkkGQ9y632zgbY5ABiwbvwQvNjdOPA5JGsIRt87A41Syw0695/8Wyu9q8tKgcMqoSM
ubelbaDUTAVmmUl0cTQGyWE2qe21J9J5PV7AkzwC8S1tUlJDS7tRNZHu09A0rxu50DdrQpSM5EnJ
tl2OWdqWVAi7RHzCr/AoSbHrEVBW6gUqFDhZfR9CqtEUpcRi9e2dOd618MBYVogv1wENxXcGmO5D
DoGP0NgGt2DxOrhE9b5wKYtPNQHnEmKaU2fJWXJ8zsDhc5HuDF4WdP5xti1dQgECLtFE1gapctTb
hDW82qvnQuyUFTQbMH5ffy9NOFbwVULTibi6tByV+d84gW7z3EfrjUzjoZlr2zc3jVKdoovq57b+
MfJLbOX2x2cCuuNolIZbOmwBOGAabASvYvajwRRIYEjRgyg8baTL61t1AmVJdBp4bQu4u3PiNx7a
zu74TLoxaJkWbhszOHrvNovPgTyUCC3osHl9K/aRBdCbwFSEHOMjxlECldzNZU73mj5I9DNhfrGf
U2PXQXsaMzJ8APyLNUdD42qP2oW2gO5bolDWetQMaoogXMBGb1couLJfvqfwzxqGD9NejoltDmUp
KzDT6mrYhV+T3ISbbaiBwlD6DdYleDEnWQvQpUwAj5Ffubb1Z0xSQjMfWjJtDHcmolYyXEivDUoM
mHN64mnVOkADC1J4lnc84AyDnIMO2NfqSIrVRvuTsWV9QU44wjI5nD7N6IrARQC2Xigx+fLMoeuQ
869bBjjtKW6GSWllvGO5gT1ZepQizEC4Mv31fGJ/tFBVb9x/aUZZ/0ma74CzrXl95L8l9EyyVgvA
WwrFMwRYRcvdQg4Pq+sdpWLZZn0YjozX7WQ9mXoUIXWiIJmm0rYB948BKq4U25QGhKecXeq5VRx8
qoGrZ7lBD35rAAyPVOFIL7iEo/YhUZ62nDJp8l9uFSSngJP2naOIUzDPPmfvunQ6oVNaHJf+ruKB
uuhd+v7hcTVVm2YqB9SJfUmAmJkgHUPe4gQn8QNJNUJD0VWTiySwVUUBEvgJxsjwBPwi0KFC1Xle
MMzwyBYPCF6P/+MU0fPTG/LQ4vMmUgjlp5USCjduK6vCMyBqa4kRDbKA+2Lx3GDkWTgi+ZR77PGW
dveagNAb7dblF6Kw3tP/uqCab2KFZ14ney664nt750GI+0z46dDMjtQ7xdkFlanXq0Y34RvqpJnN
O0kzkgGe3pLn5EioO1XQDd7q4Toe8Cx0h8/SYQ92ID6Q73gZi9Jj+XORw7o/HUCi3PiqEPSw9LlK
ogKMvXiSER25nMohkZqAxZq3Cr/N6g/RGxy6robK3gOv2UgghlFkxM0hZohddvbvvBhNgfWp1pV3
HZVMV06afUdATx22r6EhQ2tHC699L8K/O7i/cpEyynwG/E0hbiHhwVDbgVxZie+Gkw5GhXPBCc6X
FhwqUADECbjayqCl3MWox7UY0ZLYtLjdMFbs3Pjiygc8+t5M2AQhi88o2ErCiz6bZI4kxSJt0tDK
kOcfa0uMxUeBycyL3Sm3xV7lrrMJ/py0CwuYcdNAyNASlelcSBz0HO+WBmuhEx6ywTdi3Bh6bBFO
BTvSQAe48yY577vfOSUWak0ewz/zTd+cAHdOmhglQOC2PGEHwZOoalviyplPQLSs6RfPGo/l9aUG
/SOKaShfdHS8U8C3LKfQ7aaZ8uYWM5pydolE+Mg2/p7uXgiC6QkLBjLWZmJaYw8VoVkceKUNLA4u
2f6BpnnZbmZNdUbIRL46mihynY9rhx8UO9PaD3z3CJiRkVRv2aRkrUWt9Q/5Kpk85uaARVftuj4j
/l38XQ4ia/Q1xbrDHhA/KOPGEDihU8H/AXG9veyTkGeSKrTUkG3EJkqvII3CZzOHTko5rDaiTw9/
hMVnB5ldnEGJURnjCmvVamiHcakt2Sei6oyd/c4PnuCyuD44TEL42KkCwl8kMDIK6uf72oY88jm7
iXfmx1MYE/xL+7gXDUGlNN9fMqJ8Sx29Pv/Lv/MnSQAYNrg5b0ggUEY6dbzc/RmWiQ1HOX3Evnhw
MX5IMh2HJ10dqYEjjmMnzhcySuQ63a0VI5utYXU8/Lteqccr/RRLAOiRtYIS6WSd1uHECumdE4Bt
AgmszgJLS5l9AqmNXScraY4PY2dD9XyLzhT8eC6efDGZXJeGqPlb3UkESZryrgftAJuc937tpA/N
3R4EEXNW27VahaC3JEv39HvXbP+PBDk4ZepfQGtYvgcEbxwp0jgeyIgO8qgGZHytal1zZgu3f9Gg
0VdpxCFEiPOAjK36V/tH5TtG6kl9MryowdlvbNKSpkEFNO/AgTaZ7IlJ9DiqwpZ4dHOveaCF4bOI
wZ5BU5NfO66hIpljHmol3HsuZKjcl2wvu8W4WngjuUlvXDB2IAB9y4KZwjv62mxXrjNOR0UeyT6J
WAGzv9xTLMa15pR/3nBnatBFWZA7IFM4EQ/PQDA9qGSdddDH+D1s/2ib3rjQzvR/YOGXh041SF9F
wsZktLbdlcP3G99+rAzG/LdMrMrBTaautMfnWUH3PTt2289x2fx1V6B4Wb37wYK1v91yqsfsy5RU
n3No5K2qzwfeYGw/YcxLj4kkCgXfosevh90egJBBxBqfRkKELpheu2SI0pZF8olT4t6w8/CfUmJ9
f622jMH5Av+TkKWxDs+7OMmh9LN1V8ooD1G49PLZZ/E+ulloXPslHikhkZcoCvm/3+KnUzl5qGfB
NYdKIIMWo303+D4CCLKYbOM7QGyO2kuwgCwBbdHIdaUn7zGUKv77wvnwdvb8ICPmaEBG83ts+SN0
vesoQfvfdTjz3ik6Hr5QnHv5/CgKFmMXGLyFiSx1IpzLlDuo10iluLc/HomCkgUXqmeHumwGsE2S
WcRxZdvIu3x16XHaYSlB9X7oJRELWEMji+FPI5V0B0tUzUh5zSk6OptwBTAZOejzODguo1mKigTy
sPlpy0wGZVpBtRGWd/lztmi9aidyYWa6gISwtK5WBauN7n+o9l9C4Nm094rDkKPEegzpRt7eIZtJ
E+rp8Q1C5qo8oOycOdGSBf6/vTXfjOVRj5FIKQAYSfzXsK/J7hR/XLrP+tjLqbY6QzBEAoQaPi3A
QpYp+4OsP0hx5HNm4RAjTliF2awHhdohDf+rc+0bH5daYvMJ3UkvyurtsKplrjO73l5pXyyNORxU
dAZggKW9qe3/APMl403INF5CjAAcV1tsc7jGkx29pooUQxhgB353Q2RfyGTQPLAezBTSKiG8gx+8
BiN3X2RWf28OX8vbb1qhyUrGon168+DhlnpmCMYskPSN9AOeZDmjtW7P1R58m7g8OCP2Rvn6FKOn
SrXAY5L3p1bVcT5bcFZSKairqZmAzDZL31Mnr9GtqiDK3nzzZATKEqJ9BLIAsQeEsB+tOZ7bk9xy
f/YXCdWOjQGJO63hBcfSvow1V/FRxUSyTDaCZCdw2cFhpd7F249NfT2ITra0zakdD6yGzw0bzF6m
3cxgBIydHog7NgWz5w1AUkCuU4mUh0DxoLyi4wG78PlGMmefCxRqQtW+7CHqo1BQmA20+4rAPJQP
qsHU54F0Pu13e3YXfAlyv6Z7GTMlR7r5tt+hU3n9d/mB3V28W9mAXF8iK8kCTRZ5MqWjTz2qh9Uz
5uqnSGN+kdlpcm27VoEWOt5CvgiTeeOkvXRBItrHtQVYUlaxDISW/OUb8K9A+CsKUjw2lsSgU0Xq
wMVW//1nvs81DTx+0djyqhtrckHBFB29nweg0mDBOWzMy+E0L40aK/sgu6fydyDiApAtyQWD009n
M8n/RTqNBDuYfZUgyoOGRMjsQ14QHAcG3dIXSNaMFfYs/L9nbOOfwbNRs6ej+Jn6BQuA8sfZ+gl9
DghsiqbBju/ohyX1tqNf0o1MKSIO+X8tN4Tyqp4eu/Ql2wSpaN0e8zVIftsKyDxgnm6NjC4wM7/S
Hu8isZXfZKxYC/QSCraiQmwghRyQGGMga7g5tlv5NZCrOSMS06+PeWGoeWRlI/L7Hx4wp5vmxneK
QnFmXB9FMbWe8N2NY4/SWx6jTYkiBFmC08o6FBBXSFYbGkD1VaegYdRV5VN8G6iqTYmwHzkVcZOp
Jg1lIiFCbQ6D5rPb3A+HTVk4tYEdbTzkOcY4lYfIupzVXBZ8yvSZXBC5mHK3g+qpOBkZlhfhM2X6
l3r3/owHODni1GbarRPhsx5zgJXlWWwM/4zB9ThatNFD3BapXTXO/vB2cNmV1WRC2nV/2hRsNhB6
oOk+LCUpC6dqISPg1xcDi1wKqtDP/gDxxfca/WoXhmebbIepYjQMRzXK/A7aaTv+ffPsc+6JU3G7
ELwM8a/Uv3ujy+mh0Z0278LMFpD8D9JI2IlGUIx6YwUUuCKmKOYMKUNWAkCNavQE0c0WQVF6DJnn
8M/sPATlNhmQhNsNQURILCvJEYvdDWBTSKcNALzwDAUGSLdMld7jGr+m0cq3OkNg78tMZZmtKbNq
cgSJxcZG2Gwe+LHMKKvVLaBeQc0buF/KMx022PmYKPoPLr2Ca0dRv3hoxhMey4HSb9Pf79xIqeSN
TxMhZHEBBUO77hlb1+uDtoo1XK1hsxbFOmf4sHjkDZr4OMLAt+MdmdY/JrhZ6iX5hAhnFzFOHLTr
80VJjPulrKlLtMNajstpBeQhXYrid5ROH3ttFj97JsOQnE33JIyfJwyx/wrcgGX+gOpJp6qUCZc0
k8pMM4BF2z/NVyagLW86bVftJtUThpJgwzuXhtjZx9U6Y/D0EtT4/qvGq5xnvA8XoSFWi4QpO3WO
tCWBnvJybrcG7dwwvI/UX1HWuKz9TeqlnhQkEZfZzAwoX+4yCx/9wMiQPcC9D3P72lFoASa2mlDB
xXbVEwPu6eAws0LfkDZXPR6GQWB7HmkXRm9wrF7TU42t8SdIUTaeoUkcxjwHrqtMZEUIyTIqP5CU
KU114up/CMEZHd/worexTxza4RjBA+EvOiHukmOtLDxEYDqlVmZa8Xu2Ez2CQxnNIu+i7wOdvlxp
f8zD8iBqbMZx2D5p9nRLMdURyjgZHr40sjdKdda7sr/V8ROon25MSW8zAWFVuH1wIK/5Vg1yyw29
VG1upiwsV+urLhlafnuFU0TOZzIREPb9/nIzu6AVI/IksNzQExIy0IJu/X0JLRIJuT1QWWTg/qGp
eco6tazF/XY+FkCuEQGQC4BQPJAsfy0z9dlgPb6DoZJqmqp9EhId20IqZ8z/wZyzlDshP8h2lGbN
R+PBfARjIfusEll/kLZRnNN3fAX+P5wTxdbKQqDrEiGBXgcm7FUuJWJ1WN4uOOhT5LMh72yp/W9h
HWsBlyvNFSNX3HegIyIvWlgeH0HLrwekbbPPw89eS16eJYLaWpSHgRGrMcaMrOro0AOcRZoNJb1Z
T60JKN7RSWq4IJSdQvKvuvG5cBeWFFDMpGAD9Tl7b9upsGLI28Su4+nGn8r+GFkg4cu9RN05qr9l
p/Wv7ShbFL66IyJfzftk9o0yWPN8yJuBahy6S6amXaafPQEVl20W9dgg0r+oQ5OFCLjP8j+NKWvA
RCzvm9KilrAnu1RlicMsl5kdgS7f2fMfkTA2+nvnsEpX0y/n3jycaMiGmnbzHiFeWL+zd94jlvsE
3jkSPqFIUbe4WZuzLHdPR14/x8LRKycS4Xr/EJybUR6jPMNpYWLYrEAnMZf4SKtzeFoDKxLT9a0K
Wy+C7g56Wk3EYkZRKmdaabr+vqOY6cO3htcDkuMjAVa+vYof7VeVJAE2itHsWzFWvABsFr5PN3yt
EDKWxKUQTNly6CSZyO/EMLJ+0Ozsujg7WfcIDXeBoT3RItkIUF+c6ZLbkdPjWlEQJMHCfmDH+ocL
7p/LkU//gIKEDsoYzDb8zRsbC5Cm5uWxyNegFHIVj7EN8WK/5Xbd0+t0Vy4Ib9YaWt1AHyX4Glj5
cpBNkiGwLVxD7nDeoB7/AsPE2eex51y38MWPUhQq5SjMOTSkkyl34uxB50YMoIHXX8g0KmAzjGlV
qMUqlOmI6xz/nSdq5M3HxAYX4HNECo5ecvVqOqvdv68lPX03VocGOtxbQ9DNNpfDmIpPp8Y6V6me
6NbbeOQd/18YRtad8Wl5DOcOcGGwM0nSSIpmMXA0x637btrZiCVSfrgfcuU69CLUwjfoNJZIep0P
D7S7/hLEOmluKXuC8Ua/3rZDHcBahZWs1e5HINWbJD+a6da/ATwXsw8zsvJUiDK+7qP+52ZgCA3n
JIaXj1AkBbj47wLI+zksePE5XBI0no/3PwN12W1j2RnvcFkzCu2BPqOdmswZ5DEd/e0xsWgHuOQP
UCvVSer6b8ngyAWnaGHz4k/7mhYqXIyIQA8kRkWv4lnEmnmEjcCh/owFLBt6YIWg4lUodM69vR08
2Y7JTi8AZ0JDN8RbrMZqC9Jjw+PXnuzsP6CKNabt/rj2ANdqsDun0CIh88V84dATKWFeVGYitvAt
0qaFyOcP4Gn71Y1FUaCeaYOi9SMZVkUi9zIXGq6s7q7XN0oVzCc3zIKlPQXy3NtnF1Q7CJQilTCP
/STHeYze9JBZLfn/Z2EPlpNcL+u4YiqluRGQCX3caqO54wmHkE6BSTzUbHbdnYudDqq+KYG9dpWg
0GoyKFX8j/beW53cDutHW6IYgezXOQmB3jGAwoAGq7EgIeXvsUcAGF8+rjWj4m5WDlphfOEMHYQ2
iDALQep06BtZB7Xc16cHmLjkp9RGsL6gA5HmmrN8NotaicVeBJcuJqQiwHn1szIhMa9lumxBJ/pN
ssbRWd6Zr0jSvEQmG3oV6ojki6yj5dfeNMUMwhGbh1ZCQUQrSTeAqOCST5kPM2C7N+gEwBLv0VrM
31jxbosgkNtbawLbVLXgB4fdxiEGa+3d0L+MWhusqwlPnBw4rvoKuVJYh0CbKpDkbGUTTl+5SWPK
YW8dn/gzTT4sn9BybOTwvopOTpXUQShVMVDvCE82x/RdWa1XP0Lx2zmTjf1boup6h/N1xG9ximv3
nYJluQv3+HCPviRzbRcokpiQG6VPCNf6HsdyDVLMbU/cSrZzcUwsBzdLeV/l4DM/YHiJEat5ZAtm
XninkGLvNSKXB4vcXkUAHuX2/JDprH8uRHuka67jul3e7iqoFbxs6yeGnGDtvrf/VHpOsYjusFyl
JQRM0Zv3hi5XMNYt6F5xj0x/isHs+HgkT2pl0uPLPGaMuC8Be2XFOqVvuSGkQx8Xo9uiAeP4CzKR
LoTYUMblfO3JaroThucpcWIQxi86gTQrUbZdok+hn1/qJMw3KbsLtcMI1xoKAc+YZCZNOahLfX/O
PG+zu3oGL3MT/Olr9z3vfQY1X5xQrhUhCHgsA9Kxps39ScqN/MpzVvXqVKERExmZwahAhN1YVuPX
/sH2dSwibMkjYBau/IsV8TAAemSBTlF0gcETUac8fTBVLYxZIFkvLOv1hoXfYl7YPdH9GXMQ8Z/5
+qUJ+A1YI4OCkjxYjrrfR+Qaacg14br2ECH0FsyQMf9RdKcoRc7Tq5UFFojTiZFcnp5xYdAwoW33
8V/eD7cdqb7BNknHg9XJBQ+ANCLVbBgldlQ/LBHtmZJfH4jSsgUxX3idFNq1M33jKnf0NYlpV8gP
yA08eIQ9JwAQYMrTQkbFgxe+RKoSWhqp0POB+JG7fdhtV3DMdvihCak0njGadH2iBZvC/Kt+xby/
J1Kj+PYPVfoyIBqT/2ng0/JNGVJnzUorKl8fSY4HMYU/XSKHfstXZKlBoV48QLqWwon/rX3Oskk/
VED10CEZMOiN51QnZtkggam3bsgabHquN/gZPuy1SPcGcWpZf4g9Wv8lRSqbVLuYx6xS/VAmSXMH
kAyOIT2ZtywElmR5DBOTc1rxCwgSQ/4jhqTQ1NnzKoCYFyyJRC4bxyPR74rI+9CT5elWpe7rZA+a
6jsz+YyFlrmjUEUJBLggSJRAKB4XCK7vg/gu2DhZEegEzye4spt4GA8DANxtFzc78ZFSCk9ha8BS
Gpfwubo9jtFygg7EMh1B7KoS1sJ1Dnvf3zxPBYUHndpMcC0sBCjblCob5HsFJq5woWCtjshZlVa9
RHRjcQSUemI11JgVF0emYIkBPsemkwp6+xhdqoC1dxcMFdIkmhgIIvxQNwUP1ARngmdbtzLbpc1f
WIPJ/rv0DTQteXbPpuxewonOWKMudfZnXvVhk6G7hgSYsvkd/VqX1ZM6QPuOeVpSWsA17pW46ZSb
ZEIPbA+WJlj2YuAGSzDtvIXb5kcCWSqnwB8sZ0jpszMkrGSz61It72GvBwPT4MNLwQsRwu6EtP7d
kdTbyd9l6KaSLHo0kJKSLvNa7KUTl4YqWOtpEOIx6GoSF+KnxH0le0H/tUWnhmpXAkZrmiQ5/3RH
eSI+t5fO7C7X2UszFEyEqnMTFJjLBrBXLzGA1DsWYPTxLxGNPQrb76v7cFGvOFMjvLxkU9Ql7/zk
DZdcmMOZnL+XetQ2khGl+eAHusX5magFWetTv8lav4ZHSAqzEBRHB8RGd5loIauZQjQ53M6ubsLV
c7PwTvvwHCQa0R3UPzbQSmxF0N4Q5vl5ugmmXZSn6ja6uJNCZkzXapURNhL1d3C0rPInipDXdAdc
/3jXiWyXaomzPZvLRgCgGb6ErFq43uMNz5nQfDFE8y8ue4Yw6D79C+njDIRmopwwSsCqE1UpAvU0
DDJS2uduzwoLVQojUVubbLBKgxpvpyCFtqADnr0SMLN0+C6SwsMPWxSYabA+GiEKSbkQh3lmBPaM
QCNzkg8VvoK0mrEBU633s2PwyMk0yZNbpd7HjUVQinGxy0ZMK3INhC7MsWwSPAX9dJmr4FtGjngR
t2d3ZBqg3RuxPJjO+htDv0hVGo5ENdqMKeOszAeXl5s4gcvDikxaEgUUOLG3RW1Oqn9sVf1Busjb
13bZ4UWh1SKkeMV69SaaBvJqYvKfFAHqpmnrc/o7zy+UinDj8L5C1XMbFCTdWdFQyjx2696LGCFv
6LELZc6S/+wH8h8X/12jEjhsnKFEw7moi2g+S+XLoI7fTWTlE/B2WalgIAo+2J+J8Zf8T7h8EsPW
yesk2kTR4c2zDC1f9w7lW+TjPQ7Qkko1gAsAkh2iRV0SxVozFcUmPEf/SlzyZ19Eh9GUPvCXlo73
VpYdZKdQ3xkKQ0dVhgQoonlC3LptFpKVTb6tAyOxAzW7/brlcZXqMl+9uZBBm76L/NA0E33zVtsQ
B5fk2sjJJAUWWNv8KY0+dUb7M2R05WkSV+Az9r6a5M9zOlYXLKGjVNPmMxWPHAdArKSuUWf1z1FF
KdLDgIDJFOVrHc0jaj0F24uVHzcptXdDj8lau3sxsZAzT2EmqkhVjf3OOaOpXb8DEtPDsFtBdOs5
ehJAouLiKPR8e6vNmVm72rXsnJ9BUOQovAfDK6ABKoYdJyL1jmd4ru0unPHwZrzrmqpPeOdQCNoV
rdiD0orAhxaRLvWwt+n8NMCEDePjIOgEMSyjbMd+MM58QYDm9J9mIrUa6qUI5QqKYivI2P1LLEt3
IauZt68zrHoL+WIoUgcwVmeYj3T4nvURAZLjY+o0wJWEA+hBonn5Zy8908KwH5ECoWZxlaCb5siD
1cBdbxGjKRtZT+0h9GKAkBrw/PNLzhi40JWkOb2cDfltyN58MMqoRtMsdkzUdIQsRYrGcCGCijG/
Q2j/lCFBJ6ONq+MTKGxnHUjiDg2tiU6GTw8RtFPtiVhI+1KGn0qHv79iVeh424tyXzs3vPbggYaS
Hmt3f63YwoX8zK0tX1l5YnaAXDMpA718UB5gbY5dcbTcFkGetQPXVWCuOGnGEfW66aB/Ebkbam39
nFuYy4pn74deXF5ItAFVQ1F6eAFqPEwEE+ARA7KkNQDvba5dPUG0TGvg4qkcGJmseemPVtzipZio
D5j20dk9rzNRsF18QpaBzK09ntqoptAnRh7/AyNhl85BWj7NBnXXHK0/SBYEy+HKhWS8a0Yur98H
fZfCfmUgxdsKyGFNSBIiqiklyMTPViRcIRVolcNLpia1HMGUgnUxqbMeuXBZYPSIBliHxljSMDyM
1YZUgepaND1byF4cagZdM+Ns6xg/ABJksw5+UItQOzLyp8LCBSK2uJBvJi9BClR0QEvzPxDceADL
ctQEoXZ/88RSHRJJpPn/bFZnomsTRffJKE2tYVkY+jGiL/Z/Rkqo57o3OvZ8qVhMrxcq+rY8fY0s
7soEDfs/XRsNix8u2A6w+kr92aMwlxjy1xrTncXhfblTF1XLEhZhtBpXiuW0N4bN6VfkJuS/JWE1
dsWy1PFUB64m9ycq7+RhqBCF04wimTMFvYFBx9ZRnEK3Z6xds/GPGqBKAhAz4qoSpCwL486yakt/
OO1LEuwZoP6k291Wv+c/bp3arRdkFYlndlNEb1YoFjsgqx0v2yPanFhqJZHfn+rGZLuRQU1KmlRx
vzBeyL8qXW6Sqn0TKWY4r/J3xw0WAs3q8kT634Gq9/HzWQ2yS5QnDGOn+jIgb3ySYozC3345sdDZ
JGdwUvSVCa0u1SMpGLu+ubQ+AUDatOd/MJboJIBw6MsZ7fxTe75gAXnZq7naHzRY7u9BY4YhDZxi
mbsobAy/qnYAov7+FR+dSE0WqA4HD991XexDHVutGRGHJGbWVQfB7ksBHy+PHW4NNPjRshOim/MU
j0yoZU7+Zkqe+23DkCIAGYRAkiok00i6dGuNh0CCHx83Ek9Ar8tcA0cTdspyWz3Sbcigsgj1UYFN
nnhcc0GniylectyHa6nqeNWrDB2ismwY5FWAAgEVyx9V4RYIQ8QE1BIr6l0x0ufh1HWNGEW8nRC6
y9JrKymyBZ6lpXPkoCzRtGmWWswKb2QxbvdUC/tq/zQa6i4yUwU7guhu0Ow3dqA84c6bwys7Hyv7
kBi0CFy1T1qXkfO8OeAR1ur9fF0Oz2rl8DjTFfpQZNtHpJSVaO/HAY+g9YQQVMDuwAgIK232rW9W
w/HpsDb/TELYGhUkvG8+GngJWwgEP9iC4hlpi+tYN2Po1KDq9m+AYn+XrZ3hcXbzpR2fIKtzbb/i
J1YWu23La4ON+9D8hI3mLPdeVCI+vWGJmsSmCiofhb0G4P+MdX0NnFBtAP/aRrSLXAwB68+xZMsy
THsOomlY2PS3na8AaesB8p86YZK9fuulJtXeL6id6La3oM5/mBfwL+7fojnKDY06h9e+z2fJQW8D
70Zaw8pwfS71tEno0oON0aLy99Vt+0WgiYA5oYdCTe38H8/1rQ9XDKTKIJWaO0Vi4k0dWaXKWDaD
MpmevAIMRaufs7PGPt4/3JbBVP7P8mhDVrTUPhtIJXxb29sAx6CcIG+q3IaoIBv5RDOu2laqFRsc
bH5Wy5qw1LaGwYS7zP+Mg5Qy/gb5dvknvl8OLMbCstykl8f4fCx9m3LNsn29xeG81mcc0d8lpEy7
4siERAbEjwftcrVSumy8jNHzcZgUnrtUjA17KgwYHJjBURBh4QQ/uIBcpQI7/I9nq7eqOu7aX7cl
VQQTFDz19BPLXHfYnccdBxMmBVftU7/9fD+GAHf4LawxdQs4Zu7G2j/38wGNuiVpFbYF63w9d3E9
4QyRcseAABmkZ741xaoDzqv7TF8c0rJNdsBC4GW3S+JH86MZi7oyU1I1x/LzAFqtHQhF58OkqMYe
NzW+ma6o8jhUBj0HWELCiDDZJEZNpnEYK1+jK23Jseyp0TpZP2n+HwaVWbG+YgQxp1F//lnyHBxk
25INJ5S09ldy/huYO+ZJXfzRWkEwyfHB++CWVYmnYim77SKsxBOS+KP/7Z1wYWdtdYPVU64k5eTY
RPC4TFKhiaGLTk3124Pj2DQPeiLkeccyd9GRuVumsxCHYuiugM0qoKK9MNWzYw99w3DcKAwCsCln
9A3GW9MjZ9Z7S+Abb2v8/WrxbZNlcuv6gwtw6juvhFEUMSoAsJwXYpYkLCILZwPqDRlLTowYRs8V
dFj7FcFyzSDrCZLzmVimTVRwfCsSwsC7wi7P0g3dqdXVJCm+3C6bf0EUNb7yq7LgRZ2vqKG5cKVf
xYwMLRWe6Y8J0G2oukPCdXnmy4mGOlt1MtmEK0zuvePwD0c7tcc1akWW3wJBCLAZLwBbhSm2IScK
u3dn0Gj0Sl0PpCJ/opY475piqHNNo9PYOkcjRqmx65A2S/by+yaB1j05Ri9sDeS6n8mzB/yHoeRR
bcIrt8TGjjwFecFer7FXaqdXpsrbTJ3xINAumqK+Uk+gO13O0PKBH1GAp6N9DhR1aVOzIZxrqlJw
ZMQq+gADa9lfpuCuNC8xir33zVIRq2GDAMTyMHS21slPSCa+2L6npANHuk74uhxgyV5OkgqpyQbd
KOwEBXXQed6ul/eYJQ2M+hGQmXFl0noyy8V7BeXJXY3Ezt4vk0rtp3u2/wh7SHTRs5j787LJi+ov
PKfS9YmrzH1fER6JHkTR+25PPQ+v1MlF+XzCXwWFwECzAGqPTwbMzIWWGya70LRjGZbyTCrAChM7
G3Z75DzDZB8+DY8vj+pE1yoesUYtP/YUZ3vUInw/RHHznVN+D+APsvJQcz3hIMz+lDYMamO7l3Qn
OXiw0DZohwzh9OQ7VeiDpchzs3rsrLfbDCMDXmN/anRJvaKbPrw7ZUc66JzfNELigtsAdqYVCoSQ
KC++OfE7XoaFPTaJmRsGLgyNHoXkSFdLkbke78cq8z8VWBbtOUVFINGOn4T5wdLvVNaZDoioFXjm
TyYzsT8jO5N2R1/jVotKedGrvBiL4GJhgJEX1RqUU0HvwNPujKh92d8Mn8EE9OKZ54/wv9FuDaBQ
iQrhSHesC/GQ+bpkd6cZoTsX/VDYiYljGrWdePUpjCVnd0vyAt2OOqTzf4YyZdUmT6sa39EIZoVn
SxVcJ/MszcgOF+yMTzagAMFy4Fl+48S3/KODfoO4OenNYWPJOgWQukqF8viHH8FXO7J38GgfkF57
nvrQi1XtZWg10e6fcbZJFZs/sMMFn3sFi9B3d2U/kiVtln9yNtELgmjdWwYxfjks42Gq0a11ljTW
sWYaVXN3d74yxVLXBMPzVJdJO0i858LbgRphCozrzmuZc3yf+5dUZqvstXdwP049USrsYZQzbXSs
f9sYBUoMCac0xuegaLtg/bBCDv9wJHMKyE04Gb3aOQHBnuB/ZcP5W0RHXPpoJ9qF+LTFMzj5TgDc
rNY0k0w/jCjzjLbRxvuBEQQGXuvRimh8dlfENXdP5L9f6rNYrNtm1ZF+/Tuc2c4BoGiQ4H052Dzw
QKRnjD2xn4T79oQjv3m4jNPtmKi++PqjXzX0X3IdGsopnj+8gFoOu5hNkWUiWccxAcSoSUn9YdLZ
d0PaGEy0KxQF7pMvTU7AvBxkHm5GiWJ6M7Evt5Oxiv4u+/rvBND76QM7iqtjxS2FHG0Ui+BdMaRH
2W6NqHuFR7hNUtShp9PbLwvEo95dUu+XsX168yUYvXCvyfQN4vuT23nX94Q/el18CKpVndw+3m/f
31qT5K/d+x1jAQ2NbRutodypFg0EjaPLnNw1n4zZm7iuFrsUMn5BOJE0kzbWlyNNwyuTkke/y/Qx
WGgUFGehZRvNmrR6I+1yrWSYx3g+AtcPjURMeIPuiIWD6XfVS5GJN11ElTkyDQAoPeDIwpLAQdKE
8KhlwnhVPCQd8zdyTuHsiKYUu6MVwFJ9mwPiab2lcgnzcjvCakxHBIzAuVxiBzWz96aBbbW4pL0a
LkquTIgmPfhHeA4jJXH4uIa5lsuOV+FgH52auHffFqeQ2XaMFB3uPL/Uq5fJ/MhFHqmlyEKX0UDS
g4XWmzZvP2gUwOJR7ElTzD/psE6GtHEEHrO2HbD/Wo+SuaZImoXzI0oyFidh7MXxTmQV3Qwr2L0A
t35XnK1PMFvNTzF5R0gnnMc+OHvJfSH/2xljKMfznJm95ef/prZ8HcTw5zTDOOH/G9c+vZcI3BQu
LzYCwUwVcu3m6MKsJAvI1quooIDR7XgUr2rKeOn6/9SSHbypVGoFOQwuwCNwZbEcLBvW04jo4Z5F
ou1q/HCemPr02Ed8VBMmAx2RU1FrsBfyckC4eUMT0pkkCV5DO57v9JQWFvljBidgX5zVHaAJZH29
4TfX5LCcTopxPJIHiiUv9oZneqpZfoGbAOiP/XF0pnvyJxyT+tDd2CLSmzAFQzz5Z+iLRN4OejeJ
FSYwXn3CfaAQHrx5WueYYomyS9KWOVupjNLLZu56HbPSjVdWyrnxnzG8SFopw9ZfM8Ws3VjHzIH5
kSmMg85oXrwYkOREAf8RwoiOVq2BrnWcJY9CrhgOMROKVV5w9v/nsoKEpOF4btXl60G/8PikblXa
zE8eA+rkchf2i0iY4iPbv8DxJzW9zPB31UjS5ElzmEL4day6ScDz/d5Dt238Cz+WtnUvecqT7pdB
1YQiWaX4LfdqAJB8krtdKkHZWxwOwzhupiv0KJU78r6XY4P4TH/w3b1R3+A32t/z0/5pzHErbVce
8aob6C0aoETn9vnu5SIWouq/wEykgK1QMoVibG3ZwA5BJHUtMoo5eeTa+dCzlTidwqvwcA4aNwgJ
9jDhRYBNyzExhdWQcSGy6oAIQHQ7zJAfhkLDLZb6dkeKogb6cEM5Z5QG6dlRWYZ274dmovL2iGCl
fFF3+S5ofGB7ROBGy7RHlbACfTe4mgAyVE/an/uAJ559kenlDYnHzxFhlSZwG59dEDENqbsvMCu2
F1PLX+Mf9RGth4tiENrEoAUttqvNSU0A3tnOd7EsLaI6CtZkw05yHF71f/XMokH1LU4HOL+Xr4v5
f8/0tGzJvS4Cq1FBjpUoL1sd916WRHSwJ8qbcVzmfDrT/5XfF1GthycFhhBsZI+pUKjiODsiAPOi
GAX/U0KqVGUuomRf0LzWBvNoKHn2zuPoAqUOBrWX3oqFAApg6EIK6QINl4yMRFl/NZYomFGMohYH
tyW9Sn8d0bjyx3L37mG3E265mesCymJrEjuLjglpiHfRtpAAvWYCkfws98xLviI1u9p7F/sSMMR8
oCN0PA9JDLCxNCqXaX/75uTnv/zl0qMblsrJCEL0fjK2z0Z3bfHpfKRZuWaycWhl7tNu/Iai+IUA
AVWzUpEkEKrI/+a2EIuFJnxTRX/uUSwW64Hjb8ZnyvIVK+m2H02IN/Qq12TZB+IHK2mOenfJ0N6A
pivx3FZb2Hr9RJnfpvf8XaI+8IxTQPDqf3yrb5ITTb6w9/wahatSkxeZ7DoUT0FbM0fB6Jt/+mlW
XS7ASGxoFc/c01WlE8O6G0utyp8N5Jc0Ncf7edAwKWlSvawLwLPMmuJcVKhBs0Ecy+10udStuJKj
wOchR1dFSn561i5hP/MH7gXbx4EaCXKNBEbFbcxTZad+b0Bjin7cdkNiOf1/A9JCWKTQ/vas1Qw4
mB6gDE8YpT4DlVv7YVS+Ancd+TShttWjYvz40ChBRS3A4NdR/P28n95VNJFxQcb8dKrp/cxGwHuw
kl2D/rXyxfMJCKm+iNakmp/dMYAT7C+LwnFdDEat5Y1F4i9FBuBtXsUaJezYeS0n3+j6nlfbSdAx
atvcH5BOjOHjxnfnplsi1hJdi1V+9nkmaxwx1AZs0YpIMPwuBVcbBGfyRQlLq2hgxMidvFK4Nqib
f6VmLpCwmcIq7yqiJDF1eGnV+iNFiRvn+NIzcDZQaW1FacfcOGb2W5khnNnY3A+GzhemzoYS8L3L
gUlw6IPZU3h2Kw3yj2im4cTqwLA/Z5SPPRTdV9ZybxPYY4z6Umudb2rUD6Y5PlNeh5YIJjP5t0w7
1PqTAdDViF45dPTU6LQ8SXWbwJKjACVqUIUw3RRCq20glT9GOoWjKVOWgVzVCwzMEtYS5vcmRMeh
rvu/KPdXpflxu1RZoBA1Io1uf4/Q5FLRR/lu18GbZqG4HVbfJKljYBlH1oAR+OPCyyrLKx4f+Vha
ySPhU+O13j5XbLpPcrxnsInt12QcY3le9cSSYJl5A5t2+Ll9bTlrA5Q+d8fnBl8lgA7eS/P/0brJ
CuX8no0TY0fCQUUQauISmj9AcH9KPemJ0Rs2DELttsm1e2tNbebUvjQLaEDKHPcdoEYk7aDl9/Is
yFkHAx4TL4D+Ym87HhnjN6yBC2oLe6Pi/PL2ZXOa7B1iGGROzodhxVRfcpe9M3VJRpMIoG8N6gNZ
EGvv5DIm3/mwEKI/2yylq6a5/sER9Igu9G6zcHa9biECsdNnVd9JsQajYpCSGvw66E/I1FRvb5Eb
sPi00M+slEkwRb4IebH3e+NkXPWvC1eAX284NBPIO8XQi2+EUkLWETUo//jZZ8ddOUHDun6jA9lG
kr+r9JqPagydmuEIytZmskEUROzXH2JZjhLVxjh/p7oBqRz+i6LJRV6+NNO9KxOCkCRRnwUflXER
ts+mrGwVRCuBw/l4yLNuxOgde2cKcNsD1ef8iHtOpY7nuU/1pCQxkwD1PlcIn/QDsF2GiQjlfG3Q
Xa2fwnLtoJK7hDcSNTxz0wQV4fSPIESaV+6ILmi7V8dz2EZjltfoQxHPxtLI8KVirERlymiNOOeW
Yjazh3U1ihRwj3DCq19HUnAuJTtKuOEKAXnq6qdkyGbr9mB4PtYlGI39eGtyMXUpXOdKJ4z99TRZ
uaRX/cG+FhbbLLcf8qGzbecB6IbJCqJs1sM01ESczhA3aYDyDqSVBPRI5qeMIA4QVnv9kiGqtoMS
hlfnGW25CgZ56uaVNQ/M2NrgjCMeg9fojQZwWTn9Tgj14u34ZEg1QeaaP3cOhLqsJkD26dlIwW46
bCSOm3hTp6jCfU+4hF8riUy6QT9vV/6lDZmSesdi9GraMy/E+56sKMJhd4voM7cIz67eLwka3JXF
CsWs/5+x6fpeQGaIsOBSsWCdb2R6jart576fWNjXMLC8k8IeZbz/a43J1DejY5eqe8mVR9xLmZTr
FbI47KF7eZPlzI8R3sCi6ZcXINVxROrXw1/Tbdzc+uop6Cs44o8NBSUuMndVAkACdGJ0m4F7bXS2
i92UB84xWPan8oZm1jgJydjvXgJ+wTjH9l9eHnsN8bw2F/s4qPlTmR5aWJUTAi7V2uYQC7zEdmvC
BpVs8bpCBRkgGvybmXustJWgrtgz9pUbk8Uwl+2Mp1OlKJ0aZ7CU2w1puJwsu+2knPNOil5mm1RH
5USgmxrdtkm2VNfQPbPPNVEhXEeuDNl+6E4E2JtpuTdmaDGFO6kyLBbh9nA2fUUZQHvOqWYmPLe8
PJ5BaTDkZXruAY/HQPd54KhAUDL8uKBvHWmGbjxmLKX/a213s1sdQFdH9Px/xbvSVjpGVL/EN2zu
OjNoGfynLv3/FY5D7fd/0l6QeJFHVrcQazSjsltj1mZ3c10VsT4ClaaahXUl48YLkcipkjkn/mCt
vBoWcnGezOSIp3XoV3BG/Tw1QlXVDBfgj/fd0KkK5GbMiD1jjsCz07THzX0TFDrkri98O9PmtFj9
z7LGVg7SNcJOfPUJ42l8oVUKNG3ovd3LHTQo+33nDFYCthjlzZL/BKrWRmy3Fms1Z1F7gu0QkM86
XuYtaFmoYc034d+mJ/IUE+wldBecBkmV3pi6FkhQN0gxZL82xV1x6Ji2lEn6t+uAiG8dXfVIubLl
VO0zR++deinwJwRvt1Iu8xb+Zl5B01LBLMs9mrljMpoU+X1LD3+7yIPGbgEnehCMkUCzyuxfwKIk
vRMLZEDVHnlx2Tmfto1DFhK8apRJIhfCyUc4g/RhpfKrJ1FYfXvGV7vWDhs3xczCN9nSHkSP3cfm
TPixZT1rR1b059AJ7ozRw/y8kmdzmt0IfkRrLUvToqKFnKNCLqCZ8EpUemUEqVDBW56l6EgHYkB8
mNutrtmuQf5C+fARhI6RTlY4NqrKZzXvgew8+0eVSiFeR/pYMvEgyszR1mNpilQUEHvCeiTqSvGD
7kf/ZutVQIHLWkouWv8zM1uMUAGBLIN5AOGlobMquOf991h6aaBL3VruoyIBkxzxto9UD/S3LCjo
0FW0z6BVblBXKlrsgmOIdnujL5m2eg8oGhVJzTh5jK9asPyRO3D8Nli9TGX2pT1+B51Y6FLGn/ER
PvyCfZH8x3KIBJYIrpUgTSFKtvtlG6zp5KAqXPkq/IWyglrsTY8WLJdbS0Ufi+XWgv6i5X4IURyi
DeZ2Yo4lNhzrWuH6t32a63ixS8cFTJLbKSubGHFFa7DSQwg19lWxvS5AbKPrhfwnGwQNY0yn/VYF
cnLaLsLr+3VWDgxlXEwwcB1LKKVaVwlie9YJ5sVy0d0NN2582aqzM40kRCuWs1mzx0RZ8dx4dZe2
RJfORLXZbjnOAwI99A3/UnjX1Jg/Yp9PpFKnpJrGTJhhPZEbdFmNHhMX9uWfNLSbBkLEf1+5C9rX
8wTUvltAPbIKzxon9rQNF9GIXUtNaL1QjPAzIVM8fn4u/wev8y2zB2BzFuJabELWWeGtZKw7lEfD
FwcaG9F0qFz9A86zo3+hH4Qa0iWba2htFcvlA6CWnnRiCnzvz4x+tOyebrIT8/tmHc1BCmfcf4He
OSxzGi0RY8fL9MN23iwsAupJXz/yNTHwndJQR4It5GIbEDX9Myqt8A0H1Nu+2+962v2wYz69lCry
HWUJEIUjkGNgt7xYK6yVyGc4hjS/C9uC3uiWkhI1u5NPQqRDzDkoLeSYwDZpO/OoLNBlW3Vhb/CP
I06uDFrIXUujEGlXnXuJVRYg+bDliyOhpeOxnFBWhc2Cdc2GJnbkdlxv4NVpFYIQYTDzXACgQj7s
DwErfB/EhdhzJsz80g3MYroEKp2B+ZWD9rZssZoCzAp2XstV7qf98nmEyOsRq3beLCsB6X7E9bdI
gmqreYeQESJ66AUkoO2bwp1BYOilIjoD2jFvIuPowX+zgyutk4Es2rhipWTWINs+cQWV+e61gd3C
ut2gGgB83EA9ViyHSnHuy2Ni4XTGfXrC+xBD3jBG3/zwVkEEOVLXcmj1cIhJoFZp/Ek8mBq4xiPy
lUxEzpZekG/8N5Y3KfiMj/VfoaGn85HieOwtzxYYw2Ps3hNFAlFjw4zHWX62FCgK7h+w+oDxrP8w
j+ZeJepCKV1RbWte9QPvhYXmCs7yhEhitXiFVr0inP3Aez10X0EuRXbPKAyvLPrLYeYoaOLa4r5z
2YNqgwBulSC+7rYZ+z5JNhwP2czMJQ/fhCmLL2h33gpoJRAmx1ogMCk1gw8p86yruSoISADtlAsg
RtAw8Yxp/mKO3bNapJLu0iQpC2Ic2sIDFA0hC9CHHhd0Kk6cN7ZSCslFbrqPkh2nCPMGgISVDF4k
huJSFE/phRNts2OSbXwTgEnt3aO7DlP/tnMn6fDbdbfoQdm9dmX3kMVg7mqmAoO5OwVv4sxKKeU6
Pst8wVogofZ+ofaiclx1j8yrtjzYihKdnRx5DrsQGymF/c1/pXMwmHZGcWE5ebin4bYm2Jg8Qr5B
GlCwXANokgTqx4ma0zDYyihq0xhGYJR/JNMJ+y4ghVo6DUXAyPfc0MlQ3CBeTMdkki6cCllRmhS4
t0imtyfuXieotzeXj5/LfjoVyl1K3dNErvs5p5nApYJaouGofLdUl04rdQB3Hggs2NVeo6ADUAN+
8lXlAhnnhMHXP0RLMTG0FlJrX36ccOpiSXpfEAtLfH4gF8JGYV240k8pI63SKXaDAU9EoO50IM6k
mO4JD8WdWg4GH0t53j96sYFhQWBRz8d9yIBOx/gZ608WFoc0VPh4TIkQCARy7nOa8QRycrTcViWh
2ytd09PTFHwsHXU61qcPfBKnbLVSaaDuQKT37U+8spvNiboPIc6AD43lpVjlF9p5pOIENJevdPro
FRlzH2SxVH861kblywQsnVnIm0H+NTp2o1zGmPwctJJ+66myB8f7NxWsPEuCqcubeKSJGRnmGtCc
2gudKtgbiFbls4DlEuGKIMBFpVkJuEU5gDPsE67/goSl4NTVq6SUTQKMhxTLLDdvs6gPMam7cSn9
FY9eSnWbKb+ex8/6ne58+nzWwVj1hWEF8v5809oTRarzgbno0k1QCWQ5P1AR2MjlQLXAy1+Eb168
C3aDLq5jc4z1JMafzbP/9srLBKgeZxrjUHTErPuf0V4HU/m1tJVQL2mQuI8LNawMoeJDOiTH/Mh5
A4NykNg4U5NZUauE2SmpRDFNzIwI1tkL5u9suGQfMgPg6zhXzdtMb0h6IqfecO26T+/3wbqOmIEv
2eoCiWdQK809TDUYp5NujkWPYTQLS73YUDejmkidYwSAW57iaGV6SSzXxprAaSwm8o0nEWjF65sx
xaQEp7PtQEDJh6ZPbq6X+wW8BQY3nBlVdMPOGaEVPWjhpFwkwu68GaW8vX/eVHhLhcxNTKGCLGdg
Y6lqvirblv71jbDMItD3zxkWrmG9jLo4DKhyhNOhyEsQ42/S6CKlAQOvuNBG6lc9U5bLwGPuRQxx
wlP2+acsvR6GDK/iEk3kBjsElS0L/zhdqMOoyaA2MQ7l0n6r4ZZN5dQ/YqvMo4HnxgFhOcLytdVW
c86ZrgAVK/7/ph9Yrrs/BQJKn9dogwTEv4iNWicMYcrGTmgQ0oxUI9TVdpg+J1tPEeoYN0ovshTS
j2HWGDug3jyPEmgK1WOjZQaaNmwcW3ApwVcM04FT9rMgDy5L/DC2CNJgbCkx8a6qxmRU/o/qsiZO
y6nzjRr3YrE4mJBxqaNipcJ1nRcwr+HBXc4CkO+Oq+oViLqQGf5Af8xdVlLuhfgm3BkNLrks0jTc
pn8A6D5Lm3Qqy4qVRYpJrvTVHat2Sgt62f7ZUNFXXXX4TusLo7CcX5PTCzT2Kvtupqr9nClj7rem
bQHE36rTosPAUPq60E0EEONHXOCJl2ikahJW9DaNDeEtZWoKH6atswGaB4TLgy4Kwj2Zyo+BZ4d5
iN+D49Hl/DHtagIElJ35AUjL5KrULoH8cBMBHD/TAyLyVroAjVChm1t4ZbGgyMFiBsYXCY02oTwU
WGtbGpoJD74BDdWKqOGtiDseX0aoaYlxe81QngCVm819JqaBz3ePHoMqiOjwL5P7y+W/iisv1kQJ
5Q1j5qsqydATnNNngjLF6As60IpqZ9wAuzZhr9KbhoeSVxr1lfckGG1raH88UfpvIx1j00Uj/sen
xx86i/QBuiasIjRfyZZlqe9AMOWdcgOBuHy9TFmnLGtGqzK7TBEMPH8c1kg1QqWWlSt1hDYJmOxk
gU9lVhj1srIaBBIynbJos8EfN+MWC3QbZB2yfgFWPkguo5VdLXc7G3EIW8N1BGFHCeTahGsyIHtt
PDbnVdIkWJYvZ6NiiDYh0AWiezd2hfZzJis3pPRpTJp3yFXOD+xmFfPjlkpVjmF7CFwzpWs1Qq+N
68+rLYxTgAnUwl3D2e+FL6aihco/XZ7ywNLiN6JGWY7JplvVstRTsRjrZz3YU9sK7r48EUaoEfvS
xdKvW6iIMwaYyLAGT89NDXU2UxesatekmW39U3xA9Kv5GJ3S9ln5vh+PM37s5UmYyes6E+odOsFV
zV9rI0IVRousSzlmRVNXIIR0e5/ksENunwiK8lBLamT0vITou7qp4oWtaNxgY7laN2kUr/07WZXd
541dEiwEDA/2FkZbC0eCHneH5KA4l7U6K6hSRiJv21pH8mswTY0NyvAEmD1wVCqk2Od59WkY3qeJ
QbBHnaD2HnpTaNa8tFoLPGs1u2LBVMuDe48CRkIQxeoHP77/PGsT6tgtI7+GEbn+AV6aQfGBdMdd
vmGUKwSRPjvYFodTb3KwxpfJZq8yffq5tcjTvqWcB03KgVg3Z5UQj8pm89qIW+Vytm9hKGYiaO3d
UBtD4YPpm5XihxMwVKqugkPxY1NigGPZ5ATono/6zyDZDcQOkFFmwxEhRAx5PJczgORzpdbMuKr9
SSLbqZU+/wc2iXLJTXnJqg16cn/DViqGve+IrOJ6XEm4tTc+3NAlgKx/pj9gbdBzyu54GYJbUC2B
hKAU0z7t5IH88cua4eA3vEhDhnbhrAIi/OPHtYx9TfSmYxW0TgmFPFVWCQkzY1QJOFmt8+4Vyiac
ZPxLuEI2L83FSrG5EhaLKoFvpLogRAT5a0qWfwArA+pQHN0xQzTe4Htlwg0KmeXQCXanGKZhGMKg
sq34hZexrd6+RYckmPMcQkJAI2iAuhCv59NM3+aqMkoGtVLKftLoHg0vELQL7CnwkhE85KB2YxxW
lWYo2hK5Zk1mc/ZSxC4SRC0vN9AuKH1CTcWc8xx6y2M1JBBF6JS4FtN3uQcD+b0UgMl8ZjPoGlhR
suiQTFJaaZRs3L6uK3RBkPCVeVeYXa1lti7l/j9ZWJo3ST25Z5C/wokRSDthy3ZNWbD55LHdOkf1
teqJsZWBrgx4NcmN2S5K21YUWvB9UlgqdDyww5GoCc1mquhHd4v+AXyCp0xvJej+041y/PUho4TB
5VGAST5FFYlGTl2tTqvlBeaMYrYFI+vl0AXn5xPY8Urc60GvV6DdJROIEgtB6dCo0KdEWggQ0qQk
cD9GZkfxP1CAKrqjuSEEM6e0Mj1p2CxWNwmZz22LSqR6X781z+r0fA8L6VlPFCjvT1M7RxLhV0VZ
JJCJ8kyjKb/Qk6svhapVQD/F1OmmOlsRW4kc1NWCKl9tul32McVTkKSGn8lprQpD1rfQrFkJyMF9
13xfCXBH7O7ceiUEZbWTe25we6yNJc5HIAtZ3xvoqWEhExe1FM6+I4sVBSGrNLNX/9bpjKjD+6mr
Xp/OatghoAgQMU4MJQNCAJoYMJY/zfDrfVRzN9bEnsj2bDfa8PjfmipetQ7zdlfo1tiZRpgnZtA9
QVXmHJN74nGNesp6KyCleYd3ezivm5qarJpfsJ/SW2kAM+WplcQvq+YfsMht7Y/mZOfndQq5wnPi
cAfoQw9IdkZdJE3bFkfTPZeuoLuXVBg389IBn5KtA4sGQkQlKVBjXO17JmyHbvKVtuJuWPJwycwd
mEcThF1V8/z/Fz3xN/CHM35RAsD0PrAFV+mEiTYod8b1h0WnwVwuunkFQCstqmr2Jug8gFX9HMef
Vqf+sSmLFZF7eGcdGlPzuYn/zpfnWxUX7FAJWOhXf4MTW0qRMedBUgYtnG4g9zh/JFJFj3d10cre
ektLamaSwQkYVXB0sBgpyuNoA/yN/kvCn0a9kAQMNbTfS8D5SxHIEjkMiD6HNZLZcN0maEgDRlnI
d2ulZaHEcFPHZQmMqkB/cOWvSEaz+mpob4dr/LbKjb5PjgpsC4L7TpXk87n6hQEZoWVTFoTesZ3F
n7Q+c5oapzwzuK/RI4oOQhXP6LCzS9aI8Z0dEvboHbXcTvgxAQDnatINVwXkg9rn1upkWdyk73gN
ovFZd/9iLkZQWGPmZkL9+IvRq5tn2Q7MAO7IQnWkRV6ukn9/ED2Yd70nvCjNDFRgNqCSA3EPnGO5
a8LkDlYQb0f2kJK5K1jo0fwUENLuJYNEY8f+VKPZi5YNr7jxBIA/m+byHaVGQWH+zl1QeI1IgJvH
MXsJS6xLSnSfZzdb5ZtOCy3wCUtxohYLTXg//a3EDCmG2rMIPqRhkqwc1gde3NtYqlsi9/HH48st
rGSPc5BdPlpZjE9rDXw/sJakXrMc3batO0b6CnNWAf8le2nCvLr94vlPl2/q3Yd6bOzme9V2FI0L
ek1kIg3wizpbLxVp67ZTAVJSsmt8ee22PmKMdma8Uks/XoqEeHIWX6mCaEmaGfY3Bn7nSaRICDYo
cx1adtaG5oZp2phID6YlxTWt+IrMHR9HrYeoTobvRX0oUPCNPcpyebe6J0tIAML72t1GtKkTbI6W
pXjX3UuPP64TqxFCvMDBX8o6AQ3naACVdclXj9yjx3qhUU9uF69enBj13DXnoL/R2NW2p/3Fsk0t
Wu/x8lgc/6/y2DYJyQ3LTDfK0R2uRtexswqOIwkvrufEQH3i7gBMmJzENtREAOJOOhMcaZGdYxwA
JsracnK+gFw2tlkkpIsxeZtuiMo5777Wjd0H24ydjOQ/3ni9DKwZrNydbnB/Clar7OgagDENoLlb
4mH4bCM5x8dMc/0UypmbOrplc7HF4JLyt1X+Kdi9t7KPTiOgosLWKGSBjIq1db04POFQJZxKXPGz
eRTcw7hXQVpjQXQfTF5Ql8l+VozNL8/LqRYtLoMI5IkAHmiV1ft3naVkNnhOGCWBlR2DcmmsztTf
Ojmh6nCEWJXq5F5job89KG00lUoGqNcfmLgXlmIWpN4cgLhiH+VEs1GaTBuXtKOFMv2Ps3SZ23ZZ
fFnfz1NDrm32m0dLlzBC6p0YOAq8Hwe/YrE01nx0DynuZLQwuOFoeDubpo9kEIf6k1lYhGRe38Cb
K1RdqjddGTMx+E9gttq2ExVYS1HbTBKfG97Rn/V4vRO3H+7g3NHk3+LFnNOl+u4x6zR4gFONSolL
DKCF6QaxzlEyK8aNbHBGKx1OYWQs5dQzF23dAlG5OIgx6lD9HsMI+o5VbAsTofzq2a8CW5wqEyKW
zmX5mBzn45HTChb5f7cPBAfTuBjUCwKlYsy/92MxxPnfeNoeCMV36sVkYplWocN+VErE6JnqIg3b
/V8M6LblQJe6urs1u9nXp8X8GcjU6EcvV02VXxOTUe1YrLz5YUTXQH5SRBBKnh6ygcQpsVZ8H2Vt
GdYlWb4ZsAABTVwlXNOKInFlvCOg4lEO6Ou0rwTMLt/LtDTtxwiHoWl1zH5rnD3KX/nO5MwUVpnq
f7yPpQNkt8h4kAr1qm2FyETzn+JahObCgZXuAdhTc3Uk1IE1VdEhIhYx6NHaGXMDnOj7AtYB1dKA
fU4yIBFX69ldGXVx9vrC55KqT4vyGYXZfEZbzrVg7Zn/wHzN+ECVquTr29yNFDhLtr9jioxav8HQ
injuX2Ms7x47/G5xMO4cJw6D5AfbVFVu0808ww3e10QPAvf4pjqVxwgNoojttpD5cfZVrExXMAvH
eyLtdLrNzv+PIpDlFpjhqaaIhQeJGjUurpvvX0BSSvvIB1ZGx8HdwAUO3kqJM/IiFdkngIKRkHsI
tGmAotQ9VuwYPXKHb5JZQvgMqNUAGssEXLecbQhT7J82uYu7TdcrRwV9VIVsghaMBx4KyNCWCCA8
Cs41s0+3bl3r6KXs5aJiAG2zi0pjsnDcYJog4rWw2MD+RWXHWNY+h/mYAQbnPaw3QsHQ+uY/VIsm
u99QE09vn5K+juYgXxUwsUIqWlE1Eav3fhH+zCOEq6qJq7Yxfq1cJNM0YQgu47SMH8D5nfQiMGs4
OTO7FCH8jbtUnE6oBlll/vgWQLHucESDKeRX7kpXc8eTD/aqnXONTQxfJTwEdbXfz6gMchpYRJOB
EPOwzrgAo0tlXaUV1xpo4b0WfqMSaVgktkV7kj/wHn+TJSxSG+29ljfOas4kOmdszukdthnaU6Z3
C3s5+F3cwD2KfP97fGs2yBTvQHAJFEm171wZHtI2Qa06oHDcnwKCr3vo358ZMzpW17q7k/PH3D6u
Mlx8MijIZ9lbI60fKEvN15NtWoUI6r04TA+nLobIx4eRfP768PPqOGC7Ts4fOjGNbic2piHZYRJb
okGzzCywhFD4Pd/MOQmtmwO1TXubElSEj2tFm4XmsIDxdQTSvYcYNNjAgPmeeuLPhqIWb1MnaUdk
f6ytzauPqPQtWjeFOvAhQW0PMLc2I9TI2EM0ISJPlz/APxfXCYs7/EvoNgKnFVazw4qi7fz62lxt
24Hcxnq8I6s0xs4m9gst8/H0rNYDQNDFcKVhNe/4LgUxu/hZjr6Iz5UBz0QT2sntyUb/6PNVhq3Z
YZh1feLPYxFVlNy7qNOOWfzd9V2NPTiIB1E+PPfAOWUyeZhj9QfACRCsGoroX8xyROtmgKDxrLjM
wt29UVVtoFtCKdEOqnHfcgrtxGbv0SBZrRHxxFvV7g7xNo82TWKAsRmKNoir/NXBOk3fVWr8JxnT
9kkmR38rPm99Me3C9SbpPbk/xSjSFUg9JwEV8/moafLfN2frmpib2gSluLUrE25HzunDyb0vtHyn
z0zGRoZCwSwmkwENfCy3uCjqAnQRpCeK8VqItvKlHlOSPvQYbW4hHa/n5d3D7FthNSs4vnIRbzez
DCr0vIcePKeVi/zkXgPUs9nkoqxXv+wsKT18t7VwniDdwov2GEetcYLxKuoesqgHxym6H5uMhQEa
GYU+JXZylEnKO8WzK/Qx4wSC23PUl4stSUzCHdBHduhCnlGI2zkrj5rdRc5670rE7HoY2kHYADdA
aaYQiiqifkQ8kuXGxKtLx7MJecHdu83B8HGDwj4gyXZFbID8329jsiRiOkd5r/KCaX3ABJHioEY9
FYQ9y+IK1SKZf0Z9BUnmvLI4GyY+yihHmS/bSUPG6NFgT/mxkmVgh9RD+cBZnJ7L7ZhYIPprxnlC
o/Txyg2D4QFquFlvLp3JSK793pFn0VhjYpe7roBJFMVDHVeC96hMObxTLdlv4x6qwDXyB2bV9SCo
XkwvjB0v0NFTJflCAXcj1MgfuomvXkkKYqZZpJofMpGjvujMsCvdpWZetFWay/AoClGkr3oxx3Sq
MvQA7DOZza1cn6Ir8/flOJD5/kPSqHxOA5pku1Usvp7hitCc7v31cqwhzPJg7OrHg5cBWtDuuf6T
yZiRfT6FW8cm3W+2jbMTgr1i39acq6cRef0ZsoUIGBAknK3Sa0/+XV23c11+TxcE0esk25AdQPR6
9A6DxhOZYPI75GrbX5vmL4Al0KsegDKBE9TcSM8foiCXWKvPeyjzCywZa65rdCJoapRBkYZfprsv
962AYoVQ65Am4s5Df81vbesLXhNPI4SOoW5SbrnsqFXd9d3wcz/JidVsF06Sb2I5jh6WOI3GqpV8
sqspWJNyiqes3/mqoUzRgY/DJhKWJfweIqWTVYrhVovP8+m5sQbGIz+4TztgD+pqex8+wDNK6sGV
tpSwALzp8vT6WcdVnCV0uESO9dO9jay+Qqv2BQu0+LLXjtTR7FchpHNtHo9MIUdOt2343pnvCsQe
ysLW2MWZu+jsvFLqjztOS7J06ra1VT+TxV362GOWbLsKQQb7sKMDjFqTwxRmhLTsX6b565QH/hFn
4BVh/kY66FB0tZb65P22PFfHlUDK8scH8EngZmWaC54L2xCMA6vQRJkA16Cmcrp86UaGSCtIOvFn
Ob7ERPhiqD637vJxQv0E7TST+H5GqqrAwxumqIsjOialSn4+Gv6+c0RplBUWp6Rwlz3ZEZaUAbZ6
psq0+AwI6+a8NaELi2r/zkE7O/FR/cjNNuxbFnpFCCQ5V+QzDBPTBvLrEoJ6h8wkArNOALnEtAj4
zj/w+cPHTPyFx/+deuvBBBtLEf7ll9g/4Pg0YX2U1K2Va5Xr66+2kOr6FoXYd4Ni03UYGLRywwCZ
eiBd1/weXp4iFo4vrpn/p1epMCL5GM2h73px0ix4K17aUUhPnpWriftWSYhgUtNMNV7/M4a7TLW9
H+wpOZpkhEULpY1S/jxmwtOWVp9xIH4SxaRWifvaQw/EcHGk+FbaRiKzyuGnlCCmsyP7PeuNzuoK
a7QEL7WYIJhRQIr7dq8G0OrFY22/pH+wL2KDhpattUj3DR6VB3dpybcxSeuKj0M25dgxDoCEAF9W
zK75AjF3yX7Hz5b1UClgOyk1HVEtg66rXGswiCGs/QLuwBE3B7LUA9VYCvoVxE2U9BYd4e/oQh1W
8Za1K9+oUp8Pew5GBdh9tR63LZD1+yRuylPZ3qwr/8k7o+PNmrmvN6HfgQTYij41RNE/ZXxmpr3N
3Gs4e3eaP72R+Vz5gx9FTqQViJ/f//KUAe7RQyZSijcgSeXfugrGGycvKWTa0OkXKcAhoS89xYDR
y89nXC+axftJu1vmAIZSrvOsLHBJAM0sEsmdef/ulHmRYm5Qf8A8bb6/i02bmfTJPltmmS88cJ4E
l3lYM3ZjCJC3Q72T7eI3T6lrjKQaoOrnqQrfMpTl4vmad966Ffvya/x4QdPUJdJ+Qlng5F4d4RYj
Zp5xRlpOBWXVBzrbuuHQxVfJe7yPNfHBOA2Fe00GEJsOcSQDebpYVNx1XfKA0Qp5DmFEw8XeSvrj
wab9LBGrFlCZjSSK5gCUl0B1LFr72rpo3+fUY+sDmUGJyoLRntLDiSYgeYmhmh0pGz6GkqQpQlOC
U3QmoH6R0Cj/q73ZFq54H8Zmy4Md2MUV84sbZJ6A2dpt8uA3quzeP2/bfyRynHV15BT9PT5ogz0g
9TyakdroYA9E4GJifn2pWkFYWVaOPg0pzHFGT/PNlN/qqsdURRQjrkIPtX0bheE70KXXQfWgQThI
mfrTwHvAmubcg2YZI5bHKCvyy3GISLVUrcJitmLIGrpFY8efCt1NtsamlAOQFyvsm5fTKO3SPU78
qmJ8usBA+kzDNhzAqy2aDw4WaWu1p3CRs86CrZKn8erj8DoG2WtmFLmNCYZpq5r80XYCKC0Fwt6E
oZC7aQK5l/+WmBrOBD0oPiTKDhsLlVAMzTyGpriSNmrC4bvubAzSEM6ZwjCHAxnC/lO/wUxtDYtz
6qwHWo4qgMYtlUghWToMiZcVB1YX5ROnfd3QslbjqSEIpkcoZZko930kvGBAwV7RuUagc0dAHLHO
E5RP5zIQJUQq1YNyxUuKXInggVd7B4y8G4cX0rDuM3dOLEKORJ6l+ZwcfoRs5AtMiJY+uXFLH788
yw+1oDEVc85AqtM2fX03Q1oAIgpn2fsbFejd/eVFwjst125e3h2Bn0CXcDne5kJ/ZgHb7jbmdgka
CVkLAGukLRys4de03k42dacQxGtHy11ej7Bkb4m5HbF4jHo8NgqTlO9g7XEGqos36A5dF1is8IM5
EZmcH+4y30Jqd/T7qgw7xyIJT4Zos8/8os3pMGNgfhWZDAh5h/1uud2APR8EFAdu4fxlpfhfA7Hp
5iSwmL9pXuClN6Av2hBuqptZraXNqwZS8iNDHH4Hgayzci1fTFXnQPPBWRLHYWT1M4eYV+xJnVUP
Gjy+59xqIrnU7fQYcjblihIsuyRmtXhwk7t+VJyl4s+sC0mdGwoioBlN7ecazyHMiAdA7p7oGJGb
xWMUoxlW7YJ7sz7FMqA7rwjH2Oui1jmSyEhN8KeKhJoOxvWkeED8oUFKrI+d5Emsxv+O1uUSeJyg
UfuSmjsZzBieYMGS8Y0clQlPbfLK5RgI/TPZ2sT2hhu70DvkBEpjZW8PoXOCz1jtpihi/EfGk9eu
0i4s9lZyrP3gJINqFw6wifpwnTeIRZXMLZnlRwaQuUYhPRvqahRrGPfyF+uCRyW/loQpWDYwmV+O
urAgNUNttrMlUXJAKJhfiU3QJMYNhWtU4Han7xm1+NaXCo337RlxYyHVMihNWVA8wzaxikFDAezl
NozIJ2LyU8l6oV1WkPI7Igeru8Lcihpr+KOl3jmq8nSnERI7qa8sDE8tUMwSfRqA5+HIf+dK1e2N
fyB+Hr+oQN+5lgNF1b38+u+qnnhkV8bOTJD1mx3g2LZcow7F/Vdo6oOFkH3WVm0tjC7fZCSKTo7w
HRH6E3m2DgDPVs31nx1i9m/iDP0oMGN3L4JrXcOtTkygfeNaKfEIvPOg7EIJTfu8yKp5hrmZVeJ5
um6/lezm2xIZNbueQxUpB9Gc1eTMM25qTx2D5c83YaIjkBX+tJ0tqAabilPMu/nBB953MomXOXF4
QOGPGO+765osgFguaQ+Zo8FbB5Ps8e888PoL7rLeE/DhuN+hmfwHC0Ptz6mYrmesk0qz1MxkaenL
r84YMJdFtrXlqqJlufT3E85Dfk+iEI/4EceDbzixngpvSH/tPfMh8KYAyJ8cN7ujFaZYD8Tvq1D+
96UA9/LEAZfDlcvWTLYtYF/wT7nSC1MQ7HHxt36unru6Sxnybzg9cHVyeuQNdrSh7yh5CVKI9gEq
ga1m8n/vpRtF/uLgK43nlV78UToDuoMVXV3hKBQ248GgJdp/quAcx5yLcmhn/KpdUkjqWBN7BWmO
RI+DnT/16GD3KkGBmusqWK5yDOlbHdp+dU5JVOa7BjNQ+hkBrYLjk7d4vH7NNv/1fhf7y9vGtJHn
vzgy5n5VNQa1dncres2utUSvDgaTDJrqQl+GJsXwxguIjcY29eSieaVrTIkOVEKIB14S4I6ehsmt
Sk7G8//wVfX6ss5nyaQIWVMUVopg1ppLhR441lqTfAT7rpnB0Llrg3NoBXOVOp1h9eFAq1h7iKlZ
I3uDRhKBmNje4QprVnZzHGer7WW+wol6h/NpQGdZ3sobGPjb2w12U0vXVv17BLVQXklP6REOISFZ
11vw6Xapb8cvQeQvZ+awmnsIvsoXvrIpFEcRR4ovk0UkdqdrWYbuCKWl7p+4R2j99V0LlXS+T/Sl
KjkIYOoH6SLkmpsLg/c88dxe6aFspi0ykwMs/kpYKVedcQF6mSvzmEzXcfbztOsMH0QsWbsngjvU
qQPqQVMbjxvUtPmdOcGYV5cdfez/HcWe3O3hKfkRk5c0S1OVLHJralXcsabYlxDz36tg7G02LfS2
R4XZ+EOYP3Z8+z+R2dUCVsAvh2h59yhh8+8i7xuFCid4XiRCSvwtIvLqzzgPuy6OopRuCVOFYZzT
+GaYtcHk9LrS+6J7lxv8ylThdXfSQWKBxbyBFtvrSw2pT3QHW9tD9F3luYPMx+SpQ0syeNpkyKw0
Wn3Opeu0xjtdWnxuRuauN/AcIgB0k19hDlUnEwt+tHUTJ8P5+1RyAWngjE/EfR7ZqLvypTaeUUUY
3bRoNbhmMEVaQAP4lnpWq0hhYxsyNdsBpSnW2Pp4nVHHW5bz2W3z+wYINAZnuFzh+toqtqvY1PDd
pJmUBnQRxi83NnrF74RImYKSGrwsTofXuZl9xyMZyJ5Jw/+R6mly8KNymChA8hkROLngDfYTmKEU
j6jmVcTEfHZtSFT9Z53+Fe3qSDAK/X+Qx2UR+jQBPnCrUBcDz5UrU7t6fczY1GvqExYfrJztxUv0
imzXie1XE5V/2deRG8o7S0Y4GNoqn8R+CxDlY3Rh6CtThuumwkZlBOlQeQ3osF50etjT1pFd4S59
q16NfNjB0viyrUokjIdNoJrreJh5svV4N70lTu6jKJB/SHf+lZKr72vBherbResl4Y552k8hKFQU
f0Puxz1OwGsv7E81E2mRqNfK9iSILLIHpqlrrkQ4KUss0ZBtu3KpPuZwPcEo2/ftNYRlKvRCe77Q
sWlEFbTEx9Zyrztw1nAPuXu2+qlA5+9LYIyqtlvgtPuATyWmQhC5Z3x7+qDAg63YWcWATJUKBj7+
ZNMKmxgk9JmG6EUdPSlxfItKHn/j0LX6pi8FeQwWHlXkXcEHGCYaHvHnIUVPvaPWAlJs8dk6/SHq
Cx4AH7arPxfZ867JmvCMVVpcCpwn0zRJaofIvSbuYUynlG5csg9iUUik/GiyoatPgIcTEzVmB/ou
SNotWGKh8TH3qKDmrBW7eeF2yyfYv9F1M4cUjC21Dhk/BQDifgKw47wD79GCxNa+dQmDzkQhj6ZU
8+YkZccO6kl+N2i8teM4P4Gc88zPRgxIkApvI2x8m/Z9b5FaRZVJCWajGb+Ssj+9DNUdPZCZWKiP
kl36gX69bkxK/lnsfsiD4oK+1GoSRuGpyMxAuPY3/GD2cruWO0NX6YNDSd5DnA+hoayKXcnBrZMX
MAeIMifQPdcg2D/DPXLk59gIJqneHW2xmuVqA/Ey6phU4kyGbqp6WlCBmdQTNdHzIOUXuvUEMcr5
5/qaRhWDWZ+Tv3UYphDfb2Z+BNpU49k+FhN5VsJiUJ5h/ng3UYHj3qIqRKE5DbgZUlWlDFW46MTo
URoE7733cgzdTN1UyTpS3TZrWrtdkitm2B5r7NBJZMq9w0c3g98lkKvG5TEgSNCXvgpcIiZnq/H3
xOih2KjDnsh/KZkyj3+qwQofmD5U4mU2dAovEoPwwBM3hqoNB0eZ8eJUFeBznTCLq8/FeZ9yZHZC
ysk9DGCuiEqP6XdHQs47HtW80rYg0ygC1c6X9H9uwwWOmbYMOCdO1eZvl4ffpSuznfX9V+4Nf5Gr
W3qxUCE7QOCEIef1OXxMJBVUK0RSCt2GaVuL+jFI7HIL28xHYB6ZM3OBECaLgQCxzUVyzU4r7vQ8
18SqedA40ZvdQjxcUX7riwnBp3CF7RHjFP+iCpje2uJQysfmXNrsIlZqsMTXPC7vc851uGWHTdMv
R7rpAAr8Z0WLqR9iti/XqEFMT49Eg4UOy9G8y6l6dsIZh9ODQQGQDsn/T+K27U5m+iKoKz8TXJgr
H+E51PuEa4nR2VinWPd/Dg+c8+fuP6a1zfWUksMQGicJoFJlYbMALqAhNhJwm2ig0zimK249vcn2
3T7BZmxIA1nsZ6s4eGcaXlAA8HFoZS2KzL44WRxx4C2g3PgzCWxUJVqBYkh8R7ll2xswz8yGddzr
65HaFn+LxY6ffJpR+Lt/2lWa2DOy1Vs/ZooCwTAb8U3ZRTsymcu5Xph9bI4I1aRNNVVq5tV4gJfn
u4UaVxNKyg5aai5gFqrgzMClMaKSjAtk4VR2AB1DzC2pcZQziNxXHLeJwwlb2lfiE+B12frBqI5g
UMBA4buMwW7A5gcn3xaiCIbFd0JEPaedN9WdMZAnN7i0OPyjtyYSosuQWEmwOZUBgF8AS9OxLC10
cFygMtrnelITcmxLmAD5iqbhunBrZAc64pd54dSDOZtBoXTFyDhTK0sqC3U2D9x8CA15PFqdv9Qv
UVDXBdujfYTCY773xob7/BkUbzt5+fW6ZsvKlfuNLNSiSzYSnCV3QKo7kbX9NpFB8LYd9DsWs3rW
baoBiLo+EnAoNVQZa0xbFf/AnFkiZ+SXkZGlbEgGXz/2NazbZbFlKQ9ILteC61MLnUIMlraXaGFU
kSsP2xloUsH0wMJQ4F9QQjyMTkfp9QO4SZsYkVu3CTXw+XfjyfHjKDSpZcdLe0sbiJ4uMPViTKGX
lRXf3OhrxJ7UhNOfvXVbGWt/PAi6qkuxsGU4yBeukg8wAlhEKeHKN8ZHqnz8KWZhtPrjsD3R311A
aNjeou8eiP/j1LQD0hi3V4fneXL6iPsCAiDUep85eYePCnspfr4jj0ZB1J76bggL6NnENHuQ8l2S
yEPEmZbHsMxrGMPsnveGoSbzEjMs9+CtRsy0ndJI3k2RTSlCwp8uT+Lv7L+4mD01mIF9VDNjNW0c
fiyG2laANwnsRzvgi9DA8gzazGR8VKsEhEruLiL9CeiqpOUuui/npTAIPBNOGD8r/oRPKNLZwhLh
nM4/h8WGbNffvjq8m6ge4zZVmF0SXjqQrqGCkKkCUB4Bxq3eD5f4ANYoNoPex4C1Lwjp0qX9GcHi
T3V8jV9bclwd69DQYt8KHthNZFi6RJwGzRo5aC05IZHb9jwShRLjW3Xmc369f6GoGeEn2PxJPDtJ
xq3pwPLeKd8TdJ0WECbYXEUaYVI/uA8mb+mO7ckOE5xP642fA9Ouj8Z61V8+jhCcNDotLodwznCn
hiMX8PfOaFyB9WVfX/V0xyB7uUfOAn/mgGXwREdXCePTg5iOj7DBjQPogYSKg1GTmdFYaubqcSC/
axOCiXQ4y99DTuR6atD3JyRuzfcKyWozMi+ywO5ztkUccmjbaKVtSLDOqo6nlJsAEeNLW4bLaxKI
f1iXAPIirXPkuNj8AMLRJx9N3E0wK4B87jNv+wVpuf+Q938W2GpZCNVmk6SKYzSYdjfOfeRxkaaG
G+42AWoBDek8yuDgBqP+Rd455x105kmbBxOsTGVlgSORP415vQ+SgQRGAPG5FhfGZU+D/7tZShLc
esrfN4IM8txMdKUAfG9IN0eOeLl5vB3AnewaUSRrls9IrkaeGqRfW/FaJQFfPKADFibvkFGTjMzB
zHpokWqYxDLpm8r+zyWYLdf0ptlrzLbxeR4EtoHoIWDKj+Hz8FCr4SXFdtMsnT0rpOhFo9uqIFwN
JRdjSsamhcpzG92h4zBmX0iY/ckVrG1/jOUkZtkyVabtKgbizWyOf8UO9IWfs0S0fN1EHvTz5wxk
dX57Yy3PqpBeDikojmG9IRFO/axMPKbKeD9am9bHRWQ6L1Tm5cWfg5Fc1f5FPRCNLzMLTg7uE6Or
f3P78wVVXomEo2jUlmj8B0OPjZWdY2Bi5FRG3+ALDoVR4XgXidgZpnNzkQL+4XV0ZQN4+1xJVcs+
qfophb29nRYGX1rWlioyUHa9SCCufJ8OfD3R/vNodRm8U0m8o0oeOsdjN8Ndw0zOC4gy24gxRg1E
6ER3KS/52RlqndKBuVJC+5jxGyALU0IWY3ahZw/za+wI+ZXlEGxMVojqbv2kDLTwbEQxL3rqPqcV
k8Zsu6pXb/XqleGshGcBYEUY8kwJPPWKGGFAUKpGIy/WIm8vtDHTB5ARrZ/yT4fbV9qsST4v+w6T
CuPkCJJ3Jx6ftuKhKI40D5nNe2tbXDEEbq7tClbZMmzpK0mYK6cdhX/ZKtTDUZ66x6WCzUiuJ3Z9
wTB60AD39NXktFpy3MI7xl84G4dmm7pvmuNyag3qN27OQQR9yt4c3b0t5J2iDlS9MWzf/PBlopli
xlIQ0AxuTw2mtKwcDX9U9NFbt9H4oa103cWbUi1tHSxrNmWW7IrW8DnIk24pDZ7LXV6C2CXmEOec
NIxmXHftLylq8edxHDYcutZUwV6eJxvGkkReDyz2yiGPkdhg2dxarBWMFBKuuV92jk8JHA5tdURW
ExYAzzvx0AFCg+CxAlNzIe1nH2mJYcSBdFJ4Q4ON7GfZOl8QtqQo/CAz8hh4rojHuubG4HiEclzM
YoXMLMn7Lk1Vq52d20AJGkqWLP9a677fOX1jliYnD6kiBUw5yvkvVdmDqkpr1+UAMPxgLpSuxh5A
TkvpKoxz/FPap7xIieojr/HAPs5Mnt44qCcJKuJXpJS72v0x71HG8cD4LNLR44Psr+yTw2KdyX8W
+Uax2H2rQz/cRsLUYjZ5oQ7ibIQ276cEzlOqXBXpNpbdA5OiOKNi3tBlFHD7VxJ7bFfugBCjRyhL
MYqaRsijRr6IueM4kb4XepEg9UBI83a3PDeiUNgUyCVtAEPE9QmE2nj04HblSL0uVgLOSb2wghfZ
T/ScnK/GZy5U6VFmkLS1jj0HSjam20A/+Ldqg1dUQl/TQPZ7bZN23q9U5Z8/YVwbZbpIMNrUtQXC
5GXTxcgBsOc0/E9g9YOqlpWRrT7yVzBrDWycaDDAqM6KnXEHJ6t4m2+cZ7VnczVgenvgWMIiYF0l
jpJrpL7uV/8raWudyg/BglkgOJ5ZEHEiAQvR31K4dEeNduR3fdkqtclOeKqfD9ow1l3HRu/fawYU
O4vJHPljpnAZZpmSTJ9GRzbBcSe7+5Y3Lgh3xVX8Tewnh6rjIH12zHTaPY0XZsyFnPeSdqFBMasR
4zN+P4AHIiB9QdZVuEgChU+F8XtHAcCyLzjvRViKdPMtQgInXnN1KzVbf96q4VHTv62VrYeIIt7U
XhnW/Be76zn3EJlPNVfzm202pOirGhNmeaad1Dp8XhJonflw/BbaFaScoI+Jo6/167I6qzAmo5dd
8U7rOcPLgR3KrAM3RB7mjJBCbNFHKyv5bgdi0styymoMv8jTkj5M3g1zzKGsCluTBichGA62xoyb
JL9d0iZOFmqVMoGBqc5+oZmc40/xrmpXTAJ/35tDTyNDsgEuokPoZia6QtOVoTLuOlUXQWq2r1HM
zk1jrtQBolr5EXqhy0DfDcGCgBVzLnuICVFN5uAbuHlZTXv0HvboR7LSAN1zXpBxJwjsvFQVOE1q
OdJ06Sqx3dT8lj2H43vQS2dy3SIocRMpOvfDtmoXRIemIuvwIf9c+6bH4ZXU6B2wZF5x9w7anmXE
mVsgJ9eDOmuko2OSCaOiPdYq7+gxZ7SDI2dRZYj6frQ+IUdaPAL7cTk7ZZl4FfqTZ6O251YQI3UP
g0+YU+qDtVPsUq09Z74MpAnZOwO5ZHt5/sO1hxw/cYJAakOQjNOuU0XDIvlB3iGI2g8G9j4/H2eP
7cOXZKkCW9+arapl/+ESE2FEhJqnQY7ftMufqvzaqUnKTqkKbwgKp7eoFC2HRgtvsqpHWaEbSaCj
xdWlbVtvpQVqg8tOpsRxDpUnR4225DgZ/39iHKNDQBF2ww6ixsNbA9oqdRQ7B8BQGU1nacZSVUQi
thW6ywBLmRtMPtDF8YsVS/x8Ps3a7mtVb0LtslqeNCgBGrmNnIKrwzD5j5aL//m3wWGBRdv6geL8
CsYrVdReWyx3BUB6SEuwmEbniAnznaWCAI+mdWlXaBjFEDLyBx0AV9W7ZFTruxZYoi0QoU/YiLZC
ReGZg3gvsetLqNGEh66RsNfaKctyf413AlfsRrO1R9LSLlxSbXb48YS+Cqf2+aMVFLOMU3l3DBSZ
+ydsQmfkNUdhhGWaPLhygAsGATfBGQ98jCJNYh9/pmFwUVgaDVMYHUbDTeodoM1w7EjPqXKQHnln
ZDpGiGxkyAtgbaEuryD2AMaZPacikjPXBHJ4iTDDKYqi/Y6Iux3Mlgxug96BNF/oOSmC5mxZkbSi
4LfF+NPJkh7DM+hQ5JR5d7bCIafJPaelvz3zd8lCkdOC4lONyYOWQZ2Q+BQgJNv7u8Z4r9SHFqs+
n0GmbE3aTrdYrgC8+0fodFvE/araL8/XiW9as9Ng+Bs3O05KR2wcaY5yYHDzfBX5lor1UX4BEEpU
9B6ndFAJ8UmuJg3OBuEzQMppf5ZhACmv4ljh4Z62Fzf440SJ071y2RYLz4rSafxXX589a+YZg9Dc
Pt/iNr27QHUtrOL15z0J8GFzfsaf0YROg2dPpCQ7f6b//lpakbChY1Q8h07hHVGtZ+jVwpoSId7B
0dQcIqEb6lT2x2AGrIDy1cPy1Me53Zmxc+xIJUD/u94C4YavUbEltcg8S8aCfHOsi6dQhjmEeGPv
WbZyNER95xKDjbgh+AH4TCf/ABXBwtugnWFVmcFV/ExDxPfO07KidlfbvAqPUiCkfhiw8nJJ/iLb
Pw4I9wsn9KvAltMfASqjhXnsMY3EGcYWZp4INsUUpo3kSLsSEWvmLrdrZlJdi4oJJ0k1d96tYhRK
pTppsIz0frZC0vKnMcdjQHefq+N7g4Ej5MqiSXnwuJLa7IyIEfQzu2OCXM44uRXmGoup2eahR79i
W66gLL6mPpcV3SsUiJ3PW0Kls4fpVkTVsqWyZaP01s28qAMJj1eiw7CsVJ6NGuGC/CsRk8dL12Bi
mW0n5cviMC0IH/N8goqnfPo524iuEMI6mv3A/OA72F2+NTWBbOB83AG9Wm2+8ViyJzn85IPMkXLB
CSgTcuFfa61FtEOisr43dQQDTCa5LzdA6fSQb5HBIJJQ+njYYyEd0BW01qKJ4O2/powy9bGSkmxD
0JgEQ80l45e0Y+Zs3pIaYVsopRtYrc5OG+sq01LZEItP7Ebm8fXeTgD40Zd7C8ETLUScKGTVbdGO
yPJ+n32qi8kNAigkpxkdmWhaMXqLBci8pWZaWtnR7A6wi6aqLnWsS4mWS5T/rjRCHV3tKYzQY2be
xU/iS6GJGBzYYSSM/0GZm4qNz2Pw5mn5IGkqq6kv8UF23UoyXf/Q6GsGjUHTTnrv3DKeP87omIOj
3fi+wmaRO/Zm2rgk6nj4TiWfX3TDajAxFzl5SpmwqiqzTugnCnb2eBTP8sytxQOYfsUxDAboT0UQ
h1uBzd88QDdNaovelY3z9zJ09rjg7EmgBZGRlBDYJ0yUQm6R7koOzMEdezozkjlgF77U43AQ8VDV
BDJEGmCLIavVM9/sfteY3mBuAfEoDpuxQI8woPOjW+XLZrKhhs+yaw0bxLx6XMLOy2zx0eWKolzJ
tPOSNcwRelmy7LPOi6+6xHFJawCQV3NY7OSzqsmLzTOzc6GptGCS8/ltBBfWi8GkY7js/Ip8BDDL
t3kSH2cXpSuz/xhS2NaUyLMzeme4aM8IaYI1DONahM4qjcwyQtoU0YAS0C2pWfoP/dFUmQqCgZr8
RTiTzVrLTP3NODAIFnU+v1dLI+4FQLU0yZPIu16rr5RkzgrRrwjRelrXPV3FQj+300hPqIWZWL3Z
oMQUwVKhzrfMyO3G+uxuKvPxgDfHErFbw0VDQ1nJ4PLOOQuFs4d8idScosmbCdb7Vzvzlb0OW9GZ
hQhv3ta5RVs6bbsrC1nyNwyzwnCCnMMfo/2S6qbGrwdMI5/USgDhzv7daSLMKfI5BmPBXg5oECIz
b0mLJ4qJd8oi+FhPWZ9V3WpvyW57EDVpOX0XF7IWp9tnYYhBFGmrY4KiAVC7r0VZuKXxVkEO4dZE
8+VQbqmuVEF2l9m0gV/Gw8zgTSjrTH4F2x1Oy00wMBBJ2/eoLSY868veCbz3s27rKHmaRPDfR+qP
qvLk57fSE3LrJ8ftSo5Iq3IHWs3f/oYWLDIOpFuwTFgbof7m7SkgqgqQHXZEaD4uJOS2g4JuWbBB
wDPC8aLLKR1o8IyWlzwxCLKuf/s4cco9vc+PVbIob4BG7jPutSGEYN8egm7NYWduD6fX+LlgePP4
coIuHGLwiJXSGyczIfOKZRwwXlGBnKtF0CKCpcq+a555kGm0rDKmHT13rrq++Gi+skxIAV4QUFaY
yBXvYixpBrVcdX0YyJm544Ik2XMbKAyetAXvQ5KSN4q8KmTlePqxUVQz9PnnYcODaexkyQFIJf8s
sfaXJdFZH2a2yMUr3vFh4GdVPegk6esOyKy4MUQHqanZhenUyrpN7urpS7G1s/Rm9pb/3OfnXQnL
7r+dttJ6vkCCnn5wywXk/bLffFcbr5ZJK/adVvm0nVDGBGFJz6t+/iF51Zxm5IIxlko3wF3Z9SCs
xqDL8jfLQBTn6Rcjt3NbkywyHe+eHvGdMSahuG5g04x7HxlKQTAxMOjshNVI3m9zGn/ObsrligAq
SNswsJwcsz5go2QrF7C10rawGoOmFU35JpMn/tNIXthmS4U6Kaj1OAMtMa7wEQR7qHzy5TCm8UJu
m41bfgicnsKpmnABzKKBuwNYyZFKr+fYOUrfCrlFViRDhg6ziD3LFXTQ4IV6lgTww2wulc1gmiwL
/f8oeuZ1Rt2JmgWZqmosZbWNhOQRh1MlgqXIYRY1X9Qi8JPe0Niqf/TsQd7ydF4sx79CQyv2OYAG
U8OxXrcwJjR0Pa2eC5olvsCll1fXFGekySQSNFKAnwmaO7DcG+67viEywl/+vPGBijqysSEirIC7
TQy9JbF2FBWGe3b+jtcF2PPnhq58+gF1FgZ3UTOtoYDiZlU66m68OWeyAaihbBfqqffg+KtLOzBF
hSnIK4mDmnPbfGgWPstVa/l8rQcy6B3mKO63VlkUftMgXgkkhocCbc25n8+H7s4CTRV1LH8tbRXq
TimfvxvAovvA5eSXYKzYcUlyDKah3Wup9wGM8OekbmZpxhzi71DsjKWygvBa781XJdBr19JFuVfh
GqTk4eIRflXhw5/MR7tUxJuTvqwGmSobdNALcKfii+MP1ER+B01himUfV8irBTlVFztAncN7m82T
Ibn741x0yi7HF7gugn3o11GuzkZ2Ix5XXAkV25qedV3SKSqnoGFoDghnjzofaYt3TFuJ6nGqF1Eo
qxLwZqH+aTFdpRbRHz7rU6iEWb3QQQP3D/P0T8wkwKhwcc1j2dD3i0B/O/QjazsFfb+oI6GaeSfL
i2XUzXoDkOlGXBZWLnp9Jfid6TvxVUoFN49hF2tMthwVd5d3TIhEMiibLbb8nixNRoxFdL7lzE0a
U4meX34BewpA7ndqDgR3D43vCsxaF1/gpdeCDOScAPsiBRd9jDECYAGIYEuTBs9IFUFCDUYRscdd
qEJNSwyMDVkN4hKHe8AF69O1EghF+cW0QaxLBck5IqSO36HTOZyBHAqlEWu44WnuW46CRltcOzT/
PxNX8QjggOG5JlsCyrDrpEN7LEmLoYG0ONK4gxPluZJ+/i3TlOLb4YpE7sqXwbMJNa+EuALyEiW1
giTKbwSygSJ1Rauup5tEjSCV5g/xthmjvdas8ptp2qgMrJSlU/c/7Vx33DqGSKk03RTw1eo3yJWB
aj8nT0e6qpXC8hyrXB6oJsyvlqR8tzkiwIWd9WbFUaoPByS0jwlzYLfSGTMd3/+2GevjlSdT7DZe
ElwhgdJ2WCdv9n7brs2wb74ltRoDHOKX58zh6RyevJ0XmUmCmqSpcSdf4MX3PkWxMelJwpEDKb64
8mU6CFrRTQZn+8hNZr8kZc8Yj0nZf/iyUSwQLDy3G5jMdkI5o3QLwYONOzl+W82id2gU8hLdqeXH
bI0hoejl7UUNTbtTgWPVdLDgVaUQLCiniWtGWJbOdj6GkBjToRUICyXU6BwoOpb5eaFH8AmYOfvP
KFIvKsl28zaQY891QSg06JyrErIj2yhOUTVdxid+n1yZQQg0mpzOg8jBqHCJ5won8HQ7QzjvAXDo
tUPYij+lu74Qrc8kcLjvGOcgmq7PMqRgTfc5hE4RixLMs9Oeu1fieieZtzQvA5C6vy1OHdb+awIW
Mw+Q0lO08fKkzKZVdGSna+j3/UTyiSGqWbanESa8Ipx0pIwm2xArnrK9i8qygIw2GZr7hR6n36+W
cxBUse3NyX8Yhq9attUJHrQbb8azxvGfcYJUGr7imKaTy4lEqf/tzamhU0ioRtnfqkk/O0/bKI6O
mbkSE8Dgdkt5GlvtihJcQaNOkILXvuRDD9J75VchgGce46ZBLhL8GUxiNesIKbruuHOmr5LorpBP
So4imeaKG1Fe1rfhFOwOaLS8yf/DuXVSurOZBozJR+mOwFwQU4uvgtShFD6WKHskvKGdAxFT9AwP
fCGmWTUQasxWu5mdALEPyzTFnzrqs9OHZQtht3qfl3Aiv/yo6AQJ4BIkfPoOH7fYTHKokvlTSbSf
cQQ/RlkTQ6k4/YHQDR1JZYIUvdN8DTKRkwYa+uuiP0yG94Uh3u+pF8Q3Qgen8SspK7tJ+LiiXRvY
erKtLlyWfDJ5fja5pXcIBckam+d7chnlmrdXcUDQoaAh+7eEzVu/JoGZdBwv4QlgWD9rYMLf2bkW
mQVts4KQw/iae6YDrhn86c41w4nyGRCbcYI2csbD1xaJenixwQ5hRSm0Lg/4jFCEssFrfWhLWrNj
ulSdLy7FBhdxeWzYhQ2qx9PQeRL32h85Ez9OHfTuUbf1eaOLnjHR1/Ni+sCiW2s8PKbHbd6D1xYq
+poESK4n9cknXOKayImsrQIdnvrC5wvKEz6zu2w6n48Jl7zZF7+6N6tjeUwBVH3e0GY8Rzc6rEIJ
ASwCrbQxktBUHO80gHTRANs+IqoXUup3y6ltnDA3qxYGkKzxBTXe+X7u9LnV+IdtR3hq5HBk4bTk
byuF1YW9wLOoeX9kHYzh37Awx/SSeW4FCrjoowexnqvAPEcngVH2VImdSyWuTAJUF4zS24n94QeP
csiJdDl2HA0EA57g51EjoRNpNVvbt6ZZ0G2QjsNa1wWMsVPgHsYntbPs98uk6mC2N4j8b8/chzmI
tAELX7i5m1bC9H+hit5MCqANpyPjz22cx2y0/9kzDU45X7UzmU1hPq20eUlZSRLOtgJ/SlMr3xI1
i3SC79W4TVqgRB5GcMlGqq/n+67Dijn6W/33oujSkHEkBGm9il5FUWXwnFRPCvbU3S6LuB648Ljl
ptsuwVGkGsbrAwt4iw6IHIY8jfO5GlbogVtJ3CssGE4MejIlw9HEab/BnAupycLtgZdLUU8LK094
bhVYFN+nkroh1hi7yPtSF68HdI+SYjhP0K87itWXp7kXdbDNAgysl9nZpFeb4WXi3e+iDP4uju9P
4GHSFI78LT8RZPCPa0QC45TE6fXWkatNpnikqXOQ8lhwYZyxB8n5SanAM6uu/QkYX1DKMTD0AaVN
DlSIRonZ6egEyrcNCNiPl2E6Qr1y5UxhhEZNhpFg+d1ZiViwjh7e87qWq8LVhaMIVveAJ+w3PI5n
U0YYPLKNARui422VwIj6zaq+JkwWm6riQnYJEzMNAVEbkgRINpzYSszcz/3eB+IlqM4W4nzu2+2u
rr6L/OO9Mw7UIk85r34E5HpP27lg1K8mFE5vZFP4fP3S6561Xvr51XCCZG3COV6H33XCI3lmmWXd
7/opvo/eaJ4omuSZ7uPJRsujQ5qb5jhRC0UmpZlyK+9Ay9ax+fI0z7QlZAWXRMzvJWCXy0hRFZqC
2c9TRIt+W+plXFlrM615KfWRRKGKYPJV5qC9qydZNgBDIC4S1MVL+sc1TyuyHc0EnvAXf8tq+MOn
OKadF1asX68YwPF1UtStW81SWZ6rLmZKmAeL6xVERZ2pQuriGq+AXF72Tc+KZEvW/72l+c4OfbLK
/FXiFzhs2iez1SUQUIXPYrZUB1c3jInSh1T0XgRTC+DQuXLdlHH5Pn2V0JkvA2Qt9fur7CrnoNt/
k2Y+7e9VEY9eoyQBHK8XKNiiC+cr8Ve/o0hyCYWcWB/W5eH6oroh8SLnrrNJmIO70TN9RcvKMjq1
MJwd0xY/96ntU5n7rR6rC+6SYq65UgY5OYxoKpk24Qh90U9Xb+EtSM0n698+Gx2odJyHiKqt8z5T
KOblfmN5rAiqDlXIa78h4sP3pNQDaxSaykaaxRkC7k/unyux98PW0NQs04CdOJ6NxvKg1QOG+wqO
1fgGfwaPx1uowx2BKaXLxyXT0+oO1aME6q8PwWbsNfDyQ2c2rul221LcoRwAxxU9O4hregD27+qM
56CYsCnV+YNa8TRdr/VGF2XjJ45WWV28pqMdFt7FQCf48iFKvisq0G6SwAIjzZKYtMGZ/Jl1ucDx
LZrIl2IldIohufLBOOPUf9ea9izYtOpqJIn1A8QllOFm25TNhdjgMiVa2wSFtcCrV9y2KTUBFs+f
7v+T8iX5J5+fJvptaw62vAcMyLdTFjcvDrCts59WjquWEgGpkoT2e9us4E7pjYNOfQVltmVIuhIt
snJ9GwxMQ7JiV56azozyO1PXqlV5KE5mU0kg1hCX6uroKwwBM8cglj5P47wiYtdlpjYJdjD2m/SB
UpCGURl7kcx+nqrLIjKwV9XZSQ9zABGJ8Uq3IivhkcZO8+pytgpJ2RNgchJV9TWNoXQQy3BdvEV7
N0lc5Wnnsnn7Gco93zoiHDYUcON2FJnXVgYx0ujT/MEh3OJXnFxd2sZVF1/cs/fYUrZQszfGP5ta
sz5j6mc45yMR2psufL38P9yDdIMo+GvmdxPXh9mrvUVAxjkMsGAVYFieLAxX7I7AWKBdZ+nVMadu
IP013HoYDp1WCWssLp9EAPbnnTiW1d8jQHe6Heu9yV4x9B21YmGt4zeTrqIfsOu+UDrSlrzbK7iQ
LFcXFLA23NE/47FGEdc0t5swmxMtT1fUfFcMmc5MqALVU/NMMBdrnDOKDoP7SmmWu7mLpBHXqcG9
LGkUQd0pgPUhCc6hM9oEiC+hUlUyJQNemWx3yO7Puxogx8DTz7Oq9cagQHGCKkDlVvtD9NAB5TjX
nszkOnujWVInZaAghaULLtTvKW61ngFWLWwidLalTWT36t6VCb9rOQhzbh4aNc7qDx1rPtQv0wEo
lC+qzWDnJD41dJ01yUU1/Qv4W3PLJyuhMAzK09ySPD1hz4YFWbyem7GECDgFIgNZajV14yts0it1
Pg4iW1E3pV+yEBZyuO+nRmmxhF592MgPJ1r0YjBhQYkdNHa6LnViD5IE6UrWK0sEtQNp/ZQPddRh
4b5SfPx+jPpzUPaL0KJ3PmPE5RNMMXlYoiCkFRk2jiXCLN+ADoVn2UZxlG1Fmw+OWaRO6Y9lPhw9
6gig/4SDeORD5duGKNUtyCS1SqwHEExry8gyopDGQB641AwExdBrnkU4WhUWXwCXV+v45+Ogo4YK
NGqpBcpM67TkpgHDKQUKVJb0fVxSJEQk4Zu3nEMrOt/gw9xZzQE7zIQjXj/IL8MhQAtqa0AuzYaj
zTA8r/I6gKFO6qQw+9dORpReCi/KobXz0/LDtuSkuPC8cAl4A5ByhSkwqZBcUjW9LywaYT7KTM3S
s6odoaGSgrZWVDDetTSbae6ojL1lpr0R4Jp2xFHYcPA8/TH+RzDjSdj996xMKyuhkgdUdXe/XH3u
oLUk6IBIxBi4sO77CSXjtNRpiVJGwr9ik17b5fM3F2Vb07F4sMMmXm5lO5esWsD17xwP6g0YgNcq
8tS6pliQXexZhqQPb2UHYbzdfuvPXGd6dbKI9QLK555MSuiA3bbks8f8UJzJPBFSa+I4a9RIhINu
NUb7bHsUz6k1FIFx1xA8a1HeUdXKEAC5/iJj3vSJssaYQEVq/WifmZ0B05ABnIXFEChA7628fO7E
8229Bxsln+90K5jrR5DFRjhhY6HLYxcbJk6uVZ7rnkpHXgq60EuWfXgyZfsqpKOCaeR8mD4q8Xps
VFac4qaWo62RE0YCItuNnq26OBoIkL9uDxHvVvNkPLfraLBIMgGzCFJlIUz++ja1IO2/hu6HuTgz
SXThmetW3ztyewWOTqp3t+JhkwW5yF2hT7MSORwWKwOx7kIJomM6Q4g0jO+Kq/QKibriuY+jy5CJ
vwZzRzSMILkOmzCPdihrZKvw4FnqpPuI02y7GaHbUbxMUXUeSprozD11CIdmgDyov45RpmFJWcx8
y91vhzNb2SYOzI2IT64DneIpbFLdGpXqv2yzSgQB2aTN7O7DwRTETpd8jpu1l3VUezB6UCio+615
eIG+3iaFcr9CuHefCoSWaeshRJ2Crj3K90m5/Jewic3rlu4go1JDY1nIuhtTtkvLMK/1ApGS8Ltn
Rdq+I/JFeDs6druzyzVGnx6uA1lXvAJ61vc9JZ//t+7Bp/hOzQbFlcMPM9fOJle/tTo38VTxBaew
+QtneVb/8E3RoMd/3DVYkvsamtU+qjVr4vPSGgcCJ8aEPcp1oUxgOBxznR5Rs1wHnZ5xj940TteH
GNU9eKFuGdGSxA0JjOKkBOaOMPGI7a3NipceJY62HwF16SjP76nY32dJCDkXIGTELTkd8VVdeA+s
mNVhXKw3V8KMFqSaIBLukbRYj9wrA6EAjbVqLnFt2eX8HbbMCrE667FNXfMh+Zer8khipEIvizKn
E3sAn6w9uzfRYEUw7EmysuKF7XnH50CEpLtsLghcv2DmswXZ1AxBByfOzWHaXADkkRv+Zj1NRkv6
gkdIrfFJ1XJ3Ev6qqr6z2tDjLKP3ps8OwKXHnNg18EoI4nyC52sttnGS+5YWQCT9IznuLSkeCFtt
YYyvIm1qorG/ymcigD49XNBU8LEALjXJW6imkovr54YyuM8KjqLPowjSfxeA8EWrOKxwvxVS4BCF
ex9FV9JcJxymAjaQVwIqZlmSfaS+P6sGQeDQMfmDvwBeQGpPiFHaBnAjwjrQq4BeDjKNzGfOHmq1
nIv6ZfxXLEWCRNfpcF+8EMyv9Y/sjl6MAmAYwO2/R7PAPanCRzTWyStLlACziP67KCWxAU8ZBLu5
d4MMQA1MX96YevdB5nHJ7Urm5Z/p/tl4d+tf5bGUsRkobjWDYXAuTMmRMfiO76R3rDQUMJvj52Zx
D0Ta166F+VBtAOnUMzxTLLfbkwl9sl67OELFgDCuszHSKTtTt+IrXmB+MLw6pWdO9jBZ9ErtwFi3
2E96BUzTnJcEGRSEmbn9d271vHVPjdrCaA1eKxc8p2ybmpLO+4GQ0RJJ20OmyOZHXn90xH9DifUJ
F43tM+wpreTdPbWi7Ud88CYWGIL8RCZNGJQvjDCfJ8qfHMK6nqQTK+Ee+vRz4JGgbzJ/KEIIb+tS
9DAk5QVTeMc8jqtbGkCM+y1jcGPtWUZkpqgDbzzOrMGDZYMxN5yTTurXra2Ri9ThY1zsonGZYKF+
kf478+rvxqIJ83FcEwecle3LdVioD/0czS4HIHYW/VMtmTBs6DTMniU6pHcFIwfocQw5BwRheQKN
jcV5yPy1936b5wlx93U8XkGKOVG6uN/15SKbwNJ5dGhE0yJrgS4k7JLT1EZBlhObjbXtLkPFWyTR
ooTDtv/lRYBRO30jTm+IDwvwNYLQ6es4q/B8oQT6GKdRWw89fb6M4XMv3kvq1QrVIG+dqpZFlsXw
E+TfmjfmO1eHsd7/rvNthlDOfH67agWdup6q2rNXjeBhsFRb9163iZVcvzPitAKkj2Wf4tRVxHn0
f43D/Xd+1QbY+3RLNh2rD2ARlfhIFwk/Pmi7HBLo9zh9+MrGXKTAoazfQW/xMVJfoYOhlrLncWj9
jWNWyvsB5UHHR6NYLPa7i//Vy0+d7w7AAgDppRzDNPbsoVbwxtxZSp+bf3FQwTRTSzBXDiDgY9to
BXh5gtNkU7mhNZ94iw5Irv/n1lBr4iQodXtT/aGEyJp9qC2/Zm2PPucuYN8NhiNMeEKejdRx/Dro
wBtnSanWZ48fwRrXeONlto8POjjHG3cR0fCKqyCwcIvTRMC1b0wQkKonpkYWrur97TEMfUSQC3HM
EuC9EhXjOMbNEfNNKbyhYz7BzLL2GJJmQTZPVCAs8hc5oZC5WdyDkGieWglSYSFRUlpHwbW9n1aQ
utO+SfXKu7eQUASUQpQFrjBVChFiv8/ZrShFub6CFi+LV1s8hTBRQ7gI/zhvQeuGQDs4fOe0QWZO
pz7YT+eJUGwcFR90R75pYcgKDSDNW0n35DPGbslmbEv9k0bgImSTft9EhaEsWb7Mh+Q7aUJ5vKHc
BA3UnBZ3WSFZp/pYUnQwbFZUlQPvUVdDspIpCMwSUYjzo1mIQy9kKeQCF/DCxc1tfuuQHl9DVNhA
wu9L55Ekq6ENLEx9WlkPuRu2qT9ib8/0hDteJxEv1/eAJFIbHv9aj5vNUynNlKehsP8ZBZKAP2gZ
gOB/zWQ267cIUC+19UZTkql5Rw2GnnaFz5Y/4Sr68KFgfWtstegUvTVMXxXTybKxWW1nfBPKcsep
RQgfg57sFxDf4xiR1UKWmPxMcwc4rTPdXJ0RZVS4JcT3TrYp5OYj6pQKMojJ8o6j0Z3DgRKNYlD5
j9ealApj29zVKMWgbkFxffnm+T6l1oWvEl5T0UJhxSl9q5SVCjoKvyPT6EYrT/kFtlKalWvOA15M
p/kj5+ye7cn6TvcW4+3sdMRdC4VPDcQxtBvx7ARx35Dk9/aRr1SA/2m+na3NHGW5O0ZwqfwBoe82
5GMgyDdTYme1f6RsmvxGfw59YPjmAMqjtYvY9VV/iuGmMyELbKYPz5ji763F0A1lh18f2s6epu94
eXOkW1wW5GdiRbLn13Fcq73aIX/jvSc0LkI+iUFQvZC1PGNUFD5I6WyKQypW38f12cG7rnYfe/lk
hmFclYNxq8xDk9PFFH/O2/8SBpV/ALso2Fa2AHtaEpWNe2KvSVxICPYR7fwwN56Q94/jY8qltiTO
R7gEPnd08Z697qOVMPmPK7LNS7g6/ylWWKI1bSpp49YP5xaoWqzfyOtjkHQwzZHSJofPeOai6ifs
N0gWTFD3nITgLkPIsqxZyQkW8G+cT9nKjjgggaD3NQfuW/yHlZo9f+LCJ3tY2LULzxfqGtvyMSCn
GX4YhAuRsvDwXV1mNc4IvFvdH4PBxCLo+hA66xhy5sr7KC3R5sqFmvkSCCHWFp/pdAwQKocSmVfU
A3RlgIMoWkHh7gW/uekSXY146QIsP9ZTz3zOgq433/ceVzx2GdAS7uVOtULuHm72qPYKhBb8Moi4
SJPaNG0rBQM+zlD8Y8yebBw+tiUCyMdopb+UK2XV/FECEU7moqpyukh5c0Tfvqw4GYw3IBlLL5Hk
Wwb2uwLH83eSY//9JEXSDBQBVMLDCBKWKbT52EXrxIFrMsMqAvu2ptz2YRvXOflLxFqe+VpRN0qk
DGio7r2TZncwbz3bZNa53rMe/U4ul6OiPH+qj73Y9CXha3NS3082CcKbLqTbxvIZw8BvZRrPf2d3
JY89Lnt3SAtDRWnuzj7mbDBpnqWIkVOMrWH9boaf7AOqoJa+Yh39HIHYk6gcs4Ke0ouJuYODPNof
yUeWzXONdI3+gK7kZUlbY5RRfgtJnwGzzRxHmvMVRohy7o1Md/ZXmlX2lfSroQAb6+k+iNPi3SoK
A2PMazji1/60vrWxsf9nTOV9+CmwpLBEmUI83XgOxRiBp+TifrKmwGhbp0Cot9rzWHE3JNjsPkVs
I8exEtQv1QWpHPCR+gHGSAUQbx4ctOqf+lWIhLieXCnAYYDlSQMG2xAMarjSrfkM5Ey1dCqJQHeg
R2x7ziKfsvtY/+OIOa40B9JJGqqsRMJfz2d4xHNuc2dYPKRJlFyKBOWVAN/P7v3pKiWAJhjjrlE1
sSusBa0Vm/u4Pq3WibPs6UdEEoN8r/49eU6VP5/L1GvjppMbeOpvdFrIfzfClhh6RfQd//wTZZGf
cW+VRLfwpaZyoNp/tyHW3RehWNLUC1CoscmraYD6Z5Fdx7u5Q+k4P6lGFeFcNvm3PZJ17dzAla+p
fv3UmtC9zMXAgnXuBLZupd1eMPjqTixV0hMkkwF8OF9PSN1kpVK2RPcjPYT26yFz+Zc0DwgDjYxh
4JYModz8p2behG9XYdW+uCD1q7ZxQfvfJU5JgzB5fhhMa1vS5ADMzyMJtJFLxmoLXkALD12bQIIp
Kf58MQU6pY6t2WnxIex62CiC9eE/svF9Za8QJh95onbwevG5Tl2UJ9abFjPo9yM7BN8+wpPJpqtE
yEFuX6ng3Wbbned4Tm8e6l+d+lI4WIjc26lxJxCcpZAq0yLICqPwI/eDZ6CfhK6QlTZVYJkPF2Uv
UjxyN/hEJpDDL8mLdsWxQ/R3VmgqeIqcGFeb8tSTFV5eqTqwNW1459SR+uTLBJdIWXgp/QhYxk5X
9yGKw+mZARbXjB7yWQGzbMBVBTU6m8J7W38Acia4q9FHDU3GW2E+CTpzp7gWXd0pMyhKGCEa+RHe
UVG2dk2B1KO55eoQAPdvaXgFowv1eKmlGZ/lZXS+Qdv1eUkLpxx3f6LIP9XOlPZeM4J/dvhvSQA2
ywDls9gmfzrhO7xEQK2R/ZqheM8+RFwpvVvqUdwQd/FH1Hniix/z3+bW+feOlGNdksZTipw6bhOY
1V/d+J3zZ41pHhTbou424dK5w3VRBoPuEnVtkKPG/1sFJ7y/nzbyBUT9oYfbviF86oczGGfCB/mq
5UebZMcUVQAzW5OZzzvPcijRucHDnSWZ3flVc9bBxhaU/nBmUqJg+T/X+co+6kmTLJzyNI8pGtdg
dueQu63MsNq7a43b9CrIxhyEqhqs+A0045EZC0LcprcCQFCxtz3JUNGJITMxHM96MGHo3/nq1UYe
N2ltpny/YEFuEogOG/oyaKUAzpmcfLaMqxTf50WclFTChvy79bZPqviMNWZcPXCxGNuHGtYDKIin
whpjYHaWEjo+zHzWYeI0iU6pENiSQ0Z5zqnFnS2gaszBZr8UVeh4keap2AcLz8jGictXq0QmBetU
KJEvIKyns9rS2f3vmZRrTEEc8CIdIbFlw0wiFpR7kdU71Ocivz8KSymRQvIdIvbCeexUd+H//W0O
CxBTvfvL/xfi+VVMtcx2258rplDUQU+B0+JLW4pS/4x0hXaV08kKRv9eUNSYFFpKhTY74BMKfbyc
yTAYAQvdcTuVaVOOYsFR0HDDB+ISYEekRhj1cYt6KmTh6jvMhS5smAIjNR2iVH8WhiQuTanm8ddt
Hxogb2eO8t1PIh3q0n+v14BnmIsvVpzoZtjCSp/hZFb+CFX7ucbi0lFA5eILOPlqMrlD61ZZjeCR
PnxYB2exx989afS2qSmr1DB/inoh58fDUBHtQ3pg94MoEtMeaNu58EX238nLNMmuf+NWj+O+v9W5
AuXF2zmleB7SVko7y/jHsoS96KParHiaQPt6Dq462n1uH71ZwimIPM723LNItM2Eg+kjCGIADE1G
6x7RQcRINQGhKvr38qNxYZNVZZArHTER0oc9+dk3B3X35KfE8Y9/b703NlSWgHliR651wlJ5K4LE
qsDbtAPtfuZ8hvza5f7VC+UAuAYxHvmDTw8yd5/2cWTkI77aqvZ6M0Gg0QtMcW4i7KFk0lQjRpy6
XT0k/wd7ja1HZujhluTireubY0e9YACfAZQ9Th4b7hjItk+Joza5+ox+tQJ9CdBXJSuDOHckBBju
8VqPnDD4T0imUaeJlxyq88O+7f+c/rLsdEVAXo7lzi6qvDvUJ/jbEzZRKbDs6DOmOrplROkHTRa4
X+qSA49Ozr/ULD8Xlo7SNF/+PJloXB1VGJ6ENY/rFw/sylD7fDkoc+J85etYj8PBGmbLIjHJUKks
Y+DbN0M9dkXt/OSAjjh7gZf77Tt7yu8IwWN1lWM6Mf1MUOVr9TbxZ4t48mTsstLja93VzeERjku6
rVbY0d38i3U40602olp/PcQS3EHru3JAz4BrqjqXz4eeLuNJAkhJOcZOo0GWYCIsy+SUVGRBcDXr
x9DvVIICBXPU31a8TvTkgQd90BQ9KsSYmMSXH9PHOapRL/iwZasj3VSPUXgNEJ5oIEHBcTHTnM7j
GWOp0CkjQh9bur7QcxDLlZwM2oxHTuwvch+7385wZcMflW9Oq30aa/9l86epsE88UGRDiGfyklTP
81DkhyTZ1Pf6kK5eylh5JK/bEHUwtoLuiKHUGfrlsaEc64XmKFakbJcbRx9MqcA0zfJn46kRausL
JoMdbXO4GjEsBcOMZ8pIqzNfNMv611KztwI4NmAkEZLu7cNStsol7O4biJI0QMeGSwVFmDvBfhfG
iwMdg1Nrfd8ojond1NIT4LHWqDdQolRcJQM6+VWgyokD0ZEpe17Geg5w1jCcgWkWLyry0OTLAlL2
Dh+25/iS6DQfTs4i87M26YaWd5BNFGWXGdqQZsV3ov0pID2yRa7mEeDfZFj8Af7fovM1+cRfQmRo
T5eQ2HVjBekZqrSUy7bOrk3INm3YlB0Ts5XMkyMRU8VArFNUXCnXTCA3U0w8UgPNb0BDSOE0MxQM
zkApiaKjKyZMeTMmwYrBrNtEL+sMniNFEtCUjNFFr02D3xWvPvRX31dty7z1adrPQdJ8oDIWvRNP
KkqYgAO9j5tWNJhbYTptDPdzTp0oO5KJ0MWXdha+8tOg0Oo+INOfpG0/5Sq4c96mzoyw1zZAKxZy
9bj8Me0F48NI+9+c7M5tT1/GjH8eHNHhRWpJAyqPOOsz/PkAgABEiIm4/JPT0/uYiOjIV7BJcE+U
2coSfDLvPqS7+JVrLeFCGnc+kiDGRv/ufK1ctB5kA3D2NxXUVk2gbaPMnmjqLZRIJ4i7h2tP8sA5
WwFcnrjULYHUH+amy9fx/KthdoFiYRmBIBXM1tgB8TLrZH1Mo7138taaKGTsB6sT5Rs3sj8NWU4J
jNNx3D5sJbc2RYXb6oAniiBcbVyBKjNMZCPuBgT7lH7+aOjTgVosk/M2rHHzEACiONAXIZSeR/kM
+jY+TUONqMhLEfHBMOn+pmS3YY0pqorEMqBKzE4dUgtwrB7AUhw7tMjCqrNDLyfoBkhbm8u+QPk+
NTtzi91QFDEHUMNJqjMObFx9iaGQBy4WNAbVRQChWJRXLd0zOHZ3DTmPq+LFwng8C9V22HdgOUos
b4pOheGikmcmlqwEU2hTmCY5yT3O88nAJb0h6z62rMqMMsgJ+RPHbuMvSgD/25cXUQF6bclSbKBM
hjmBbdtluV3KhZRSkHYxNGAnKxlUUjP5gxGvVJaUUdU4fHwLMqXymDCyBHRhUO0Go7E7My3cdUrY
uwn5t2IADb2PRifVtGg6vWtntVKXuDSZDiqk4e3tVd1uoFYbC3PSHcdVuN0mWbY4OeunBjfmnJC1
SnI7JK8wPLTVV0zwbPwFT1RV8GBR0xRfe7GsJ+O7z4576YwkN0p4vwpQYdTZAgrcB5g8Zj4fHma2
X7nAi/y3Dc+w7ZFH86ovq28bjq3m6YIU4o3TmGyfh3rJYEPsElR079JnIS+RaiIwM2y14Boe/O9v
ciORPQS1nhst/S/WMLcqdB0fX2ne49Ery/L7W7mec75ASb9ggLUmE7fevcSFLLKlD0y29E4EW5+v
RL+lp2TM7rDdDbXtjeWx5MSzguuIN5mRyv3algyosOF/NkfIkDoWhieLOvsojPejgTA6NKvIWG45
zP8wMefAlih7+BkYzhEVoCQojNnHrD3dSKAXQ9Lsh9ZiTK/d/RbOkN7IsBg2qBDQXRQ9Sqod3oY3
qjkkbjOAMsNmYUnM/ABj9JgB2yp+urqYqtyOPB/tDJY52i1repjgUsvhmlDn3k/9bvdOXYxySUxA
gi09Fngmwdl8BUlEYZLn2bLPOz++WPbSvXJklv4rPYhRwqBInFdlV+SAJcFkQCPwOXVbzrKx7mmv
fM2G60f3nS2JG3+luWbyPm6RK85B66suh50AeP2m2LPEIwIW+1fqzghMD2z9AjQ0LzrmxrP3BrYl
OfvtLtAFsEPf0zaKr8OfQO/qiumumvPYmhKMXjg24+pUS2zlVW67CoiPkQj3u8lhm0a89NrwFr5W
7k58Do+MEu7dGLZBure8SKna1YsS6NGhGYMyQYjwZpUSnRV/DpISYT4/4xS14vrcmeS7yEgD0DPe
vlSVIXGtOmC4+5Bcne1RgDR0sicilEiA0i7A5y8ixcD3bqzTAwzHPN5GJ0QUj5W5u2oxQxgext/5
/v4cuylz8irY/p6U+pT5oowEKvYkcRqh6na1Ayh8a2AtQxD/WczJMNEAJOsqLpuhD6W6M1VrUt/C
ar1fEY9wY91vmazQOx5T7GDNjTxz7jBe7cdUaMxFwQO77hYbNvSvxmb7DoalIR3ew8i8af+2iXb0
Wv8l4d4X6oHLJO9l+/FZwpRwuIW5x5Nog3QKxSPemF2cjKKw67mpbiZyLwnN4eH6QQCIgW3pr08R
c9SA5IKbjud8q59V6KCHgw12A3RZ1Kw30EsVsxbIoCsZFNoocZ/zuGXagOOi9ziDKEs3DNmv0wBj
zaoRzNWZiBuHraTM0L8aDtYjWWrlDCQ2bOPF6Kya398BHhjwbIZFHyxYKfrJoYQ8ZYG9DtK9gvAA
KLf9LUbU0w6rQbt+bToCEMZbnp4zwo83z1rY6SpxvOayFp9OGvJjAXGCzENoCqXn70Kwtv+viE0f
6ImUF83My8I0l7vgy6o/yIT8vXT5IhjpGg/B8eNxUT5pLI16pw1S1ZzFnRcjVA995R3xFpv2vdEs
M4BUZg52oSn7YqK4KoTkxRzBnz7iLiEVp+nJhLaXokBuzaItQbJNmSFpIqKKuggIflh29l4RAmnT
m+/QvX16ioi2SS7DAYmhictr1VKakEyvyMcDOCRaT0YqJyCcPNnoIMeuGcKE664JmGotWAvkCH8c
0buzpxDQPqyYwwQaYEyyQ8ssf9nwpchw4OXd1QBo8jjTc65nwrZouc7qZXBO99rEQjiJM+9xMFJw
9TRXQumrkHrpgheNHKnrDmH6drsTzG3xYx4t/c8Fs4OSobfqkfkhqCqrLiWPdqpzzLhITqT0ZyyC
dYwZkgpVFPeFm+ITDOQWMcAPAIfm7iQgK4Sdg/531nCetVO/8awGw9sMZnYL3u0mOHy4fP7DJjNb
GaybnMlAwHDczOzMrRNHMcqm9TKOhrdTud4e05DAbiRmtr+3+9BzOYWiBS3CPrcZFvcI6PKIUB82
tQ35Tdj5RluXGmZQ+EsrfI0AVlAudPiIDvhmSXJaSaq357UVsw0B0au9Ke1a036K351bN/AmQ6Au
ZKhahmM5IKuWS+lFDh9EtwGiEq5U6SZPCSo/eTSGIdByMLy+zFS0va/V5bS1mK4TJ3xAuV1s/VP4
HN9hfBlIVNxnEKbQ6RNcwDUTnOSZIlwNHb/7x33w9cz6PIACop0E1Eya190lfiD8UyTYfr9ZyScf
tQ+ybd9r9LvRbJeC3B3+SkrfzZ7qjJLEm+TUIvdEh1fRcZPTChLZRQ3Jv0EExoGcZ187iSrZA+YU
DJ5sSCcRLJ9h+hSunv3S69hV9OLLXbytMkdN9K9B1IzvewsXFxoulsjTnv95Kc36HhfcByElqY3N
jMnwHs3Dj7csjx/ro0jrLh0OTm1irCFJC+i20lX2e5AG4bW0qbwe2AW041uwyBWf035+zWOVCF/3
WjgqkYZcLvYG2HP3PYxuS8kCfEAgq4/1xl1WpJuRSOxhM/Gwi1TMp57yULt/ZzwcD2DTzm2nOlBC
cXjSIV6eT1gFbviL5wuX8UqcWCXL7OPC9emrjL1x2UHYUbja2uYREqJho4wZWN8Ik8dQFg3qeiLA
eKPc7WD1zmlsJSjr8w4NTtVFsDdgOgd0dX2kuwbGM/qGgXsNMFJEof1LfXcSL55HUuSL64nWB8PM
G0BVE/D9b7m07KbxNLSuWWeEzcufbCSF+hCHjZ/9Mp/kLtf438tHicjDVW5CmC848x5F0ml2SHnw
QwyXltc8YboWG0MA7Jb14sodOiMGCW1tJ+ql//CZsJ7bf61fIUPB+OugE3nx+ObgaYuK/COcbkbS
ycd2henm+96K05074jYr5sWuWmcgDVg/YCtIVoZWOQNdYFw7tKcngiR5nchK4tK/oZ7GI9jZGok/
67lrGpjg6hLheSE/5BLQWBof8qlNXVPm7wVZjcKXi9mk5kTUuHlI5btHE9oWU9QGUkH16lyKwyJZ
GBoGTQEBHyCHUU3iaCXVKkUTCZhn4uOjeyqa+VpLibLGJ77+u/Ja3tzlGhqTos8z7ETitguP+fff
ibHcOw4322/JHaIiYu/ycslvNoCeYrhx6y0SizsxouNlFgj2R2Ql1GIG9NqWtjM1esAGft3guejG
4K5nwnDi51wfFdeNBLeLE2CXA8B5VUHo5lE/DGbHmF3IAbpvauhzZ6cbg/JUdHy5UgGlLGoOVKfW
5LcjCjCQ6m+RxwtmrysYwmVoqiGQuWDBxpOmu5vD47dh3KuZPYXZ
`pragma protect end_protected


endmodule
