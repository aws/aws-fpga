`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2024.1"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2023_11", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
BdLMkrBowDA8e10h+B94E6qIVj1d7WJjEOG/CJTJZ62FfMPToxzYV5ySTi/3wvQzqBMT2Sqdm1s4
aprTg4FlOE0w4X5TT06nXMCYhdAsNBTDtqHXcfPMdkFocZxBq8AIMt+d10gWsa1vAXkCFfzuZrGj
8yJmPPoCOvRX6+Cp8q6vXY4AI2FDMEc/w38UrSrvprB0PWk0V3G5yGEnSD+nvCwaU6arKuaqQ2fu
w9ysUaE/wDULsz/6KjyGPf8aN4EXVzSxIAb9vwmHnPrX58a7faurk4/HOek/Cedm7xcFVhrog+zb
+429j70QPRqJF6BcyIFzS4FUJNnIP8bTHGCQrg==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
Xp5WSp+yhGUniwy/jF7Em96RdRmeoHo7zW+9LPlehDw4cn6Sm2torQ5pLOd/cRXuajDHo/ZpSZSc
5dS+k9MQpn/QCXLF64qR4w6HHK9RY8HsE1ITXEpGGeJte5tul4obcd1gHc9MCmbfSEYsgKhtdkhn
Ss2PTfjcsAag2vsG430=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
JtVfUKjt+FmrD+G+L1bj1kr2bQ0dfq2IB3LMhPemI77Im6JH3RSTad2jGVf0mQ5+ToKmx1McOtr6
VFcxV2NyztybN+lJNffJ4aQ69yDrL8G/IsOZVB4dOSU53nIqaIElnrH53YrurGf3M4k6dmF6kZ4p
XZ4uARR/0mczprM74bQ=

`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
YHAr+MBd/X3uZPbN7yJxf0tsc1J2tp0a857w9ObaZV9IFq4916cra11kvd3rZWwObdzofw553xDx
QrfphoeQYA==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6304)
`pragma protect data_block
+zpjtILdugUS85yH7qK6xi+Olub+UGcoGwMueW+esfJqKe6Tzjd5SArLr5qvXIfIydTmMIy3BDj0
AAiXOM/lW1c+jOPO/xdf+D3VTmjEhBAzeXp1+JRQt8Ikjg6zUA2+5+PMGJy560OTa0OqcaOCXScX
dx++ArHe4ZjPBDLAcsSNc9l8UMTlsoE6NGHgT6zY1QR/UUtTSlYOHHfSwEt6ikVZNb5nM1zWYGRL
XNM/I/3uz+zkkp1H5SQyE6dC9vQRgfPP42UFHmy0ZvppeyUHd62ZCtg9ZjYoAmmc/ttLHEA7DFPl
hkW8newsGMPnFeKCr4r2ETKgsaPszoHSDnxWmE0HKfTzSYI/yWFTux6+sJcG1f2cLF6mELBW8y/e
FJ3sKiDSswzwaEJvVvVVqwWz3NMzNS2nIJib59Fhep0xkM09IXjERoxVG5lwGeFsvIKRFADzwOHr
16jBe2tZVS5t+X0seBwwuLFzcy/mzxIjolkpw7X+LoACjLHKuDfi1YJLjG7jVSNwPNY3OrLTXPd9
lc61jv8oqvcY+ekeRLXJhX8LhBfpjbNb2206IrKoQdxkyMil18XqyBK5djKW2gsZ9kk4LqsA1+lO
wvQamNX33Wq5k2hAHCQxlvinlQ4V67qmOS0JmV2xQd9c5vZjOFEySk7Hdmy7VkaKgNPRhPrcQYgj
tWAr0NMjEH463gu4PUqkAxJdkDKMi90LbPWplpF9ljjjCo5AyawAVWm5m/kuqhbAbeeBr0eFO/up
bJRp3ABS95TRd+4fKnZP0z2XXzHKFUaHj9QrF1y6coWvA5kbH8uNq6ucGpJS2Z1sJOE/P0r2nGmZ
P0IG06msF54pqVy0yTKnIW9jOorvw7f/xbVfCUzkC+IOtD4ClmE4cbU8rfEydkdCjEizmzf6cjpo
eLP7WMApbaQXk3w3S+LOtVOVosebeYs9smGmG2pF3N+SpZjpMqAVSl4SQoFutmbsD6o7/T4fqQ3l
kxHsjRkw2CR5AlihSrt88EGxVCsIuVHaCCVhs1UapxN9ZZJV4Jr+VHv66wg8QalntLMlf+xzKf6Y
sEMz8bMc9FDIOEfPWeLdHr+o4E/vFspF2UAUYPAwPuHKlxzCgvwY1gZAPUWZFJcgCkfWNgG/MpYc
1csWYBAJxr2qDPple+VkiORS0xSRafHGBD40xMtfsghjhMHIl8ojVKoB7IDykb+9T2MvLCoCPY4Q
PEzI9fyarxd3DeDATtixQSUfX7BfapKWlRWwHrNzTIClQ8Jv/S39WK5SfYDUB6BRXqNmFwMM/mQ1
p+tMC1cwKrTXzeYBehEXbsVpoSxKAfa0MQb6V3uaaOMGOnMAUb61NlhQS8ZUXPGAbKpr2nbV4MvN
o3UcojpVoNGx6Nik9I3J6tCT/R4yCuSJC6QjYXvEH7RhAB0FNqDhBnTPlYwIGtEvaDjHhWGhQ8hu
eXh6DBegbFPnBYcQDgWIDEgAvHWlHNk1eKby3/bsBkHV+jp8opBKYTNZrm9d75who4zTpcvsnSOp
urmUcIsD35Q50EOrFD/e3WAaH709Pw3vhE29senDDRvV9NI4sWF+b8nh10tif8APpX0a1GGMmNCr
If/rFSNhArzWnUGHezQIT7aLE6z0Nu8ISa0J7AQuuLLEKxDlNnZvshRO4K8sJRfZ9KDhi680lsP1
jmrJJt2LZ1H0yL/GijAJOAmqEnm0yICZ5y9I9GbobS9Z3xaOqKw23lCraBUBscAWu2cWu0gw8odr
WXBdrFeWWm6DRDhrpge3hGRmSWxCuh95cTbe9i51MfsQeQD5C/WiGLTH52loJlvew1YsYHmv7L84
pzZC1Jzlj2D4JNDUvH2Mj8oW9mUoSBx5dNJi9psKZXNQW8wGvV6af/hLn7342YEGp3cwn8AOPpt7
5dpJ+afNuRzT4l+/umMPCpzB1Q9JxM+pR1a8iJr9AmKY1rXIM06Y/tiKT8pCNWKQ8TkbZXqjGNZL
ySBPuQmuWoqIfSI+8Wh31+ice/g3EIwuNzchjPPVWkFU1qvr4ihuStyNGiLf+9530ZdB9mJE9TOD
fT006kOVRGjbum4ydkKXyb04MOuuIa/hxJ1SypSVKI51lukZjCiAOMtvPTCHTLkLT4kVb6RoeYY3
/ykZ+AYg2yTIUvMHcq9X9a1FzohdREPID2fFU0caB5S2NB3F3YAEpCBxAw6ulZ2uE+lJ3p6IoWD+
s4x1b/2OQbSiGluFKtX3n9SPlcDEya2e6AalYaTBYxSnsDL0XRgPsl6DTzDVvkRZgb+Y2xOyrq9/
48ZfytU9B5Ba2uutAHR2uXU/qOqJXFzBUGHpd4cp/teW6ZkE5hwExDTAMsUYKQo6feeXNiazM9D9
GKQvHbxKVaF9WGc+5oQnxTaMoCFkubqFfu26htQ94A33npT7M0lv5JRxbxzGN6oBm+VizYhE9HOX
4JSC22Kt5CpgeyYXMJmXBHxP4w1MVxHSkavCtx9vhk24JZ+y9N/OhASFz3FVRaA8kKK1Tc/0FlYq
nc3bisLkg3+JVNeSkHdRIwG++L18pOOV90QfuHPqOND3u/UKAh5kbc4AUijgnspUuVBn+mUEihXM
LwpfNHeXz9l3OLADtOdjPYh4t9xeTvI7/8VpBs7z0ymjMOlbtU85Fnqre54NDFrImQ3FPu8YuH+1
2mvnMW4yg/qmOJDtnTqnk9JMVI5AHkqlV/wWooz5YcOQehfdz1Rpg+am4x8hbqtRJSESDdl1ryp8
1imyZzpC0HgKDmqz61AJLX6C/afJ2OlGWQg2DW4c/s8sdWgpGpa3CDPXK4DR3qWmPi+C1J7bNSWB
eEUjmHUPXVPUBuFHtiqiCvrFA/JfmZSPOGKYdN5JliDZZYjAv5SzD+FQghBK/z3E1Ub+NDHl54vi
g9PGXVFBZVdULJC+BmhcBwG4c7v7GU7SrBUp2/p1D8IXTtUnISDwBsdqezWpGOVWWzzeCy/ji1ba
/59Gua06duokV2cH5m2HdNmGQ2i3su6L/7Rge57M7FGt4mlNgQr5pUQ5WNRPW9OyrVzAErLXUJvn
43aCjMK2gMWV6nJLM4JQZu56kmz7yL4FQLT/Ln5rZP9SK3V3C3PEnYB5UUG+62yyqduy+x82DFny
je2FN39n5vWEhBnkXsIRPajHJAnPMVTB3NCr5txfLZFeKrVjEan/y3zEQFPfjoTIx2E6NXvn7fCs
0SUx6pNotDprxlqP7qL6DwN3fLGcwA+Vejjph1v0WAzLm1UOt23vbQG2DX8/hZLe5j7z+tGvJfxj
fDEdrzbozDt1QJkA5Hmz/gI6fk2WTe38OBl2LlQ2FMdbWmmsfq/gc8ZlvFRkjiyE650loIGESQB2
/aEk/cQ5DC/1ZWFbmtUZRLav4a6Ps5XbpxKcTIYHVEibAfe4vlmNTWu2cadV8lJw+iXKqnAS207T
A9uYolG28ea62c3EzeM/W8cI1amc/zcAkle8qO6fxAOOnnFJ7Hbz3Dpvhznl9jdAcixgiWyPOYrj
AHMn9kkAkGjTu0aN95eGw4HwsC9DhQYB+cbYaT/Oy5ZPmqxtwM9yus9WluuK7zKUZbwLH69bmlxI
4k2Ais17T+woOZnERqu3C4iFjlBZpaIL6fNwRF9HvA0Am2e3xnJ1EXgbyMjWhgRiew4DEP/RnBfB
2V50U9IExh0VS33iY58uxbQpNux8j/mOhsMDXkOOlDAeJrfv8H411uOIBrUwm7xm0h8zBDsxA8hh
UbZQTae1fbq/XPMZxZi7a+CAOH+SayZNAhyLr35xertqRbKVQrf0M6j+Eq4f4GhWTCYbR/rYk643
E12bWRfDgK2sHS0vwBT9pUSPUy4yDe38Kr2zVTV14afPNizGPlMjOP3Wj047czOm+vCyzopJvXK1
SeIUYABKVJazylaB5Zgcxya7hojfD9AYXTQYnVVR4RN4Vd6MKXmj+lqif7hwYx5Fhlogm2rx90iC
ThxlsPCKyOrjj2O8r6Dq3oNIdvMMKITh4mYF9t7twTz7mgZNi+bZnbYXVj7zAE1MHB/X9JgeExTl
oZk87AAqwA+pzFC8KfXSEG7w0MyaVs/Iath4ufmve/3efVPk2SPuOi4FxwvovACTQxUFhOOkAUAZ
cJ2OvAMSTY63rRg60lYkWC92eJ3WXmCJ3FYiwTsdkgxDf4ijkXNeCnokrnUHBZJGaSNzdmDnMLK4
NRTwHWOQ1j+1v7d6YNxf+Cl6tiKXzTM89c+LgmHTCmx0ju6ggurVvwmHl9u/LRx8p+IxLJHUred3
J9pZh7yuQUCk0EVtIdZoQ6ougyItlMhQcq9IfeoPEhqg3rCErRTNMDgxyUzVPOkpdkY7sL6xsi+S
eOTFJOV8XhLMbzA2fR9ue+t8v2O4OQBSgXfXiQ7yWmjwE2KFNLVrtxlJi+460yDKBvlCADI5+AS/
c1df/ycKqJjnM+5iJ7inTPok9Mek5YNiRHG8UgYHKrSaRv8Ff0dbgraoifrfzICzlG+lujqIWSEF
nxt7ROe2Q6+4BXb0bgJmADSpi0RL6CJsY3rtvDNCJzFdZAQZ4uhTtKbAWhmrP/J7YxIccscWOcbO
2Tv7XBMpwouAVlDE7AZ7hty9p85cNj/5yrT0RMjkl0iP1sOUpAYaPk63Vhs50JDLPUnKBq/lkzOV
v1fj3iUMGkiQ8nBfAqMnonqHBKb7vVzQrD3XKGjMTmH+XLTbjVCRisQynFzAPRD/0rGqziT+oGT2
N88R/AK1DYKGjv06pIxCjIphgN0OFKMLUjHFH+7HIXRokhh6CSeomgrxSiebwYBbr19RLdoaUQOC
TpGvdRbF1FESPYrr4nnpoYPEBW/cew6Og5OL1Ib7dMlEFB3blOENiw+314zuy5DBC542cuwF1Dch
6uedr9cfEy/4mU/Q325shhdz9Mb4qmdD5uB8XroeYbAKbC9eia8XsiYx4kQkHKs86fqHGT14R5hF
zk2nW/Dx6+8J/ELW/rOiyd7E7GrVNSSrvUMX0MYlwj4ghjaqhga8goQmahIWIhGV2+ASuvYxVWq3
gycjQXSNckjh3tC+L3vvL391wJWlQL8jNTzTCzMzuuU8xL6H2x660rgc7OvFauZF4DcDEPGjCc9f
62ii4WfTGyh0ra077AFrZvdGU8z3dz24I7HscgpC8YsomPp+7ezrDAa7HPQ3fH0WOxrrf+BdPb99
1IJP8wW728wF2eypgLfub6axjTJN87ER+d61LNqU1DhLo8r+YDKlRtYEdwqPFGTDe5O/tzVSgYBr
56a8u9RY3wtzzJjhV3ahn5uXeXXyLxNnuDczMuyUBxWOobhU5frxjWoULo1TAaTvIDFhVr8lON/1
WwxJkrne1af/xWlvkz7xV8GPhZCtgWTkcD2PMQIMCf1kc0Wb/yIqckryp6KWPuz8ognz+AgQT1Ry
uQjMp6YK4dgj1ckdgQHNQ0dYrcTygpFGoEgC58OoEBQ6t5cDK3Y2EKSUXhhruwS64ikDHoxqbrjR
CGa0dvTxJTvtTQCuGqmuA55COuSjHWI66AtXGtY7MIhI3llvuZ++x0bUYIisjfVUkhYW1cN6+ukt
PsbXf/EQ1Bz4MubU7KWvfxvoiuEPcPhVPH1QCI4FtFZfYzM1shOszp80AGmWTQMUlW0iYKoRHEM6
uD8Thcht1mdQv/hZfc/AZQX7TOfybyCO5syb3gl9+n+bflr4/Od3s5JlFv6okTB2GJFbLSBsSwRh
dHyuPfmYRgxCVX6fZUXcvmTTk1QUNUb04HnLwATyR7BK8v4CDCt9Nm6FwhRv1L5nQrcWy/Ddu6VY
zPEc+iuiecObbejRCZhjbTnctxGeK+4YxbUB0JgLP4YqR6SBddEFTMSgsSBEJgv3Jyw9WGJ1Gh2X
q81WNSt2670XPXlTc2/iwIqOVeaSKkS/g3QmKA5V+9aledons9h4J9tvvkPMg68YqAmgi8nz2t9d
q/0AgZKX3yL4S6qLztqY5MBJFthZLNE7Ywa6TxfghbKDoa6jmn75UGQpn1mnItJeV16jFjuHHKJs
X68gZYIfjuOvzADk3RlCirW/aJF8w2sPkgmQ75HnWK0AyOaIYxRrz2PIm9jNvGRFumfTBaRzq8FT
GTfaV2n9bDnsIJjwAGizlKQ0xQjgeg61cRq/JZybHAgXlQFBeZmytDQ86XWIH1K26CNIhHSzyKaZ
rhMexW38ahEYeJ+CUrzOF8dMH6RyHY8qbYEamjvSgvDyNV81slMoV+8tR1IYb5NAieeYNaxbYDsS
gqEV9TzFYOm5y662Qzp9johIyBgtFzOePyUSJqePapyLWvZ6IJvIpEe7xXUfFHcWypNKOUGxztEL
pxXg8Z+Pmw4qBfodW1rFqfUezvIiJuD6xTWLV73TYHUW4gw3qWBSl4CIXfN/xEElcv6Vsfg5IqCw
70rqFXcKFeHZskZNSBMkmYqaShzhqteCkH2c1p32lX97+Ih1n62ymQKxUF2fYhZM9WqQPnhsiadK
kXOINwB1hQVh5X6QYJXrnQPKKZppqTeCvnCUVs0kQY/gowyEgUNFgj8mw6D9WOBRCZrSTNU4mZXf
5nuE+wPfFTuks9CMNxCepVdDKl6NF87puYe5FXgo7agE6hTsES0B27h442kSblucCXbrq6sBLOhD
Amyjemyq+/vpWhXcKtxvTkqIqkTBUjjJpwh/RuwjlU3Q1wIZZoNF7IKaW5nXNMx8lbSLkfG82mHI
gQnPJJZq1BhYxsd+J4lB317Y2HL3dgzVnvbbZPzoEVa4plPX/W/kbrxBdypTVtX82CqB/dnov2go
QVY/gMQLXClTN7qz29vUwc8fl5bpc90lbyyLlvQ6JhOOp3AjucOSJL7RFcbZYHimqDMrIFh3wCan
wCwDe19bcyfP0hiT/uvBhBvB4j0Dt8sUqaBdPBHqoKiDEF+02VU0DGgykHveDe7wXydW1UImFaBy
eDxT1o6+FHzBmvLgeemoBN3lNONaGVidNpczkjKayVbBrtXxqetTpj+yUbTP/4lihRhxzvpWhmm+
Yemy6gg5gK1Y8UedZ1aW3Sh7fTTTkUvVunGdp37iaYPAo+JYF+xAgqHBm0fq9LRvIF7XbdDW23EI
lPrTxkftgyAxT9dUY9TTEy/u8QVKkk00n47Zjhyou17dTRbWq2m9k+I2DGk5TlebOWUzhdq6OAzk
ZNgPy+GJL0e/7v4NuS/WedaixeitwwF28YGNQzTOA8yfa+0zk5n2ENvDXYuEGfw2t6mUX+xwR5gv
0zRS0LIvLNZ1sTgSDrpjQ/zlmhaukhytoo2odxlLMwEc3o75dkIBqZOgy5RQFfgD3bQKrJ1dD7w3
1ir8RcOcnTi6FowfPY2jA8TM4sp+/h9NxNdZUdwJ6WgyO+fbE7ywQUAZ0wJdNXQZoovrYpt7otq4
BhG/WuS3WGH4AbK6dlKAmq0XVsRz8Kjvhrjkcp5ke5DRz4Ug8z3M+lKipr4xWSu2nBtNQHiPMls0
TE+FGfjvN5glKOe0JMUngkMjiyriNaX7ze2ie5RldEWqQZwwenIj/69UPQEPFHQZ+E6jUZHR56WN
ginQCK42by0uFEbhJuoeZJ2In25+MiZgf9x5RuIhhEiHUclJ7gXq90gP4pha00yqVYJdPZ2zWuyI
Az7GD3v0ZNFWpxBXbT8tikiTDfBBAdrS0FoyE2Vl7vCr7pSl5dIDqYgCS6CMVQT4jD1WRJuhOz90
n+/zgorAturER0DswAjLm+UjCIdp65iMnIpAiwtaRCF6p4ZDr2aGWydKUOgs3OzwyE2ejkx05sZR
+1CxTUBZ/1XGvZEZihM+gXD343sBRA3dsx4FrQiN6rFs5kdUIGWi3JAo5wGEECXcw/9+pRVjMxsm
REeVttEjUcN4Fd5+zDiCe0BK8BMFydrDeTz8R+sT6C4JopRlwz1Aje1GEQkGciokwfOxfB3xcMU7
zLpalDewVZxA88mPyTeR7rjd9p4gNAenug7PUeZfLU9eAvgyiU+c3oGQXRM52JzYIO5XrlqAdYc2
rOpoPwAs1RW7dSLaLV8C8vYXf905oNTGmsXtlW6l7Dl1yD4Qx4Jwnr0UJyGIY4Ef71TOPnjW3Vur
rh3XjQgtS5EMJddhQxrAskGr9JC2tzblECOuAiPa2Lq7RhKRYSIdFVRCKwuijPWiuKb9LSnMHhqN
FRSM59jwItQJ0sTRR45pgwCXpnvgthSTAD+fEXWOfcJq2c6ARnPPOrSpDlMpFcQSYbnUjLQ6JPBK
lkBx8YAK+49I588LI+hLVko1LRqMZgbI37VsVy7PCDbxWoW149FTzvO4MjB/DDnDJgwocWtdpTUs
kmiZGesLgAH1kmXLqKZPd1Xq7M0SDB2eeFh6zUxYD5jKw+paV3FqnagkaJ/6L7B1V4taIdZyUjQK
1q91vBfTA0R7/MGdbxMIIuGMys96DiIlA/4KbMUtuKBRtA==
`pragma protect end_protected
