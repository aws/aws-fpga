`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2024.1"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2023_11", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
k31BtE0mli2q86FQAozbvCuaVnrA1qPYotLn9gvbOF2WSTBN7r68U8SGqWke0AqjlpSxK/cu2cJp
bOn+bS68hIRvWOkHR869yaJz2cD1VHMX6g1jfW1o2F+/7jEOLLER5J5MTYEbL4RT0NZCHtOVEajE
UCLAB5yqUAwh6c7jpRuiZ+Y2CiqVMaBI2OuNLvUVhR0wq+WtL+QUlmike8MKOsIz5Re6klF2EXPH
S0XlljlqPeqJZDO5OidDtnbE0FBVe4JdLoljgjxFLMLuuSnGh9lGUe33fh08zq/jv/qG9/tEywzv
Pf4AQe1KhWvvVHcLDwDe3sKXbASwM78eMHZvuw==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
p7E0UfmMBbr7TLaDDWB26yDKz84ghhYE5m6uPs5064JcniiojiA0HuDQQhSzEZSfLMW9N9Y1PIf2
sckE9YJhba1Lbsy2xrOfF5belpqvJ2om5lxQ355QHLAOFXcnBLEsXiN9YNaH+vwmGwp7NP3d8Bn+
bMHB+2uS7Xoao9TOtWA=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
dd9ycREIjKheskezwU8l+8KOahXm5iqGNCRO0fTjPtPjPwZGIKkVIAVh7aYOgQtyNejBHnYq1Rzm
c+9dx8VX5OSeyvcvtXOKNm48r9ZLkC9CwO18nG6Jaew5r0BknbYHL2+CI8693UnTpoBNnE61puRa
gzKZ8fx4e+LP62NsoV0=

`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
Gas2ladCjOtkhakWq6MtiVu9bVTbx8zn3nlHQlRz7au1QaEWA87rOoCvrwBpcP/cdurGYEwl9kZU
AMCPPnZHvQ==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3504)
`pragma protect data_block
1VN4mB4QgZYDt9ywLVUSgMpLlHxCESCtmNvvbt6kuxglt4t7sLPm7VwY4xryl8rFkGGh4HsRuUDm
Y0OMnJwue52n6gUoLzQDd/GobGnbQPTNd3/w1RM4AjyT/RtV97Q93umYijq60K4Cwpr1bPoAzAUV
lSBp2lFN8EkTn320VGQ49+ofK4vUtNbrW1Fk5zpzSPDTIIu7WzfjPnZV9Z3rh2P75Xbu6h5VQhGv
g3yHrtXknb6v5pI/Q8pguKAwJlfbqBLw5xECVPCaz1HP6+ilp5ilEIEbAhZD4Glbx8vRZtSDtTJ5
0OjQfWEGwuq0Mqwbmf8Hzz9zCuGjEYKKjL/Mhs5b1N8JuTYQQ7uh/RvyZZqaWhFoVlnarj/iG0Gq
pLAMIUHESeJxsaEPk9Q+1Jzn3zPi0r11YiVWYzHlTbV5y29xXkPDsq2IBbbykDBzpfS8jUwqWhZ2
nqfC/0sUYjxVin6x1dML/XdEXwem1gjteZqgSn6TMWfKuTwIA0RsKCGbB74bB+4vXo4VDrn2arFx
/qmxUJ60DZo5O4r4+IS4jXCFsKc2wzUN8+FKxPQfu37z1GnGBbPerpCsiB9urv9flA3O67egksr5
hjYeLDGyWCkHMbcJ2M0ji5nt2VaQbCZ0dBjTjXxvro+yU8gA1M0cmBwa+K8OE3LVI3bW8+AE/kwC
4SFCebxk83OwbIVyUqiMA8oTkmtIub9e36nq75TdGu2GtFAMDFPrtaheaCZ331gwlIrhxxlLguCa
2p8bHWjJThvds288NpWSo1eTLzyNiZqujQKGiaIGAkRbHqJfQUq14TtBo6ILdD6m3XAOBVESz5X+
eqisecH7onY52VJXHGDdU/aBm6xjkLaKdQu4NbagP/r/1OmIidnXn9B1Wfy1PyHKknhr6G3HI8I9
idsxCKzxi6Z4t2wq1yRd5RB0c9xcSSStnFCJBqSAF37sMODyk2Wt4qrSgRrt0LXtIDj/fA2UwF/q
oEFTDy4BiL7pLquM+faH7O26EZs77x/n53zBMDPu4dz4QirjcgyL4hSUMag3mBy1pIPcuaFfuoaC
Ute/XAdM1Ahx4mZGkZDWQDm3/Cp5f8XNpDO+hSC6AOEth+8P7ZqXISRlWO1D1dQk/uIl1ZprZ1hY
WVC+d79VKV9S27HYvlN9NoJC1sA3ilUhb8BFryQG2axOrYuhdWSCtp1h/vBEwm0HR8v6RBRXw+44
rWe71fHUt4z7NCKcYrJ9GlZOCEFTT4awn3bH6gMXddsZvOwV4qFATkmoS7E8wEihYe1B6z1ZhQDd
Qiu8VcxIJz3QdbDCM+8MWOFrQsm36FafJSB2a4kKMARlYHs+tGPCUqKBiw4LaJeQZm9YzmtA69bF
vlkqOlRIFG+GnIwmqhGOv+duFzFZoqalKELnK2ajABDKY+CXx8MsPInOYpEgIhQ8DQrw02jIvyMV
yYUQMo/iWPo0DT2q3eSCqVwCzJVIGiBuyND50IM4DYc5SqQTLLZ0lfjAUwAsye1FlxID5r+z9nzo
OC2nfQ+dl3X0psNNEzFcApdg7OG0eTlS1y/aiYTaZAQI2LZ4GNGjTUrCKkKNiFTGSUYQlAqqPfjW
hUBdSnf5EPH/Ahtoen+pSvEtx1bn4iuqxKKdUn/QLy+9718gy07G/l4PkUTPpaqSIFzb10Q7qoOa
JNHNm1rCmc5XJLfa1f+/B/TaKZE/yTFOlySYxl/RsTiFeF24G9W5uy7mPQNlF9Sbm8qQYJQ5or/d
dK5/WzMXythqM9ScCuhZLqvDPfCyxn2RGmFMry0lfqMDw3wKknNVpYMjWsI9/qMzWtNssqtiFPBJ
wEGN5CYsQ59pbarLoS/HvhoPnl3c5tM44h/gfaC830PzLpQEKo3z6bx35BSZ9gOMerbw3LsjNO07
cO56mbHjPa6DPe+RwsGQhzEiDUvUsEQ221Ict34JBomVJmNI43XPraNMKQ80H337ZPaAkpTddsu/
T1a1l7bDXbNEuNd6rlYyIHEZki52oTehEzEwL+zy0f94HbZK/FhNQ1Pl/yoZOOQuZBWmgxvLEpMR
loUgn2Jyzs1TSRrynQvRudPSYHoEkW8uOJO3yMBB2MHbta6sfN9NKV1y+r95D3/6fsO1MLQ0O0d5
ok8sT7lOt5pLnnbpfpwucPk5vMdhvuT21LVNaHLgiqvesJSxYfY3ZeT7vJF2ac5N2PWzUeEkJqsv
ODInsnesEFRwh3oCuWCMgBjPRgpmAZzY13xkMcVYC57FL2yZ4cbMXr4KeVNuvefT8O1a/0wqZjJB
iDjO/sRQCXq84I4YmRqdAlOU2Jn76eLBuHpb8isF6ro3m7jwYtP8ZvTR4uxQNNipx8rl+zSlc/I5
Mkfu9SA1016xDFFT5mw+Ex+ZLQEK7qoh0UitUQzrA0J8XAGVpKucjhgBBJBgXO++6WsvjW714R71
QZQXLhAIlFyoHwTMB8mI7X75CHpt0mxQvrXyGJCgJ6z1ArpteAJLQ73/BekDYlMv661tCuG22jc7
nK2U7Dn1Nv1Bd5YADLNJtFjkWapEW/h99lIRDWhvm1W89tTaTnarc1yr/vKLf26SvBqthPcS5gsn
sFfoL4TFwAVRgZ0Wv3uzPvWk9XiZ5lQWDozVh7RJTdGhOCyY6N3JPIVt1c8rkowyd6vTa+CmIixJ
wIUlzD0hvHJlYBepz7W4fhVHpRbVbThoxSyNC1gZ7oJk813OfV/VXDz+am3VoUPOA00x6nu10Gq1
Y/MRKY/d25z7150Ff4aZz7zckpyQ1vctGEGxSgM1kfD/lE1LsCKFPwt7E38Tvg1xSo4W+S/lHpZE
UeHGR+TlxiDJ7JO1Yy+PDliilPFJKaynsFFhvZGUhtaV5R5HHcJNmZF9vsApnF7K7c16AwXbfuPV
jr1ndfCtOexKFiAuqz5p3xJgoGmU4SWqCGef1By6sw275jxv3XfVA3fMNSir2pbwT1QtBtpNyV/n
ryDiru0N3VI19punwLxdC1B+9gBuiM42DVoestp1FXlOi+ff/JDDaRvE5doFqIZuwokWYYNRAxVg
gb9UpwWAY7JBEEekCEEXL2Byl8Ad0vC4z08sR0AD+5wHMAuURrIUCa1lpCyM3ExqHRJlXGh0262N
b8ytUN/MHe+uJT4rUuSLOIsTVaPfERPWNzGBkzrP4hSWU0ov6Jq4vemqyW4euCBNq5yVOjftG3p0
vUn4RuKHp7ebMJ8u89nan2LDXJTFWCZTD4fyav6jagR8puFI/l+twXpRAIFib/wPp4HFTYXC09G5
1sJnmjYO9aIP+EjHWejddSqb7BO5QCftw8B1dVaBktT8Edf/2+5dUofzHvm5BxNiKORYxdguZarJ
G/6yqtD5WI95nOzzJ1ErUbOGFr0aCwoL05mSixgEm+1jH/7f154kA6ELisiJ+andqcwHxP63ONy8
6X4DjMiBrFlO+0Zm2ReepqLXUOmmTNjJifjcitUJgQPqr4V1/pp6NArz7/L6LfoFJmo5ZpvKKOux
mW5w9JXrIPuCd7lrOZsd9tjSaxjweM9l+HsSv3oO63kkImhT2qI7zZTq3IhkXQzpsHovde6CxIt3
dqSV0SyKElNHn3u25aLMSbX+5rEuz9euNJYQKC+D1WBLz+4d9zS42TsPEn/rm8klQdRHPbln7LQW
Wc3PR5KsRuQOBrPPicZvqEiEtm4fhKadNcIMVK8YvQMV980GFbdZptqsVwwwFaKVaEsGovi8wOoB
VcrsZ9ZVAy4TdLl50/cv5khZ+SN7diX/YyspyqdErO7UVOmtfYnuVF35B/MGtITovVyLw31u8tVf
YuAzqRqCdSsT75VaLwA2Nvz0OVViUl22kQca2CMOEwyU2u+FBlA7gOch35YCKmwV21S7NpZJ/49Z
Ek2izKJHQdhR49fYhFn6p/dqHSTkAzjUUCZGKo7AHsYD3U/BkPoSxBIPmWt+W9OGN4IbZmEvn0VQ
f4CQWMn6r+vPxEdPb6nQkUGueht3x9koj03ghd8nEd0hZkk/gMywiVz6u7h5h6/NfXWukV8VbzLX
kq+geARrc3C+SaSR8oEC+jYtg9FKhjoEJaeZiIg7rDqm2ismiB0Qh6Nc9/GQIp/uO4m+BJeDnGGn
YKUwWK+MRwXyK2zeaTEv+QMGP7+2tJWHZEFQ/6Y+CrFIxOv08rcbGyGPYG6MNREaIbWffvv0i3O+
3FZbQP6rnbMLgYOcga+PHmlKurOfgSC+EOoJ3+/HaWu0MrHGqzNDB3YB5Pjmwfsh8+HMqTcMNJaL
pVCIBhYY5h/9g1BEKPgKm+WScVV4z7n4oHcwpfUbFBnUmg2yUwEPA7fkML0rUshedatYzytdEHOR
7aGpiTr5RJ7CT1WNf5EUQHnMKfEOTfNXHiqd3756MNXq0A8rtDiitFC7vGASlzVANvU3dEWfuKtG
kQ/s0wVgBkijiXF8Xt+kX01ZI0MBdFXxU89AFS3v7uFRsk5fT8McZoGWs05IO2IorK4p6d3/11Tl
lGuAE0q8AqgjHTILmosW6Mz891Zdc1LSfRe9pMgZwM8kEWDxEQQM6qdq023BwwtbUppSknni7B1e
9XwtIl5HJqfEhczkBr5Igb6avPU/X8QNHx6R/IjilvmqBEQejhcQwBKu7xElRtoAmRBI/WDLxYk4
3AWEMIzt0/OoReuQufRVta4F/HH9RZrVlP0W
`pragma protect end_protected
