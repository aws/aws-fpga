`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
rbSnzE3A6NMcajBzhPp0QKPkaxazGZQEVPGqFHa1SoTdeehiuR2yjSR3BTpl0zyINgowAYd1RBXo
G994kg/QwJdE+tJwyisfGcoXXQYFxbFXNXsN/0jLLsJhMlgIt3UYdyPYZ7BdtL8Q+x1WTD9wES+j
ge26tOxAQGfkA6EXBHyB/7e08se/TwsGhONQelcn5EjbqFxciJVnbi+C9lbT7ie2GlwqbYdlSYVd
xjxjFiWyblkIV3Tr2o27ApokqwjDFemNHGpgezkVPijZo/bQtp7hP0QWYdtbVhgE3BGddPlUegM2
LTKcdY1UOlbfn4k+1aG6ikMxjaadWkS5w1QrOg==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
sKiAyNDsUEe6ubgOc2qjZytA6O6iLGWNowCWnIwCsND7N8Vjde8NyPxZWJVuA1XlyBED2T0WDNjO
/8HEfR8tv7RwQkuHPN3gReZXzmlPCXNt9cZJSUq2ERkYvjMc6+hy6EtguLb2RilxfoYxDcVFmpv1
4W9ZHkVipqzKOa1YEtc=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
osd7NIJGGKqxJxWBmj/Yo697UFCqvFXD4SOgAPUAIOJrR7WVOVG0jRj7LZor/z2QJ3Ld909B3ei5
lARexGgVAK+aBZGmBkWeTMolAV+IhRdohUZNCafnlOmNrRLvcOXVeGsxiKXIqwhYd2QZatL1T9Of
a+aR4oHyrZHRsqddO+k=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11520)
`pragma protect data_block
dptqAUtRXzrLfclJecbajy9fn8qVidVcUyVztgVK+jCeLWOWs7alRbFxMTmZO+ZIIFeJHDGaC6Y4
jIgiN0kzuNgOrLMcK7oHgdt5tp/6nNVmir7NujVJEFyY8I9fq0MNlxEqYAxzX3KITpC1XHHC5/rA
a+uFr9z6hfWcQNPRl4QINuyAXJ9G6qUIGFymbrenPi5fuzgEACYhAZcLmGccVlnjydLLb7/3uTQr
Uzh1vxs7KWuTNj/9BlTHGzxZcMWBZbaf7ygWcZw8dJlrPq6iPqtpfrbBefseJUjtnVfR060IXlbV
dbJgkPfXKO9tLEftczNsh3uE7p/V20dsGSDFvq4ClrVCcgPp6EaZvToSE6f2cDz0kst9n9vrtwJK
w5mQoK9l7ntWEPJWca27uPElKidOjlrc5sBSbjsL4BRG6g20SYTwYYDeQmuiNlbvr5xZGn0/9kpu
aex4N6vXLKtVeX46f35FUzly6mpjgCYXOcbAD5CASvGcPPG44UavPkKnD7m2ayRfW+ZgBzInEf2z
aF60BLgfOREI60ZFdBkI8oh1H/hHeKu8v2kInn78VWAD/nixywm3UDZBxt8RJQDmvcx2WMWws/gU
/xQVvs4H3PZOppUY1E/6EcxrI36R5mUaTjnvQWBX4go7jNIL5GgOvLEJjr6LQmoYKcubUdddlpCU
uT/0I5OAoYwYw2nWv/OnmvktSJ+3yk0C42AQmBB7q/ji3Jvjtn9cFG1OvH4mSr7osKU7hSCGWSCo
C1jU98U76k/2E/L7OKgy2OAJhSnjFe1qWIBD9zjAK3UsezJahpsisq96rn+/q1OpT0pnHkdnRpe9
LSg7cGLzgm/xf6DtEE3Ouq9/cDQZB7JWYxuqxkBTBkyI4yIwXhvuR6EKA4C2Sy9q7m44FAmTukPT
Svt7RNT8qsFysDd54cuP+eUmnQQ1+K17Zznd50AbJhNnKjE5FuzOHsEvT0dhRJ4kSsdEkL/PcROI
O+JstzQXr6DDocH8TqHiqaYh/dISnIq6tYRPZP8Fc5t0pK0XgVvoWAXPYs+D667Atf+Hco/iF9Zg
30INKkoWkxSLXqE6trlWlMj9oBMocIpMuCi+FbiiXu4Ur1KyZDUuMX9bWxrkL3TOlUG98vPTf/7U
pxFRnzG7G8Ikab5QXa32+lijxthC8Vkk9dI04FidYbyD/7TZ2uN5taciXIZsdP3ujxhiRqRCMjDa
f1NuwdjtNP2QTdT+2AW/U6EfIIcpB/PllgAL0hnuQ8ZM3B21XCxWAyxIWVJqMo4YScDYaaa4m020
cJUyGaZ5s7v5Ehjx/h8H+VwMCmYJLxYcJZ9JkXdP8MktHny6kBfEVcICm24IeSVxmiZazpMAItTo
2eCkXOYTTKz+5+omR0YooSh7x3GoxFcMnqe9JlajJUQDeWfSJv8R5RKXVpwZMiUckLj5y4jtdZx1
1CT4Uf2X2C2YSM8cZwuX7TOqSOEAbOvfq8/vpstF24P8K9YlCP6PxemBKbkevJt98VpiCoo+sHUU
7oCkdGVtxOd16tHctrmHeVVEhezqVbddcjr1336N7hmhiF7jQQXshPXFCYekzbcVAc5RZavBAzgE
+gpH5pde0eQCzuSMcHd+jVfN9VLclXxuFjfn10IXcaIT+Tf19lgbrW867gwdZMqL0pLrubI3m60y
FpwXgAqi9s72DeqGW46VDaGnW9KXoi3Ro39ErF3jG1KLx77sLuMb2VqNCw+qQc3ZZcmneWMNzUuD
154XFnVrbYFMXv+gO09GlattSRqzlDQ6bpPLiK6UlD/M7nSb976DGK1wQYaXMxhfUp1Mx9WkUil3
2sJMxRCzxGIggGCNR6ZPXRt5BJMfewp2qnrLAykJ/jZGvzEZeMre3apuw778GIBiKHhYRATTcfcH
ndawQP2SjM14D+UF29YcYIm+DOiEAeqaJB0Iag2LiyLm4gFkjO8wi/mGEvCg0kVQj4dzIz0uJaRs
QPajjbhq2RXjavtDd4LDRrKw5WtKRW8JeTEy7CJ1/EoxW04o0x6PF3prVgYsDXfjLauuBONKj7ra
S2bpDACsGR2Iky+3ATCC83denDQxGaB+aPQ8zR9mG+liHL0YLI9Is2aU2MOvnAAKdCgE1cdsdnKP
IlHBoa+myvLbre7llOI/JQVA2bKFSlUAEnan9FxYr4nDEnvtgjQDpV0b/iIaH04MrgPKuVjnqDuq
mW8wAT5x5IuTCyeVUK8PM8BZPqFn4goBoM7zKvZ1UbiClNWHMtvHYCbgmGu2QVI+6Gyl1GkBcRvU
Vhd0jtJbuke9X20UrSh92Rb+KfgfQpS8Jk/cANLxsxKBiwB18endM4nerkEE/mnKR2Ib+kHP2ZpC
Qj5aNOQrmOqgzawcKIW69TlClwZrfYc27+2Q/FrQmSs5E1iTFLMQE2NtA1Su/I3yPNd0tvhyPt/u
8jXOSJr2X0PYHs+bYTb2VMCpottfCRukG6NyrHuMTnzYbNVQ+fKWXeicpsckiArs5804I8Fa9u95
bxgpwzw8km1iJMFF8M0ac7L57/yjNL8JureYVnp7VIwqDmqEyVSm1tMh9NVKE+BMYcTCmUte6XuL
43ZjtO2oCi43oNrI+dwkNz8k6kExwptAdS45HSoXBsQBDyYo5+MSy4Q4p4ReBotJKUqf55g5daaY
hKUr1oSCeeOwG2FelxldQKBEFk7xQ5mFlP3Ocol6ikC9fbVz2TknnqvjpxAqTnbbKZurpIKpxSbS
iFZndyYaym4+kPYXteWCm9OJUgL0g+Lt1+16wthkcH7DzK8x7L+WBsl1OnnhW1SG410Zw2oQAS7J
1Cju3LS57BsuBHARnrajLzgmsBFNVDK6wE9of+jFdZ3THJMhz2RhVVNIpwPNXfjvwfn5HKsdmVap
TYqaTI6rwQULSYt+Y2YpfmuFrxtkWb7ss+pgyX1khw4gc/EWT3lnQVBlpWtuQRsClUb32c8icW4+
MoY0goPfopC5XDpbijKAbNKHNh+lWDpLAkG3YUdAo6Sg7k9Ox9po2X/S6hotIMBmKaePq5KP0aMn
u3YTT9mz8J37aLYnYiOEA5TaBhyJESErXjHgqc7GUy165f5PuEA7fckdDI385cnvo3CCh6+DAr2R
OThv322mqgDb5MNDWD32MdUNiGMhmSE8+9bn82w6bzEmjUjn8sQXSq3F8j7q8QN3SQ8f1tIGmIUR
qErcD60m/abcjvbB2psOZy9xG0P47X2YZfODPhUp2ldGlSuSFTu/L1lv++X+6jrkGBy08BZ7ZoYl
fhG2eS/w/v+dg61MY5PxS0+Ynky5uu8e4DC2AvQ+WsdCBp+4VLnuwRvTuY5U6iUpdfiTXeWnQFqG
It3GWP9lHDsg4QZmVJs8RR3/01GEeIRCEJpdq9ewmX6UPEV3BbdKEzdRqPUJDCqIWc0jcKb+TOs4
+joXSrGdk2ND/kHZZdzqZzj9AZve7w+iZ5OcbykuhZly6wmtfDHm4ZfNfWPvZ7yULYyHmPZrdlja
5p5tOwMuU2KDZJfqZk18/HUy5nFedqL9l6Syqlqm2fjBixgumToJUErcZjLf/lq3G1FBWlkwJdbD
KQIhvquWaJ8GQ0+3zZFxpFocj6enUA30mp/lk87j+M/1l2NyJTyQx753moLOKqslma2haFr8o69x
xi3KjnxZMi/w+hLjXHp4N4Ev3rIKbY1aPIoU2V9RbYP1UIK/Ogtt4lwM+CH7MBi+6rjqPt3PxUWW
+mpo4HHx0vGUGdtNmq2bTDdBhta6i7sxmCTLNq3LrJzvBytvZdKp9/mLYJmdUDr2KOFK+PrdP8hQ
HMnPS+/i8UoFaynRgYYWgo+LNYdH59XsvlEnNUZgpHkrBjVhRqhGbjGUbf+rAHLMegx79C2hRPDM
Vud+2AQvPakHIUuLUndBQrh6GfwS+Cd18BNN2co5gQE3L8mLulP31CydXd3FF74Rl3qYnHHHK+ks
TeJMq2KYTzL8NEX9iUP9tZ+K9+Xjz7TxaLZ6Wqbg6eEL1NT3/hNfcqElNNDR/vB61lF2NafCwTpV
KplsfSY7ljEzEYf9Vp+tltY1eSf7Zjjvf7y3nxvJLknBYrJundYQbHBJhqGAnnLAUc2N6bwMdF3b
hup5ThXSdFBI9JQRjMErz/Wisd0Ox3MRCzROxY8Yt23o+pOYNlsQ9hAfalC3Bz9v9V1QTZI9VGIA
9CPo84q4O+RrEJPnDG+BtuG1qi/LDALjhEv4Jb+VKSxylovxt9hGuumZYIznuC5KUZmYvx1Rptd8
PtsNF98VigMtYUo26jptqZDq+aSt3Lu/gcMLOYhb3h1SJAicISdMhXD8xeGzZq8pBRXCHhm7XLZs
rEkgCtDlLYOseygiVveVim+aKopXePOzGzlrYVROlkTtl/g1Utr1DxCl2EzBTMXgp4ZeAX+162f3
s9lzy/0z82K9ekLBKL7jCIrbcHVZYfzMVWSVeyX2PpTLWOPKqYRij5NxABxx2LkPoqIIy1sPt6zO
TQiCVEMP7T+rJTayBbw67D7Q8md35z1dboSKPJIRbUH25M0RNQOEO0um0bj3wmPo2bWLBYljVnVj
zTa3dAm0SRgJcL/Ho9Cs9zC0tp8Q5+U6okU2QhRanLI/572O9QOVvCIB6JUoejxuduRlZzGRwxUc
RfH1NEqBMae2DgauaY7tRZPwEQ1LYk/QVXhof/kgRDdOg4o8pjJiuuZfTWFfR5hKVpRJ1GgGajnL
t77EPmnsrdHW2MT3+TyAJdDJKoSXZ28z2a/cBEt31aQ1daOgNzV9JvzLO4UFzrm3VjBHozsNT+Tn
rEoX266WELrPGCYGgnlB8TiYo+EIgYpGZFReZDSiaqLwIOsmhcjfMiw+c/4j2PxxcTCH5oUgpAAp
ubKPaeQmVZXyFqmaKkVuafiS62pAuwQ0x7C5RWWE7TY0ZACaDoxKY4pwPLUAEzSBBrRt1Kw/6mte
SNZrg2fjc/pAAbrL6incUufTloUYkZ8PEJ8CDuZwGSmV1oNWK144SrgagkaRTLEpMncbY9bG5Ina
PL79LONuHjLOMFvGHZzIUD3nxr1zxFPay7s77lrKb73j2NOjjkrD1ej6ppYVtLrllkAqMNtVyWBz
gKxyvDPX18grsvxwazjvAWuYQgMrtq6wpCf7xoYWtJy7Elmpa6oaWMgEkQQHGuzj0CRyzqeAVNyz
W9svpD8djlrYZ87V/486Ke1Xhzzq9NPMpf+gSiW/6holJduBlZFtIz+BqH/+kczJCs5Lsiedqwea
8FR+NT+8I7WjeGZvfipLQxJFMm1Qm2W+5rAkJChey8ZkZIxF2YIJUrQienBA8X5HPCa2nV97m0VA
B5I2Orj6svd9CZedafxREf+1FBQ/VQ9sJsUal9/7jqPkyElNfRgNBBo12UeCei44vZcfSEi0iFwk
IeqISu+4gRaV9lCh3PJEt/cI49g3LQdHfkO/LSErQwLV8SwXowU2DNHbiFLJVMFtm82HG9K19TaB
62htcMipoAqvayiCEVAE1mLbLKOf1qeHAMJM7EX3HekfoJTqbL4VcuvT/zMrWXgdqeb2Pb6naypj
Dye2acHYvpDfCCxubdRJ+ZqHBb3FtcnUZg7z9o3DfWE6D9oQYruvkJTO1P8Jb7RteXK2GF45/A2h
z4RK9X1gBEdWqxCSZwIaLjfmCahur2DbOGLkrQ9dXmpXo2uTrK244vbQMI5fzN7isAMy/AGGcOAs
HyB2t6KesLUmMVUxud2XG64LxIoitlTJBKKTUcB9gAkiqFna4ZwxdKuREqRJn45iLpOLk1XqpqNm
UE956CFPWiJmS+bwPvKcUKWuXabx1cZKR/4KdS+XlaOp9uGBOqVsAvacWi47b4h6mgtg4Lz5SlBm
LohL9GsLUEQFZec0PiClz3sLXMqCaIMptygjHxeUZEixz1BNAjMkXafg1Rw/DZMXD5+SCFkZ7Gnk
jTdFXYRbPJMPmhazNC6EqUa038vcXDKaqdk3vA+tqyAnfB61o9PNkFFk/6a3OKPp+Iz3TYRfMLhD
qXrZRhqLfgPa3uDxPsL2wMrLxKTrmiriTT+wCvOIsHXPanuR/kxpKLn775Aow4OCAJICTci6gvGd
tbJMyKyYuRGSKnCrkYEqT3rYbugxKwO68lHsh272d+VFcO5x22CDZDpX/DEXMK485jxeM96WXibs
Ul3rfxptueGxv04yR3OXZIcQYP484SpmutaphW9gQUxA0/c0wgN7WxKcJEQDgti4H/6ThYokLJcB
QU1u/vLyREVZ21ZClgGbe4afsZOCAwXq7lIjJzZ4caskUc+nwDAkcfI6gsSBmO2sZ+axkyVHwzr7
qwRLWak97Il1/lazbff66bQjorDBTsVSg1M9NU3zrJmwF/m1yLxsBFUw9cyKNnerxNDZ4xqqsVQa
GpHriWMWZMtcCMPn252JF60hY7cRRWu1nfgrpj+ZqQozcbl4gBDV8BCCPHfMYAv0IECcjQPGTWld
IsZPZc6uy+t85mFozmXPjKmlNiw/tFaeeIWM9IpXFdZbFSV6ZQrKzvNWi46b+aO9KtUYx7rgFhqN
q/Fibfo6LG9kGN2GtmIEO09MC+e4/52Z8BW+hTXAwvYujTfvB/OpA6gDtTxJynSAXjDRX/GOJwEQ
lo0jmgqB9RHhZqVcq/vIG+Hs6MgD47Xtqwiaxb211ar6uMqzGrnzzt3zGHfKWh7irGIG7yCOIrfb
vUZj3K4m6bMlbdwpqhkny+Fg0IW+1hhnrZ1+NJOet2dQR4mM9nh6D9nViMuMD+ns5zYpZyc8tByz
t5AnMYyuKYPDnTAdxst4cWVQ1aQ4lwuwOorbQ6FdUkZ0+SYrWcm3KMgFR0se9kN7pjnoffVksNPn
oRem4R8D3WQtLv8jgdFCMMPEWWlKxERkM9dpSvFWghc6eX8MoLeDJaoRuaqWOcw4jGzE3FpAVCbw
2bBq8zxoSp6jJHrkzCroFPxdo/7ythYevlGgGsWRVayuf7WCfdwxnqZ5xyphqH8VlKXWpBCnapT5
QWDrn7U8HHRyV/IK0+WYQtObqwFFcm6QRkvF5fqFPKsdaZCITrg6UzFMlV67JwkMs4lp2DuQBbBc
Cg5jfH7zkFg7TkleaPZ0YWyeQKgpOvnvVxam8jZvGNjPCz0ohy5/H2WQWh2g9/1REhQc44GEfSYm
2bRUnhbIW6psF5104VE8DHH7xfLAxetkxMaKNw2l8MtqMn54Mor2l5kXlYhR0Hqtpp5GKV7P6XXz
flXC5pq1Ehii8+5xMcThklo9k4wNcju3x6imy2FYMJCI8GBYqBeMrMd9g+i+hoeBV+bBtLzAT3yZ
0sQ01Ncc2Nvc6joKiJR7Zjj0oveI3URwNfXHcuBiHN4us/ViHIodQJUwYPZbc4tigVzmyeV+tEtD
zs2x5891WCRqxwk8RQCck91/mzfmUVjuBFpieERBi6E6EF97/PfLdBODg5dxrdTX1/t3dvapaoJG
/mDMVTpriGM10hAht2bCeeB86/uLvCmdC9/Dhi95TCphg7oVeg+gZQVKuijLTmSbuJFmon5W01St
ISagi5u/EcPFhVT423h6Xxmm7TSowW+viP7YnuZ9UhCynV2d4UGC4FvGS/mbUv/RI1qP/nkHZW/I
JqFOjw4/DFhzyyhImNfURMRToZU8y5OEGHrR5tpw5wUeEZkXAY7WQWsVBwc89RAjMto8rFVJ2p/L
FC64SG9BT6/uq/zoNeUMKWDGNaZdFYDItxkL1vmYWzc0c7n+bTKLcHSVrz64mYyDYiQ1Ufj1W29U
RkyZUyJ8eZIHh6Ea27jvE5LJaJYyHzbFKzlm7n/r3Bscz7wKvA+PWpJYHZhrI8KTnVHCAhS2XO+8
wO6jL7nRp3jUX9xZFEN4/NIPt1oxcVeYRb1Bpeyh4+l2cqZAW3eQ/CpUr5RqBz1hz7exLB2I9Ryd
GlvLMIKf33nHXM523B4fVEmCOXxLfPAX7f9U42KcKk5ikg1pNM0Sv3jpWhuGTWSSYlZWTTdU3ODb
3x0JLQCsdlLkHgubMC42x/D5F12CVWHFnmQyV5gfC7TI2dqpivqGe+KEoz48iNEvvTNajamY0N98
CiNSNrsLdG63StTB/Wyt1ZIs1yUSpaM5jyZBok8CkUNykPtTO05Y+oFIetWzz7E/4MjQzyhG9YsV
DiaL8ZYBOnd9iBzPIdcPq9L8Ti7C2JsLP/2DFzeGo79o+/YSiWPy01cmNhOrYXqjod1LCAq6EIbl
LngH/AnfEg9BDxNmELESWcCeL5mXBjmQ7VFbrIYqtxCtXJq0c+Nv9L0ev5/tVu7+TuW/lCvonrqW
Nfl18fo2QCLLgPCcLFPXu/F3mxaCYoRA1twsCc7iJyt/zXSH9gVgSu80ah25w+ArLFwaBthBzITx
ILR6d52o2WG80Nbda2ilhZUkQwzaAtYmwN1qJeni2uu0scLil64cySxEPhPenxiCPkWWGY7dG7WG
g35JWOb2Q27zB8/PnHyONR8yjcDXRaeHx8RpKPAsmlOuLb45NVJuUx0iAlynKtoJlBn6rBftsK2D
y/ophyKBWRTLNkHU0SRICDlX7wxBzSY85Syrdt6EycXg5PhAuY9xnF2/bjy4mul3LXEoz5tygaQU
m3YXZeYYAdjDhF5hhPT/MOYrdreewjyE8y+keAm8JHTL05BasdAejZQILDCyrMi5NwOc9N96fBZR
OGw8/cO9NiaWPMyd0+HN+fpVemxB894kjne8KTYy3+TGT1o1ztxi1PC0n5CwOO3RxfrkceVI+UUJ
3w8xP3eWz3pjmgNDyV7xBzNo2FivIqLUfJSD3wRAd1/oXZoN/Eb/Kl13QhRGO1dMZj45I4jmfZmD
lKFKPCwLhktxrnR/CZojbeySBeclq21l00yctSdO2IudjhmRVaqlj5Dv8CtYyOZMRR1lrid63xKf
em6lM45MuM9XvLvq6cYkZxhgbfi6TkevzILVnfkNW/ier1juwxiIPjdqiBXw3tYPxFAKZDzDNrzm
4GwSJFpDew1FAN5cV5IsipEOLI6YV1bNV4Xh4MiF61om6YQ156V6WhXkKPQed57d4VVaJ4uNvEgf
Fy4MhGGsjxgql+3ACUFfYXtpzqQbS4DOBodKPqibWSIvNQuKnXWHomPUu93s6B8Xx1l2HQS6lOPo
AvOhb8rPOv6yT+qhDhWp71fwrqFxnzOsiBKIFE9zUICBrw6phxud++52yigtvVCeaxelbAzrVZqQ
Y1hSPSOe6CT5N3IVbqBjbDVkF+YQAv75PFHIJx9LhL+yGSWqJruPGdrrPu2T5ry08aU/J6S6rK7C
tbcDPAV+8U4rWXXmSAJsjo8CirlfCqTnuSJGqGxsF9XSI6nJg3H0r31XvmwyN6qEJeE0twa9banR
ryScypnxZ8cJkfiNJQ0PMNZAAPiQYV0PJyycZkDzMpA4EJduTW8Xak2cjA5NK7ZNQ7gF6712LD2t
q1esB9hk04tKZOLMdMaz3mWuAoxXml9omPjWEbyn8Y06nEdueG5ES8ws5DBPW4i5xru6mOn94GeP
h+fWWrzpysMq8woX5MuEGl94USE0QTT2iHL3raOpJKJHp4O5QkhQB0/Uf3bTW5mWnwOmgeGPHjdr
YueYMh5T8MoLSvm+c4EVdv+cR55YoeQ5adk4C6Ou7aGZh+/S5VW2EwEbuT5CErOJiSIk8C9JIWYK
/0aGMmhxJo/TEMQwdpE7pLgjInID6i/YcTlLVGaYq0qUIyrF9lSenaCV+vy/5KTDHRhvZ5pWY8/S
lfMzQIoyywpP3QRrj5cqmhdc6O1w7n3t42IBTCHLy1/+5AiZCgMqLJJ1lCl6E0FqPfGH4WLsOobp
ux4goWp2JBvfQqg3ayK8Au3erG807Q1hnekVPvryO37csCFQUMxOkbbYCt2DUs6TapShxG/B5Z/l
ZSFXJP90dcgISN5uK9p2RK023eiGcfN1HPS+D7Ddzw+N7uEBofCTTgOGooadA+blqdslURoqvWO/
nAZjZX2bANXZa6nfq1n0R1Ulcpzh3+RhY30tB7GFaxriMaVZ+uVGUXxawmDPClS+c7Y7yILRTBpR
c3gXQWOKC7yz8hcaqS+QIej3INHWB5JYL2ee/TD7jIRTlFr+G1Z1AOMdrbgrZnjB05M1tr7dtnh4
px5uLIibcn+438PtdPvAKmU3WxEZQ27M2I3E3svCdHsKTeYuA6hnZ08/DnI8i7lO8VihuQW/4UX1
oBpOuO8cM1N14YEDUfNHy+JKiIxVC2aNUGN+xQGKEgfIIi9rJGGQAuraqC+D7P+zpcZWmYqK3SqX
fPh69vsWSPs0vtPVv3BHuFpLlHbIGNUiq3rNoRTmueLs6+gxWNtTsP648ghU+KDEA0oLtfSspdLU
tfFMO3Xg2kJccuPtqsJThpRhVjEDyLQ6SIiWOVSCWGWQ14BbqulMMmWJVa1gVgZfFTBiH9exCJQL
b3U+4UQauYFrEEkFR1os7lL6ir5QoRCvv5QSrPiwKeOjUoULJNGaSwAj8F/FiyLb6ZZSIgeMvDjH
eTgPHGRkyy9YpcES0pjLxviWcUI68Sf+TSWnNHgWtzs08in01BYQAsTESrewWLJ3y1UE65Hrzl7C
YsBgxv4CzAYrez7wVXEwbf1wqbfk5LWGXlzs/uZyyoVUh0oRuUtJb+dXCIwTheEjWVDAPDIjgV5m
kDqoAyMtwSOug0/9I0zXnRU8UMagufBf7Aj3AVsnt1RMGzlYqwbivssVmt6+sMOGGrak44QCikjY
CdNqpVBgsQJN9RxfJdSlO2JpdcZx2R5tMjIia3kZwBbl0+qgxnrq8epG/+8kqNUdl6d4AZ8NoBJa
ib1deYY3Yv35cDoSMRhHiTTFDhleCUa0HOOazwHYOBfJiJ+/dhCt3SYrOtmlAx55NVBwR554zyDr
+hdGltpR7rS3LttCT4y2gE9WKqIT9mz4DC79KS6XgIjlOAG59I56kp9lgFGMV+eKvKbqcO+d9zud
MxybXiXf+OPeVH/mQtl3wk5Jpac+Jnn291E44ho+ULRq0kSHbcWA77RjrOe7xFTPGZW4yMVP2dlO
6+fpb/KSJoFBE78XW5Rx297duDk4eJ+4ASY2DlvGmVO/7ycUxk11QBEcwoWc9+Z1Uf1IbICcxiHB
TWX5Q6ZXPwJiRl5xQaN16JFo3ONvBrL5cVvr5aNKX1iBsG3H2OCjJxz+h+VzMOwzIrPkDC0QMCTu
Xp+CGONmnNuNDeSMzHCYs1s/ucTH1BXsrzO0W2wleqEukSdk9djKCP1LhaIEWR0irQ2lDMQJw7hf
YlOIZxN/eMa8gKiakcF7bbSCdZyPTK42NnxR0WVlQmqG5D1Q5W+UEfH/D4FZh0SCMmz9aLSBjVzW
W2Xe9GGtalmYY02LrD2+Jmd4bSwhZktbskkog1uDr3Rw3mM33nUGa0OgBXWtbOxBjODvuRJPAwKz
JADTouatG3gJv8pPwCNGNU4BsU45OmOIrOZhHgETP4dZOQQUB0c8QZGPyHbq02g6XE83TGwfCeJw
yv9vLRinIgA2uyiEfiB50LXJY2Trn0ELrqN34Vfq7oTi3fdotHJJKDc1OMwX4JtswHfFB2bZX/rQ
/eTQGErwxo4yYnBQc7eStq261nrzkI+PJ4IsZnbx6wxzzdDSKg9m+RJUWB8GX95txI4O+rckdfDS
k81iyRRenaEt2BjSWCEqAWlRejqQsSJBnKLvDceG2OD83m1fSYIIbqpPGRO4Pazz1WJ2YkO3ixdh
6NFO093U8NUAb1lqPzsX+UXgb10jFIDCP54vlX/As3kS2qHeBKse3oXzf156KoF0lM0WijVFvNXk
9h2B42WhCOpwbD4dH9C6UgFf0ZwRGyCnO3gUZJMhIaApHyZJnGlFqK1hb05c2edqqAinnt6N1bJc
OtYhivLt3cekLF/0Htf7aJy2Wr7nnE/34JcyTuw5aXgV596QsnGT+mwwy2kU6PzDjongKgxheLB7
g/Hbj93n5wKhoi/QIl2iREGSRxSSnu3JddVin2qGT0MIKfn8/URCoidy3TxLTOjKOupRepztHFfr
92bdgOm4SBXfFaPVH5rfnaE63w6Ot0Oyr9SJjZnIOA71Yc6LEvUaUee5WV/UktE0jwyLIN7pZchh
p2eBBz2QJFZ7D/0GmoHCVs3aNJh5O0HoQvp4T5ZOEzE8U+jLzX5PrI+mAu3f+gmTO39/Zl3UqDfU
UlStLLf0fV03JJ5oUsYo/TZrhLSKVt2IHeBxSUvJ8Aujpx84z/Rw7dQa63Lh5El3j0jfzw0SWQr6
vRM8LP5OOb6zJEM1OkdT7zH2HhPS7bN7hjRKGCdBleKrEPUVcpXyEDyAYrr+l23ftwsNXpclTjLy
qvU/JvMx5PSA2XgFhsCWQS4unmcARacaNWOMRa4+aiTu8G1SVst57owXruV4hE1JSIkxOt1NdRxY
C5/fHlBVpDBwh4oN/3nBqM02uhgEFl5uMhzxpjXRHNVr0MDxBhNMWNrxXH5PKtGQhGbDl+IaP0+a
6K5TLv4G6/YGraYdRe3hsrfobv7PGXwkLrCVzEMomwOp2FhA2+nxCXXGZ7ngYX2nR+MBf8w0GI6+
n8ErNZI/WKRPKyLIbWaP/7yv+Yeo8Ztsi2PJT5sDmQlgY6ok1B/mWyte6y/cxGQeDNO8O1g2KCG1
UEU/DlxsPzWvrkpKgSct1DTRW/fUF7HWa6ivaMKcgXlr9lEy8JeVWW77doyxJtZqKLMt5PJsupth
SRXhOfMwPjlJOvvA8Ty1yOWPMox1fJn4+CULGEpr2Caj7pmJL+2u9rHFfzf/8B1+J5HokjuzDesv
0ygTERmKOuMKRkUVwoyK4tS0f9HtsPLTVMjdOOksV4x243rvwUv2XeX+4K778d/VoMscqIMPjhdr
JFUt53y6jVZRoiIbxB2i1u+QFoqdd1upf4dgb/d4jjkxq3nI6zHnDEalJjAzG3CA98JJnR9+/lvJ
pEcIWnJPgPqiNygjwx6+Na94p7fJodWR6thKDkDlQwMuyHgij8rw834Fe5u+DwSdqEezNfbYt2yX
JlUiFg3FJs5FulI5rlm+8pM2qz+kqJ9/xjSfLn/mkUh5IOmWmO+Fqssvw69rIzGkltv4bC2OHixU
8YP+P2YmpLS8b0/fmbrlx2JHnLJ04vDF5tgxyV7jWoaXgOwFA8uwJyd+MNRPzgacn0BAK/uGyump
LAFYvGw4pWmlx9+XSdZnMFSn6MkHLaiGymKfAHPQFfpUtTV2tVicFTqENqOCL82i47SlRUfcIPNS
/IurThEedSUYMATAmDIv1t4o8545J8xGNaL45PV4C9iXCu0uFU4cSl1hmFf6mwdbGf8pgOpvvBAb
ZsQ1XLc38i9vDn9s4S9Wijoru8kT7ZnCmZe0LccRwOs8GcI+lZY5IP8KDPruyCBdzNG9OsMfsb5T
wal3DUzIEP74LowU3Hut/KXOHEs4eqmUXEqQjMo3nnuGDIOdXoOojSZAdhIcnZD6jHk0SCS7pD2Z
57BcEQSRfV22t7/BuOTGeYnpamQK8dPGPsayS5WdOV6MPd8NpmiYA1L9KzmHNAs4is8Ep3DPre7I
VL7dzmjaTE1DdQs2P+mzt+sUPBEN7rnfOBwRbvfsjPlplxlj0r0Kman6/WTcHEGSpkyie8DyDgog
wambvQZ7MaS0S8SenaxoPBq+AOPWAGXwePTr1EJWMQRzCO4THYRi1MArU+rTpir/yMtrXvZT60oK
wAjJWtRH89UOZtduXa/tdpJvEcIAX0HdnscE4ofwjjILAQOXCCa92Y8hrtQKdS1I0tsNpQ/NHSMB
HuSmJSd5AWbN+1q8UNt+uIl2fAfLHotUjeboYRlHjOvE1XSoFBoo5BqlzVpULNJqjr5T3vaJEO+c
/RpUNHZ0KFgZxW3TxC5UL94sKfALzX6+x5FEG5mDrxy2fwGGL7ISRcO6Ec3JdQzwMlvbvbYhWwCq
Vc+z0IGJWuwN1+ZLPjLf6R6dGwvWDhcXTJ1AxxITbjme3QjhQolRo9TULTiN4Jo9IjkZA2uYfgXp
jvX7h3Vv810AaaHZbl73pPNlsUM5VNzVhjJ+FEKFmjyy4CHLeHJW0SzmLFyJYiJ/8ruX586tRFC3
Al4lqey0elDPZMnWL5X7bpz8ID1eqGpofVJ+Z2JKt5FRHTrirK3SO10RZ7uVy7hS/tleuMvE/xk6
NDSRuhcGtv7IDlEjc4t+2X2Y9WrAaM3+Q2Zs/MvuEuWizJ9fpy9IC0an6xIrVXOuCH8GHyfWnLUM
9SBR5Ck/jr6FEdRdN/52Zh/WF687NYxNadCrCpDy3esP7EPhBeXgsMGue/yBOrT2NZ5R27wvz7Z/
ARZeSdJ9LMCF2fmFP5elJ40ZahuoEZeu/jGIIZ7VBQ1nNwgREnvaEFzlPobjYGQAoCKMkfMKx01u
XMpQyJGCfV+Z8Zf5WLlSSwwubSRyz9yGiTccOGFStGP+kxgv0MHGT5sCe012B+ut6YwctkFW3tY9
xAbu1f4qT1yqsuv5VHVgGXPP5osYpVXQLTeih1Xlo62h4OSl54fE5RBb/Ezq0Gf+tti3AD6TsAH6
e/QHE+0qhWsNxUh4Xkq/mGcB79Tr4IUNGLMXafgbFZwmHYjFGrvVK6y7P9NLlJuv5pMaVftcFY3Y
nOjM8PRX1hqZJ0UMZFgMGVufsBwKA3MDROcWmSSlTWVx17sC1lUSqnb2N4sPIlyTZo6ugg3Zfd1v
jdW3RILW15/SF7RqstpPUicxmuJrmEzv0Aez6UWds1jzz+O8F+vuVNWlJMD5qtia0mVvH2FBQJau
91v06w36kbSn1iIpgybn8glcH456z6E7V3Ucqi++kChY8+Hf1C1lFtF5ggCSzV+IoUizg+11OrVc
2XLz0ARhRdkWlORqNSCVjMUgbroVzF48eKle88SSeUvAwEBk8AYT6qgrYbPP1o1lQ4XmuvulUBdC
5jFcnDq+m5kX/wxnIHjJW39hc2Z5GJ5m78/tZpw7PO8c3BJU7uOzt8gPg+2D6BKUgNUPNAO1AI2t
nVE3pBAP4OK6hLmLSF5BqwJ4D7jpdVkCfEoXpPegokrlfyLUFeurYTaBx/eDnfoYuk+mFQsCqvEr
CxY641DvhkpcK7qDb7RZZb4JquDfykfm3QWNRbVGg3IDgkMttV0U8PYp2M94991nWooRVxhRDeJD
ktZZhnVl8StA5Ae0n1eyAxprDa1dvy3+eYrgcysQMXb/86ihBsVcucWhnVHTpgXRwzWcyOmq6V1Q
wuGoIUmkc3Zbr+TKnjW9cUbhNM2WkLJ49WAlpA6Qu5L11aBRG4QqaL5OzQCguvylokn93MaI24bW
SHSEUsVbQCfQRkTTYDHEuBv1x27H7nWCGlGEIgWE9d/kujW7lpQiWLV+tdlwnmbwfhSlCakuzBv1
t62kPIWw
`pragma protect end_protected
