// ============================================================================
// Amazon FPGA Hardware Development Kit
//
// Copyright 2024 Amazon.com, Inc. or its affiliates. All Rights Reserved.
//
// Licensed under the Amazon Software License (the "License"). You may not use
// this file except in compliance with the License. A copy of the License is
// located at
//
//    http://aws.amazon.com/asl/
//
// or in the "license" file accompanying this file. This file is distributed on
// an "AS IS" BASIS, WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, express or
// implied. See the License for the specific language governing permissions and
// limitations under the License.
// ============================================================================


`ifndef CL_ID_DEFINES
`define CL_ID_DEFINES

  // This file is required for all CL designs in order to generate the proper manifest file for AFI creation

  // CL_SH_ID0
  // - PCIe Vendor/Device ID Values
  //    31:16: PCIe Device ID
  //    15: 0: PCIe Vendor ID
  //    - A Vendor ID value of 0x8086 is not valid.
  //    - If using a Vendor ID value of 0x1D0F (Amazon) then valid
  //      values for Device ID's are in the range of 0xF000 - 0xF0FF.
  //    - A Vendor/Device ID of 0 (zero) is not valid.
  `define CL_SH_ID0       32'hF010_1D0F

  // CL_SH_ID1
  // - PCIe Subsystem/Subsystem Vendor ID Values
  //    31:16: PCIe Subsystem ID
  //    15: 0: PCIe Subsystem Vendor ID
  // - A PCIe Subsystem/Subsystem Vendor ID of 0 (zero) is not valid
  `define CL_SH_ID1       32'h1D51_FEDC


`endif
