`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
aJzqDB1fzprIDzuflIiv5AxvIWzZTbteP7xwl8wJM3VUkUPU8yRX6OAC/x/S7SOL0ADDAifZe0IR
axltt1Oxav8QyIoloWYIPHnhz0wYia0m2Z+tipoD99zObiH7mAWFmLGRCbzhVpXIp6bpjSt8lN+E
C2Y2GiHRhswSKK/PquVsEcWWUFOzs2reI9fR7YSzL9sDkhV04fZ/v9SFgpD1O97AJqrpyIUZsfTi
K+4t5B2mU3SCAUsMZiI9nu5K+I1q9Usqc1T9v8zMy+c8j4GW0Hf8eoXdzrUHnCtqt1PKc78oTFOb
g2HNQ6EyO9ZnIrOlh0ztafPMfcV0y/SViLOgOw==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
CAKfHbjQ+UvOYLyPsP6I795+j3j2kz5xKDt5SNnsJq53Gphm2ZmEQkNmZky59IYKLAozoafqEqCD
GGkKMgml/xqe8ixIs3BaQur2QbKJ9veU69jhpAYZklY/lTAhggBaWPV8ORsbAW3fp2b+LybUQMhD
VeownLIBf6ccx4x5ENw=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
YZAWdqIkhjaUYnTrXgVTSzMeDt2YFe2CY3vrDyJMtpdFzeYD3FB3pE/RX8QXT/FAK4IR0R6OruH7
HMDPhlCUnMvuvR2q43z7wnDYtfG4XLtkHuS+wtOiBC06gXw5+2iqM86aRjSuptiQ/3pdJRZbk+hJ
SwuzWVO/9TF6ufYtd0k=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3488)
`pragma protect data_block
vcp1Af8EO9OXsxrJyW+jmSmWMcjPD3Q6dLRC5oO8k9giAorbED1CbO2Vi53sTxKKpXlqFbbWVK6K
dq6D7VoFMpSW+5MS+MA7lKxva4pz3VU8xYuHzCQLUGFMxNw4zNyUMHgYP3E6Vry7cehfo2xthFZo
dJJtXIjiW5czMyntAItjR4pBlXMVg48NUOyYUGgVCpFHzDawEXPBcECIVwkRLFeBw7gmMvK2gvbw
/NuMCx2zA9ZFOk5gj9xRcvwvdAgfFkercSozmZm1SaAU+426YiI0HkMSlGaFTYG1qmJqSCSQWj5c
p8gtLwix0inJtbRXb4J6El2kPQrjoj/4X8hCYa7lbXt0ylGEfmKdodkA8zZBfPLu2oq3xHIE/ins
1Y6fJcJUh4hGrqXvRoz+zGa2gJCbTnOyJiD3vt5yn3pBtr2gfh8FwYcpBwGbGn4J2ems+wRoXHoK
c1Hh/8sciQw/PAyKfKdZbC6hde5KcrXqTJAuiWEoSTSox2xgms0hDetMTlwevCf1bpAAmUNQ/v2x
amjazLX4IlqsRAra1z6n34e284XINxHXkouRKHduFQTvZ+3UtmsEDz81tP9vF6ktMeCCOhUXa8Zn
ZTaR06j5x7dtziTTpUTcRTZ6VtytCLdv1UdZp1pXBKFGNIDHu9mpUoE99juzuFSR1Tv+UXhuh5Ey
o2dgXmLf2FE2Gj0TbhZu5EPHAV1Vxlg3PDWACsDYfnoJNHhw8dto49y2uW5VO+BPIZFX5P1DaNx0
2gy20U8sMK8JJIj1JbyFFBoEXz9kLIILrGFXyomiYXaQGK3YRSuGrsYte+oJhRieyPPKA0hE4gsd
C32qhLXf+TW0hiZ8EvXzA+JGGBaRwtAFXuAIPCqJhLSeMdu2ap6glqj6vAe+MowXMh9Zj+rXVeV1
A5hyPvtmChrXqGo0LXC0e1ozuIDUTIcRRk//6HofcY5bUFbXQI1+/7PR4yALojQ0HaNqm4VNIDjx
yC8sFP8NMiT4Blmoq/KG4caR0HE6lPKNsA8hOgYXCpMJQf+yIgD1bKB6PxiFruXtm8peNebCTIWJ
EpANQIYONWQ1Gdf9oeWFRVvPSOc0B8oxTAXplGRCHUsMJo6z+c9vRyvWlcze19cmpI1sT5a7WsRO
OF2ENV0XUAqpIxqSxnwHWcmfgbuw1FaWR0qnVvv8iKofwoA4gFfcRJycFLXpsFmQxjP5lRSIxxqI
X7qRtmNKJWalnW7HvfdLTdy4LvP7v/hmxC+CSdT82wjvWAH3huFnJDlGg36ggwQPUxuxKDCQCcSg
upVAEtw0WvV1FUKCleLmpxugy/xlNi8t/deYp9bVMWunoMtss4oAJn6jET0ti3QLjnnHOwKsNH47
Ux5xjF9gEoAJ0XYak9alxhRfoqKICX3ZHTuyL/0rt+BZQKkhDQulP2rWwfXwMc0OkbsQt+PiR0qH
qgN+OZPkxe5sO+hNk8cQV0rhgllRLsqzH6QkqL01Veq4vOuc5vUMQlxwPKUdBO0r/Kg5fRC74EvB
x+Jk+6RzzOMBUeRVLc2e5jTJ5IcnNA5DBb1srBqxcu8SVsGQwC0Dhbgz0xnn4P+PuYPwZpKZLrpy
iqqARiDMBp+7Gqh80SaulK1qzngnMeiQwVaJYXnQKi5KSsYj+b32CBWGcm6ZJ04DUwY/O053yonI
E5rNRtQZLBxMekVgV8M6OaKLPaEEokKMKye8w+oSapHq7WoqK9+cNANVywe1+Y85r0iH55x6KE1Q
Pl8cDitneGvsiqt/naO2MqFcL5LE9Rpc6cvX5nZXMO5AqdkgLP8/62r6wNa8otAAEiMct3HEOCcz
jrEMb4VfCBWTAvydpcpbij/aPTdNDdx2dc7jOHGa9stnuhH4oV4FBwM3sWXttQGsVqwcGOL/wRHz
jSgati90YweE9WNhIVVbTpqMy2sM9Pfx7qDta5YNSEMD8xjIDm7H+lVi4MxVczBBhkAtePQwR4Wr
RanUANSzcLBtvb3eCuwIjqCtlkakQzHF0sFYDHi8ymvC87qgBlQh7jgFhd1VQRtx5HGfFyq5UdAw
yiYetHWLgSXTX2OJ3OkxHewpAtKw6dC3T/If8PLgtRChLEw7rlLjMJS+xsKIkx0g79feS+1cGow0
7Za8Wt+Nu//a83ZDHrA1IOjNB2w6VE3jPv3FvC0T6mRHZM1AWrcmLsdqHtQf5n62Zbfvr/+fF6b6
hayyuFsLs+pPuHJYKJIuMM+6SBkwmympuquQFt1bzWoI177Zw0YSV6i3L+5rDVgipEaQwJa9K9w3
o6Wn5jH2+0nXg718QQStsyhp+xAcq6pHJBVxiN/sQjSLgxgZ2+VimC2sPB1QUvIaCdKGPSYfJsS5
kOgOt/Y6+UfnJFPERLixmQPPF7Q3ad7l0a7KxgXrvJbc7XRxEj5Z7DubLGGWBb+z/7MAnPJz2KPl
cfdi2/4U70j5sfJbd4bI6Yrd71+02l/zO6GkPZNSVMV6g6curJP2PDLf60bDmKxRh9SIUGs0nZq0
PIWisiicRWFM5RH3NYtr8L4tUvcUEc7LWnjOR4dJcQstz3Yg0joNbNLGjKUy/woFD70eWIzR2HGP
7MRSIpp7dYNxcHZJjCPnZy0aFSY2P5XtAvZuDwLbarCHTaPAFCF80qVDvMywFVCw7Yn0+YxPzvVz
sIgfIs46uU/ZKPN+tIhb/47KQj0KZJTSAqwVXG4mzcDR9rgnAYRm77FDg6uPM5Frh3uh9ctMqTU0
xttdTrho2eb5Qe1ZyZsyByHMs1hjSoLtXV7fzRlLndYfP31dK4OzXmkIqivkMuDG5elSE253iEuq
0hc7+Z4s1tk0Qut8bxJ7IbC48uliUPuKFD5w7unS1FaNbmb410rgSeR788ZoPa2sWhPoSgVgYvN5
ZBONXsNeuiI8nrHjdkeS7AIgO5h/6hM600ZSSbYihln1CTSQFKI6zCkQGCyk/JB8prfUnFrnEpI3
7nWAuvtGVjz9noszc/a1CBgXGUkI1GILnFwoz3PlYYN1w9UePSgeNkbsuZMO9FsUl/4lzaWNMIur
8QLztidH/cZXwOdWHiUIj6mw1LHxo6cpgvnusYLi2/JKYzjAV7cAIZo+YkcbtpwmLZOhuOaWNkJH
1OkD56hZujaON3lZSG1EPRTTMkGKESH3bgl1ChnHn0x+lfYGFiQ0K4c3D/W061Ey15D/qEM0KSDS
KljZYloppDvUHnygjBAFte5BjAYGN7irpiRig37rjaGYbBrFXgQgMXoUfe8tqJfi+ynqybpek3UC
hxpHj3uoVzSh5d8frsQLcUMBjRGAmJSVmGmvIPxuv+oiK1iTRPTjo+qJivhK2Q8c9xLLMA7XXBaO
68EIlMEUDFLragf6gMyFUQIyGIoLU2LC4XusWi6RQ/92VeK5wR1htPpIeLA4blkugdYru26Gd30s
vBy4hZ/phG1YYQzzBsgFN9Qx9EyLOwqOhbyIlRPh1xlwhZ4VxIUuLEJgbnqeNi68q/jlSRwGDg/T
kSlqJODJ0x8RMTuAV0Zqm85zKb3BatNVVmS0MgZS/VHxPgcduYRLMs1ndHco30AI44H3kLhM3+GO
no/GzlOESa+ueCD+UuJZHiKM/aEykDxnF2wg/md/rwLLUwyioHiAkQ2jcaH9P57bdojew2Zd3ZXV
jxe6JFc+nkUtgWV9v+kKmEQxOJcM3IYnYau6mgsI1DXFGkvABfT38OU381Go4h3YkscYjb4iIxnp
Mu/JIs+Ys/yjn4FhSMEufMMh7FXj5ZBNVXgfyUVoHkUy/PeQBTD+afA2jsRdjtmzCsmg8CFnJS4L
1hQl1x00eVgnaZG0CPfb7C5DPvlPFyuwGXvFjwFktSSQEA1V5cqOWE4MohA6lvNTiu345nS6ktm5
NKQK/l2/jNnC67yK+eg8ENqPMuYWkp0a/lW/stZ/x2gmxvUBJxq2+84ERDIVGdWcoZdGTTOy1iYT
Spqt+Lc+nMhwQuS9AoIYMnfe2Kmqsh76oSrtlW6fd4+CUgq1xpD47Rh0Smwo9vrFhVQNjdqFMmv8
Ys5/foBiKWePvgZYQvLN23vyzb2KAQQZWC8RymzVne9kQ1SPsAnvO7KPYkJFgSvXj8QXz3z/4lZU
4PrSed9jAmac4CuWUAbTu0ypKQKygBmsbLvzuSDZdTYFBkcmMO/Iai3K7Hc0ZcY2gszBvaB/PW7t
15Tlm4wbZwRdR+7kDtX74xVAZ/G/GAtljg13Dp0PeM+2AudXxiMOG5GthO+IjWhRSw9TV0ZJXzI9
H/d4XSF7X5Afn984Wnpp9PgUM8IZX8CRGv2aWBhOoETl71/OpdeWizytdQhFawNbxFBtl9NDN3SN
AY665JLKiyODvxAOAepcHGJDHG9z2sdHs56UqJc61GBUporVma0uDLqi+d7K3gyLTx+93mE5xwHM
bgbqzfoprAodniSdcgwCC2idXR1VQ8m2FLLHhV3urmc9bB1LvYJ6AXpxUxUXQ6yr8JjaN8M6RSg6
h3+CDp+Y1aIswslS/lXKkVy+6O9AKyTwoSGOlIEWteajJLxw7tV9iKnLWb+JtJ3hRKA+v2j9hDWp
XGhaBddc8eeQcURQ3qawl6R7Ucyz7WFgmwdCExwb+HmpW1y5JRFNXKUS5NVrhWrYPILtjKvIts47
oGqUflaliXTG4Ak=
`pragma protect end_protected
