`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
ANb2zWjJ2NcmSpRc8TMtVcYwA7BXlywMRXSObmltrpAFxDMyNxq4B9fWjz/08GVZ2v5JgDbUoQcl
CNLiIEdVjf4m+4iNct9x18EkkUOMgI7ttSa8YOMPWwfUqnCuFcA/XcztzwpW5SIThgdzYiL6jn6j
ParH0mI8aRKCuvDKX4PPmtSSXyBFu+IWkLkHwFFru6Iuj5oJ24uMiQ7DC9LEQoZhge6R/KV5LcNs
kcy8tCVib1rIEYq49OYm8S/C+xr2RiUXCokvNNBUPfiVZ+5RZUs3oPB0JTmAa7OKggYRTv9FdbnE
n0xaDJV/viQhC4tgJX6ZSl1ZwNorFbfxNopSjw==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
hY//EbHblwixnRtZF8oEe6d9MQQDegLIN/dRQFrtEsIculLHRjk8JcJSSurTRaC+6Nf2s0xcwmBA
TRnwqdY/1c5KX92kAGYO5EvN1Lppzupy6vOTkiqj2YW76ST5KYWFjWN4AM93i7T4QU6XCHSH6g26
rI1RseD93dhIZzm5d1Q=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
EdDYLf1SEM6M2s3SvEDNmLea1X81d/8ul/hsu2Z3n/9J8NuHlv0RvuZPQTWcbYg0+B1lOCysiYkW
6sa5qpWeNeqZo8ZejtmT+cgJ02xYM7F6yfJ0VsAR8eB62JzoXMLUPiCZ+/mviTMBRY+NDCmCym+U
3iwT8QiUqzDyPergW+Y=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2160)
`pragma protect data_block
sA3Benc2IRHfUBSr0WPyA2e0pdu2W7O0QAibJfHgBCee5dfbEx7Oqv6XjVShdZfI5bGgWdLA3i9O
Lsw/A2rEv+gcT95AHpjpUIjxOCHphcTrRxpVK/qQFzvaefMGfxEnbDjHk+CACfPMUotLXRiUYDAH
7ksYF33R5zjscJ0MHl5MEitkQRMHfyTLOnQmN5Fsyrlm5/BoSOg7jCgJz3E/r5kPyTDJj8vFQEUD
1hncLfzZ975Ue+MuX+jGjHFpZCZR3cLKQYFv1+NTSsuEDnA59iSVtdKhVtfPE+ZbztLqswG81IeJ
3lQc4RWGHoGWHxooWgLT3heHKiBMju0ZsKpur57TyE1yIJ/OIWmF6VGe0DA9DplAYKyrkvlzddrr
2S/+ipdIzXlQt3y8jXcAjNiu60DyIP/AJz6A3MJKbl0+1GSxHtNkgGLskJxMFphcw2kYZLbujf9S
vssYIFPZj5sZnTlsJJkXD6hEkpLvOjpHSiMN03Yx7t2m9toOBP09JLa1sYeCSWtWBQ7tO10PFjGT
Kyl46bVaJakfwwo5amt3P1RoOTOWxgYE+kGC8/AXp2dhOfXmdW5wYo7Ri2P2EdbTWWWok+p6oX+L
GVBfGivWp3mHKAyHDBltGLWKKILunT5sv2ik8utjJoOQMuqc9/F5WIklceIMX7IuIsLtcSSpBg8B
nC0O1yFzv4aOFzbuK2gPwOitqA6hzWGtE6QNT+sKPIenREdW78bD0SGNVizRRUGs6WKPumeFxv2i
ZPDQXdKowNF/fxH2vJ6zYVpf+PEA/LapW/sxf7QylIDHhNw6KcvCfsvua8Zk5fBFTTl/dMr/gAuT
ZoANGiIgQ12UColcqbaBc7lxCtzimUes+b1qn8PBXEcHNdHzsCCbUKAS/8KGkTcRStjwjM3R6K4H
JPwSjQZtu4fy8V0opEwENTRRdgJv+qZC76gDXE6G1Rg+SHk95R+7vUXeU3y/HTeIPzRAsfhBQ8wl
7cT6fu9n413UWf4lrYkl49rQTXPxBcFwNcMs4k5JnYH1I4q3J8OZbQ9DliSFwWE/B/o+NY3A5fsv
TeV4cTEHaNZjrUIyXVzA3T6h0GZqvRB5aEJ/JbpdyEbg32msK6OcB/s4gKJv65BbYmcMntXxoSRn
0M/DfKmjJhdzA/cTg+/lP6TZ7LEDe27hITBrk4H5adJ0IrBDGorBOWSFKf43vVpOxvCaKDYYKsaI
3xz6YHjGg5lsbXzYsc9oCUJ0CLsxIr7PSF3EjkuugvVnxH+eZHg3+/14oT+NflZuZ+XsbI9OmFRn
Z3diLTOlwWNxo5b8g9wHepFeRxPsrfmzxeiktDtn1sNKGPH80K1DwuFFIcDgk3Y0Z6fdgOP19Drs
vXA+YkwEVFgMzMzy3Gzaciq2LZsCes3jd3TEhTPqORPrVfkG6nTUj7dXYme64NSlIMmz/xcjax/k
zPFoa98GhgblbAGJ2uSVvh1DyQ+OAYpew57XYi97RMraGl073bLg+yhA3JJV0xh3UQHsTvKU+0Cs
Sk0tuFbgowqUcciHw5Hh7ACEYYOEmpdzUDkfhIFil6DZOSob+colU2Erhr+28NIOb7BM0y9ilWAv
EIiW6HxW3Lb67DnDJh8WYF7mx0gCyMs+M8NwK2UdRE3uYH5FysZnyRDJWvAcwUI22zH2vEX5RbmK
RFWaWfllgDf5gW1JmECiVn9HszuL3wGe6qbFwEO8k2clSg2enT41Ry6JVyK346xkXtXFZL0uJJWT
S/c1aRZ47ZCDC4yu4/7+rimZjhl1p8lpNOv/1dQwW8H/1A5Tb9NcTxg4x/YoEQ4uYjadrTYlbncw
qEGCVn95h8M36LvhxqMeR3rS7M0ZXX7/JSMWQV2kXBbE6WRoI6DjAYdRm60srA6eAKI4hdf1ILX3
7t4co58KXUXLRE5Ti6Z7FVR5nts3b+B+XagVUi+xUvXJcv8aTJkEhm0c5vBfIrDq9H/YQW5qRaP5
sxEYLXpnNfty+Z7LW6DE7VTVr1Zbz+3Rs18m3dCueWX+279H9OZzYBRtzdOR1+Yh2ue5ENMdLRfh
45nwkrtIYbf4UWWYMNLJ6DiNwQACLVjvG0iDm48KnmbW7tAV+eijYORP65GIKbaix/6609o0D1Zy
J7EOwDmrrNUgQbYqUFwcyGRgTu76pI+fu8/4Eybz8CH8dBoCHy9q/NyBgPkn+HhvWPPWpJfk+KZZ
6nsvVa15z9AXaGPiJN2rt5giKHgtt6+ERe/lr21VQBmnOcS7vnTPvkgaWI2VMlnAS3DUin2QTGDC
DxO+sTLykzyGyJlvzKiVIgXGElgmnnA5qrOGzZokXpc5zj411xIozweqH2BYJC1OkeTHDBjdMHjL
OC4LmRxxsrKbpkVcGcqgR2x3kitRje71Vk9JCQiwCOsib+d/gVAMT+0Oz+D4Pk1aRHVS8BfVczLI
yUvxYSXGegd7bcfd5KtCdGHLuIEMKeJ/HLLG2Y63VCUo7zM0Jz7EYRrmf2bIlqqorWCnvHc/jfi9
nLirAP/T/6YsKVESLkMJXgz8qTyXouxexACuXB0cv5GBv2Usr5+o6F7BJrg4haIZLX/lNXb6d0wx
vp/vA0V2FxmmoR3AwrLd0nmHZQz/EWozJX8qNxNy3LzXh4yk/cXgri7N0strum/ooFYqsaZVXdoS
g1ZxVzoCxsImfNJulmiqQ/2WUvo7x3Dn3zPW6JsOrRAWu8PSfY5Xejlx2D/y9lthFy1bS3DoaNRu
JTVy4QDy4ym/hxWq1Z8AVXjsOm33p4dCXgm0A8FCZZAQMEG8lwDCNV6oZ3AYvdBjF6HMghxNjEFU
zWwaOGXG6mWYYhAnvj3Son9JSh6mOwQk1ALNisO72xyrHDbU0h0ZecBzHB/7swjgCuK2
`pragma protect end_protected
