`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2024.1"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2023_11", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
qM3NLSP5NvsKtk0Lp9uS4aUiJneQOh8vU0nd1efdgzY9Auq61yJTJzcoGHk9G5LUfQomCjNti6tS
f/ARdQcGNdK3PxmJZdFK1Bwvuq8F/HV5CDlgNtL22MBHyZjTQDKo+EmepQ8GcT2BwnER8qj1WllB
bujVyOp/SbuKWJNKv/fL2ZIXoBmPzu6+giEmnERgo+lLkv6IEVcWkbtH2wX4x/vmUordFi9ifcOK
ceZKL7mU2xwVUwIBbD+TCMS7Vl6+Js5Pju4+XEQX7sbhZRjxBv13Z2nHzk0CG1pKiGMgffinCiRz
yJE25S5uYggVkUe1TLAkHFQH2dTuRrfjkLOECg==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
lIlmUpT3kYIhSrLBeok3FIamWg+BbMZFMzejN1VqgpiIFh3OJYn0BQ9yxw0F3iRRMT/EumCueMlJ
2OCJetEjInAYBs+t/hfgwcO4ip8n8ajYApnfZiH2G9QJmG7KoADTV+XYtgeSlkrj3a+udrBu4NTh
I0zVNQLOKss1vb/0MeI=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
RmhhnHFGVPJI7oxx4JJJXWsOz5sVdQ6FYdbWV7AT5D8jYTnhjzsn3i7StIq7sKuXQYBTdCDNsUy1
XXvd/kr/r9VVokUucMJCCZENJ1wPYkmWs981d5QN88mZ9sCMJP6lcww9ES0a7EWz8PVSacaiQ+b/
qkhGc4yYpQBFqFhzemk=

`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
WVTE3eICZATh3yUxe0p8Rck00P/eqNbSoVvpiXthq1LExKR7+CeJnxlSewPJ0vPNSBI86Gmq8anx
6d8E14/owQ==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 81424)
`pragma protect data_block
QT/ODwBDxiL3LUrihg2ldK5hoPa/BPUj+6MUVtW4ie3TWHefSXcwIhat22K5xVMffZrjrEZXekFS
fHnFUiS95OxKfESP5nGHExwc6zVq6D6h800eeVzajVIAJXNYVW6pO2ZFShku1w0eSQzihbrJsNUp
/xuzLTp8YKqMP1Npb4OEO/iaZLvbApFdklhKhhl7WnmCBQRYMXtOX0MGtJygw6cM945SVK0dtPLV
dwI/pfWssH2L7FQGu+Ro5bkPDgLZGn6n5iXhVpDP8tgN1BGAbAnhMy3lldJznv9GFdHlNRTdFPuF
ttSdV8A0bokJDqMTRehT66Fki9hQg6YKcVDengVUoBf9g3nT00HMguJrSp6jbDkwLLVrfv33PaeP
Xobqfoe4LsTm6wMhD+Q5H01tY9xnLdH5MLH+3I79Xl2cEhOntVKt30ppvlvqGGmvthfnocFfVDjb
d15eFkaaNCWuETE8fL4a4/7Mx+ljeUXZYGStAsOjYaMvIGSHN9LK2R/Sie++hIMsv6afQJSIGVM0
FjBA/7KD+KdjT9GTxRRYi79OETTBoPEyrQ5Z9YadPyHVtmKnkmHFuFMhMGsuaS4DT7cfd1TsCGAR
Yl2wYSJ/vbzBEQcpV7nq7tIwpJbiRFRHKTYsZBcIGdN9G2H8NbJrQrQ/iuAiMDhKLByONCUf12ka
l+FCmphaq8hxA4KOsLhlU2cGycBW1DKy7nkBmWekhwaq7VHZ3FXm/r8EjrxjlDLOa1J+ZmPtkyYQ
MJdsSgKnUXvZqBb6l0lWEnAtQhGBF+NNPYfoxXIR1Qv2zSRve81RoC/nzUg2rEnT/G+/bAbGKfoJ
wFiiCS8Yf50tcu7+6JDazY2dtllFYt9JyLUQ1eNs9Nr01HriFxihERZ/HWjYE0O5XjcWQ4ynat4C
s8FF+WeUs7wQEWJdlEr1vF8tFtzhoOfvcXIgqzEMZXTWN/aF/Sz20pjEkHpw92tMyJGPhiA+Zf34
lVsOxiv/cHlSe+SFwncAJ7besPbXpBHqeYV3Jg55ICIqdb4kEsZ5yCmYddjWNsafuTE++83kolPl
o0FBswSH9UDKW8+ND199rryf32nF8GBtgYAppSismQw6srwDZpTSsNxzfMnftGaq7V/KEz/BXgVI
Kl9nCJz5DtQtyvxzoa1cnNTVmio+6QQ1E7DI7CaiZ6H6nWZu6idHOlozIXZpmUdm+DPrk88+TDbP
fmyHpIm8cD93QpNQevhIVcGq0tj6WC6RDvVh4Trwt0p6wlWwsUtcl/v6mINsDyYSgtsKRExbm4RH
CJkiWyQi+60zOQfZGyTHKaO9PzXoOYUIKANRvZ0QPl2FlQD/XJnkD84Ah2uyjwTqRr+lxurvfcXE
sPN8cOASzgjdlPkqcD5ui2SMqa7zbpIYDCME1wtsyJdLkKR+Ca8VxPsjk+uGkmocvuyoBPA4hHGG
xPWZfDjXKiUYB+VFyDKr6Xo8hvtbNCr3kS1qx2IdFu0MK9itO/X3/BSCXA32z4MGuBF77g1nyOta
HUTl0CVfK8HBPLU1JV68vwebFC/bwa1eK8gMZ6i0tfaEkCWHFXRXqBc55lN6ThBD/598ussmQ7Bq
53hN7uzAzkN6y/WQPmKNL8Kh2NnKmrFvzpUNVYPBKTMksnbViIFp4eGaAZ2gpclZHVSC1LthfrAZ
TVLQ3de7mhoC2kM+ExmARlJpej7sT/TKtTUZckBB9TvwOM181ehUSNMwhKgZLWI6cziDIOvK45Zo
XcL/60JxymnBSDcIsTw9yOrz9CN+s9gY+C/LkKEvUXk5oWcwMTp+DYYU8hK69Nc9YuM2eAjIeXKH
SBxeRIigcFlwf9UHVWKjQIlQSO4d5CdFfSQvHa5gtpVnC1JsbvGJJJZZtxCA92uyD9n+QtXXrQht
mWJyCmPK6DtAeZWokDlz5jpUz8MOvH1aFUJ23ZxRBZPh+RriMgFhpwQwT15HULyP/YEmhjlKfmit
wN7GJwbIr0zSjDP1OnWylQLtTNwV5fHbb71wI2G20xnluurLfubSWedZPPt/OShpI4U27SXP8114
TBPDxkl2Si1fZG0A/gazGQXORdYDS7Ok7Kw2/37y/8iOW1eFzO1abmbjCHEzjmuvQYipTmkaHJGE
Z8TLo0WGk75OxpRjvr2QyNEDq2MQ7pmhtqxvcKSjFGsqYZv4KrJa6jBZVKXrebHR3EjPIowo8Mt+
us8WA+VqFYZTkIYIwY9WZRsS1XWlVwilmY+9iPEnhGelM/2KGa1lZ7ldwSVGBGB+FspPk2pHTUby
LjGDqX+OmXMtwtz/mnxaNVtS8/tCGoyU0eFeQXAG83GyglpxzT3Kha/goN92obxw30LzDXoiNasg
IS4zYciz8qISyhcDQuVf/pynvJgq3bOfrOLUTuh4kIEZZUEeospSOn9ysH5+deoeY7+nH6yyBpFF
7CEhT6sJ+XO9hwnJ0bwnG0PGpS1gFsvbW+JKa0im3NNd3LTe650rY9MJWXjsCRXdrwG96ryVzNKg
Anqvp1imNOGzXOqtmjmD83lMs700dVe8PEzuU+vcvb37CBttgEnIXSFSXZM5fHVIfyb3VFM+EAIy
+OZBrYiyuW1QvXqWCr75P5yA6liaJIozFzqPw25aGbz7ZJAJQyp2qn/rfgSew5uEv6eeBRla3JWI
6ctxNsLIJWbokSRqV5dMtJXkGuq+wnOlKBTkjnYtyZXkbYm//RqDpuzfBPKrufhqCuoZoDj5M/cc
EbsNLhlEZB/nB3A5btV/iGDzcMGKuH0vKaJv5qJks17SkCOyyV7ySmuollwW0SlPU8PK9pFA2blN
jALL0Mua2Baz5zRc1UDTSUyCajoLu6OQBEMKQd4C1n/f5ZfGKrQY/cYemxxak+niGH5Cps1Z2AKd
IpLWFbk1GmPAheviYPVthpJGoDU7aXtnZ1grKjfrQbSKB+dKFbI/iMiZxoOUGGfZ+/Ku3x+XxNOJ
f6mNc1Me4LbdUaiCxDObwSPfUCLuuot7fJmghlrbTm+shbc6MP2vDmcPZPnF8MtH083aR4uqW7r+
JwEs67vwIQFAVkgKn01w0Z7txiXOfYHjXbQNP/ULd4jEpTjQr/81xgaeAIk2+ic+VT2HnHKFJISH
jAzxTOjBM54vxCFtk6ECGwZI2kiakv/aZ/p8Zyg9c5uTzO3CCn3424SKW2c3u95AZTz970OlfuCM
gxjZDxYsmmJ88YZKBacmATEdfDSQXAuD3EYEGDp//GFMSUCqSeS1BujGAsUk/sDC6oeiGD+31QZg
FqyfC9GeP5B6usWR5DNEch0YePUfWjOu+pHgrMgOe0EVV15qXV4OlfY3ONe8ZLcAfk+Dzgg9dGTp
MGYk4EIUl0YbPawGXtQDlMzrahFtWOJS3QsneG+ZvhhPJ2fsjUfdLkMtSQ+br0hPjlEAW8lZhTAr
C7uwdgFBeDeabcvdozeXz6FPKG6JufWG2ZxAdx0RQdJj6hA336kRRnwsK1xy61HjNmPdXJjfRowV
rSstXF4F5ciCQPPzxTm2FjwCjh6ADJH4RJWn+Il6+5GiHPfBrvUVdd9JVcRf+KorNuEwfrqe8Rms
rQBsX9Ddzec1nMBxfPtWw9VztbDEoxNsPyWOJ3bknrm/AtEKDAlRTVvYuBnfq1RfhgxdFpj0TD2M
2/I8jkiINBCtubXZLHwnnhTV/NiA0RcQIEIZwthbOgzd1mCmbmEqzKZ37TGmHmk4wSEbkCnRFVHg
efwfPwtTnD16EL9dgAMcrfBZW4hdF9VhguUU12BjmgT7yetqTHXIXTZfPHwnB6cQM549XIc8gcs4
ts4BSvJ+1GxvK6YtFfH5C+jl2H+ctLjccgHeopDnQFKYIkHMG8LxYiSMgYobrFijDOqS+jpEpH0r
qYBes822fm+xvHIqiaLmRbv647xPmtyIz/7VbynXGCc/xMLZ7yKECNDPDjCsf+tIoXFF5YvGs6YB
kaT5py0Kz8rDBc+Rpc1r4ptF/5xn+OpSQdRU511Ay3pWPwDhYxdUO4Sa/bVClnwlWtjdk1qrd1aA
O7l1DhfdwF8/Okh/00MHkRBQy6LkZVJ3Uz/YP8UHHL1K7ts0EKNNirAOWw9UM1ULK2Nfo7D+ra+7
1i6a26dhNOpcKkIqM7prm9Szfd1J2uEp7117uTtquHLeRU+o8j4Y2pewM/nW5UjX8bEC82LxZ3LM
vRjHQBJR764c8JCVUwzs+jFfwNPHw8xEWS2U+SbJReu7JaHtj9xcQkx1z4b6tCWgPubTIRwq6/Aa
Sl6B+mqwj+rU+e+P2MR9yeoG7hAlbYnAZJoZOFX3XYBnwa9BPNWSm/BEXOTzs2SO0z3SNPQJBwgI
E80MELo/JRhI4CUlguTpyB9saMuUv25l4FYKn8fhjtMuxK15uQCrYhR9DDiIVLNOvHZ2dtVqbT98
MwsnUItQvVLBGBjLRhKENDhu3IKlye+9VAMV8agqyz6gU3fsb+fqh7CtY7I/1/oh6i8J2E1eaeC1
bbieAYBHQE02/KZaUgBdWSnxNNhYkWZgnCl/K9i/9jvzA4hs0qFR71SWeERcmXb5a+y7VQy+1FHw
MuiVcGvBynYPKT+73nYukyoVY0fS8YbwofaVDB1vxwDlZrgD4BePO6GN6V6Hwu+lL3MvOjBNOEZ5
rymtQmJ7/UFXNocjAi8sG8qhS0ufCPACRiI4U1Lpjfn11ph1T9+c7CPzRTGdWhdX8iORMgxdUyDP
CHszYO4XNJifD9DkyLbphPfqPHtYPfoI+jfO2oK24m/hnck5KvXnVcbIgihPxa4mTS2uEASeOrrg
aBz/Gx2Mj1cjY54pNycTVEl4BorcYSGbMTHfJYb8d9kF14Oa6SZNcH9JpmpYnYdVcITy1vVpcbNp
/1czBKeL3d2l5f5WwrEwUffnM8pELyw0keFn9JYJIkdPYMr4yXvj8aBVspWRiMrbFTIL14ZAGgZ0
fU3zePaJT8+mVSNFSRuAiyWHOHFmaBuPOLcOd+PyRu39E6nG8maGg4rmSrONz/y31h91796088ow
knsku6vsJJ1MX2IYzjgJKTeWV8aA6736Ujzw01gVh85ugL1J4a+7uhowBL4egRI80r7zilzwLn2/
aLPfCHUsYpRH8eGyUJA1UVSJfUZGTgW/IJoKxhtmtrBwX6e1viluXOrhOUnpq1/CPIIiTz0Husji
WVHA3fKYdUsioGEcUbvq6VXbAFhw+3CKITBe6WPKT/tmpEoYhAWXH4PD8m5F3K8m0GXkXbFPQrL7
VKPlVD4Cv2D7SYIvxaYruYKrhdwCyIsTewVsIJ2mcer+4S7cBHvyuWsccytL69UFfrkiLomE8K4y
kUxJI3np3yLrOUhaZGg/T/26iuIwH741RUp+1kKsZBzn7DMNLUkLr1J7KJxesnzGpjYi7k0A1jR7
W9FJ96BK8SFJzAskZqPcajN8v7BenFXuhF5tGclyZYYEfE3hdJ6rmb86JILhDcac8JWTXq7oqejJ
kcp4hNiTfJrguc/pKnc3sibAwH3M9ogdyxdeJW7J438jHGLZpYVVvFtXRLdx5Yju92GeLM6zehS3
LaW/JqVsWvKRdKOLqTJvY6vPdsHIiO/IkUG43uPIvY1Y8G1NsETQtxW5EhlKr+dKnYzctf/DxQFT
wuGaWXrJ2usjXSN4y5+UXEEzKDzt5TusxBnLn42THfass7QBZUzI9av9IS7q3jJjnL4EUmtRxOdc
QY35zbH2TkxOzXbJ1y701orZ8i8qN3KmLvviXEh3mreA1sNoYpctXDVzavQd8Yd+Z3y3AsKqC6fP
Zj6zR3w3RVIU4MwbDEVYE6p9Z2aGoWCqjSDM/h/yKoRoXRqyj1PilPu2NDuET1GNT1/nSKGWpEns
fuLO5BsUCF/ywAvbJP6w2uMS0hpy2mcQL1Ow09caMXr3RyxuZIKf38/o1X/FILao3huE4iwbETBp
gRjDKLVxoLVYJBtAMZkZrt/0jRiJ71vJWdK5Ec+BpDeDxFPoTD161vzF0t5zqJTBf4K1HIHyyWuk
Gu1nYRmBn7GVWuXExbNcwVoqi7hAoFkmPZ4z2kjGi5va2z+9XsEqdRooyWwffnt74VgtyzCVq37w
enEEiKWuXni4dQ42GNxh0edglTjt1V1eAfu75VSasMnpIpTow8E2K3yoLaioROptb2TUd+qaBYa9
u71eAYQGNrz4hAk96a13HYUp9FaJjlZrmaN1PW9gcmZFjDEPyeenANawjezaQXcjkax8ONHtwxzJ
NRqvxn3rtllIuDL6uVB6DPxmb91rVwf8dzhMvS7n5f8saFjNfnO1NV+GcyXdbdZQ4YzSvisVRcOZ
aR2SUynGOpx3b4Si/k9aVkNAU4occIYIh9rzufkdtNZWueGXfwgWLN6u4tRdDTDqrGLz1/Mu77KW
Y1n7bBEtPTYG1ZQtY6n6jMJaHtApS3ctnRchp/A+0LPxTbM8/ISUprROsWqe+DAhwylAsCW6uWCJ
UXOq2XOVnee/VenSgp3S2EKXGfrYT6MepF0qVfxvr2zd6U/AHZAwklABx8zVVfsbOuBlWRzM0wDC
HOWnaL192YrZIT46LMvn/oXQsMgrKwcC0D0mUOIeQZh3sC+ILTTGeGA2n2oTuCoL9Yuc8trKeJz/
1w82zfC3U3VjU4MjYvXphlm2CO+8v38vUZ7AtLk5hZFWPH/MrzK+yYUXpBITLYEcxtkAqB9hUgIv
bZTv7Cqydilb3JceL1xGD3P0V+CFJqrGRoOEvYzXS0XtHGfHLnGLQclGjZ1R0OODZS0CWZvBwI5A
GklmnaEEa7XOYc1dw98f35s6NdVmeEyhsNr2PadmliNpL57yyabsYN52IU8oZbdgw7HRnwsEj8yJ
Cii1yusEZWO2vc+9wdEyDjNOSBoYFRa890ta94U255JLARvZUXTyXk+abPtT7Hqpy8Njmk0RzdPy
F4fKvXL0oOzpgDLZf5AMoskNhuXOmnpBNoOf56ntRt5SAOEGGxpalQ9KOepJbRPHl1EgzYdQpy05
eXiDZ+WXojkFWjJ97ATeURnh0kzo8Z+nj70WUTK9nzvsqMq9B9SwlTyH9sp4aAqSVrR89e/sA+aQ
Zmi6cEEDoYe29XbNc8eETL8QezwWfYMOMLUEMd0ddbJfnP9P1zf6HQ7JYExrRAGR3rAvapBcb5Kv
jieK7R7g0kheARUB5XPFLVJECSLy6psbyC9sC7G6e0kPnOy6P+wNLDanqScd0ptMGpTP8mSEmBMC
f4evP2dsXx3ZG/du2/AGdzdLnk8VC5Ygl6zFQ5TCdGZEpPs8jL9+qlSFVp++4n3AU/95WzRkYPhH
hJTJyRbrkSROkLcb0MXGjj1/rAf373l5FPx0/YdzEgF8aIdlMgqdqtaJ9azJmhUuFmX8ISNy0Jcw
iLdIraTrNBE8zKFucOJeQAO9+MvgNugjkYoQyfur3aScEhVI8nAkXU/YTtnPrLNAsR7vKO4RN+zi
RTQ67fTeKrjSuUypdrA810k0nd4TfFyvOS4Uwo5IkuN3O+P+3zdmdbz5e4Mnwhoy0y6wR1F18WLN
aacXlOO07troI0iYd3NvjrcjDzk39Xd6y1b+3hhnIMat6U2ciNbAMxyddUBLgpNZlIYXWZZ5DkYc
MJzNIo4Mlb7bzFYHhp8SdpoUeOE4PkwUTmrqsoJDrJROo1YB9SqL6C4kD7eOUpDauKg4amwSV6tK
7DpaLIeXqW1trV6uV0LrqevBCw4hT9twrE80ifgvfEvZ92we5Xrma8Z601IQ4XMCCsEmQq8jHBH1
cvnOYdDrDmn7lxUSVrHyZTyh7CHNxLzgXb0DIildoJ1LiNur1yC6d5gt1/9PQIQnIxKKQiNrLli1
CxuoSzSX9PuaSMcpJa4uw9Hc2G+r6zFHlZcHiQkdy6jtfAf5uW+b0lL9vFU4v6GzqI6FiPiwN5VM
gDpgENbEGCw3ybSFAAVWjKJlhe5zF/Bswmx0uTAKSJtVT6JZnjJ1w34r57tzgcgZyfqnT0XvJDzU
UWIwNGLaboZmvIYtRqFQ/XWeQGZX0nctFoxfAp+K2LnL1jU7BNDfkk5933mLzUpzK06ZHRa63V/4
Zc1eJsxqN1PokD23ysKn5S622WV6w2fT+hymMJNhYQ5Za77iFHBT4BBCUVlMxP4e+sBskDlVFsHR
yYKsfznCwjl0nz1B02kfPoAM9F8l2lOl3MO0CVUrco2UOMVAqAH/U1InA15x3hsD/zk8OP/7+3Vz
5xoeuWexYIBnm5WdHWg8k1yH8BqEuy1zz2D6uF0qCK+L3AXRfPMMMVsxHmLJ4pbfsjxNZBy/CFJ8
EQhuRJc45Y8lO20iiLC0rUGQ47RiVy2+kGYKa/LhzyohfEe+gO1GGzFFXctr9H0ISQOCgOp62Ftn
ht+5tYfhcgdyRlU6zZ0Lst1cJgmUXeowuYK5TwPNqprjcd3G34sd71eScHtomBOxZzSmuhF5yXhi
ZfzT3wpWV+WDFFioAlLn1+CehmvDqnhpD27StMpPoZiiERKec4U/SHYL+HXy+j88kqETuHHatm9f
bkJhUaFELHOAkzRripE5YMuXyPF9sVMhfUBiDbizVg+uaV3Hi8qDUe1+ScdNBX8NOM/1cJGexIcE
UXKu1euawe2JwYJBgTm1sW+UwN/YZCWmW1Ak2phj5uxcHb9M2HK9qTQyNQw4eLblHPRbexJNeAi8
PsgMqCL1ch5RD2XMK20e9dp8BuEGPiaWzMnupWHgWp4ap3KIdQzO6xBImXm4bi/3PDuJ/eB/vDnq
H3EdqKF1C/t7+eR7+cAoUVo68L2KSCoCtU26njnUVvXJAMJ9WodsUby4HApcwWLkT4jaG7PygdsE
ozXvO489xss7JnEOSRKTT6nuywNbWSXzOY8dPelxcLhccjqWZ0sdXv14RkQV5vbKkmLbI5Wp8Tel
gjAfnY6/8qm76ZZhG3oxS/sTBTw2TTGQTvZwxJ5LjfkRer6+84jJlLZhMHnMJSSM/PwufCOmKz1X
2yU2jT/OCu4b5Y7v4vk3dpx+DQmJQJ3dM2JGPkt6Su9CHOgkwZV2EKHoggGBqcKg/8Rch76CyWMu
ZIfyaJkzgZRReG8cGHyYO1fRNZmV92CNJfT1eA8Ih0jUSZTdtIdVnsajA2A8qOq6HM3Bq1qn1sTA
QSAcYQfGxBZ4G1Rg8E4WxBp4s3w4lzegJtsWuXdflYwQbFgG0PqN12nc9pVGGEtAX11zPSSKb0b+
S+OKO+Xf/5Bg1Bl7QNIvyEB+oMkqXjlz6ZcLyPGouveITsd69e9rkat1HKW/MoIEnPuCK6S9Krpz
P4f3adR4NBs+85rJI2b90imc2jZ8lT0Pb4Ea7gMDThLymuHUkvaMXhb5flmhBLo43fdAxGL6D35Y
E7KVi0B+zIFa/YS3Sra4DfUU5s02S5F8UgeG+pWAFTVA8NuWpIYHenwKW1kNlNAG4PMJkx24+E34
HcGdA4EYujiWphN4+1fDdCMdRtTt3OT8fR+OAy3fb+B/X9nC4lftLcfC4MRPQvGU32/8V2cE+a6I
JMhp/abLvl7eHNoINEKzhOw0foSmHH7/4lJxtYS8XluTopVvH2UAyGKEXECO6GpsqB+FYDjC6mIi
q4KKitV8tLdPtTLs9dhCDSoXGkd8jcmLHKKHhE9NY36srn+Vlm86a7la6ck6xTKyg74vNWIh9VdZ
ZIN5517KWO3+f9xDDyiZnftclYf+ysPlS8jMf8Zda42tzG9g8v6GsunfBQOQHQnoYPFzE5AzxKgQ
6r2iqOVNsiY5SZfdRxLv9d1LwtJdIabtzS1AucvA/xxzEewVOsFhi0WtSXCI1y/XS+xxtXVkdKip
ctvV0y1WvXPX5Uy2Jfb86TFJ32vZrGh6sk4+0KEYwfvuLdEk/VAm1+UKVAs+RdvzkkBwBmsQPeev
k3iRGFVo4GayxJRoeTC/wTLhw5p6/Ju5HEz1iveqktO4N6+LxYKMV09b2fBVERn47JtYwMwMc4uX
LDNu1xAFTFH0qFl7VstO8ZGDIdc6UCAFolv+qPW09dVZKF4yTZ1gPVLtAg+gfi5LSTsJOS+JvwdB
uZC4S0CGnGp2VXDgNGOEnjUmIyiCQeo0kXTCZVej9ZTg3Q75aW7AwMnN35H1TdWcMMs0qi9mCjmQ
MeSuXhM5fvLBUF/GaU2FAc69wNe7N8QT7KtAhF5KMuUXKa7fFn3hRtMRgu/QBMlDLNXnPMHEeDmH
E6KriA9eZ8dYYPJbZJ03dq3/S5p3Ayd0M79LiEKLqivPnUkYO6tc3C0r6OIFCd/uLG9D6lFFmyyB
lWHJIc7YoKxwYBpaaeBEer21OuKK1wPhlDjOmRcFzTelFZVo11p+OJgrJn4bKtSgJdA9EhnnInMN
rgcBiyyqhJzQSuAocCrmVJsJ4yTV79Czc/tYrHjMfasmIBENbse6hatzxxkgIynksFNBl3MVevgb
vlIxwXxYeH/8Kx50b/RaEeWa3OXNCA5zx6SgleRHBrwx3Bjo4G3z7vuZPTczNdTMhTfSlO4BUzGX
AkSlrRWyLRR63Q26BT0mnI9/RWMLr3vKwjHOGAiuew1BCz1AFBt2WMj+lS8/KDUsUOE1h0MOd3xW
vx2uyULdH/uWD86QgItiX/V9aAQNAy5fVkFa1Z1hyIzMdI1ACXakmYr4hSuhNUVgZhLI/wdaPaDH
Y/xgJn+mUWiRgFzRMmcTv9l9oLG5r+i9ZuBQH1icWPX9RXr3UB0Qc4aCxLP13dwVhrGr7zTTVQ8j
2GMeo/b0qmQujp2JUYtJMgIhiUC1yapWHOT6JR3cAb0/dIpVKj2scozuwhgq8+UAZy6mlGOCmvJE
+JnChr4K87uwMc4ShThhI2vFRmIk3frlv88hKmrUTHCiDhkzIB9twwvzefZL4E8SW5DNP9MGT7ZW
gEPmdl63lpx8D/i0rMYcuO2x3FGXrlQARtQ9shCnTPb1SzipUlOnxG3l/yiFVidSRsgYznve68wF
m0cgRuWcJ49PsxxpiLAQR+yMLGHgyHBkgJZ/HQ5+JfB4cWkzQt4UrbIOmJJ09w79ha3H0U5D+9Q/
Kw/XcO1FIYDRp3v21pGzMxoh+05co4HU7EoHGoPptTUbc/LMcokv+FtSMHbrTcGoLGV21KPUQtV0
7PdHD5+28RVSvZC7xOvB9uPgwPKv+8eHoSADVGF32qnCKRCB1ymDSgffGr+3rJXTUYzO4GnA1/mI
tpIMZZ7aGCff8c/oAd24zJiyQc08fLJvYNqsUZDXz/mZexmwXunlFIIBo4GT/Ou+P+r5/0vvLjUo
E6nm2/j7DcYJVHJSs4OJkyMzM/Wx4tuUbssHVad/wV2sTwjedWStPEQsdoQbDEcbLSJ2xoApYpu+
ITfJYweGQkKtNXNUe8SjusiYUTFfvvbEMLHwsPD8IiA+ERdqzpvxtXYzKj0lcQYQHvvR9aISxslG
WHN4BzQTSgUBIlmEIk+k7QA2QEwg/hkqA3AqUzXeNe0Diwyg48T2l4hXMUCDXX8mqhIYDOEnHq3U
SLz9cTulWHVVYR5yOX7zJDtahjFxF80a2TRkYeEz4TuBROv8+FNIx71vfUUzIpMtCFTkqJAW8TVa
eOAJoB7xGL2QtGKvtFEu0u8qdLzjOM2rSgR+Fnh0u/TOG+szPjGVWTCg01QBmfsHX2A7LX6BkPMd
elQF7l9JqsEJhSo2YC/g0SKd6ddSEAJEN4yDEeGZibdeTW3lu6ucfUiR6TSPVJiNbMN/+B1XaQqA
x1FoEQrRfaQL8UIc3WQKUjD7ft8ley0N36wiEHRUEK6LnBYEE00OERbQQCUveKp6DjP8BkViKYkD
H303J2barLUWf0sKu2QUmZocMrl0jOBSaeWORYCHfUmwIuFplnvyH7rmHUpyeWQMDeNDe3pYIRJG
NoPv0xE9lWm3EeSG+LTy8SwqOEK8VzGBZamgMS9qhmpQf86cWhVWmNO/Yz0vngvgpY0/Hd04w297
UDFRlXFov1SPGSywf36/eN3ADdb5U9SJb+U1AKGYchvSse+uQqpm5zlPsTxtW2JMowlA5O5axhhg
+ldVXFllG3qXxgY/2+0MkrO2+bJSvzxMIlfNUQqpXrlm6CYdoL7uQdoO043RETsiwa/Rwr794s6d
fjFBdCHI6tfz4USw//j9VFkjS3gNdmKZYgNJU7EwCFnmy8DDu+WKKQHcM04OvTIkMQXDfgD+tjiX
ijwtRSJMNw86a6nEgUHKcDj/C/x7aZi+n7xAV10BKsTristuAmzshvqO2F98hQvQpVtBa1Ohsk2D
QvvsxXVAit55M3/RkVDf+ziqdJOalXS0jAK5IQydCfFxy6DmXHueV/aLX80Y3HM58/zgBt8grnkZ
tWJQoPelhkrAeCr5dPvBPlXPQgIBWdJBq4u3gFonbKvVHdt7marI7q5gXUO9t1cajgDo3JpoP9Qf
Luxtd+9IPMZsmfCcVc1xo+QzptWM5fSwUeyj1Rcp2gOUuIFFf6XPp794dqzBbnVfELPUBxNPAjsn
331XrDo1fbxGVQUQNP94T3Q2xmUXCRGDDKBk6qR/zjhWXh6RremK9mD3lOva7viTz60C8OmITszl
YpJhmV96cxE8lTaupGGQAVdfVPLg38HAUuULalXA0YuPsHOrKh3H+L0ZHXZtmcwOJReD0JuiIKaI
x/AdBq+z6/jApcfNtrwcLPKyy7La+q2d+IJr41TjJjhUZ8vp36vMivB7UqnyuCGxkOzu1Wvg/brM
CZ5agFMmYlPvkbf/Pmm32C1KiguuTeXVrPnA+WPkUvQsSlKue+nVM91ioWW4qCo6vxuvx3QcGCPs
oAn1+zdsvSia+aecAn1ejL8d9V1O+2brr5gQK56Fvz7toMdW6P9jmR+W1FrIOR7jciE1WHCxUQ07
50A07idSpb30hnRh4JXKBHFIEvjk3Ja/hLnf2rUifPfeijy76v4SA9TxYQUWQPFz79XR6/yL+sFm
xOfM35FtYCMKSU9hOZ/rbIAoypLsa2cLsecP9/UWwFqQ/J/ZWjUFc9CxAvBIbJ4A064A/Hf8i5Z4
W5T0OrVzkw16yFNGOXx7S6KkkNHtPpd5k9511sNRNwWwOWiDJH1k6oFqM50H66ixybK6+nmM1Jwt
XKULnQFhlSqK7Z23O2o4IAkJfPE7aCP3qHa2y4HxgXbgvoqDUaYAzUEoBQp+iEu9ELkcQ4p2ZDd1
vwanywNZIZByzRJh2ABq58QTNLjKIrWApL1P+ST/hazE1+C+DPHK7J0zcKLdP/AZRwxovSoRwk77
p5MgNwOf5vchkYlK+hZoKv7HkHAF2Gr8qAKGeuxF3jRlQBtPZX5VIfIAQ6jRVqJpfRqpbhvmsiUb
rakSn3PWzIwcF5rL+tNfCviX2uu/DLWqVE6sLLvyCkmWTefd6aaBz5T0FOhnzNIFHBMd6QEkX+Mg
m1VxhD9Ng4I8I5hv2qSIsh4vXntgYCaNiE1CE9PeWbCVg6t0qS/MsFrMu5ObCLaCyMI/3xrX1H8t
5qnQ4Jth1D6crilqspbmQF0yHt5TEgdbTK+b89iafuJYNGYgVKQ+GBSHYkVgpFj/C7k5fsCgok6U
/4MhXc/wVDOlaPjxMda7DoRp8ylk8vcERiOk2RwbRZ2CoOSoUUZ3sMV2CaGDvvYR9+JVF3BxlfWk
o2HiskGNyBoAzDf9+nijMvJygJiVgXfx/iXpU7u29O+9Lfvq3vtFCI1Mu5LQ+XMev6aS65zzpfg7
0jLDD3N2xJx3T/WDux1rX0HNC2Q0ZeDeHMQFTKuSgegFFK+2ocC7m0Mr3tLH4dD6+yCG3r/oVYNE
bWV/YYeAhBiu/7kDc1b4cx7MzJ4DZueMAot2fj7A9fxiITze6pt4e6qnp/HT2e9fHxAYYag4+aIG
k2r2211lOS5C3UGiesl6bvEcnrkNpZTjHIVBwOZCF4gDdjL8L2B0sRnhPKt5VxI82Q2S9TbqYDYK
MZAPfy6DLRkLbteNXJ/SpJJoePRVjduby/b03Idx/I1YqBbI0DnWd7hFp/wyRU/B6OZCarUxFIWT
3alXOHvxmXJf+xUf0hBeNVpxqxjcfyzERRZU3mrorpsGdUruuh1ztvMlCpdccLv7dBBN+dWSG+t5
mz+8sNlohK5KJGfg12WtGWaWri2drdanCdCfjxnl8r98vfgwdJyOrTuh12/fcP6VJhbnTfUanvM1
yQbSPGjesEMlKyxMvRFPmmIbrrNSjEL5AQZc8CCkmKYaWKcT4Cu2jHosYbyy6zNIO4X3VKeWKkhP
qJgj7AYxAhSLaHEO8+aQbUw5ydtArxI5j6DZYmTX0fQq55acIV+T3vG1CaZeJaa7AD/CqT9Mybbc
97uWgXcC5cJErlhSEelOI00AdoYIWnbqhXTXJaB8yCNsMPvuyalCCCeFH4NQvfDc4s40AD0a0qWf
xbpAh6ofehGNiLO1lrheUxK7M8GgqOV5I/troMlUGA2CzR5uNJnU0xnA1Gz1J43fXtffwL6kZGh7
2AY67QHK/0IbXt0ruCkOfFccTOMylEEZsKhuL6GuA6aMZEDgPByOOFZQyPLEEUCWamQC6nITPTc8
f1w8VBh0ZcVx3uAZAqfXcjMOqaElObQ0xSrdgPA1BByYhwJ0hKb6WAXB1LBTNj+bJe90h1dJxKur
2DKR1cF+1LZIiEs0v0BU0p3TZBt4dSgf1RYqnOaMtgSeweEUe1U/160msoh4W30XSYg/FYCQBTNo
SqGkXuxleZWuWHPvrZsFixk/+qnTjtgxiqKXJDWL/4vVBzUpc6N6OKORoIwvJoCZgnGOjxDt+3XA
CX9diG2c952Gee4A3wNhDtg72djP01mXc+pQUubZHPlX0tKPKLI3FQdi9XTRyEYhEcSMt1rBtvCU
Cq1ksHzywJnnnqnEMOZEcdpPSIEWgkS0I5U+pntOgkacDebD8aGVXbXC57ygyp0Oty7ljoY44Zv5
rsHY/UOlwsW6a1vxCWJU12r217kIiIWDHHZCUp4KshM4G4i2SxKi8dYTVRatl2LibKjbjT8qoU4U
GqQR68+2AwbT+GsuxyLOLP22b1py0hZuzmf7U7jOPcAv083X7Ym+O4t6vKZ3vQLFaAdzV9Zpwsj2
/JmcJIQf3TaG+shq+nu3zx5ZBpKZtS0eKRxwqyb7rVSV8653A6L1B4SzXikMOHUUm97qms3lbYGe
kUYdL/FXf3GYfefzwlf+yscG7EpNyWAY4tTAtWcEUS1DNFs6XHlZQl4SYV4fiGn54YV+e7gFtekk
5RiccdeL86TMeu2zEx7QboWxMKAeIOHwJAIWt57Nj5ihks3ur3jsehUngltIZuEVN9Qje4oci/zJ
+n4pfmMEBU97awWezC36eCnpA7iAnBYYPt8Laf6xnAp2D4LyhpVg/KxUk4Ra+gWmYZc0hFi96+BO
0QWvE5+f8712f5gqqe0v9zqLu/B+vxH4908EmM8m6laEWXwzxTq/9CqCY532tVv07hIYonIXLRxr
jedE6bZ0Z/vOjUOjlTrM35eDTYdtRCeVYXJB3bP9wjSV3KGj+BAcp+Xi8gvMUuPU7X04duJ1GIm1
duIf8OVig+FucpZJZ+pVwA0iUuSoDZVsU8tRJn84WItemhiuyMzNThFjas7rTDiLsCaljhRsl/XF
E8kQWfsSlEDjR9rtn3Ab7v0mQnUbaY1lPs9SOD1RXt0Kpw14heQTuxW9RGXm4woXCNOJybYfmcMu
9Hmy8uAf/7Z+jp7YJhxOss2gZZIBwbPUuywyopMKhDljetWU000vGHKclFZkZPTFFOtkNFUgozIU
C4Xt4/FsVkWzbK4m5yO8CoQDf4YJso5aTXbLuqKt5MClcpewWHJVDvM6H/vIDc0qHp8PciHNnHx8
clPvXnzdUdqQVXH7HwztuQL6hdMWOINc683/Ss3mrAUMATuYaSd14bCD5+u8cD/OvVExGP7zs64P
R28YvaOKfxjk84e42SydiDPgcdhKo9fUWh5Vzc9jt7hOWPqgBIyibMH3t8ZW5VluDVnNVO+ey4du
OvZYCytBeUmAEc1IX3viXSFTkqAeCraL+KN1iKlCY8tIGBwmfG3t2jjVaAs8RYPL0c4kt2hfSyKr
x/c3qUraKeZlqoUX9VuK1kLCLXJmlv9+LugBkRIqUaXVm5e2wIUXoKckY1Xd4vjH151yhOAbcKoS
UTY72YjEQudDfK1kDgqfF+8rN5iF4EydIvYdaqhozcDU9LTjed9o+vtkcDWXd+46KoF7DCK5y5uQ
9G7lvJsLxZ68/B8tsCEqvgkmjqqn2hMoGz0t2C2nKBJF47APDgP7GBjKiQzaXSBm90hRCBDpAf0U
02W+YwllAVIQvqYJxLcykY43afurV4ps8VOtl3vg5rwPrhH3Cw8opSnjcnnSnf/q9F6LwL3H5gdj
x3D4IuUqq6uqvAKjFPBF9XW1oovDduc9a0PSyXJ6hDMeeZ//jEeWxjkC8JyTnuATYPvhWBYPlsDk
HnRqoUTYbBkjuDo/a0bD+hxAZtnKgsmV5jrqVpiUk2AtEKHlY7D9NFCVt5ELfhmGiJWvDwOeDJln
IJkKCSBKJH8xlegSNIVdeFT4jbEEK14LLEWC8Kc4kMGFnY9tAO2y+s/xlVN14mqVip3qLox6EFpa
eTDa5rsGHO98dtBl96MEGM9Olcb5ovuGbA4F4XOUCB9PoYpZiDEo01niUrpVCc9e97a2yT7/Ao6Z
IQTSGdLa4mdt3M0RHd5BKzGHP7TsyUWQWEygJi7eHaJXrYUe83RtgL6fzqdKNWrmwLZTCE1wkSCA
EWXwe2PNC58M/+Gblcx29QyzH1F2yWljIbgu9OsprWhTdVv4tS7habwFFqBMCh8NzxK45C7I8DV/
0hVLLpXgTtMx8F/LuUuDAj1zBzBXBoWQbM6jzlODa26X0qW0TaVoY2hu8a35cSw2VdipBIWGQFsK
1fZzNZ3hIX/Y/TdsBRvaADI82pZcdsAv4kpOKhqEDm1XQGaNMBzypN2+wYIMAkApQ9xedXNKgCEV
2XmkE26BRuO1uoMFYHU3bn7RLiXDcy5EsthISPtDMVpf5MiloxIHdDsMTap5DxJ+cprImLzQIpY6
+ATYDh79Na2f+x1AsiyUGn1+i9ePb1nRpdnIEugpF0kGsFPpoEmzEYBedReVmp7W3ProdDKECpQO
0HDo3qwLraVsDQofEtC7Wod8mEp1Nk5gMHPBk+Bha1+qFrbT0dRTp3TJMq9sRZObc8xxCeyuAU3y
Edw/t6fl6bbKFdbDYrImpBQI5zQUYXIQtLqyNjsv49K1IWD7mbyWIpHwfmMfHTfupAlMvX/VPlsW
2sAQ31t4TuBdpoz4dYT5w/eZzQkwhoZvkygoNhxpiD0I8ckQUa2l7gzdqdsNuGBtqkNAwj1Mjtp4
eVGsuN+ZDMbYbA6kKIVNvhHAeE5FuOS0n67r4fuzs7QVAFrb9uz2M2e1ZFhdRS6L1XaKh3rbO/H8
cZsmQgFlOy9TBgTJL4OLBcKNAxjRU6CLGFfGNioCkgrCdmq6sxt+AAPe3+35hHpP2llHmy3XQ7bF
JQbDVz7bRxuzDJkwYCb9HrGOxRJijmReZNdtWtRFboOIs0cvgrlR4l+82C19lz2PUOv7sMqoPABX
Hxbwi4PTjne63x/1UBT4EZJVIjEVuXirIwxQ8XdN+ipA5hG51Pqq/TJCev5upOYEBtWOEGWaiFQ4
cyUKnovHdgmjyR6KIn62pebJcvO6zTIA9NYnxWuNKymc3Z5LW/fLNPaAU9mHyXZI7FyQ/wNv0vVC
GbBn8Y7otmqQNej4T1WqsrCJV0YlKOIx9xNrMZjlOR1sc7pT2q6JtVPbw2hZSdfmBuisqJYedF55
6RGS02qBCWSK3cb2LVggKADMAzrkkK6OSn+DEksR7KxpFbzH7VN3F+vB9yxpScEo/JcVb2f0BHtI
WciIzPoxyXowjSIq20xPrcdXONT08xY5cmmcE01x58YbsK5wHjfNQMSOlylrGBd3x1y5P4KR8phP
FJ7RrJhqyURI3ezEiq/Y8VKQrGe58xClxLbVihKVz4nBgDze7ID5T8zBRL8pXDB9p22xr1nLAYzz
E4C1hL4SRWY895ieqUuycCglLUNVrEzpIICBpm8/5UW/bbMS7//Iv9NVeN+JyzunMh0OF4szZdAO
FFJ2djEX6KqIA1oG5LX5ar2Rp9Gg5Wk73Rxi6Z/jeh9+pxz3xMATvnOcOw7yFhU32qYKru7I6QWj
uzJv/mVaKO+FHiNPdZXeBJeQTgUvhhIRKZJo2XoI3pOHnfvloZwe1Eg+UBHrZc4b8eOH4Y630G73
x4y6gaIEte2DFgXlXF9K14b8br+OncWqzKFtbgNrNaRvramTPNoSStRPMonWUnUKzBGooDzjrAAU
4+V0e/WN7DJYHzCSUquSiWWWqU3C4lvHYEopVF7C6eGd17LLpFpuDpxwZq3X7MNr5rhUhdajC5jz
Ws8x40wJ8rPDUjBTFhiRp8s9Tj1l+caZo/4+av8Ns/fthZgP9PuPRtoUdmPUFj+YbVHas3wFlGtL
hEetdmk1stoJlUb78QkWMXh+iaA2cbLhri5lP/B4maTeM173M6FtxuLS+7sAujZlH5QWOx/fHFGB
y7vchblAjC/C+VnZPYJXcSccvTTvJKGv3qWV0ttT52UlC2cvRB9Z/CCeSeGWs7J06BHlnCz94g4V
AgO0vuidTd8aVOOQptIfIMd1ZeiJYJz4GcnUVfbE9Txni8tQXqtFsvxsQ2S6qseuiPPvBn6ZRzw+
r+y2r6mYdqPHf+bDUqwpjmmAR/IavzMXptGodqEKtSy1Vzz34yDGvRVGp0+zQ5XKU6IxAyLJj3Fz
NqWujHyyEcnb+foKPmhUus+vUec7jvqhH2GkHztANQKXaPyJSATVo1Wjc41azXtplmaa699rt5mk
S+xS2JdwYalktWj091LZjqnKYagM4BkXuW6xaEfWkXT4uUmOBK0A6mrw2Ygr1zumyjZF76zvTllI
EzHKR6C8eWvKXpaLrgkg4TJw7ywU9znFCKL/9i4+bdCgljaKlm3Pu2uJmWBeAkNHqu8HF9aJTH/v
vFGCtU3wS3mvCa2FjefmRUV39jme/OWA/ygE+V7YFm6f2r0LbbFfB6uW/QI2+aqDokSDXoVpcAUm
nAoeJQENFoXZYO4mNEsNqMJ0JmJV2g2BcbIYEySsTVFwqrzy9ANE0+FuOAnxG7GONQKALRZKL+Ir
/2RW0rC4G3AeGBrPJ9Ptt8XZF2ThfKWwx3AS1D2dgS9sdtZMJ+Dytb58zLDo43wjoXoQhndj4KKj
nIKFXdXl8oBoJTvy2TP7tEcvoWkl6z4kqUozvzMRPR0sxv7mSrdPk9keWKFvAMr49s6Um630YA+Y
CzRyBQ7x0+4PtGgT0sg/t65C7T8kS4KyhMxOujIu4xSUo8NvDKcJAdg/oSU8JzZGJLQ2BMRPevye
pGDBHxakdzCgpUTXHPH32xlv+lWg/NHxqQWTweqNePAfunCPc65eKgubunhNHiy/4CjBB0pJQDjy
VMQ075egW3JcLw/DPTAdvnYftMcQA/HzjFMR2+cZCu490PhdgbZ2ryMpJqnRcGENB37qcB0Io6Du
98/euJXlzCq1uvVqldHZX5obXwwXWNeSn8IrDAmLtvyrvXdG9Xi8KQ2VklTU8pw8OBJJKmgVX+lL
TjDrS+mjNKpWAwmNj+BHEXl3zL3euSlQTWxsIYDprOSJTXOASfmwKkNuReKZWjmjyNY3Ea7gB9uy
P3jL4rS4zZauHhhJ0uDRGkKNFU/PXELNMmjdCbK/gTMQVy7Z1PQ6tSgqtdpul7pA+YBFMNKjySZt
Z9TM5lIMFU39jrkOtzaXmxy94RGhjGWblOGXWQRpoS/5Hq31t9R9JpHdvG4f+fcPKz+h30GWB+VM
3kGL6GVwjWgvBVXexSTcu9QaDliQd9OoVlGzooW4+syyj7ewYsXU9eoMViswoMSaI2RyIM/HlVVk
iFQalGISs8DKG2DiNNyMTbhwUBg5MYHYXi34qPcunfEmhrAS624VP+lkvhu0kBgg3gJFKcWB76FG
yJB4i67H1TCcLSu7RxIo9itXY0/P3s9FICF4aYwhpugnTUVSt5CgDSHJJlaxqF3pS6o955p4RCZ5
1DVdnR/dHxYIQiawzGfWH0OWuCdh/SH+DBJAWeRmXp0uCXXspWIbyL5AGzNWMgYRnZlcbKF5lk26
N8rhP0jaUpP2Dtg6GT5oVpd00DPuf7/LyCsOe7q3/9U5/9hv+AsIZ8QWg5Y4pOu8mzXOgrhrsjw0
TbZIzGVsakbPPJ6IHdMYcgoGgLcs7o+xrp3X+qA9SLur5UM65zf3gOrpLDI1hQxtFAMZ1Dp4JfPZ
UEpP0zqU1ARI3DiCVossPNTyVRG9u8gqjHfeqLGIlgUW3tKUhYL89WD/5NRSEVuLWZLDk4XjJLjh
EMSrtKDFBsI/mAXhCgPiuhCvdd8ytwkElrBT7CfueNR9Y6WLK5tMN2shyIvjeUiPFK4nb4Rc60D9
iz10KYQlRD/wk9b34dk6vMXk1NFT/YH1OQfOQ3Li+JV5FW6hmINcowKt9sYFISR1jB2U6TCKdkny
Ik6ls4lxs/JTAJzvY4M5uX6WaAVwiVvDmAAaav+E/9nuJNzURys1uJiJE5jwZ7PWY5CTJBi7j2Be
e9KeBnSSoByxLx/AlNETWMJ6631AUtaZ9xe1sPfBdYyIEQWdbFNRjydg/M95knkRm0l+Lxf5hXuk
ZprawhF0gvlIEoWKdjxIvLqTpshQHVD7oCl0w+yDScHJxRoYHX8TYst8KQk4f0m44/ZmtvD5DEha
01qEDRrSXUMQBRU3FuSU16cBpE0VOjtClv5zAW2KSdgDaURiHiLL5rdzfUYy+8QAk92ztWPqml1s
ExmxgJ2hjw7K8xJTxGNS58TwlE53WTxWNvxGkbOEgWDW9FirHHrQJyChYEcN0YtA/wmh76wLc7k4
JcxSBRSXibhIkLV5UmzsPeLDhqhtt4pMA2oMdXye1WYxaJuLAP4hNe+qYlLk9fgemZSHry0zR82O
ZfYsQWlKRD+5H+QOFv0ITADQPDg/EUddSt3ZUxmzW0WiRS7ikLXSLqVQ5cJQdHQPQ23sGLLNc7DY
A2/SM+RMsRMxaeH3L88VFcm8RwVCpqzRPE6SJrqJ2DogzlVoT8p01nZHp6PGIchFceISfPn6IPwW
5i/eNxOlI22vwA2jRbXv2hVhWOo+zyGpTSPP3YjcCZ4MsxmRwM6iuQZxF+8Q2U+yq18bF4c3QCyc
QqmSxrlnym7SeMZQMTS9JpMbJFmceiR2rC5lA2DsmJ0G4YIUFGafe83KTsmmtg/QN835jf4gw3jr
y2RjtxmdvQGqOU3AJ5r9Pj91gzW4mJk5v5Pz5giNe1ne5Ivx3c/P2zgbND7NscovXY5ktkySacT2
/ZUfwEQzMZ/pUrncOi1qX2lYVa9ZniPb3oWXGkI3RE9sfhUkS3Kt5HOXtjALkiDD6Io0qXjhOXRr
VmeSkSQPCfi551sEOfjwzjluxeO0WoEDZLMKk8BRZ0cLkFpJD6D7Q3Tc1K1psGgIO6kK9XXYRdCf
bJdTKDLMvxWQErwaIWQYDs+1FKFA1ywZYRItp4uxhvwkoQ/GcyJlOmGz/mOInzFcY/tJGgmky1w2
7AW7S4Q/eU2ar45/QZEfVybr8AdrDHkNQaqhARzP47E3XEP7K/+Bk5QoeFUgTV94rlojYc6OR7IT
ttQD5ajHu38Z2XzYe6mHDVUrSiS71PfaL+y/VLsQ9qAk8sck/9VldAvuBjukKPkuDSL7XJsK5x6r
UJ+80mD0HcAlyaNoLC9+ERDvk4UtEl7Sw6x0QFckuGOKgfr/ta1QxOAezNPUAs3nDtOqjBdHs08j
02JrBJMFSmPbwOK5OCtsS27yp4BAKTDHNW7+y4ZVZjOS4wgFUweJpOqHApXe3zXHNMrLLmMImNji
NwtmHKsNYkoVywqETIful66NyDtT3m33lVgQBfY3iMG58jkrzHvxJkryOsUg/mZ+DXYemWP/Nyhb
6Hr8WWh6CWjgxSjY/yhC3Ewa4szYux+GmACTV/ERDklPq/9yrjL+dL7ERyBPKqfRSyVYEqODdv+p
/k0aO9dGyP5MjQBK6xib7M7JfvZA1dZBygYe0+bc+f24A5S/Qlv15LYk2ECFHFbqJX+R3o35WALl
/6zRmFVBROeZwZdrHc90mFV9t/eBzpgmOLsGBcfdBGSX5YgR5EVC+Gn+T3WUVdLHlLX5oVm6gcbW
oR412ZYVcXbmnVyDsmc3z4vDxkcioINwNXONRVhS+GZnBaONUnLn56fNPGapwuxu3y03533WeZyR
9TavL7/3+BJsvQlj5ePwxuC++GlxIbZnwfgDYzyFWxtzoABPPsl28NgoFxCkB0cZCELtDumpWRr0
cPu9AMKc/qF83/Jcs2zxE+JBoch13ZbsounzZe37EeDhJmm33N1uOSPNTgUfeOsXivTY9Z/LP3aI
Q5+B5Z9nhDTEYDhKxbcmhK+5zQZrLSxVc91yRt495RhttEcuR3tg3kk0ImhutbHzuae+9yPrEPCi
apUCzhE5+nHlaCy4fBBGjZt0Jq4YlcdjKJpi0GqIse3invUytCBasJUMmeVNEMIEM0uEHwFCWhnf
i8MkyldX3TGa1eS6N3b2jmP9+W+PpgWLXFIhTzC+kV5ZEdg6vMG8IRPA47v1watme8COrYcLLyLd
rzEg6RlNKQ1G11SnkiARuk9pHRsK3SSxewkV068YQmMtAPDo4TGUONHEomJq46FV5KPBGweQgaCa
2zjLaT6wPO/d/EEIlyTgKkP5xAB7PQYmXAHP0TwGr5ykwVko3mBLtldNXGaYOa8J5LOhxeTL5SI/
nl3oIh1l8X/7gPAo9/KaJi0r24irlxL97Qrr8vGWpHMff9I22f5GRsBGeffBLsSb948pNX50jFtj
SvGdP25BIQxTAEcLIwV+ltCiyNHRRDJ8NFCwNV3VCBwSsbCwInlc8/KL+sN9KeOKStkrUpRnCWX3
wBO19AwWv/DjZGVaJJa88uU0msemzeQxFmITHkHhRVjoCuQ1BV4GnDdI/FCmZZ7rTuD3rUQ9Fb2O
slQ//u0GDIOx4muMlj7/c2E+mRPmY40Q5HjwH+O1rtrdceGWjsccWc33VicXKtXS/R8tsmuf9gNo
fRVnD+fKjkp9j17w2hmVz7xLu+Mt3xC4BLT8erphaTlmm1Aug6lMLqRUoDFbUKNqnaLujkc5/HJe
pc5F1YHLwKrtWnrUPNwrzGTNYalRvnOFe+7y/NeqmBdjNq0TReIXO2wSbr6k+D5SQp7J1qoEqheH
49EwrNjH2ZWIwKovoDNI/TBDcKboUVPqSc9oUFF3CXU1a/YJsI68i+w5to8GcXgkhh2AqF590/fS
jpwIBpkRD7i4FGmqzJzzozJT0SC2FG7xxodN2l7xolm6xEJPObd+DuxuGUdacAtnBH/RfjQBnsXF
nBNPawe4jOVQMO8sA65/brgkpsuz4B7xpOo1/jArMp1Xl8iD02KTmBU02fiqxtAgBdHHJ2cTozaM
Ip1tdwE6pEVjGMq7nUTAAqSsWtu5Udr/m+RdGBJlUqMmf+pDIt0SDFyDajzsa3BDG84hOYAZMPQ3
795CrHoNVYazZlMvVwMI5EnaAT7SisLHQWvdyFdqg/2Yq5z6Cz4YGDQ78rP2oMvh7nNGYICmKDSc
VPUjQv4J2+Y4Aujuzg/IOAlwT36W4Bpp80QSo+2KLXDVTQGy7uyReZvIbNRL58nxnpvquukqZPJu
hLVnq/oPsuUOOx4IOpdI6riAmlWA7M/rcBYxErSHT7/5oXI5W3j0A9E1SZood/Ktvi/srOBuR3Jh
CzXCiwjZaiVv/Zd7UvVP+r0Zny/B4/NKFLTkjIm8aYJUdM9H9KF0MSwLcgrv5eiga68js1SwER6q
K4tLx/119igZ+NMbzNaI7BS2zdXgYwD9BBifO5EGtmjnnxnSMcTH7P9kGBsFh2oxHANC4M9/W/W+
olcECNM+yLJKBYqmACER2rj3myMNMzxuwCOI99HUrykArMgU3ONQY6RmDSnpu/qh6devJD5L6XUn
L+TPMOYCuPFIZtNKw0XW8e9icNByLtIdE31aLaj6SwzVHL/eAxMoWJ5D96FEawCoGbxfHFFdbSC+
rkbTk+x3X+RwRmmBFlcKCMANH4SlkWPeCKZnk4RWX0cJVj9qUEql9US8DYTfIjWEneuDW8Nt8d67
xQ6nm9rG1C8zuuS71jFrRe1uErxXrIjwALAv6DPjt8E+ZGe5VvCfqar+tg0iKI2DWG1ce4U3spIi
cmywZO63PGxZK5obPNYBsRsqASe2sQyMRA51NzmLAVSLfCuY8SzR+hYlU+vEeBeu7d+ru31HtplK
8KZ+9tNm4f6pJXbYZKxbfLVqdaTRfOhPd+Hv94O0HzYUuMJ0Mi2gkRAgJmr0m/1s/42GjOBZjlao
C0otpF7zyTpvH7FxfgWz8PVjytGP4E3xjd6OwCgYfSETSxsvz/y9omdIKWqx78QAY9O2aPeIq5DB
ybSbTvGgCW0Y80ZGE9OvjpxcfwsDLxiEmMi4snbCRup65TIw0trabeMZyJCKyxn+yj4FLZvkhwbD
ytUOZ/tl2XXelgtvWf6KPfej9IHmR6P/KUrruUBIq0N/+i3Noh8jb4bJRjNm8J3sWEg8re3/+3vb
+WANQ0CZtP2W8CqfChCprq1C2C88IJuoWH/x8r1Xz6seiXu1J+2cg3P4g/SCWFPKeeyDC+geCphp
mvOEgzWZ4n4KKl1lr9y94l5G7/NEVSLvugmG1sI3DceX6hQoQqM3jZlCphQDKBdwIvQUhZaLSQs0
YoM7iJ4BxY9Nen3WkCbQzvnP6BCrtaaGklyaKEQpX86uHaQBGTOWDQIA1PWeLnDWOW3MzFkoJX3H
QSXs4dpg6iIq9W1Wt4D0aIg0geJPqmVXp138biGbzp3RRPE8dlu2nBDPjpXHkjfPg0ZlYoujUHiS
A0m1N47iuNHPjwXgYz2h6hHOQ08wjlV3Ynob96lVgXCDtu4y7EY6D1aPiuP3wTOyvADH8oLroF5V
VYhMMdddo5qhtOogcUfaVvpHEEG0RXZvdfFn6hOgUIazISGKyij51vWadOWwKVIHv5KySfiD9ks8
fWTtEvaRzXjB5aUyeaXGCP61ARYn7/royNeyHWJ7jnEMM9FyIzb22v76QmpWlYAqd3VVinlo8TeF
J57/9hY0E/6Ec4PfznNNGSF3m1AcuTC3RDCfFazQGL9S0rLloTG+QCKVFJBk+YpWafS5Wo2cNCCB
010cYPKjidE+gcxphNqUoe9I21JCgS3C83dYMUHWh4N8928mppC5SmvZCsDOBUJJxeZ+xg5bM7Vn
vEZ6DWDUAFLGQFRQybHTgeXOyuUXZLel8ycq7UfwlvKzmtrsmGV2jmfKClhFYCZUaydOE49PJXC0
E7oP/H2XRLmcs8FWmTNiW9nxYSNxwke6MANAv50gz98dryvFXdpv3AFHzHK0tZFYdZGo8tubtLjM
Wmme2l91sgqhnHo8avkfXpt8MHs5rAnLrpEakAVl6k+n1QibIPnIhwgob+jx5Sht/KEg6nyhq/MZ
IaE3aSY7FXfVo9pcFx+7p2rjGarfqZPbFBxGWOvjrNJ1X6YO186RcgoUnOGb5DiyIc46ajB2Qnfm
lOBp+jH+83dOMrhNJjQwv+54IB18ekfbo4W+QsZuIUbQCSopUPb44jCEaGpOeVoqT60IDAip+NOX
MF0iIh7LC3hqmabivbI+GhoNoPrHFYOp96x/Gotb5lwlCenGE4RaYtCHG7MaagfFF4Cl3OAYKUM4
IdTxI10cPPXiB407McUoGvswPzw07jbNfwaKpKR9jneT8lbnZO/G7tNNBIB9NaLOaYHomnbV4a78
uFm9qMjEQl87uuP7JFPQxXbRG1EF/SORkY/lrZoJDIlQMo+E0o37jl4wnyko6nbVAVdUKVy3OlI2
yLNjKlMmvNM33frhNlsLc5QWBSqbyAVhK6RJ2/fX03e/jlPlotinUOUpt6PZ4T3eYBk8StUVhKFN
zELAe3P57/aBlpKAzZXjK+GTLP2pIfE6VOc94wDFTsQYZu0stAjf7I47Tcky5Yl8roW2Z49ypK/b
sfpySrFHsWSXN/gufyhqu7D8RBczBV3+jz84ZFh49Z0bbjM1ls96PqfxVhaow5vQxt2u6AArp1sB
TqkCz8xNF/QE8kpo28qRbbfzM7jkwG4f+YfpZtWYI0pbzNdo+FVp4NHH2gGnTBwLavs/AswTcH67
P/RtKa/bRQoYWJByqOK7O/Yi32kgXr0Ufp09F4gJTeQenJSV9beMZe+qqpXY5kohA+PpT16iUSgy
YVS5AaGY90mQe9vlo1QLH6UUvAWzAsWtcSViiScabLWf4dz9ZdPlqEv7crfhth7m8/t/h77A2Iot
zq86I7/YuuxkmxmASERbWcvhBk/zT2CVlb1Sl5PW34VJpuMGtYKONABbMkf9hBfBl6N5u063D1Ny
Dt5+O//wrQuozfjatr4xtLDc20MecD9og0Xyqz6KuVYkaQCnjECNw/DD3+Yhuj28wx4XiJCZPU63
mmT4JiOWlCCkFYn4Bxbq8UyUtiUvLk7TY8bycHfo3SSfR+hvbt4lqhYpKrEkXm3guWYqjUrONziD
n/4oadDSRnvWroONc07FGu87oBHj39s8JqhlWHp5lNqdTyWOPXKMLX6mB0NkgWYZEL1Z18zuUyEQ
dXqWrS5YIzH8VUlrEo+k9uEf64cL1xWj3itWwiQZuOA4wO1QIIMyzlCa1kV0RN/NzgHQMiWkuMcW
OZveEg59gxatG9CKit4Cpq1xWTl58AyMONdtqbnk6/pHGM045pCUrxfHLSs61Jz8kKE/zNo2sNlr
73Y2eWasXpwuarJmc7KzEdJ9xJu8/PP9N4Ky5HyHs8KXfA5zcH0P5WQ+dllM7gAg9JD4YMFbnjDC
E5obu2HovJv0rxaMVKKjI2+L0Hl11qLUdlGKDdi3wmFcP7xvvGeYoZv4ipDjFpY7hmNzGo0Ir1fL
2s4Y+E1MfihHHdFPJv+qIRIiXrNAb4pzyiCBjtSH38aJktawa93vva6HSM7hr4egishyZdnCYJ5+
N+R0ij7/f/Y8wI8PhZgOreA4Nugmh/kwIvo2s9Wfez+DyEyqsfLUcY8aReH7jTQiDN7+rRL45HGJ
w8kn/tgG4iUia8BT7kQBV2zqb1WAbJdY+WQHbZ6mS/xMp0tYJ3YKv9gt8BamYaWi1YQIRP7eaYbu
wiZ1xCHDrZSbSkhXzKMmNDfjI22joaZ6bcgRWVfCqRiPkuGGQ6WZe8T9CQYWC+W88u0p0aopTs3X
ZOT6ZOQ+mKyv40dvPdaDwY9Vs2gJO8QzHzQPiFndA1hO4fn9yqaHebOis0powXbMjbe2n24LZolz
jpsF2DKO5fbpJhjnhGUynByDJN8rlmZWMEaLvO+3UddHEHaKKh6BRpWQlfTEmpNaC7JAGiRHhP3T
Y/OgKQP5fWkFugbz+n8zoLKmLNPU/hnhYCNGMP1tY27aDCxv0jY7+HAyTeSRVwPu1L6pHm0FgPfQ
K0BN4hLtS45lx1x9nkPzchPUu2sbJiAiYSK1UgBy42glDeap8ILhWRmByiULer+nDzjqNEEC7VLl
YZrsF1NbTDdMCsYVQtY1Zs3caTp0w/6UY89HJfhzjt3egtdzskAvZTic8r9jts6ugyBZCEi6XPqz
lMOE3Y2ciqUFqAnv3KE7RfOcaq8rJFgI+hWUpOIme1JyFf7WdDM1jwCuiI29dqf6MsfkANhetBCh
J3K3Xwx4bgwM4PB5ae6EQZSEBC43O/RaqfOVNEOq2P9sBjPo74Cgz+oSFQfVEBOQSq2o15Lz2PgE
+ngvrYUnh+8SZ3DtdKZYmLtJzhtXKyYAMGFkc5PD2N1Z88vnymkXw1OIKMrvUaBtPEVsGUW5ue7i
4it+2a6SMW6zRqR7MNWIIJnjMZrrhNKb7nkpQq+rIgCirnVSRqOsqbFOeUcJyjysm8ABWHhTJnVL
9j7KijCmW4KOwbKM/nVgnaXSN61T1TZEn5PDnsKMu/8qX0HJqRzjB0+4LwNSSWuS6xp3UKoOh0vH
MgTKMEZZUm/HJCsDtgQXIlR1Wp05JvH6D4FK7+3vOBWhcuBzxK2FKeUNqHaGrevTfwWm75z3pUjC
cEFz36Ni4QRqShLi+LSRbjdXObxKEwpFBSuZNMoFG6gKop22QBdpZyS6P4aMDp6WSZZP6Hj9eCsm
YI3qKqeQt9M+Ig0Mt7ucWO45ptoKaq7E4WEHGXhzGVneTLnyDYGabvn2ERrIEkx8LNcE+sCc469H
VKQn+rkhLvs7z9qdRExpHCJl1PN2mwwzHgmMWl1dYUXFJ1oieEjyu6mfLu+ATGqjReXIvjDqxIHb
wg8vDaRJ9WVs1594XBqsW6of79Z+weTutWGRBgQymeRGvM5I8/DANkY0LRDFfhpnmdFjDbifEwrY
MFzzwBHml4Cm5uk7t0PU/aMqXFTR+hAmTlGOd72tbOBhIPIIHWszwSkvGh7P/Cmj8XQ+vHWoGvKk
d2t+hKdjfbMk67O5Ikpta7B9TqS8WatEugfhx1j3Ie2lxcxGQZpjzjFmZnBAd/vV0+XEdBglG6//
iQQ7/GkOLQtPzUf/Q3eH7d6Re4udnaWbyQ1ylSA5d3NaPYmQTjPNjkRMkSzuHVfikm8KDlsVEn7D
G6nGfrOWJiEge2bTVqixZCjp6wxS3kR0N9ANEJ9afieqTWlIoGhMkMNylFBwc4/CXMnj2Hjd7a9+
0jP77C9lK1IaLUNMN2aP3gsHFrIvB4bU2YZ3Frr5o4PWtf4aNSyEKzS3EIqwJtbgZTYz4Qp1ybxS
pwyx9TDLldXU23rUIDj7GKY1n+1MQsphpSUcXJAN3PmFXsJeKCvV4jxZSs0QJEcJeqktgZyDpPmi
GGanB35zmj6mQjuCHxDirJINAeSLClzs2wsQ+WyssldNUXoNfFHbCYmN/CPAQmjZkoMJmG26aQ+F
3hV0FOOcKolWUFgn3eXnJLjK0CVxiXpjR6w3NIrxi0ZvpygJs3IJQawv7d1JiCHCw/UsUSeBxvX3
KCGO8AkEOStv40dOj5x65fbmcOMeDIEs2T/vhAuRtuHRdcUmp+YVTJDPOQPgdWOi+jAae6rQIC2R
8Cn3Igu8AuMdZU9+LrleNQUIXl7DcJZ0BG091UTDEiaIgB/PPrJgtrb8Rpy1eGfm47nM4JZp+M7u
nhhwARBEf9HfBOJ1VepdDHjjqPrNzODY6gmsv+C7Pn43YqQ0mlndHPkgl81n4XvgQoPx46EsUhG/
Hq1POehJY04MoDzp0aCk115Xzf1BP/klNlo1wyNpU+iCq07DakxEA53spKM89Z/sbMUQQueZxsiH
NJW6hOMRmivhr9k/gTfjMSXvTcqn++JXPuXouSl3xLuHBW2ligmWcz4akL9o3hNEBel9tidSuU/O
1MgvgRbb41nkN9EYYylsnjEabTzvIJ2Pur3g2IbJod5pp3rPSmhG3eiIj4erC9KoxIARih98zbEk
D5qoC9obu0MqwJK3lNpJtW+BKSQfLUFhdCP2b6c8z/CLaxf3t3xP4JsIffhCYlGXoMxpPYAWtoP6
96IPeJ5Yxqi6nH+pLlWihScm0FNrPq4pB/3P0W5J7cfqoylO9vAp1Qm4ZWSEPLqlLfv+yJ+6pbFn
DugR0/m6+KJxjB8CXjujrYKpSQwF8X3K3stwU0O3F+SFVZTyZjsEwjaQ0kmQ+acuvH4MWKXqsY++
+bDUL6IIwmTzk0LCgvkgSItvb15jp1pLAGmkokBl3xZbrDJTbrxdGK+NNSUuPJmvBvjBPAt+q0yU
tR059nFJlSghMLRi+09WC/pD+lJinA2x3UKDpI29J0H1gFX34C+sBmN/SHDETpc8QTSxkFf9QWSj
M2XbcTDZQfpvziwInsqE5h+IHdIHENc1Lt4f17ZaEnXVi7XE3RNRf7v0q+EOdjGnge3xl270RRRR
ViTje+PmZcQxngHxh2Fihcfum1aDlmO6lvJDKXJBWp5qY/TdHrdKiUrcjjSqIpsyvhdP+8/G9nlh
V6JqeNVHKu10yteheqQ91dU5i+RwDXfCHcI6+2Lk6Skt0okFKtHV4c+c6immKqw8JP8NcZ7mWJKf
Y1v1iAYnFQskCg1M7WqBubgzFfqPzEVVu6Bzun7xMYoXxMasngPZw4GTzFHOJd7Cz00KCeM57GHD
iYD+kmuAIbrfMVO3oHJlJWxmKDtpPzJ5n4NM8iDMh+5ayw5L4vKCNw0Ghcq/fbC46c49hV4rBpMl
jWPN6bV9L2FX2ACeMP3Ma3SYSfU1TSma0zoHSogk7HvJFSRSz6jV9U2A7fBIm0/25uTdCzBxfY2b
V1s77m6RgwVDn+pf4IV1m41uFw0xK2wLkQmy/dFvOIDOmqWZ9yh4EvZ239WD7MJVyVAYQ41g6Lp3
NsyeHQ5h6QblJMvirYPlfeigiVhUADNo1VsAuTZx+IeciOQtXP6TYoDHREW9yLq/9HZuuIrdjCcj
EqTS0cI84QBG7SBB5RcHYaz6VFvJNY22fN7pgCDuLQBFUiITnbAwIEzuUEzIcjk4c1a76L8+L64e
PKVaR1tUbspndXT3QdE6TqN/WT0NXnBj4RwVxnAu9akKlShf2iUOla/+xRefV2JksVa7q9jJo6DB
R3lwgv1IryfG0RBQueZ369FRszqlHGbUxkZCGGL6crPwvTLGHl+VTViEcgZldU8b6UqX6sKq8VPQ
zSz93y7NI/axG6saommvrgaLwUygBA6p9AaXG48f+7Oil3GoRt/0BzZPrO4mTanvLleNA+1yMfFh
PhnoRLbuwt2p12yGUE/4qXDrB9nRFhRBRH1Z2GOHOKdGxTh0zIgtl4yLLZw2jTltIZPNyoivyUkg
28Xx79AWZxLuRpN7yn0AVZZgKzpVzis1UFFDDOnKQWDPxB986dr8U0F2KoGrhOJDnfMeKESSfW+Z
uXSSL60GGWCbaig6bPTmV6yiYGPmNtHl6kWlYKeOFThsuLmEnN9RcL/07lN/ywMQqYc/eLea8eRn
vtLtTxVIRbLTJR7vqv7lXEmFR3QCkMe0uXkh1Av05Iu3B0S0c4lgUbNkBodBj6Q9ejcn14uwa9sF
0NTLVjzWTcZ2IwkmKoKKC8RG+VVPP5Cqk7D6lNjCZna1hRXM8+ymVn9MDawkRBRQKr4LY6QcStiK
g+GuDgMnguAN2CbXgDRRr7tI3ScdvGfFw8i5Sshc+u7K9JE9ea/U/xrQ4jTKn7bVDywOu1P72jTT
a5MHTz8q5fzo2Lpw89W/PGn6fDOzGpgcZABAglNamUrvIxMU6mwuryuD3qtcvTNTi7YsWhJWBmCD
lamxHfQrpwNEk1/ZDCJRlCyP8SkGVzLqeWKHBeK38L2ce8MQ8//S7QfGbVVx5Aw/u15Why1VsjpA
V7HTVEed9nx4sYoDy8s8D/L5HqUNzStqXxnhPSdYENLETmwvOsYlIkP4rNpqSyAd2wKyEli5GK5X
bggUuPMdZOfqkQppHUet4PHul3wvs1DFlaD9ioBQF6HunTWemqht/sqANTslQi7GveungmCm44N5
qPbzrp1SbTaL55gZcKNntkq656numR3VFRaaeuQgytRCdSLQQI2CLB4Ex8lAI2ju6KRk6SZL5LXJ
hi9UBitRxq15OxSoRpxKUyhG1wZVGxbZRVm0rAEj11wgpuMX6vfxoT63/xeCB7jvCqSBJ6wPDoVp
3XP3uaZJ/PYrNKosCX7j6kRHMBuYDRzlXkFRToKc+z5ZboO0jaj9A1+HOH3G7XkZ6gvo5jXrqiZr
swsSAUCsNycKaajaKOvg3wwfahoax5Yl+SpuskX1NJC8IWNp180TTITpw9P+EQrdhEBkHCW+56uU
lQuyUKCCNHIdFERdqq42iRdFh5isicYx69ZwXJJ2L5V+f3wqDGHmngHiavOaKRjZUNLOK51PFRvh
cjhx+RDX/4vaqObWdqx1viVQ+JPhINd3cci8UNV/heDtQ0w8WP6ZFDg/LJ2LmjI853Y8DlPXNGc1
/sGK0zWs5xnu8kjfbRnOspUuxxGGKzvC/UUFOvzPph55tOYddg4oePKcLLq4BL1cie7dSpFkSRkZ
iyIWhpfzJhAPGPAvhE23EaESMMvB19yIOSKqpCDrRuZJFxn0733H+T4VEXuWHF/LMVsEEgIeYB+z
lBdkeaa+soJBaDfGVxgXd2+tG5UXB7LVa/fP1sFBy/zWPWYfD7LqqFeDPiqkugvGctcmcn+RbRGY
CQ5T1952diis/EG7NS2S8Ihzqwg01727EWToUQyX3P8cHQzCkX3489cnnPdZw4P+314L45eRLny3
7WL67dtEtx+sPH29HW6xr8jfqrDWtuJQpuIeO9HDMY8AYvsTS24tCnDJRmp6MtwHdjY/d6Ej3Fqy
xBv65+4gLdRcwSJuDP/dZ+YXYDc1LzsdJIxQz7ShQ3rbvsMlVFvE1tKqEjrs7VRfEENXrQkp44ev
qH+zIzztu3k/Jf+hYlKG3GMP8UwOl28nfYA276GOo+dBsurMxdFVTni55dlIl+J0Why5pleQfpMc
WK8Usim2NNo3+qzFOFIZTsaYHiYJcDBMUvKdrhHwnLClbyoKtTfhUx7cW3hQTmsaSAt8UOpA1zp3
i2GpnyFn3i1DB5L6B7wATgz9u44L/ljCzdXUciXI4amq7csdYYfSAC61kHNou1IDFmje5T8LQDyJ
NI6TlYxMJcunvpEOtKu6gadoJ7XWS7gCqVYbVI6Ghd7BmnBxqlpPy7ztOL5+H1DyJWE1dhW5h2F/
uNjLbC5FiSKiyIoFSSbKNHZs51vMub7/LkvyuTHfhLa9cKT/xvXxir4d3BoS0qdOzZVY1CMOyuxc
u9kzGXbbyCwztZ3zDOc8NVCpADx3rlpGFTiVGgRdJkpRPom6Rkiwjbgu/RsFP6dQSKxFZc602IDr
4Az4Fj3woihJi9CCxUqNqUtdpmuXux9BpVLAftpevwtsyX+C04eqHd6184yW0dvdx3xdWNaWUTci
YpraPR64H9cLZBVaUrIpE75NSCs8cYtDBD/OpB2oKbGN3hdNEWm9/WBQs9UueTkjdmcYzGb2lxjJ
OewSwEOGHrgFWDxZf5ar4S+Ak3DQL6Xsq+gBlr2UHfT4l6jX34mjIB/j8a/VIY89lAQo61vz/VY1
tMZttICTSWEKjmdLxDO3TiIjtRoEOQry+3jX+FJmlfegYrNnP4Eh6Ch+EZYPvJGPlZDvykIahoDM
vbdY2y8wx74nb47EN2EGBdilHZK/MUMzwGOBDfgFcY0b7NVWG5kQezFQlL4jsZhpCExm2H2RViac
taa6VSbihGUQGp1LjyaWxySMmKW3Px+h42otLJX7OZoweDHZlOzSr0VAeB+XA340YdYCpDg9YOw8
kUij6AUxlz5NDl2aGbZgoQ1sTLGbM1uKcFidZd4jhuQMO9ZSOC+3S7vethtfu3RJv1XArIgpLfgz
nZws93dCYEGY2rNWcuEivl2Q8neAHJafPvefxY5tbygOKXg23EZiwoqBR0uskyvBeJBjaHtXPR63
L12QgYlbGFH3q32oHOvio0WPkkBBlQQxWuiKdfZBNDIAg/667XupoJQvFCPSq37f3pu1kRien0yG
xOwFwBc0tzvrspsAz3T50pLB90D/4CKKKtMgYnk9+ckzkFQB9opptq5zmS9aVSJi7aMl4/wMf8ak
pARlo7um442owzm/uI23WDuskY+c2gqgkgEPBQdrhVx4VV9xGvu5j0nZTr7w0eDnxHuX7YXlhMdV
bBjJfn5QtoE+j7XvuLlv5HgJW2fVmI8gIdpOOmGXsftha6+e3wym0lDuLHfljkZ+6fY+1XQopOJI
ncZj8LivPaChYLKSbiysEFYDGa/xv0HjZpw+vrQuCeLXJLrWhnI2C7yxPNBJ+HWXrpEc9dOyXkl2
seotAkog+hAbKtrOQgkPDJ+x+xKvXMONUyXb8iCyQ+nEBcq2H9x0yhHB0Qxht0FVjCyBDYN+lBxX
PzPcSpCIPSi64JeIWa0XLT6MAJ6fsGNf04efLLdFBejw7p/1/ivgCxLeTCP3hKK6JrDqhCq1Reg9
ZM5oZrojy481wuGcm3kT2g5Nzu4ERoyN9ChOwbNCbzRYwrSRV38obuzw0IAHA+xbvH/fqALnPzge
d4pOAqw9e+4Ic7xCuWF7ElnXb8S/FFDZ0q+sNmCa7qLubYWB7wzoiEO4r1joDs9RKrMtyQTC1/k3
OiOjP41Bh43Qbc7EzO7A2VRKYIzx+jBSOmbdzrrL4Nw8MitqRQU8AUbwBCQtguIOgOisbixNhv6R
Pb/8S6aLAR6yUKG18Kh+vofLn4ikKMohsYchrsP19p2KK7jHSXajWb5x2ZhUOTweldyiWWFFtZSt
0T9zIvhDXo77jRwsjtBmLiMeA7BfpuGY8SiNNabLyyr1FHSK8hqBkQB6bDkRy2ztxYAfHlw+iM2h
Jsz/pEYFLpOGEE0FRLkLsbWAGGP4Fr6bXS+3O96bvwiiSPcGQCFCt/1Nl5bnVf0F8NhRAmTdIY4q
Kkv8O9NkS0c7sc03dBdcYK3it/4FRSBC+ixWB8pXg2UO5jAAGqK0SkvwivM7+XSLooG8r8z51TAG
DjjJzI258OhDQ8WIu4SYbroCwE1AhLCXNOqR9kzdyb4XaqHQ5Qc3XruiDlkUCyUOEkADvrfmtTWJ
Hnp2/9ZaJ4LWr1UfktfM8uiwGDem0DiZy5rwwFP7FlrlQsojkdxjovHOOr/TqY3KRKHCZRz4ivlB
hFyTmcDowtNVTKHLC1MPddSMtKr9Zan5iucNvJI9/QWqv5cARwg2kRZxSMLOEQOXh6nSk70aH30m
MGxcTJO65aRwd7/16ljdLjIea9JYmpehpNOPW8Mi3KbWAdG9cl66M3Uac3omnHAWPrmd2U8pv64g
dQb6Q0YDrwwvwAqqJV8j68s6reYOcdMeMCp5G4QLBeUTZc9CUiFBGBeCtTidht0BrF6dZ+zN2vPu
uPPT3cfBokHDsHEQMPbbIlUOkdP/SVV+fNandh95jZpYFKUHSMcF56Gcyr8VMmVpMwRZxMODOcQ1
3VjXaEm7RvFJgVCssZpvj0yFmy6oEA2eWwBvW+GNyx30yWIPfEv8+Xm/JwPuUjf6xd2txSmP4str
W2kRv6IlrG/TBvontyZ5WI+KwE1QO0+1GWgky5O7Z8ZRxRdEv4DgrWVZ+kWawpXiEHtVukBR09K3
86eMnpPGpCOs/uPBXLOOrcPcb7PD1gyAOQhTTrfvqiB/KwIRj3ThlOwD1RAnTYqS1QIQGr9MBRVF
K31Bfd40vsl3iEtJ2Pa+2E8pxIY2TeKmNdHBQhlaNpNCEneIGZW/xKay2smM68zXUt/k80QTjhQ/
J9ioy3Z0uZuVGxJUloDnYN8q4PLWsSbaznKn6Zo10bf41NtUVdnbozsKfmWrsCa3nQth1W8kNiLm
IdzX4Aw/u7bnjODsBkWii/FLJShUCqp5Qg7uq0X/vFWKsV/m5tK2yjjrl8Q93jTlFXkuDKlBWD2f
AoEpZoC3lmlzfk6LKfhwOzHdQuK5pDVPwkWGsIyihzEVf4IOhkoX9cT8c+UV57fW3D68A6w0bWhx
zoSIVIblOLz5zYUc/7YSJOz/5JUjDjUo1JDXAdWajfeS+2oKj6BpN3Bo1aBiSGsRQTSAv0fIUyFa
Y9aM2rXEmTKgjGiOsVgCtQCYPdGQKoeBgXK+sOAKpzv/Yx3jhWw6OWPvP1+d/MalUlyxUOnNLebj
d8y32l/bWfPdX14uY4Xi4BJVnhcAVYcc3otxAmPEGX+Yl2rRd9jRY+Cq6ZTxvrbgb6bYBFZ6tHyX
/iE39LsdWDyniqSqKIgqRqIuAONeuYoV5BvMZkn6IEft76Nv0Pjkf6iNVyuLUyResL0ljMX/6VsE
shX22q7chg+5j8h6nR9fLNE+eIuRkdINU3rXg5q9pou8NNC4/JK2L+1LSwzosnkoukq85zUutyp0
jfD1VNlxRtIiAG/jVByB5mEbXGdvDvo589OCEZnCpz9eHAggTRn99BucGJGsBvSAuFXMwMJCuQoc
p9LWhZpI9a4cYGuTDGBQ1b2WlX2D6TEzOqMKBFKyKyBhWhCXPRqjoc59fzG+wyp75aICE5Hxifuk
Wv9xbDxyXG6ChKBNKR/1v6Sm8SEgmy8Z3GLAj6Mpk8x9mlABsa2ECc5BKuezOCiDmD80mlGfxAHe
sCUYbk9mC8fGy7863y+i2C4ORaV0PHhfqRLhmm8jvNTIB2p9G/xoigccvsLgrmw5yxB8sqfwfaSN
Qf0YzzAGiM0rMjTk3g7GE4pzoyKr0cSVs7M2XWfwaiU+psLHfIOVBCBqGmMbnyKf9vE7vRAUQB/B
e8dABlithm2xwLhoI84MZJ2x4KtHhJg8G6fuC3UbeaQmXn9D1/c1npPnK6mwbRNLYcEpJ62vGvAB
bTGdLTfak934jm+CD1hr/W2ctX9Ot4HD6o3/5e4XzketO5TCDlMy6Wk8QekwIEj++3+im85t8DYF
wbGmbzeg4DXfnSP6EzNolP3lzRm9PMYrxRGzrYfHqk3A/CfYtGhgNiVV5GVO96OJp4AR9KIc6Tzy
xMdCJhVi9CsSUU+3UpjYM1XBofJ0Fcw4FfXFFXN6Eqq+Ba1fnQAfrsS+g7WQPyq+RDqbDhKB/7NR
EzmPpdGigLhFhhwpIBUJPrw6Dbwit9QpImVffGRVP+Xi2rVTERrTF74J5dRA5QIRtG6KAa3Qq9tc
gPhAnoS5MZpl9P/LS6GghDcfyY8l6gZIOJp4SQkSyLORpXB+LKEJYptFKjslUpUHGGNZdG4geVtw
MkEFzc9QLKmEMUFa1gga7cs3pE71W2YIQWh52VrMgwNq9ZsviMPI4KTEQatDBX2PSCVIN3IDOUUQ
r/Oafm4xiNYomv05YapKOQwBE/GBGk0D2LrSI19sx7l2g9WLcn7DemjH9A6C9qlK4FEog04mMIV2
jUJaJLxrzLcjS6wOlRTUMa4RLupynrTvxsI5IJaxSBZzsD3/Djbx2Z1NTg3ddoqynksqbUPMslT5
wS0GlWcQ23E+7UEb49GvWyYkSoWbVtfXj/ULfOZEt6ZuywBXQLyDKRQysizTdEUZeML4k5RtT3os
iFatwhHkB4oy4a8wn7QYQAEYIda1GM9apcXablz+8zWiAjXUb5LCf6JpWRvDZATfGJWGov0MQhah
WI/7cfUt82pZ15/g0O/DNPsLAaqfzH/S7Z7mo+AYrfIDN92wji5Brl/IS743k0eXb42ymXvXhfk2
f23+WzvHC5bGFyu3jdPRj8OILyt28u7Bv5IJCdqgwkVPbu1ob776VJ247uTMdRJDsu75SXOkNrU2
Z4DBQRvDKOgm6oM9N177eUkKEuVlLzm/q4TEMEI08k7Sr+YPN70wLvjAHU80ySZdyyaAT/5hQQj5
bhA3faR2lV+0+A3h5pehWC9WJEOSlwgHaCvUikIzOkZBYe1c1lR8Ntz03ZlELDkVAfJ6lA3PBxg8
YZTR+menHrs+9NvMsGOWyD5FuxH7FPXCi7N23sJjPjVaRBGoqbo1u0DPbuN8g13ruYQ176dCmbrs
GSOU6srEtSSv0DNd5gUnaSXy77gJCho8TaJba+pCPDo9HLMzJ1tB1lMW/EUkjhi5WM6X8gXa0/GQ
OqywtnmBCxF8XcS9xlztuYXeZMyPJIT5vNjX13BaP2crMNHoNNIBP/1gkGu8Pp00ekUvsucGc7P0
/yJYexmjHv3/fK0ARB1WEfUY//WXs3aCazzG1lPIU5sG5c+7hI5yuq7gcLMt3AbJlLGxr/hCuLvT
y+W6afqqmTCKsOAjVWK3Kr6lgvOFWA7zYdhtR1UdE4sUMjEC1rtRh3K2RXbO1BYVZNWqk6NFMLJD
Q5b98obwfxPs1/7hK7Ir7P2XbscljIEhabaXIwopbdltr78WxEBq1B6V6Pl9ULm7W9tsBXdADfC3
8VsD9lj6JRRro7m2+Fi75zILBXPzmmgHdRekzR1JJYB0ArZKCPs/jJ0558ZLiXJrHROTcnNsIBXe
zBjp+oTlcCUukSLN49x7rTCovvGg5kV6dm89uSQkNcW7zZY6UHIH//pcEhTU4Z+EoB4OZf/7U1g7
QGBalw+I4P0CbZjf0WKf3FVXjB5p1mCvtVuIttKip4r4iJ8thuOVwczPw3FxdHKz/bwjm16e8qP7
P0Bvj+Rx2msRunCWLXU9SPiN/FQVJ147JHvvVmnaztEnVvG7a6opqC/DVCgBlhdcGWZ1MMf/S09R
f55nzpJ5qAWbUnsk+2HzvDqRd7FTslfDQIHRRwHmfdhFadH9yz2LbuYDR+vEd5VvXHFBfiyz3d3O
k4qhHDuJKeXphes5FndPOjAhCpUICKib10kwTscTLKl4oNL6JWS1EzQLZeQBuNIn9K5LEV46qjDZ
/JNUSRqmpQpd64OLzs1O7jH82av/Mp7T/jogww9GBZ6ghJPeTgAau6PFsE8RG8UZO7wAd0MXLBST
x4FMmGl8SvJd46baZFqydupvGPSjc2y+w+WOjxpoIykeX4wcvmRi07cjoKWar9I7T/ffEA8Kw3QK
+sXRSkn7BaDkuPZ4yfhUTBkl9fvvoQKJITx0vAQDKu+vwYu2Y6EPzBNGXEU6n5ZlcvpXNEMeGN+3
9Ks0I7enAlg719SKghyEiKk9bD8XhxHsoL2cz89YwwLVwseG4G4I2CDkV4F0R6BS44XBWoY+tUAx
Xfpd0urp5fnJXlQoW97BhyI1F/0zKq3NTl1rpgKzDYObfb/egd9Ufd3lhWhcXdwvb5ex/Jvsflzp
fauXIvE5kNo0TwSbJyp7xndsUnuxmgh4hou8JBY9ThY4M4gbDu9/uHnfzr2Pg8KMCy9D8fKTaZIO
QgOlE214XwIvS2zImwBo2RiKrwjiJMNitBmMTqv6QS8mS84EOJx+yMPXoOCsibcU4aOokK25bWpA
LL+VUjalH3AKdbgzCkbtA8YT2O6fXqpr706q2UQINiFd9zpW2CnHwc+HjQhnAfFaixuH0YRxJBKQ
WzfUGH+76ineawX8HFqTpYlAoyeVtulUQt8zRGbQkaZQJYr6WYd0QgG87wiMrRCDp281O9hmRQi7
qkz8uz4uhORsPqrgGU6I0RemQ6akwGXy/87YNhKJlmS5hG029Ow9sLX4lU5VoS4k/PSvvOrtzDwO
FRQFsRjC4IXKJAVg4iLRHRgZ7YU1jlg5KjM3delhvfYFg1mzuv3ZxhGgheFLlPV00diVasr+UDDS
0tVkCbE3YIxakId5p/oteR1vxBpXXjuM84DQc+FThxkwkFnqu66QEcQ2YPum346SlujxUrabFSuU
Dc6wBga+NXGnRDHn1Y8xXjuJDr6EG34cyyU7ZtpTj6JHhm9Duluv/DlnSa26t1MV9fkbTBaRixKd
a5BpjS8awX5wlGm5d47ceGTEr5kc0+OOjUujwgjGSrB3OG2uFFNBX+d5aGVY5anW1DB1DOGkW8SQ
isc4t3rnT+k9Gu+owd0TNTQtTNEM8FW2yOEpG3NxIjnSyVS3BpLShehG0gSDZKJ+lVU1nSym2Xcg
cug7td7RMBukVpeyl3yocRcI1QfTSljY6UhgIOBKkn1pFTg1Gpd32nzYusXigfV1gP/Hq0hla1aY
9QaF6W8n713Sr7Qszrj7nse0MxOI/6gL2ZQSPMdnMgjpRjCYthS899SYZaNo4E8MDHlTnBkbDW41
ilCOQcXE7qKwPRItJfBWuOHNyh2fxJmL91o3CCvH6uzlN/Ccqahg+4nlfrjQzS2pyUp9X2NKVUOG
gs9E5VJ1vK2H7Kqr4NJcF7ss1kD9EQCRf29GG0O/onARd5W5b8cpt3nZNJL/nvrBVgAYvKkMsz25
0TEKR32fiTh01dcia6kDN1Hrb3Ifv+/zNC1yH96NqgmsgomaA76GGEILXi33B7DMVbvWybeylrVM
T17tyRfoXtn22fwprJuBa3RacxYsfUHatJyIbztCDD3z++oy+E1gtjllymFbH9lrzHXdTCEAYc5r
TmDGAqWDSOg3hcPE9b97IJuSoIUFutLfU/9FG+Bc07sv8qVnr77eTzrtuYUnNxzCUvdRFLXpjxF3
JNowkM2eyfz/k8eLjVAfvQXy/6JWP/5+Unr2UCeHvND/rKG6kVvpVCcH1M9fshWMAMcnCFVL5UkU
AA03RlVVd4Ul8VjYQ6/0+0m+73FZoYcCFwXeJ4VJjCj1IfTPUVrlHFmiA//Qoow8cMklZg/W8hKC
iNFOqtDWLJBo9p2llamroVauIvuXI/Qs7/hnxAAajHRRhzh4hWRs+uM0XcRAThcTI1ACL7nFPFEq
JcI71iZ70+lZsrxQane2j6vLH9nhFG/cxhpkdLrkKkDZMtj/CSGYFqQAx66tTenhqXO2uP2VgAKd
/sINCTAGCbzc4dsN+j41G5YDCVKc/jhdulMLOHpKII3+ZavJDEV3qVl+fPN6fKnDGpFvghcbaa4E
rdB/qSh72hYQ4RPpve3c+uo+t4LOXnLsH+hI6J4MuWClUwksq1+te1fBz+dCSsrqBEa97vJkEZPS
I+yS0ALx58bZb31hXZn78o0fhMhBHoYpSUP1ZWyQMo6g+IutFu2YD+7qWQ04FlkNQEVvOUhowhpp
TD7LnZeOesWGVyyB/oJb8cYaY/S23uL9DYBa6LlT4BxSO0mIIlbNkDV57G0MJo2+7yvETFjxEDT1
sPk33BGAzc6XVnfK5+Gpl90h50skQDbmYO3xvnZqEf1cEc1RPVBx6ZBX5O3hupDFeT9dAArvZtre
dnGLauJx/NwPFJhHHdBVkNMY0OFh27fLBVD9A+WQ4/mgV0w91O8TxfoEGd1FmQG3kWTKZxEWRUyB
UrxNsz5MGYJq0Q31fihTqCs3XjZ5WXPFwPwh3CUoemk+En8MP5kS/Bvmn7uNg3b5LeCELOkSNiuY
J54IqVtVH+h63fg9UtaH+NR0Jo+BDpfqqGwJXwMAQd9sLTuKYwoZC43RB/oFIKvRjE66P/vO4Ava
8+7QMDs1PLyBJ7tWrJKzpFbuZEfF3B/TMRuXhWvU39oVu6Q5+M0fIpgP7A2RwYOxIx55ZQEK2apb
eXnV+7qKUkcW09tZCAN6jIjTZ9JWacq92y7kwdSxRvCDnTb9Vm8+yV84fUzQ2Ytzrt0NyNFlDIYM
XVeY0IDvZM2vRSH03ztW0W3KsTIoDrXcxZQ49W5KgBpSK32srb2S3VEVTVva8k1qjuCl6jaVvCcj
o4t10zWUuHVCP93RyD1QvKMQOmiZFoIy/Mxp85aKUDlZHSl+J20GhWdpCki/220O0O7wRw6bSyfR
kMQpAfjcDkjMCP20kld9rAkSC6cvmqNRiFy+tO72WdaFLe8iH0Y9IsqT5jtgdtsAcyWCEO379j3v
GXmuNCCH7cDMsxhw/LTPEn7Lu1t0e7wxZ/REongFaP7ffzWp7yShZozoD9XQq4JRliufBHmH0q+l
IFUegZ49MYPCdx10URwHcaLWBtrqSpl3xhqVJUSnY7tdpcCtXcCE9yvR+qjhTJ3/f3JEo26HDC9u
8xBaHncmJ1gBmrhCMAISFIra1+gNAJwJiHidjRPvYZW04drWZ2VXPOGQahJRXmFj4b53KTwSDPzl
tnmbHNymn6ub0r9YGRs6dW10oLNMGP8R+c1c+k9JqkUQggU9zrotN1/KD2TjMyQz4ts+WWasLolH
FpaHlrWf8y2RyuIYwhrZkpKTnOx2CS6VZg3Kjbgbsltu43CLPctla4lZ/BQeziaIPTjLBMIgxBeJ
59a2iXlHz52LBDjW07YjnW7RMIKIyzWOQrdI9EGI1OjZLHy6E2fhyTmkl6X7ChhZSoP3oZkeInmM
HMrMSyuSJDOqDRBDd1RZR9463UWNrT+NngZq7i/8vOJLDd72gNTdsr8NoTKJTfIaktSiuMjnexSk
0/9Ywzu/Po7dwdP4a1w3GmqTlEsC6scfnzf7KelOZ58N/i4uvYeQGxks5q1/TbPgEoh9W1lEfiBC
sEJ/8SHWMZad5S+KQfFlu2Yr5AOaQiUvAZKEgjLLt0MHFQ3ZcdPQJawrVax1KIrBWz1QWKY0YMwL
oXL9OVXSs7bw3zNZZ+4/D/4a7eMG2JuRdkJaIPAEQZlyqFhv+Gza1Myb4Vp7Y9x/dBFmwfxW8Tg7
rd50p/ip6TSqWX4kKiah7FQ2VH3lFASfhXwy+/ZcxSjbF58gv3baMddPvaz38SPqmOB2hJImPhJT
DzLJ/tWM01GcpEEZ9tPW9DaBoQKOYgFGyPmnhTzwWrpy3nnP1szoAhaOPjlqL3dH2FCbXCsUssoA
48jcApmqKYE0OY+mOHaZMFvM3nLc0aNNQSPDS5+klTyV5PXQ2kmqGd8KAiN+LUrHNZBOr5t/IYMh
RSs/RdlWxNEVwkZX8k4zh94oC4FoCZECkaqBUuFSXcrSfeEJTKRQKmLTFr7WRNF1MRlPYu3nUPaf
/09ZQgqSvRmlbMK+csV6mPrFz8FJJvj7HfYZPoUEbksEqijtw1JU3BgHKYs7KqBUFz1dvyjONsGZ
HQgWtyTYhsJf7yESvjsTQ0oQJI7EhfAm+2wcpUT/ZIFJVmLI5phCj0j5xONgYB0HHFKEQnBAC/MR
3Avby+T64Jutoqh/yaTOwjkhsljKHlfR5HUiAuFJm7BW5HXDMaazQx/ihE59vq3Fzr+9NxT0hD1l
LpMZeEb/vdWgCGn/Edv0xr4TZ5cwTHjR9UnFAZg0H0OMb2ANKoystiVl2Y/YbDRl2y0IBu03RbqW
G1kt+YLfsWd6HpuZdRN1TKR2z3rGhZUIxLMcqFFGbt8B8Bjeb+UyEpS9Z2rqomKXM8NrIZwCCT2D
Eh1qmKn3ZHnFL0lh8N7Qc33Zba5OzHfeYUOEX1Ad5i8dx7XIuaTItOqhi/8Ty/AaesYPwwpOLcO8
13+fkswHECGaJ5hs8+khNLFuNXrCTsN4qdHE0n0zGZ2KGF4b6o3AjYgtF07S7VIcZqugMs2P8Xt0
z6XmZu8lQ54EZpAh1RnBunWL+zuSIFhGU1ncJTLCyontq9jPGQwwA2zt5N+UFqfDtH8s0IqXINQl
yGpUwuhi7hFa/dXqxfBdEO2lHz22Fq9QqXhKPlL4kdZ/jjhQB4OEEdybDnwibrdMzk6KzueUO5mW
LoTOxHIwkDCC52eMehF6vUpitCVNaQ4/c92JlQL6QF7rnVj7+FO5/AF3DfFZ0tnzd6CDLHpmNH3F
KQ7Vdh7ibaz77TVo5srhaO4rIMkh6PYhXqKggmdd6mtf1ON1BJCO/XfmD6LRffWPiA26/FQEm0Z6
P9gPv+1ERi8OnD/rkYwkokgDDWXBBXIb9gRzY6eETeqm5dM220xY5rILz5kzioEtYG5vggGQrsfR
9HqM/645b3n0DKKXyM+WHNJiyJrUVDu/B8+J2ya06NGWTWwnBCeNE6Lqi5LPCVE4wOtvHlxnv7Dq
nlAKspgvoDoqoEoci1TyU1bgX16T7j0bHFLZrzR0Icy8/jw8K01nTudekzZJ4xvcFB5gIxyXdZTf
du6diUJ3liKi0MoxNaOZjHuYRGqpgTd5aO086eaPCzNkljjTq+BPcSM8vTXdKQcePitI4z1OfPQ5
o2mvev7aU5h4NbRIJ9UWgF0ngKsNWCyyKOV2bqIrta74Oewqc96WXz/SYBQ3x4MhEhi9okhg5XM4
Y12LaLxesblNLzIqYLcELCa2skNdnnmpWx+X+NoB2X4KJOb+O4f8CcduD8fTTB8NSikf+AWF/KcD
+g4ApVpp9d/GZzcJiTqsHdjxWGW+Mqlr3ZWKJkO2+Qz8ywpqjpiWAXWF95xyWyVrJ60+hG3qdSrh
Gr9HPV2MFAvuCCXK1IqtmBOg/nW43h42QuqAQfMbauv+QK6jlwNQ+MLnNxXQ6GM/vD7jNueeqqAF
yEnFS4znr3t3Dom6DwGxKhxJ3ChFxgysNgBszUWk/O5+RKaXt/fsquNwrBGbbFvz2FQIphmFLSaF
u+j0OO0PCxw1mUtZidlhGDhNWkv+fef4puB5ygwjeI7jHT5FU2qy8yzPMr0qOqFCJC/Q1U8MnfD1
2NhspTr9JTEXJ2Xsd5fd53FbbS2J+aqeHF2X9Te7BC3b9fr/sy4BgA5tpQ0jB8aPSKRLwHQSzlrl
xbLOgTZOKoMmTpSmp5k72eq1LJ5lIqRKhd1SDKUME/G6oIMrjaYvwAszvzl9wiHNGi4rkSDoraCC
rLH8hvS58jHVOrjLSK0X67LClUnoKivUxJqUAIvg+jECT3ZiwpzhmTJ4RCva2io/1HTgifJ4I1Fz
1dy77IHxLFbZ/Eu/jmim+swqJj8v1Y6Xb8bhXVDCVfqAp3jtZ6H0nPDr3RFo0FLI5YoQyKY34vgM
mKncqoBOmP8zEjI8wECcvf2VO7KjZhLqA9Ed4V6C1AzlX1f9/y2Q7lKxEBccPK5BKJqNGKRpOVEK
7bn76Ky/JEaAmwZxkkKZDxm/J2vzRlmt//PYGeycCoXqCJN+TmfTDCNW3M3XDlPAeidh9tiRmFad
/dicQRqkoseBHrdd8wsrwg5ItdQIgJ/P7/nCIUj00XIcmCtzBKU+yaKc5z/aYWCI9KhyxxD/KwP3
fgdJMBi6KSDFTAc0I2v24xr705Olfu4HPcZSV5oAxGLUxWV7mJyvtm3jpleLh+p8IPO1A9p0XOdQ
Ss4FEsX3hGFRbVN2i0qsCJwKSS2MgEO9uzo0BatupeO7kMZf4V/3tVHW/csKTcHMkF9hcj0sfmDQ
t9bnJHAV8ACNgN+VkIQWTcUONR7p0ZS7HlXQ0JZ9oLqAuiguU42e0LbhNPRqkG5M0Ia6LkQvT+rp
aDkEwrM8o0JCYahjpp8LM8cd150E+sieBw3SPObliHZmD3NxXHkALBIfo2cis+xl4KkpPU07nolI
PB+KseFibejlFYt1YoIhF9EpKHI6c57KSr/wXio3Szmu2yV4E6N0/6ffp6QDc85L/C4ZrTCnESlX
koVjjMzlU5j5chnMpHFAgSqMxzaEo02+QO2704/wdxquDLlk/8ZUbMj1oe8elIh8KUfQXHuNDPhh
cP9dtpLQTUut8SZfTw+ne3Xf6D6+wvL7HD2R0OQ+vXqZPxymD8HR1bqN+3TTHNz9KJP6qN1TB5nF
55LBSj9fbs9/O5miuI3I4OPsVeya2c0EJjQG3Q5kfeVWgoLUcRc0409/IaVSsEh1R+3OGbvV6kyX
BsLc9xgKO437wVyq4zTPH83zN9EijPhTwJn1hKdCx1P+ufFsxkXL1N02KzEibsdMWPAvJy9MG81B
l93sDpOeWbQoKUwDxa0DjelAoXJnYmJ2ZxbpIAwCqEyZJxmxs2mbf27aYESTa6dXZUaYDp3R7w5t
IjEzxt9k8uIDTe/uY91Vg6vS/CM2aZzk62Io4goLVM7nvw9PYzv75pl1LHcSATrUNT7Wuc89v6wK
fiRAg3Ahyq/ehCHvLHeB/PWFyU0W6TvuhqprYm/Qr2bd3zFh71MYRD7aq1F23f0lNZjPVCUckhxC
mQEr/hytO81w/05ha6E+2I5NDmTgF2NsaAfB2cmXImh05E79cGjZPFhRcX4/Sbi+2fiYRM02FaO+
ZtZYvdOwrMcG3qeuIxaRo2iL6pVy9hfozKiQQHVzXVnqMaszvpw31XhI0DDD0tOwrKKILMitZ48B
atLRnil7oqKaaCj2z85jYm/Swv00+IEVnOifrnUwRBdSAZwoL3/W3dyn0T11OAysCc/cE18/OhbJ
E4A1WJ1YJLH79bok9ssPi2tB0cKcNKo+KyV8Rf1L6Cg6ex5KikQM0K3XyOHm7wD3NXddiKI8fTAb
K53WqlvP7zGcbdaLp1ha/GmKqSnoCSYxlTs9LmXEAyZEam4uPEFFOnn8S91lbRsidtXwjiKR/xxX
d6HiH+QG2zJJ3iJn4LE3z2TeO4bntmLOJZrWspfFPktyBk3GC4+iVtiKwZYFt259ez6VmT+apXpT
oRXomPscH63NLfezTFSSK0ppxa3OPoAfukqDkx7LLDC6omZrj86E5xRvjgi7V0cYd4uuawu9RzKC
Dk4I24iMmOQoVBGH35AF24kFhmK0/gsH4XU22iKsDznUnPoUZaoTo2+oHJW9p+6mFIML1hLtrJvQ
GmcDOb1oX1aIrW1uRjief03GLTPIg0YMyOiLAFPCqIB6vNYntDNHKAuFSArMBJrIsWYsZ5Y8DtRC
+1eix61Knk87Lt0+6KNR2qEQ4rozl3bBfI0EIsyoDpLh/4ot00k9F8zy6qjA7VlWlPk0cMHKCZV9
jpOOuUM5mIJuTaqxSQNRRRUByrOqaRQNqVWQubMyJwMtYfI0y3//m1tLhb+YvucCPvjHddsi1dQe
xQC220/gZCBwYITzZ8PoBVqlZNwoDBJCKkJuVUA0a2x7PspgDHtL5X9Lj2MkboUKup59c9OzR/B4
3DvwUPdKtYeoFUDVnPk51fz/V3fQC6JeyVKoqXy+MsCBnParq077vyWFW2uP4/CXKqc3BWEC9Rog
YqBm+EPwzOav6yqMIbgtWpNk800qFCn46hStDr1SfsWv662WT3q9dzXNztmvPuTail6FxaWfQyK3
2UlFPXILKJnc/7BzigaBaxK1ob1b1KNu8XNbk/0Ava75zepD9+9Gz7f5TR9vqBAlahjF70scz0xY
J91dlLjV2c0cZ7Ug861zghl7XakSFVPZMucSOaYHLPK9nXp1ZtqL6Hqk12ZCUHCawXGqh/U0SWZS
rF03R+LlOu8zn7x06+uq+ApvX/Lhk4GVZGyQ8JlGihdHLyHyAUcJUmo4H/l5fMDq24/DFAOmS6lV
5ocfVLBcjOvftMIb2ZoY9FM12940c2PfoGdDCqSctYes5g2nk35vYX0my2bR+iEI5UUQIXYhSxlX
IE3EWdcP7c+WMkDfgujKjiu5pFHnibGsuwv3bB0m8nwae79x8vRxCrqJS09rMZgUVuIQeFE509Ou
ZsIimJAAJ7iyQ4R4+fwVGEmCSsE2kXfyJwRiMXosAUT94RRS07pKP5TjnzoOfDCcRoGKdsg63/QW
efiOMRAexiDVCRnGflqDwYWLBaE1RYRg3cYxfymP/4nbWXyr1xfq1FzKv6IFHt6m/Euj0OOFVllw
hp+qsTGCUp1mzcCusJ4VO7ZTdtTQwSLZ5LRYgF8p0WkS8i7VvGptLb5IZr7A8PG3GoZZz/X61qCt
oRUhJWCeki7ENRSZuZZLNVOVDZ4z6L23ZyKBS5YzyH+kCDqTTNI64e2qbyQaxBzUl9SEQJ4ZsuNK
0oejuwnoT7zIb3kdmXYX7oGxfIEYavLp9v2MwFbisl5FNL2/DiaKfczagWrM3dgVoTRXNIL+OF3y
Lc6S9D1lDlYdb97vgiaPdGOyhW+4OkagDCn3/pHk/8lIApEQuqHq/vOM0+IF+QLZNBhZpHE/gN+P
E2DcUhg7dX+nVe4zjCY6jeToSLZ0vdVVFh9mwTh3mnWzNv4pWmifjuJVPc9P4FXZI7HFvRQUMhAV
IoHtpR0OIvJD1xhjvsb2Mq9P/vW1Cpx1xd2lx/vzO23vcpzGVPTvPt3QivHpkEW/V3SMRPHTdw1t
xy1nPWRFQ39XIdCYqXGpmBnbzvQNTsz4gCChewRH7tvvny43Sb4lMGYrUNdxnBGyst0fGx+TM85f
HYXscw4xyBPg063lZI9LJ9pKC7Lvw1cmqzyFafDOFSsFesD9i35lNUZILO+vSyxJtv27t8go3t2P
vNSHfwxrh4T2D/b79uD32oTNTSX4x9q4Bj8Sbseo5dnqZWQDGZYhaLhyZdTODHcbyX7esiFrfZU7
AmVK4Qe4oGsBdA5/zLVxskrMdgALEe2sZDffS+v8qT8K/Mu8tfoP6EneJMQAlZkI584wY86GtlfQ
XrqvnopGn3Jf52nTLtsIaao3VpJdtBBf7kRx4Rg5WUOFd8tVltGsXvAlLX+zzVQpQImIBFzqJ8yg
Rtr2vJQt8RMUwNMeuYxzTyyqR31lzPiwx/FYp26D9FoHLZcmclFc/B3PEdGmO+cXISE6ZjNTAEh1
+zszMAWowVqLqKdKFoeHJA3Ykr9kw3yK+xocsBdnnhUhGNZlEomSvTUH/CZXATrLrvnd9dgv/JYU
dbHYatakp0fqV0k3TLelOECuhReAC9WVPRRa7zfNIeyHn5y+qIDLS3AqAnY2S3+t5XGMOszZWJib
P91kSuavKpcarDDtRwF3VbUtZ6Toe7yEtXf1xMNClJIv5SN1lmYgxHmSjcUXAbt1BLZkkk5rSutR
kNpNBjsrhdRZZDItxkR3k9ZptEu3AFX91IV/b+Il6Tehr/YF3MsA+HUYw7+RwihqEj4/JikyuLAB
iy2JvO2iL8ce7qcH/XawahiHw733+ydKeJAQyJ9xEgV6fGTJJMltXGINVS8bPyBi+UIWS0sKuzk6
n0SnHXSO6eaSe1+KtvC5lfePR6Ob6qSoQp2OI2e2wmvSNgcGdwYTRd2TidZSOJgzj0fkBDFtSbmZ
zD/ATZv1VJtLAMijz8Xo2/WgwCFLohHUXlJlXcSFofCWsLF/AK8azwFFTqp7HHMkJNJvzFxkmCmn
7b78a/JRC2K/cKvqwr0cXf+usSKqJjXRnOpv7h2ynYcUEN/RR3xdFLnMj5BdKXcoQIjXy/il2Kor
GO+ugZXpDkW0kBhXtdOQo0jku79uxuHeHQZDO28Mb/TTT9qjbKIU1xZ6z0Zib8/ms54wE1nngYQg
UFtTScAHuRTl1EbtPhHTYg0/DNNeD/nTGiuM0zTCsv21XgCa/JG4cRMDEKuh5Qk8imAqtfuyNdQF
/UoKfHyIldOMZlru3ryylnegBIf9rOXJQB0jWrHf9ley1cfAu7R388+I6/lH6Q4IWbNr2uA8dBOx
Zo0HRv0pQ32Phs1J4z9/Fa8vSLfZdZ45ABf5+4prHpuMutRFLLIhzvL1Fuowdn6N9979PCNlGXLx
X16c4mNj/F/taPq5bOoqrwuWs9DghcMO0C3ttFYjh41xjeivFqOnym41Por0MfUvfujU6rk7NDZU
RftdCFRFSCYeTX0iIkBJYCBWOYZOvGTblcI9RCmV9bZhdplW30J5CohMQkKn/9YqmcXzZJJkmXqH
3e+xarShPgkgVR+cf17DrZ3TFQKuPoSs2Wo21VyPbYWM33IXYTyk50KyvZz+n6Sg5ZrUZqwCQPdl
9yrvkYNUMBBPYPTZBupDufdVdszB2EXL2zwYWrqzOCb3Ubs8jouvmXpO4wqOUT/uXneIM/q3lxrA
ptbeBxX8vNPN/V2D7gt1aF+/HvIvgIp17oknzKceeJ+8CuGGwixjY6JHihKGlabzwfNja0oa3LQA
63RMeB6+8WE7TKmqErnZOLcMC7RyvAa36/hMo40V2Jlh2h6NzBrP2jSk1pgC83ITRPi6oSCmqwpi
XP/cJvXKeplJ58ffQf8IScBTPGbWC0Lf/oX0P4Cwkl5bYbwI9BtbdEINa11AUNE+raRteu7nt4Hv
aA38ndqSBHqZWjkcHMFCgy043CacFpJ+7WC6xHUkHqsiBUD8KM2wcceBSNgc/evwhEfF4jk/QmZt
PWCZZb4KXcyydbZNPqRmcv/W9/YDX5H1wIIie1H5l/27fhNz270xKq1boR6t29wwXLOcZ5WBdQe7
b98xO6c3nqtuaQCLnq1P8oxfcFzOvp1j4BdRJLKzz/k40jEX0viMMd/jv3uUxedTZ1s6k6AfICok
BUDs0vwhSegre1OcjwR1uCN/rs0wo1B88iyTMRqSSfOd7y0d55UC/temO0ZQ3yO05gLgXH9j3gLG
9h86Bmi3cpUy19sqS3CVzfPkR3CZhQcJpNvnTVoldOgSY6zfy5jVL6fZLv3ro5YE4F3nuso1rqSB
KIK4t8bg07qZ5tsx9hnoazsKz+lPwDhiXgSyiY11rfh015jdiX9Ex5cmBZ719cd8AdTioeojVuTW
LwISzM3AYam6FTd6vKjHzEfamFHL0WcW6o/IuQYObjgZPAP3zdrRPjbrJD1HeBl+SLASdYFFLS9Z
xvF4aSl0vNpylhOdQICIoKCDkNcuUlhgX41HDmwVm/Yf+fVF+DBpMiQ1E2Et23qpyn3XWbmrRUHi
Dy2c6EuihQ6Hph++Kpksp4kzEC86CFg2wl+LeRIJujW8hsS1U/tr3jUE8WIzDCI0r+NAis29J8T1
uRIQQYJ8ZVAUieFC3W02ZHHgPf5v8107+GDW/Vuas8D0m2yoAlArJFhDvAPd3EgdH8KyfHGPkXRO
PkfJ7V23jpc84Fxa9g+EwAg6VZIui7FC0Njb5rXSCLzvp9lACZutbZJVnT0Yc10QbK3qlCNDJ51N
7CiOEcptOm1surNkp8OcTsfG9f0/WyWUofqiUCpl98pBw6sLaZOxc8gmyqom+ALEXJuUGQlqaPZY
Zse8jXlCZbKyw/6g2Ni60+MtC+O4H1kVL7qQYFcOR862T4XKxkcejbPA/4GHxjWZhH2hDBroeMKg
fxnIJI6dnrRnmp2Lsjfz6NHkEnGnEwWrPUL4gYDpYEeTRdjYuGXXR4jgSPKm1ohRWIHYyQ+mQvJL
RdGq9EjTQg1+hQD6SE3rqyxODDoW94lzGHa4X5L90Pgm8mVqwC0uHlVYYVXmVj1zITgtwuZnGPhE
FsRO1Df16KYo39C0dq28UXW8YGTf+/n0YTmve59MfX8GhrppVG9gxNAITyqq01fcBRZKATRNjYD8
A/T+RERr1+DvG3meg7qiy6rGT5e+tNfiJ/7hg+LAE1ByxTiIhdTFv9WRKRGs9MIHesVviToJ6bJv
0hqr1tG+xY1wLYbzBtcRBKJBhsDttlLuGyIgFQfV+ossEGN4lgvtxF8VmqGgP5LOyUkaNw+oR2gR
edsbJuWwLff6s+m3W1N3lDy89tUc3wBjmT/VBilYaXd4n8C8T7urMfz5+xWgCqjYXJlzb4CQr66X
awa4ZXGAEJ+G39oKTJ2W87FKldjggkEDV80zgy4bPl2o+3YRYy5RUqHmQeR8665m88n+TkVFaGt6
pK6XuzaiQqMzLnn9HH7nYi67B+r3PzLfDr6SCYqtG9Gewkj1x9c/Qi3a/+c+Qp5ayg6UtxuSlTlx
RxRjLKCuGzYzioXhxExomXVqjY1ocEpgdlYE2JDJ6Ks2i/N8dyd4tigKUC5oX6DTcBMGNLR1f3gg
3fgZc9CADl+BYqPKLxPWS9ZKKU3eRX1CKBETkBvXvokH4zluTyM73Ej+nLXY9LNrEFlsOpFH5k+u
u3PTeJnyWgbbb82pLQKFAJeQsLJCwV6eqVJlsurdrYPrtsklA8GeO2G1bZv7KxB7dK2jO6Ps2BmG
tohBFtit03lWSajSbd6farmHJayCq2AOj9UIJHsuq3YzPHgYG7By7V6usV+u/VLpAPv06WP6EZrY
pJ2Ux3qHJVSDmCtJyOrGuRhmZGZt+rPhacyGVvoifCIjT50cubwxkPntFk4MZMZzqwzOHxZs2MID
xFIJaD+znv6tCQaBBiRLtLc7vndsgGeQan/6nsRPIkE657oP+lxAmzFVNUAOy9E1y6kGs9ejETHR
/WbEEIOzyfACdE1C1ywCMLHDsKxdduMwFBeYXE51kAJ0npMIbhp2JxCXxeNL0zi9fS3xvBJUQ3ZL
8Ac1naU9CM7GbGAB5R191qEiHe/oJMDekEKS1cEbQlrlC64I5yR/jhta5/nwbxxrVHtAuZ+ygD3v
xkkOjEJe51ttoil5AUgS5oLmRK9Q1ahadBRPaQELaiAjtyLy9wxOd7+eUCjCS2jIAwKtnosdyL33
XMMxxQtWhzhUQAxs+OE29VUnDR5M5G/GQzjY4UrcSxUrLWopJURcnHYS5NeqGqRHRIN+TnHAfu+Y
+cxQN6jyPQ0QEAHdJBTFUOBiurBC5x8dvRVBEKOk5VHrSBC/TE6Jnc9hTQyHVuresfqYH+1qXfpS
+8bBi0ASxe/QZG/tFIXemPG2lL201e/ZB4xVEkbWfsBrRxIADd8yzl94J404WfP2RlRIheZttTG0
7fIezcLQzly+13w1u1kguVyUzNtCu8gtZqc7T8f+H+Ykvt2oJIoyEU/XyCVReIetHwzIMCSDaFDW
I98FNDZnsWcLoiTlccxuWMbcr5Dkw/QiIng7P9aDhNQS57vBK8VdZjJ31zsyJ5i+1yI/cxQnVCb5
KeFPutlw4jAYUqPTP5j5CJJlBq6pG4j0dZX9Jsficxdl+36GZXPNkaiHVWfqStoGpNZhEMhxpjhG
sGqduy8i9oUWuff3VwruYDQeXpySZGk3tfeEHa+rZ2DzZ5lObBLp2LfDXIVaWBe5Oc6TEVz62/UA
qV2XmKLNKL0MF8/1FOxd/vLQyqU3nt4X5HnREPlCiG5zynSN5HoNxWXhYPx2InAy9kjnp5SRiEQK
+Lv3tv9FYsLisu9uL+qGpSHkYfDPZ89W8OphSaiCROYxba/dl/H9uyRhwdbhn446vdSH6EvC+yH4
V2roQ1P7OSn0Ve2p0osGbi25i31hPIc4KYQs1pD4d9tjUSbm+X3VmeN/gxywn8+G7LeIZdajSUMC
Y8SrizD75YoFtoPo1F2riP2F+p9MfUfL03o1ip67mF4mOYQSXo225WmV01L9g189bIkVvP/R5URX
gi1RSlQnIIVJnSKKHMheqnBh5SNRkf4qGXM+Zb60YKaXMMVtDHCQJYxSyCdFeXC406AWr0xpZgCq
OOEjsh2pO5NIXFXYR/beZH53kjNT/hdaTZHyyJCwyw4w0VPrQlV+TtZMU6T/avVxlABLU8L5MsFH
5piPPjU3skMwyUshhBlkwcpYczEzQZqkMXtpF7b1uouAfXm2Mul7GGN5jFKaF8YOS5yHPlhNjpjz
lwnP9IjmS9khsS9FVSBf96hgzpzNUakz+4A3i9Cpd5ZWvvnnKHWhO389acXflfIHrfoetjM36VYr
inXhCqFtjGBbr7GCceXoMjj3BjCz8ZMeflBXemoB+c10nUVMriyH11ez3f3fEiZ0HQ2TESnAsDix
uN3r4TsacQZq7Ueug+SEMzWvrX6xfdi9MwLUuGzz6Z54UhMbZRNWT/q/QHXKFAD6GT+v5FwGQTJW
rj8XJvYjDmaxyl2vnqvJuvVlB4FjkTEoAIUGwWuDgp1Xc6iNvSf91eO79dKEmiYzxoKLrIAoWSmL
BVvmKfmYjWXelx+qu5jGEJ3e8phNVOHLO+TKMarM5RqCO8o6QNEqZ4Ps9b2B0ZOJ6cb0Rzys3rY8
Rx16kQMXwCX6TBME0/e8hzlDW+wimcYWsds9pihp++A82COjTWUPd2QlhCQEvZHYaFYgLhWOURQ7
pnhAwRjMVBcB0fewIU3ITRX+GiWyO+Yin5VBlDDaGqIBMM/b3Ni4QaJhjB7zuqVNGbNdmUitNucb
eSlcE5+fAL5etHmmUG3S8Yk9UgIbLrCzNHL2EoVJcjF/v8c8quaGJsxJZUtyWUtqzAa9SSmDknav
PhB5wW4paknVdMAB0MO4mo86cjMiBkFn3koKAM1R7qFccaxgg6RgAV5Ws8e50hffTrok6O0stxRA
iXjWBtM7XH+3V9e54OE14JnDY4fuMC8HjHcVf/+Gv0kEHd4Qkz4Wl6ZszfaFiCBBCDSZFqlpwTaV
sNK74uyHVe1L7f1oY/cEMu6sp2CZxP+8xonXA0GCgx5W6zAhS+YHnw75+sxMlz2+NnuV7TOJuIEG
2nxOKDHO47WC66nrrqLAI6Zpw6s+hoQM7f98mh2RQZ/27IOufYAXoy+AeCgir9F/w8LfC8pPQi0P
x4LP10HU5c/5CxAa6//HIlFqPf29ed4wI68REcVvcE8YjmzCFir0KDPObLhsRuDyxn1Mqs+OcHdv
/ua8IzaCUmYCF9txhk9N/M61x4AgxLZILAFq79H24G6ZzDb73i/fhdEpE9NiQXDKDy8DmW4Ve33S
p67G01eCmlvBO5tZhOZn1WR8CP9X1tMWgpcsSPZcwWpsuvPDDIqAfnS+CBJIMECCuUHpz9eFnoTO
g9JZ2lGj/FjsdLgl6oCmlN6m2qqHC5wv1+xkn7Vizt88Pg04wa8WFcaZor7BU6U6+EucgWORmaBx
C3KYFCQtD9Fa/jFIdWl24SAXKZiX5dbxPPoj9svqf7r0Ewrs+leT8mRSnjm5kwiQjHJQFsb4TUOu
EUIEzGpsTdjlc8ROO8GLoFwG61psJ+f+gc7AIKI3261AjUc6JLU4gUxULUKYUx26CAryB1WQp1zF
oMF81peLuG2/4FiMG23ZV6R4acyZoCMWLFG0a/btZ1FJ3USZU1ZF+PqqS09IHl5UK4XuckoYp8i0
DD4rYahlQCPiMM/oC0M+mfZ/NYdd+TPFouj9qo1xrhzDUlvBUaUyKxmUUGxwTTH5G1H7Pj0ZkUet
yQnI1+fQaeOt4PzVeWM0kgnqnJfb3WwCGc2x/PMpnvR/sXnPfPo+hs1yTxGyZzwLhaWldpiC8mxp
2FuyycEsxdv+lDEgWEs3COZtvhtqQ7KfDpxLfjcFUPUJdKVsxQthP8vujd9UWrE/giKuVinTLmjr
a+zwNok089DVfzJ9iczIYFq8Z46DOq+5Mnd18FV1ieC2JilkxwifMGTjDQznz7EJWjE9P5XL4cts
86D8s5LXhO/t3lQfTODoRV5d1k8C+UvJkJX3K5RCTh3tkE/NADS2KKMEbezggpRaYa3id617U+sy
hzTTcFRon7y87r5tyM0x5cgA/1Z4vhEVzhd5AK6tPWm1zmjV6+j5osn7Js05LCXm2hwiGOfqe6FN
XNvlQQNoT8zu9JoaIfLbwA8/heWPrtolUhAJ9/AjcWBvle1b2vT8WHDAbhYjS1sAb9hQbu57SwYT
25sxj1fJd12OsbyQOa3EUArNVInloFJpIO6NYZ0+BUKDqJG2pGWrAXUYYLWKIGB0J1Lripkg6/pF
yeFDHsZreBYlyn7p0lQRHm7WdSXa7kXLBkGTImYdD9ppG/e1FX7fsg6jXPS9IHoqZa+ozAnJbwnU
UQPDThSzoeNZb8/g+GvpoH0/CdwcfdLIomLhpAYPzPng55NaBiNg5iwq/siM7isZoycLZU1Lz8xY
epPu1HhMwgw8jD6ZRw1ZcuqxMOKxdYKi3+HEt2l94BrYOU5qS5ImptGiXOGLlcf7fwM0Oux9v2lT
RctGDlUy4E9ZNnLortYu8egboGq0aJerMKdtzLESDYVXPX9ZD3QNZ9yDC1z0HjvBQLBGSqMrl1rT
jSPU/x7oTh0rkBjVtV436XVxfRQnGNqJYVvspbS0mAEgZM6CbyjnJ5/osqqLmYAm7uq75F2DUVvJ
ZahqUC80hccO2m8tY5KpU8n4rqLOpvBePlq9AsFx4AC5YY/C0TncMNSCuLEr+59b5s9NyDB+TOOw
E+k8z5QDcnvLR8EPU55T16TMMU7i+uNecFW6DHoGQhdylBenB56ja0IVgQ2WyK3rK8NmrhEn29cW
mA8xBPkLOJCGge4st+zIinA6+l7/4WVByio8AVSGZc0w4lhyuN0L10C+pR21Y8OLWn99nbJga6NW
CN51k7Mce5EJOsD8IV6q742BichQwwOXbzVINg9BP4qjbxqzz1GXTKXwhiMyKEgYBuzU8BxYwq2X
/91dfRiuxWDkTWLHj6KOWOAVRwfbJe1kwIN2lzsRUeptqASXhNVHy2So9zClIMLWSCSWEFIF0YOG
IcLudeHtUQNI9V6A9rPqcqC5w+QU94jJkXdQ0XZxXx2hae9yd+jflSqwzikrH27Ex00PIpy+eSzf
WjnsFq+v2mimjWeVhxf5hZYNxUW8YGNSbwBH72mApyZ9Ium3IaxI1QfQ+k3AXH7cvoJlEPKjv1xq
YH6gfXaA4hwzH+nggj37/TdjJpZFTcqvAgkR54vmK+fN0SrARiN1t+hiPIqgal78lq58wTAKr0Vv
eWgNajRjx0BItH+cnLUioFdroRPj8iGOlruuMjY4gbyJ3XXjdsTTmuqJjDxEiW0mGlNQOZOcwBxd
VrY1AX6dEh96NyYNYWvTWDv3AhluEAfSxNwl21k1Fcp7RqnQ4lNoawQYB8DxKwjoVOmE00oSesVk
m2P84/r9ufcG8yKkYD6/+RxWevnsJp84LR1NUgpCRiFZyh78kfUgYi7NsGWyvA4nSw+ab3B/PKOG
AgyWNa3U/MmO19nPvkLMsvjYojBKiEwTJfLw2KT1mxLNFajiDOFNtGW9R8ngH58lI/LrS49/5hs6
iKhVhLw83X/jjsM86IlEy1X+LLjOzzlQrk/p5MwEMVFoTCtRssGEpR5Zy3SptWq1obnLh0ZTdok0
vxRw3Lp5ORFFLrcT6ngm2lURt9VppK3KqCoTJr4L7A6lv+41uTBPpI+exCozfWgGAs9PYVRFd+nh
3lU2QrEw7V/7cUoxLIEeFog60YejPuwveyVajNok9iOn8xZIdfWFSdBpGJf0XvqOTp2+qvgmWmY6
6PFnV/N3LFZmeIncPvB533ns86ns/4BYbqeNHwIGKBWtG5Hyqpik3FORqMwAZjfBGKl9xjhy999Y
9GYmBwM4rV9OuskYtEOB9nDcKEXHyVSGHB7ZUhvUyfUodHqV0dDRCrhupD18ha6rsB5bu2s1v61t
wdc2uQVsp25iITiUZspvA6WRohd74zIxaPASvDwUBAcd7DyV6eTapmvSCv3fBOi2Xu6K0f+umKyp
jOkY30i4LJtPMefysuiQ+TRou+uwUQTV+akazxoG8LapVWmg67/+3OTQUY16+nzuvojkV79KK9Yo
5AEJqdEMcpu7w6ulqo2yvfE6SYR/LUIHmcAJjZ3XlrOTS1pzdVc+4dWGv4z0TKOMcEmG9I9WOBWq
FBaR/eC3VNhFL0thiXevELJy3PCa6KU6vpDyR+PRzh3oriCE1oi7DVB/rd+KKl4qqI5T5vNBRpPQ
kSoFwjxHZ+FSHhi50/aUQbqdvGYYygy3rKzQqcCh/L2+gN1Xqr0zMf/c9vBI1mFejWu7ccha122d
3+rc5PJ9Nhjel6S7uA8DO0eLEMjdMfMxcKWBwowxRehWsylMULJ2+U/Kp4PzDTylTncnxDdSFkMx
Ra88zG5XhfddkDavzFMxLRtTRIkN0+kWLjlYrB4pfq0cf5HICeabsyBHBOQn9HepavgW7ygMPTlX
m4KFzp8TpLUG/b4zjtdETRuMX9dP0Ep1KSGFmgM8hsMbaM4Mdk8SUdC0wma8+LKlJo11NhzGv547
NP4T2iGL0dotF1wpZj26h65srgkQMgEfVk4/FP9nut2bcaIB5sXS1CYidnxv3AJtv2ZTFodnW65y
92rzYSsxayivdqMEmDkIctmX1EtGEFxjhI0zrckUkLGKaAR94fFGnbFl5paDq9Ne0aSfR8Zr5gtl
xLWEHPdWC51FTzAMPvBfiOI053f0+z61jk+k3LIRUFOjzD7wM51BRpEr+1MQUP/2ZPNxH6Wtagmm
UTuMsFz7yCKsseYoSDEUwblSO1ySjL82/wsO9aOiB6rpNmyCjpA6JUv1QyzX1kYAzSsd3FVL+OUB
UHEcK3ti+xmmEarbAR0dUttC12eCMLZJqr3idXmMLy3puoTeRT3AFrO9MYIXPK4K75uvwh/is5Wd
BO5agNuDW6n6jXZlApspqm+3n3ZNDXHSPYIsMsMioHTRRXD9oUFt2PeX87b9B7M6rxDjCkEApbFW
PQc3sDe4IvwMl8LZ+/n6rAQuNW8tRx30QwZN3A2A/b4N0TxewisjSyKySbF0Lrf0pRtQxfJrYWt0
DYsUuZ1K4ezZRigCV2891f6/vTdfEtQnaYCUWnlycb0Xmrvgu3AzPfY/zIOKJUcW/TxDVF83y4YS
iJ3U5iRi+QJZWvyM8yB03ZBGUfz2EMPrYSDTnyGDB9anHp28H/gjw0EMfq+QDMxfLI+qyStk0v1m
Yv5NVZH0oUM0xZRaTo97J+EDQV7WlGypkVVspzUKfcoxIa6uvLR2PvN7ro9WR8Fi70eTPHzBqJo/
CiS8al0XtSJKcHyJzPRUz2Hh45mTT6GFZ+ogD42XHTnCcmRBZl2IRg6UI5Pbfvzpm5qHyRB0b8sr
SOZ6sEtXZmE3sR5M2Ik50/Pp+tnNmTJlSDT2B/7BBpVKWVSweJYEDxlir8suof5t8rR8FCIHs1AO
Mdj9Q5EXhwG/FVIXWEPhHKEc86CfI8C4DfVyzfZ4JGzHBaX2l8yA6P/YSoFtAcfJO4MdSFyr0JlH
TOdeXyjjR1zdlZCIHaD5mqKUJU2fAlZMgFo30kMSskGYEwwS9Ytok/TEYpkb2F7jf2foFr13eu2Q
dEshQ93WqHuISojDdwR+ItCnC0fyhPMe3NG6/Tj8+hH5FdX1pBqyrvepnXd9mD+WLD3NmmiOVRbj
ShL+Kia+sem2o3Y9GvdHHy92fx0IGGOC0ZKgyJ4nNqFsKZJTtOn1tpc/qYFW1hnFrDiMFAj4JtcI
l09v5puzts4TlK9QOpVioW+S9LnRdRA0UPkNUdYrZZ74i8BFnLMKGu9fJVCifuuGgZqVHgacQfid
dE5HWIJqpyOpfK6F8/z1YDn1PBRlK3P2tdBBkzEJ7yUdSwcUGO9MugsGP+d2k7LJBIhk8TgglAny
YLCu8P/25++qKVClEAbUueA4kNwfSpzgaXB0vu6tfggk/QE8yG9h8NOjViznxNXBTjrUjyzGHn8Q
rWn3X+RYB+6dPRHwsCleI/JmPxwbH2/vBvn/reqL0O0O+A5t9zKznvB1M0VH9ADANZRr2gYJTeM3
8Pa4p6nCTroVr6DZFZeO1BMrRMXQlpvGKksSNvKiYEDZdcnrjuluIODSgm9hYtvb4MNaXFHOH5zc
4VhYhCxfc9XiDhLdvP+ri4horprmFwKToWriDqmW5UCw9tds9iiVOcIu18kCNNsZljVQ2PLz0KRp
0WG+p3RXpranTRnrPfmkDvSr4D3aA+VZQYTrjctWWokoud0a4o6+fBBU42oRMyeWC/FnkkXgiVPK
DSFNKOvU2jXdvO0/t61/YE1Gz3HxVpkNDsPp2Liv11Lb3nuk/fuQnRgX83arCRr8MOpxgZK3sq5m
y4Oy9jfSCTfQilBafCZYy40y80DwYbxGjIMIydROQeujGKnotEEJJ89+94kl2Wm60rsjQ/pKjGXM
cNLsJZiRmp07JVuvwmIC5zOvRi9lCxklx3T+gC39p7M97h3TpOJiZVrUX+1L/ZN3owq9XwaDxQ5A
bBFdwT+GZp7bjuRqjOY7cflVDUmXUrFS+tRPZjEud78le/7XUwVrN6ZOEIqk9aBs2GdJWh4qR3oy
ECDfcVmqZuuJtm0SlfnjcA/8pfrCGL+ft7o8fQ4rYu34u28yIXrFe4bJ4RBAAirsxAx1dlyi1+7f
tR3fWtQZRq7Jooz5FAWZyPqlC4aHCWrome8/fsPBfb5gjhseTRNuHU1AfAIJfSZt4otc/8Zeq1Pp
3JmC6BLs4qBNKniJWQvGZIxkMstMGYDXQrlneKiU+YhWVzffwPruRsxSycgnWVTqQw5sdEo+x5ml
21ZkbxOG/h555Yaq503Kj2SwZuhreX5lacgo1TaQ0sGzKtb475B+RRsQgFZW7/05F8o2v0U8KzIc
wysNAPAR4EIPXlw6oj3QRYpiNMlMbbIOfrSj31wnTAwvLkaEZOd9VuVn4o6kVjyF88rM9bX0oMWD
whWCtuRdK6Flaoc2e0K2Bqwqo+BNxMQnVqUW2ihHDu6IY+I3PKl1jdwBpOicPQXB6B35C3lisxt0
aZKlQJdTU4dpSYvDFjDJs5OMBC6eOpXLBA5KELl2Z44NeFR/b+zOMifH1KK9l109nb6/wdrwijJM
ivBQ3AjH6KjjrAPrfKhHViMDqjLtnuRVoe5Sm3/IV/6sa4PQJYgwiLVGrZSzMuoxZIq3pwlylkuD
qF6OKVcM04q1J8qlR3AbTNBg6I0bzv9zdoIJbdMFpqFC6RPHBNZXx+1zEeYRur1f1d6MHz7yeshX
sdugrS0rr+pQrgph3kLoW/UJcrvjO08Zvmd3y0FZt/YmR1yb/vLoqzKxVzZ8ra9Wn51QI5CE4wDr
uJmavrDwpECf8OPGNO2dhhfMlpe43pOazzgluIPpc/piPXliFIsHtSZMGT54EZ9r4NT9EQ8WzCc8
gluf05QcOf78nXc65dExzB/PU1iJsVvQq/nRrMp+g38FZu8J9ipLuiFc4KfMoTmIzFQJ1y9mRXVu
OBi0orcYu9VvT0r+/PLcUXUc/OsvoDtYGSRk4Mr+F6KYPXoSmFEO9CfRtRk9DSy/XOkMquNoSrFW
8LcCpayw4AeifCzyS0V+hzNuHWzqvry8Ma2/H7MsMuy+tCTjYdJ81npFYxmZLfOPIsUFSH6LzPNR
3WS0DPMTSyK5JGW0lpkA87CWnfNI4InHvu5XA2NWNlJDESyoQrfozgrY7VzcNFjriCfAUFc63SQS
sKONtLR/oKX67YHsgWmLAGer/NBIZnI4qDS1YH5vy7yRvP6jWTG+lDOUWY/gno/Y7Z3Pxjf8j3ML
EA+Nay5UbJU327pLTQdcGh0pHyeSqeA79jVOJsQYbzidGMUJUdnfhGNdwoNb0RNaFw1BWSeuC/kN
Bp9SaKYB2EA9pircvhLTCh9Ij2B85TVJ4VgTpNND8llNGBn24Aar0w3oL7kqS/0qNL0byXaQK+7S
QFhYqLNXhogGmllMH2Ui6rk6T/rtE0WVF/g6aSF1xI9BhcjBjqMIXVsn/qzOQDVM483uGj5uphlv
HIBj9NGp5vUsZZ1/5mqlioN8usqmX13oWyNhobkcWQXP4mtw22C5ArwVI0RhJ2vZCg+qKlwrQQEt
pxjrbKEsAQqK/PPid74LPaZptWSZ5ibJiwZCNrV4meIqipjTBwTvfWXMj/YWPf4BGqRxPwnxNKvn
Z5GCMjUzGOw5kdBfA+O14dCCQGdFEzX3jWVEfKSAdLd+qhOlrVTrmqoa39N+gS5ozzBt9IbkDgXX
VloHymmwyvI0vlP5+9fS2nAuP6F5OMtxNJZ460MXU9fZgikM6CBeZtPeIYTEoV3pKnYPdP3oOqoF
0OR2fEO5djLjnN3R0LAuSn3UtkoTACAnqLyEcKXM7AP2dtW36bt201QjEwK8gvoi7QJ+zEzP6j1X
knDd0TFKKzBL2zAP4r3/I/0ph5BGiA9p4jtjnZ8flXIiP51Z1znox4u+y3elSUdIO30QcEnEysn5
YSxRypMpsafku06B1l9lg7uKn350RTYxUNlOQ6WW3dmnSKhYK9f4OXFEvzjsafUq3ANzbHui5knQ
jtLVJ8/HXg11tvwJ+KKH5LgSWgqE+jyqp9DNk0pK+dIea6PYE0qk8RvrpC+9orjTmGNeBLoknAb3
tzucfm8CRthBiNPHO68r0c8syJTSARJyY1QAEXaKQPVIGaHJi9l4pm/lqCKg+19SM0Q5f7n5PmSP
VCRXp1CZHgh/DG0TPweDPKgpkwZz7F0rS6A2lC083WuuFK3mFTPGpTLGvOdgAmjalRlAuTqfUIps
gSjarI4b/WtflAS6/fcijf8362ogW3rydkzjDQe8yIYSZQmO3vzZDAo6U7pEMMK9NoVbb9VnKHZ+
UO4MaiI+l/JqB/JMy0GGG/HyLnrb6uN3n8bOM0/4Ke7TDUhpimPtWDW+b1lIIxxxx/+y7ekTaIsv
2vHCpGcsNZDxmaIXAW90DehPKPNZ5/Imcd5OrUOp4g+qU9dHDbbugzoD9tfoNLXo50SAnTamD5Cm
u3ywckgZDXhCQ0Wj4JtvMuV2fcBHhWwQ/DBI/fHVjFEl/w+5FTFF2RYXbfuPxpp6n2v5AdmByhWc
XiBU0+FaTu9XSkb0lLBN2Kljt109pxzv+4zCzVPNbqgiVWncDAAP4bPhrWNRnqiuaqmyiTGlIuvP
SxVSRGLmyDulEIbt30+EmihskhA8fO0tyT0izmKJUkju389Zycnuyvck1Bqz8GeRHhhkZDRZTHb1
PSBVS6tzIJh2AsGZZ5LDgiGAHvg7PzGQkC0mRyWW3AfkT7zBJ//3xc3LZZSpdCdSyYXyHKb2IGca
gCTmI0VtzOiyptVPj02gBQN54JQ4ayicQc8aZ0MHMXxK5gwjVBu+GAclR9Kcox2hc8OulG3OPUoh
Z6rTzHtuJqrTQLxpOOK+kVKR1AcuABUL2zBqhIvXkqsreWvjZQvQ0rR9COwMRL/KOi2ubjDqPbXb
CG2ji361e3rVeZ0vgVZcP41gvbi49/KsHhlSmcAy/tVmFxlK6vfxtc2K2VFydVdsT8WdZSb0ZQgQ
bYdW3kQ8UqGuXLIo2DUK7MztuNFlZlf+rm4YCxBVm8pkfyfSbnPq6wmUmu7G4qth1PCXbKz7i0Ci
P6rlyUqAprsDM2m1mwvM1e6vF/zrzadDLEwt6ojA1ZFYbWgxr12e1NrsqF+Cq543yVYdrAcQLbUd
4tMeo/wzR9l/+xZjhJ8/fmHXw5JVX7nN766ZeGtkLAA/AmIrnLZMMF1WS0a7rz+Ir41V/V6eQ4rQ
nQHs81rdPQJaxdMJGZcV7lx2heN3LBJjw8tad75yEOtvedg2tjLmDNJ6UomO9InFHh/QWTHD7uPW
17ufyW47NW0vhC35QajMytCsyhLQ/kVRJcaWeuZBoAnKftz3zeocPnZmrAQC2wAfArO/GU8JI4zs
BrhrtLGq1hZrKRWCWdUbT/v2LCbu5SanCtpA/lKeAfFd27O7IhdtgECfjsRrwTju3deBl1zc7CbF
c0D3LHXAO8PBiYPdw81VBlAkhfGa+pRiwA2FAVAX/DaD4aF95fKQQHC14JllQiT0HFidf5HppSSY
mgPag87FQtlcTggJqXmUJlz2tjFnWaqtfMXy0NisEzdIkRULI6z1qLv2y8RWAt3m/KNwLeLqoLtE
JhKUhObLH3XWTTxRkA6lN8uberywZPiKFBg7dvNNWMCb3g6oUy5pJslXalSjyDmYe6DrVWpbwXZd
1Z/aF2h+IIsRXhjJdHAsidGB5lpobdN8nByF0I82AcWkVZkxkzzLhjR2Idl7JZL6R3ze60e/hBTp
qn4TpIWCc+DCJq6ebs5xaCCvhRWyp+iqFc/jWKCXIWWgdjpVBnJfb9Ndmv4FGFKwYNQvVqzlkg5F
NvZWkYHxI+EdePNSb3kAjYeFwU6xMlkU56TeimKz7ab6JMvQuWmGcc2C25EH3yosYPbIBEP9TfrZ
PnPiBjnqhvaPE1xFytgBEuFK1Ba9DMTKEfJKxIUQ8of+OqYfb47kiYqqqUP2o3S/9QtWewpCQIEa
gqMomaWbnio3QPMW5EqYNoM2utdqIMg1AEj+nX14HEX3nGnR+QALnfaDV+KDoVP7EJpp2O3yZMbB
PpOTnPc49rsCtQCkqCc5N1tOYY5iMxWKFb3tZc2rkqfSB8aERFy86qh1HB2EvbwpQTQgFyionIgu
et7S0K63UGfDbFkVuoyF6sp3SLUfhku7QLWZU2i5lnk0XEw6ROi1gSPQmMF0PurznYTSrs1byH5u
u07A7SCwGi78WaP4cDPagQtbEqe5D913cHfZdKkaRjElMC7hLt5OOSUToZEP8Mr4jOqVO37O527C
C49tgFbuYPzZTOrnEhArPvx8lLomDXe75J1za7RYURYfMsk1a+LFMHkqSogNMU8sIWqHH5dSeGyh
Hn7uxRnG4CX15UKQLcsuNGB6Lklf4B8ePCPfGhtdhsAVwy5LV+mqGCdkcrrIP9T/bOHm/AhVIvOX
zgTGulS2uOIIz4jjCt7+NhiWYkao5K8ClBCmCuKB6+YUnk4jHnvYoRYDb+GNqnik3Q53sTgXPS/W
Ih4N2ErgLB62LRDOamR4rGP0ciT7cSodaxoGNkkq1zyMOX2MBQ8XxFFvF6bEf+8bdUz5TH6BMVvA
QPq10+CNq7bd2i6ikSaPJNMPhooKEjyyZV/95yPt4xWeP5LptzhbWO6qHEppqW7kE4Fhz92wp39i
NFCYjzwSaD2OmMjcZNHk4tTFb3wt+GSR8kJoAybleqp6+ILmbIQDbGbhYWydEzGlzlNsppww1SNU
GccJEHOtZoiQ5/PTsFRu6nXfsnrsM/3F7RBLiYr72lu6lJ/H58rJV3X+rUcZPTmRTihQMMzZAvLu
uiL91zuePO78UFBljBY725caCw/HBBo5TJYI4RVMUJXWoXXxBKEkbOPhA74Uf79q21CgNoydFXCZ
afrkNI6cXVKvCLfRIKjpxOrJzahyiHYa+M80e9Mbw2s2/taCJfM07VI24JCJzRaB9EnU7+ySu0Ls
j0ro5Xydo00VOsvEB7dQZ6Hf21bKavmGpJ5k3v5Uryen92FBTOKjNh2nfOh9ogoGFqQaNNZB4CeF
YXIg24YdPrCWrirAKMB55gS/Kv9/z3w+BMrMPn6B/tUhOLh1Sg6CzTXQSjNjDCKvXJUj8dyhSIwx
pUfPOe7PkE0fOUTuELjnQ10oCI4toy0J5VTwZ5iWegxEtghJc59PPPJS9e+LEBF4dOgDDK0VJndE
4npvmnKlr2ETgqbVCWzVHmx3hiuPFQddsz/zMapYcGkrmd1Qdgg+3FvbK699gwkXkQE1pMJ5lQ+G
reRbdrGomc1jhvZ/5a+/dDE5sQplx4+78uEyOQN2Il2gpptf9lBUQEqpgF/fcHbGoZbSyD0demFK
Mwnvfj2qq5y7W+7pRHFnEIHghjWKMyOK1JH/rbZIPojFqfTRP8ouM8zo1rParjxPsXB4mWdFhOKj
q7toWmikjFjzeSjixK3tVm/wYKIjHyDluODYurt5ettZjLzMbwu9QYirXXRW5BP0eGVnJmRRNoTN
PCIgSwCGZ3f9IX30YmDNWlSsLlZWEa7GIF4xYrQehLmOXV1Lh0K04UuZ27QfBTd6ulv4m3+Xzo8B
ZMmMXfMZvQpNHZN00GIjizSQD7UqinYxKhGAJwd9iKbEBYeni3DgnGVEhbTJFb1/WhLkRKqaA+1u
//EyIxrstW0HDWWpMhh1FEMJRumA2wyv64qvPaoeuiPUWmg2z9/t/u2HJPmtHW47Wc4DDuuoFe9w
GYF17DCFrUO9cSoCu43tLkanTLTisb5SbiplcaFQ5VvBg+STDUt0zSMu8Db59GhkdCGxz8l0XR8F
e5woXSwsQdXQCNP2JVdzdhMIAaAdnjnIL9/DGAgNYWnm+ukmw7I4Vky89NP+JRw4+FGBc1m95WU6
UM1iXtSkclkdCSKrgbgWxRVQrQWbkPR1UGHUP09CIQuCjBn8oXgqmndgPcSqA5N2GXWyGDy+m2VR
+HSM8qzQSF2DT+WRgK3WsYZoLM2FdzVIr+K57JoYp6Tcwh/va9AGxy71EZKBa6yikp3czK4Cm0TP
MNu3xfwfnHXWALdol7qQwp0FkeLPYjS5c5X+yuEGUCoEyxOdJ9kjoUAxtQwrqx2iTKnVMCxe9Mul
JTX5i66ztRElzNztAj3KVQ126VZA4TEGbV9uZwwTg+VRLY+WsE+il+un5/brucDtvbDcrEumTQwt
1QTP7db2z7PXWUZEwA9l1P7mVC1meS3iErKxtlVwVQxSKvR9E6iSWG3deWzYuklrvM7+tz8hPUCR
/iBNB6UPFRDyNJbWdaBWqYEDOdBxRK8SVCH28Y53kPXr4/bAD/4OZ4H6eMawxWSeSga3iKRUReaB
k7Fso61ihuACg9010e75mRpDDfpOtQLwMH0eYeHd1LgoDEb3CB8I6aYWYAlgxEOuJawDV8PWYQik
nLIwm5fKWnmgPpTrlFbTcCrY5efNdUbc3Q0mNh6qgYTwCKJhIkMxsm1RWIaKEau+bxJFehAyy3I7
0dZkjsm6MXdMaGOnAMhiwwqEpv2P3XDGjT0eo7NbNBsVI4pnvDKLCPGns2YK+Fm7T54S4pIhsbaY
4tq22SsIc98kDPJ26XzfkmPLiddpK37IX5prym8M9PsyyJbEyaCnnbpu+Cm1E/9WWenZCe+d9XDk
a63cTi7ULn2ZfmgJwfbsHFFgZhOyzEWfKNtW+i19xmUe4FUXuuqfY8MN/mvD9PWygBYY1CpzJqxz
5TzXLbn/NSETaWMeFrORHzolyTvMTb6VpKmwFuGiWmSeDDjAXk2AgHwjhwOzXEx1dE8opSaNlj/2
RPO2ZOpBRIhFb12H8KxPQEeHZKuSZmHx6ALPuHErd64VkaFKpiccD6QIBgut1mmYKnikSQU9JYAw
EzAT9yNzsota2eHMp7wVDertBu4FmfuuEb3ZmHLJf+bukBzMyZMjr31+uxEqVGnnLdvdkCqBgeyo
oOlW5nCC+RtIr9bb4h05RgrDfBllEJxA+kG217mPGMm9tMn5mEZiQOEVXaxyuX6b8VKHCR+Sd9jC
pWPry81XIBMW9X857/qj7LQI2nz7eQkJE0mplEms6qQEA/NhtKUyOR7N7gyJKNuoxGFvm9nKMQOm
eUNf6tt6SAZDX0uxrQG2DdO2MwGIiNYKNH0XD7L3+5SQELPegPKbpZg2TAUMOubOdK04sGRhwd3w
c/QGbfUHn+mNthwRp4PagH9y3fzors2U/m0sxw4bG74apAdrcYc9Gb1JJpWSME+A5oM+NgbE9cnT
ov1PeFKm2O+YcZhpa7oqFP8qIhhcPT9OA8ajL9z9L9NK2DgK7O7yimG9WLYnHK7H/SR43fwsF8vT
1XvVtGv9326fXSv9ZlxD/yNh9TiO9cnyXMKCbg3fxfaY+i1jwUXm4paobqKu9J1/l2nw/r3Vbhch
b3k7R8enJGjm5asYF0/M1b0BtfmkYvAmiRSRDCo4upZ/EftWox/9G/B9lCT8Av4rgrxCaJyX+cKT
EvKIqPnhdXlDIvnYhO+hCRvgNynfQlNrXemLZ9oXiETcqsZrURj9d4oA0L4MCSHu1EtY61k/tXOe
21DMB6CvKbnr+k2yf6S/dD1jo+soL0bY+Fvm6yrCzYH50jYgUvBnHfEVrSkZHdpOOqnuAQfBMEMR
5A5SY3xkt2N8GE7e+tZ5Iaz81KYMCgIbJJnoAJeSRDo0I/Gir1pvzvmF+257H8GjUXj1q8Q0UGqZ
pej/gqRdb+SBUcDdxWxTd3/hKDnkj+CaofAKY8iXO2sc3qCX6lGwnAmQTlzJNN/Y4L7Z0ets/XL3
J8VH+/cnz6NwJdQJ1FyO/hZt+4tdWePKC8AeQXOvXrsXP7sM96bV/KgL+qCmjG84JjfjpezVQMhl
5crELFKxcA08fBfXh+wM7Iz/Iai+mYcetrHUakfdmWMi9x0PkXpZ2NC9sZonvH3FdjgX01nvLPj4
K6mRySEVLsq+CxgnMM/RFBXhgg3ROxlH1Puyl7l3S4nSLsFZWKdSHUHuSzQVOz3yF3bBhkA+Ta+F
E7uUTy9nTrVPddh6240C6PzyO65us9jxnCa43BR9H03Vay2QiUYoOQVhDlE2xfAa5is6bBU+mFC1
k+TGAh3AI8uukUGuLVlZmMuEsduZ8ZFQ1vQ4nTC2xKelBRBWxdviiw4UIQSglZr8cpgy1ZA9mKHY
ZYlRd9m/ySMt4bOOX/xPDrKxlQNXS+kwxMMmwHfSSHLWDSkU4lLxaPyTmMASE1SPOxLcP6+tCa1L
geKRjZp5VFNBsoITB8bU5thfr2KZhu1wOoh2lZyEp9m45sbrtFOCmtBHMV7u/2Gj4tKha5Shpdsc
IvHDVQvE2hSWRdY0wk8ptfH87Qe6Z0rhQnl08ElGmSODv/Gk2+cXWRzWYMnfQ2BsEkJqaTdh11gu
8B+lAotRQNTLt49O4oNV0LlROEE6rxZs0WCUL3hAR/46d+qsLeHXKKlBPbQD0/0eFzyUX6zF2J//
8IieCtspXWdH3rXVjsJyxiDUDtdHt/3Sx38YWnHfzpDZwWCuCOnYkOo6X4zyRq1YfVrFoXVWEuSO
m3vLuFQissBf4i5HkRyiyC093pI6jD1UpYy7zl0QuFLju7g66HRKRiR38IgTS71AMFobELLBxiLf
kGQn3/npKd9UT9Vb904JmDh+Tr4Udr+vKq7iVtZIiNBNyLs1X/e5i7lJSjOsuYCay4nilSjmy+ke
YRD/PfOunBZ+Wx5rUAkOJRlV4U3Tq2h/T3UXtkGBmtHCCiB0pbWJCyCvcusWa9PDuP0bRZqEXjkC
U4ACXLcfcfRBOcrLBChyGChqCuzRBYtyC57yL1n7OlhSApuQN7hZVuX+TfpGdCLzvcLDCfo6P+xm
gc1arPoTn2vzs72GkjAA+oN6rOHKYe2XmpAQasiHg1NMkze34MDVQYywvXVb7HMWz8lySGjf4EJN
BMm25N2Uf1Pu5pWrdv2j0z0gcEM3n/91b8ZxaxJFD5E6UwiuOW+V2knffXr/agUqY/3sEdRZaEZP
7QlN0jLU/GdLZCEnaS2gQP/FoTKLwNE70zAFKyKbO75vil9rYGyMeB1SoYDXk/7F8f1YkQg9/wDj
6K2ehbzWu0CI6c0G8KKnMU5AYVXMeTnZGpj1sYIXAnAwnPKXpiiZtRDsMKMCdP8q+RYKLKfCBlT8
1wifLHXHfu9+8WPE72UVMfiVStysHBF5vSJlxdnbr8JQ6NxAmlagkVs5xEEaKaqpsRE95cj4jtkl
zxKieW8EKodg8OJLXr7L+AlHbmQ1X6iU2HSZbpYyXBfjrvLx3LehKyjBxY6tSc7O4usEr2WhHxVv
1BYIg8cePgqrJTPBttmSt8GH/R5rZPw/vj/WOR2YxXhFwblJQ0tfU/3IlZSk7fRutwhjd8CYsFbA
VaqH1ElxgBTm40RazbMCG7txdByZG9WqZ5uKhT5r3wDg0bskITsHzVGa1BIlQB7mdmZY2OSopfqB
X3zEz2XRoQy4g1MvyTXB1EZICBQxGsvQbK7k1ZiCo5B95VrcLP4Zl4BLj6eZMpyc+WiNrnT+4Cfh
OGzI3XBOmBxGfgbXOaRvUd4zcoWnC2PEhX1y8JYjqeZyeJYcScuoQKkOh0ja9UmGMW8iNiX1Fsyo
i8oBSf6IS//w3D3dsSKim56IzJjGwQEO1zOBNFgT2+bTqlSjQ7yme8dB4UPmbe/lDlhqXY8ZOnQM
oQ9wcaERre2p8MwAmHa/MZSPsigoPxGCHUG+5kosbbOZEVMSMVqYCy19fal7BtqY4cVrIhcWYere
jS8VdToHzcZ1NHR2oW+73IRMUgUlv+yooOcziVbZAloDpT+O/8aOR9pGRbmIbK7eew8XT55QRKlJ
Cby2RXaODcqewYxMl0KdT03ieynU8pUmySILRdbixb+cgtUWQLE6K5trIrr7Oh0zmR4akpBySFLt
TeaOLKAONByHWnZ31oqzWdExPnLc1OOqhSnbFNtbDv/6a/z/S42Xo6c8+atnj5NKQaQ+YMHMlvQg
a+O3NE6OGmbNE0ugC+8Ro/t8aS79U+R0MyYw4t0mmj+Y7BfHgLrX7JEeSKUt1jIaV78zU1GXfYuE
MKdlEZg1UhU44dICoUAgMGMYXT+bZInSW+Sy5mjA75ifF/yftbzboB3ON8qZtbJybrOuIowITdpO
/Low+4t0knmLt3Iblwv2aq0zW69FwLuYiyZQX5SZZHeIzhBOAvIwYx7HT6xtGcTaPgCBtAQN9wHd
XyiubZ5jxlcK+/vFcZ4DKr0y4xnsh37Npvr/SyRLRS4fDB+ZZMkq7Er3cV7gr40Im68vewhofJ7C
DRuVY0CYIrLKPAx7c9BYmjrc471gwHAw4H1j+Hk1DVdfXyAPIDjSt5DzK+JsmD2lzQNOQsE9yy0e
jzUN00iYR6drUl5VyuTeLsrjx1I4ex5sLvaGFcdv5xYSGZlyUymBysGzQqvBsR3EN3BBkMRmKVNJ
/485HQHiBCi8NeoxpihAdMpSdnsxg8LFQb6ta644tf3S0l0ou2lLRdTtFY0JN3SQTyLlXJ1fW0Ar
JvvxMs8PAWI4EsiWVlxyahQVUuiohcmKTDPeDquqo0UPFOWb4+rx0MpQwQUbUnO0ocVZsF+gNW63
UthJOE5Zv5weqV78TxMGS81ZmN4ICy8wlaoa2Vmln1Tf/CJBo8WEYZExVRtOg8Am2vZZ5qOd64HY
ttAbh75POUSwPCNg1KHjTsVoJtUXGmtjHA45Zy3djTFKJbwxGv5EPFFgAzSvX6H1gH6apwL0fAZa
hOSsW26tVwQpIBrOQDXHPh1bjXig+aDlW94nFdg37/1ZliDzHisCMj9aCllQw1Nomvtkea9le2xk
afntRdOJOgC4p+IpgnaRmPOhAAozUkrPaVyeWJ5cQRXOoRS1Q4JQpjeKgCBec+lAvZl6HpAAzRMl
q7v9xeMWF251meXuOMl6Cr+GHq5ufGojYVJQsXgyOy1yAl0YWcgXmKDPEZMC+7CH1yj7PIvghfbm
nS0Ii6R+kIXNywn0HC7dpb1+62c6Sr8mxzPkcDSwbEMzRF7UKE6XfrFn9LXbuLcj7t49upU+ZHkY
bF/GRdk1h0fqdbpnjIfSA8/uPkEwcwm8BdroxPhkoos1PcxBT/w24Ak1j8XiInb9Q0+2pYO8hDTO
etSo0+iJqWI6znHbRVxJfpuDHOrH18pGtqleKDJv0SYSND4UJm0sKB1Nmx91a6FYlIdttpTJgf72
eGsY9bTMML9xlz+rfxiDe8BhTUwrhqyEAAn/JQI00PAGVz2UwjdEdH2cQeDRJ1xblUQQc+zQqBT5
NXv9rfHxHixdiMpZGdBsqQL1zSrvKSCOLwWB2VM4u/R86Hv1cOlXgiP0YZRUjjdJqUK48s+9Nhj1
zOBaEDSUbY5q8kkP62JsAf2i398AZENigcR6QfybYkp9vA/fbMV0CUMFg+OkqXAAL5Pp6OF6R+FY
jN6JWx5BhwCMnkMZiUGVvudWdbYJ5nNmg/hoPsoU7kLU3bo12VbRjt8sn06NqnGY4hnpQJzwRpS4
KUL5a8SiK37Pho8qDy6VcJ+q4I2q5SKlvqJBxIbRs8UJRKe1NPAyO3yurUx5ntcosMZ06g/s/R3b
Su9RsyytfvUeA2F7RRfBwdv8Pqatd/bYHUurkDvKNCwmS0OsLOEYACppHTwrqfziGAsFdrsIGl81
T8OepbZmPmVzKNOWkLoCHDjYlv26DMcLgT8QEUY7JRHEiMSKWaVTsAq/7ZBiBeIfAl7wBYbpeIh8
je+EyDKHsDeEd6nxtcvnlMOVx3e2uSQMVwgAqHYlrcvJkEGNe7t4fA+BkVDkQ8V/fFccY3gZrntC
OTvMDbnoO3qjIivsmYeGautPZ+1YUKIpoZFn+uGhq6Swt7Iy/fNM28856QNy/hCV0NixA1OlmLcc
NA4bYTnH5N+1hnsPdzETucOyDn9tjUlBOKPJF7/CQ8bPaV2XDU5iGGFwpDMPsMr8ECBLXntCQBpb
wUDlOkwvJcyrweSsrmpsLqKRh3KbDoQQfC8tTcIboKhv+ChfHH//0ElP+A1trwwWEztsgKAlmQN8
e7x58hBklqU6zveeVr4v/IsV39dqXx39HwevgEBdNUkXmQlY1i5TAoUv6iPMsmntmgvbbsD6Edtr
rjUNR7zBs9YG7m6UNCO466Fw+Q+6NbZfUfhSyWjD3/QNZbQTs4hVJ5sXRrVjTrFHQie8KqXzdWuB
Y7UVffnAvPw9YaYRttoA3L0INDbNQFjeOUIxo3Ol3JbElUnJ2FwC5Y3MTx1Egkzc/gOrO4PpErUP
cBu48KCwE6+2Xk0kiD4pyx6cc3iE0QUK4Ui44ecMZ+Ypj88joeRUZdaWH/6IN5pZfiDpWBkDl4mz
fiOXKH9BVMnybD7M8YsM3jhjfgTE9K8q05wfActw4b+4M47+eBTJU7MtCXC4s2rl3Gkr0iaeO1X3
nB/P4F07b0Mo7b/QyNRvuiNGFfEbgDFvzmkWU42x4t6vHvXchf9bY4VIvLXGUmtmvdfGtTJg81f2
mZYybXB7PXPy4co8FMiM4VappIsftJFin9zgXjPLKslPX8dVRgjtOvD/JFEFWzI3+y0HNdUj0L/a
z678HezEYbDIHz//NcliDcLycyaPJCy8rAxdbUnDe4I7GliMv2tT0oVWcQ0rw+I8W86Mym56/tX6
azJzZO2Ia5rROGzaTdgGf/ThFG7xSbGmNKssaiAIADOwMRqTgm6kfb1Ht3Hs2XrwxSAYHu+sQ3f2
WYdfXaFQquDfUiQdXbr4cEgsztyWfdWtHdvV8Ja7iMqLl3HqlRyMv/eYmbcvEZnE8wa1vH1q05RR
gla10MFcv2nLk8NBrMCZGedC7o0mDEs1ntgPxO8sGILVar5BAUY5Nysx1pz6Kb9R9HctFt9Gt5wX
/nzPr+emub896AsikhjDxX27ALIwj5abYBnez1dxqKwu/tZuaWjJMhOWiig5iWkJpJdXfFFmGfIg
IVY/oC8NzxzVYCCghmKnZkl59kQ0iMl4m4jp+0Rys7+Gx6g6dgVqCCGkLRmxHs2wmKxBJaKjsmgH
CJylZMzueBha44k1m+cReg+Dj539YSVhMTQJg2nMHw5EJ9hktUmwPQAv5zmDY/0T8EK1d3Y6uL+P
dlt3avtlhyky8WRJUsGxUNZSVUURghPeL3PhrjgFPw6e5m2+cBQNL/3548BptiLephwuz1nkYoo/
SGYCboz7Kmv/B75cHCGO4cS6faNHblWBFYIodL+KZYQdeZE8/rMpIOZ7iW656N4MR8Cay0PSK0f+
i4kO/UTUSThEp6RsVoSFctdScvrvTO6iCPy7oIhDmCesG0uD52KoqkOAndeyAZ0omZp1seoMx4a4
xT+SwOOjjTpzVycnq1zFfIPMB+tumVCqvjsCEYJKASPhtPy2+WUaTUJ+QjuU06e18RPqQ8Q1a4+A
0zp8eSdhQJKaP9ure3gGfATuXmWuZHICh5rZ3L6NK/SB7FErjcV89GJWvku67D2EQIRdsPv2jAS/
KXL4Jn0+Gt4g39986JZQRUEC01opef4VVB/vbf162Ws/LLT1UT7yyuaDC78gKLBmnEMsMtmwD/9o
HOn1FN0NxtssSSrxWEysCtINVCuvxSWYJzRM5kaObchCLPD7e7ZYEgBN5BvSxQYReH8l9p5DUEV9
P4DhCdlsHVfoUryU3v8iYTd95cj8DpT/P7DU0Bws6ZHk00ArIc0s0iQcfJNl46ADqwoaN4mCNDtS
lb2sdeZydxgKN9ZuftjJmo6qyVISRvMC7llGt2GNhVzrN6E8NimQFmcUCS/7Yfq3HPkhN8lhiztV
evb6OPcjioOJQnTai3a4T3Aaq9LPkjcLnzRLoLxD7YGSvIvLJE2LN7JnOMBN+pxFOefdcwJyHTti
A+lzweaToVjm8OMsiIHxD+zDNWmmR2VIuL14DkWBpMRzJaw3dQDER0P7gp6kF4d/qDaaMT/DQjRy
DYN228ZP8iMqlrbTxFxu+8iJ+ki0E/BtFR1+B55X5dMPJjq45z7e7qfafZPsY39KNuq4uoIJNfV7
m4GlhHq2MRjJ720FrKDgxdGYvliIFdhGCCXbtFodI9y1oA/HN7G+BuCkXbsKGzodCFx7osA0JL7V
86zAAXC6x71OQ+7VQgmWXXSh3GJymmfkkqOwSb+QXdbqi9GAtkbwXXa8WBSxde94qHfU8lqLnUt3
kjcOwuzGX1lcYMU2TmDLTBcj8pscPrNPQp3UH1vST635vEy9vMfHysI/9+UZ5SjWaiIXB4QP+Fhg
vo66qxujno/B5tr6EMq799+MetloaO9LYFrM/fhxD7gsfLM7liz0ddEmxXfv2h8//zv15tVg70NP
UqSsW0AjLMKNHI+VjpHh2qvT1dJemLdbamxH5I7hg4joTq4RXJFaMk6kE+oxP+nh4F3+clPm3Lqs
vWg6y4ZuazTr6tHu2hHJ/v8RF93Dgtcf4BhGZwaHtsqMrKLtHX10Bn/lXv6Vqtwuc1qYc0QrZzJW
0qKj9u41ylkmZNjZNG/o4LnwVMzTkjISMiUAHZs2EcBTYs2U+pQ4azu9+zhGgz7NuOkWrVio2lXX
LGxge8CjtcGMzauDfAKKPswqHcWS5pn2GHfkElPfl5x9yI2ozx1LZ25DP1jRIlZ+u3UhRWb/BYPA
0sA7qlbHTejEYflIuCfUHzTjGjYRIzuMV4HYs/wWDrHJiysJJMaGIiPEPmc0ewMefPBxryU2rCc9
aTAOIyqwRDMUekCqsouN90MjCT09kY1FpKmkauNfXTQ2ZnhcOy2ZKmDdhXcxwOLdQmrrISoe/6Ne
zUkcsqijDdeZZisFaSSnHzfLY6NhACFjzrs14ZnHJs0yK2mK3ZhzHim/bRTGpOtBQZLLvT8X4uUc
pAMHraUzD7zxbpFOEteIZtSWCVmNbi2nAaLegC9nErx0n4TVhA5q9RvOMW9tAsDdNNl7wTwoDA4k
WhZWsQIGRR0dUfOr5Xhw1DhFU7pgEBKCO06EXu/fxCLRvKjjSq4oNENMEanfhVyPydE/7K61Bgyd
4x2CuxOAi/RjG9y08qBEcKoNPjsJvcZaBJhx3tkXcwKCAQ/C7SYaB3y+pTw+gQc3omlfo+rKwN5P
vFCkMpBITNjEensoAeic6IUCqYX0iLIDuRnVw3KUCztEiyw+w+0+LBvNthBpcr5jN1vHdpBpDDi6
/j9d2w7JjHfvQ5CALGHJ3cHE4mESczO09f/+hpGz21+dynofYVaW0xWgzzaltsUVeNIIU8OGPpyi
O7Sk+ziWNNlTe92W+piaiwF7MVIZyi92Nqj2b95+pNnPVqlnjHm4ifX7NnXLOEn55Eo+HSga2RCp
9N8Il43Cd/vgsheQlWvvIR/zMSEw06EndABk2UJk0Ntn81Um2h4C3oaLZNNJ4k98WLiz6dGIlCCO
7K9OHBxuqpjjDCo8O9+UE8VO2VB2RUqXvsk7UoyvJZ07OR9TmoUvrIgHQ+uClwxjCy/oeMcoAwiD
NHtUbq3PLeYmtG7QXh20bACeWbBnRl0NZZQtkLZ0vTsLOiE7wt7NqqiKnVUznBzrhzisTTf1Rf34
/+dhn2ZVH0tABBoZN5IWVU0PFpOpBGJdY3/9VOZsaGGzlTpSZnF7M6CVfE/fogwpB10eCdQ49ynp
H38XT9rQUywepVeDwdzHWscXrvWoLet8YtZXpqhXePocYUyZtYkhuTIkuyUfFASjRj4pq7NsKx1N
/l97dh2A1yCslLjnRxYpKdkvo4LKKrbVVoFDbd2EDZ3tw7RHxate+w9htCD06ilJac8qMobCL+Jv
0NFuvGWrjPnywdPsIxy8PFB/5s8z5QkOW4SS2ddcCf0RYWaVaY1a25IXExhjFjd408kw9tYUuotl
U1vZC7OrVT/Wc1JbDJU5L2dFRzkjnqZegV+AbAQzq9c/h1evHQDi7gZ86fUk0Lx3DFKIr92DXAGM
NQogoVSYiT/HSq7/R6TW7ZfOzkKsZeMJqudsRddDFiAEjFJXqMEbfGMb6lkl5qK7urSet2Lg7DHY
dJCCCYYgtRqvQQ+qOqXdxKW4kBpwvFNFCb7EnQHVvKQq3Nel0NIzkKl3hIFLGibkilNsVDNWAfA1
xd+aV+vfaDUiRVcWHFi7H2WDsYh2Qg6FbNsOUfMLdgS7Vq42Nz2DGMMhk6+uyGzzdNh5fp3fsehO
ukxdGvNK5ZKFSIMID90N9rhah2NwE9bB261jLZq5gjc+TzbHirryb4tlxoyVEZ+9LDN7Lh2LTxYj
WANICrSkVZQ/ysIYXs3n74toYMFpid0UIfPcGJy9VRRl2MNIydWbK55P3u8yfZdNrJ+yjJYFogKi
KvxphTkPBXPRyLU33BbQz6gAWJgE8QDxtq5b7qyp25uvEoc/kxb5qABDlO7XIlG4Mm8u+4c6c85G
bCO11u03go6b2Fsr4tr/Qh339UdfvAB0JOj9kE3hfKmf7Lv601su18B361RX2tg8ySf4Vk48CId/
hifj5+6ehfiIYGRpg8fqSfBkPp+Ou+qmFj0yHTPfNTR9SKhKllDEGmyS1z0loPyxGT4V3lACYnvS
ye0vwGxs8t2Ef22ZHtWoM5D0EZN6FOD1iuYnQ+Cz7a2UiFvaiKK63UdnXxF125csh49qTD82wUXY
pAlMTa0oeoCLBi1fWb1UGIMWceoK7X5+ev/tyDxHCaLscqzQJYjDdXeJKISUB3DTMBMsXnsR9Yr5
AA7OTQybqvL+FGEH7DBPWYKfP8PjB8Utl7blG6oJy1bxLsn6nR43Y3eI/D6J0NKv7nFipgc8T6XI
/nuUO9wfj8aynBF2wPSqT4+z3sMObiAovks5JDUXvww/3XpoaVF0PUJmNt0fs2B9xZF8x9zCtOrN
CNBhShYQw8+1nRtwDtS8wTUX+eF2kSvz+jbd4moBH4h+u6mwXystUPWIM/x53brXnM9cKzEPE9jN
Oymxd3U9ab+60EhRODzNGH9ta4Rvw+lUUduSScb/HosG/LSraEiVHdDsQKA0c4d6JGUzLOkyoxIU
gL9Xf6IzQCHvC17EcHUHtMYbYjSHsoYnnCtC+iMsYMoAqRURCnBaYzrhcD8xaJQ8mbzNgRSHvzgS
7Nw0eOvXiVilR5HKR/TO/+D1EKGS6xVlMjtrxndKoEPQQfAzMUhZJLH/bV62Ms2F6tMKtg7xEOMW
9ZFLuWzPEw2L5jVqZzIA5VOeBV6YAZ8CC06o2Mmgz+wPbzmokISsF6BhtvTyqv4U3RwKUbMWYb6L
23bbn+6DmSu2Jpj9A6mhiy5yYCFAXbh0mwu3amHqnFXKb0JWiKLqxfLxuuWvNtcwfDLUs15scR+2
PszbgKBHugYagGbiL2oWVofgmaUYJs4eno+tQlBCvWIER8hKR/Gl01FlGG6l8tU4O8EQV28CtCv4
/H1sK2qx9q3bZM2v16tAMCPGJmGg6B3BbdpOMn4aYlj0eXJe4M6jjGYkC6kwoLk3ojzNRvc5pto2
DySkgEn4Qp6A8IZ3CzHvrwl15We2+nFstanITNDTVNXUjdqbYDDe+28jz4BsyWLIdM1MfWpAu4Xf
ev7tpkIh18QTKosMPMX53yHShmcRG0h2Hh27bdrh3Fgv2r74gAz2oo2ROp2ZAe9Xy9TDf/ioI8JU
k8nO/yMkWFcG+ZFmd58dmYSwCfdNg2Gv3xLTqeInQFTS2HZZK35SJls0iy+YS7ZHa4k2QfWaVwnk
mnI1R95MGI7g/ETaWzrYt7wKKpBi9nf4YTzaezRGs6nZQeXXqdPv0Sqfc8hf3+sJBFZ4X/Jp3hQ8
Slr7mlJKcO7pr/PtHtPRUILmqtV+2MwQrfFBvusLMxwYAnVoJZy2nIBNIFaONRhJYpcbvRwZUvWn
Z95Kcn8kFRkCUYEnvklGMwKcw2urmDNEQ3SXd+KiIZiZ+DLbpK9Geo4i35Nk7VIGqNjkM5snpZgs
KrwU+R089c+I6xyx7w1nIWZO5nrXHDrpSv6XoETzjoCD2ba4qnu8nvwsSJKaT5I0CxcUNXWV+0Nh
r2J0nE9Gdl9NVFk83rsh1S3oYET2/htpTihB1V1aQt9NfMpcq7Jzi7/oj1ku6s35I3PnSWy/zjRT
PnYNImTVGJVZ0gNI5ys6jvzdEsE+odu0mNXvRzT4mYoCGe1kt8rTdtFc4dTVxn/2nZXPpvl/1js0
9kH6PR8S0G6HwilJHjsJy6uyjIZj6UeLrDNkmt85pHOVriQS8m7x0N/R6UH1mRpkXDfyPgGkTWID
9CGY85nKuh0qIl0QE9g/96qwtMBZTEgCfvy70iwife2kVAHCv1inRPyjW/l0hkfHTFIR6dsrsiGO
Bdi3AWq0YkeJkjZaB7+eRdkfTLmntglNWD1K7IsvfuDBiob9myaZdup1hl4F4xLMx/L0VuMjexUh
UPPopBOkTT+f3qWfpEiVT4lIJxmGaSWAIoRF0Ksgg44VLkEY0PsCeH9k2s4EVYi7Sh/nNcu5f+G3
vQCXzxP8dMJaKmdQgDlULdH2h5CgX3si3aFjAW86hhhc/MZIOpuUfbyFYWXihmCS+dBzUUNAKyZT
OqcpWc+wXZmhEQpJcWKychrfvCjxCJHwNH6qaSBjP/s2c7k8TsEZpTsNkYfbwgV7mNKUWj9QteBs
9ZVlLk98X7ft0B6NRD6ECKo/eyfplu7H0t9sq0v4Y2Y9pyH2YBFhfJe8r7J+X4KGLFPnKO8fbyW4
7hpMrQipceuQhnzAKHo7sBb0UBtwoDHgyjBxRzuB8UaVhN/htA04zGHaiRFzbshQIzi1VIJTAkl4
O0IrtqNuDKDd7xigdiU1NFKeC7OqmXj/5sCrfoY0yYECpKZl7Y7UfgnTGIyTPJo0ZAKhsDLpFdAi
Z+NLIRqDvCqo/c/ajKgwAF+UFmlWCVX2C8Qb/MuQuizsR6egagx2/S/hgvkR+yJt/QyYZGui2RiA
PCrLKAMkMg8lRSQa8mYh/lt1A2TugCxUgKNr/zyQBBJH6EQ7QcCFTvRMKnPJntbAMnuY4cUsVMNJ
JhNsoBCLEGpLuBrbo/oadPwklTNWB8uNi/BHNcmxu3C1lFZ9G+bxvBo7X46eT5+aoe+6YdN32GrM
WF+4b+i0cZl1O07+rRJHN0djAsC73gak6VnI+4r9y0u1e11+u7uBjmxkYJ1zr4lPa95jMN3D4DpP
K2Lr6sVvfBMmpPvYj7PTc74AimPszTLzimEjsZP/+DuN7iaIUYB2PXofiz+Z15E+7RP506C7tYzi
aOwI2y+SPjM5zERJJqNPgc40QLG40OmneUb6ZkveM77UFkAUaeXqB2BoP1FQZFVyDQPO8slSxm4k
vJ/FZtGcp6uqOLEGQDfaVqhPTs+7yB4bbj+rYK7cjL/kbpSRKmLXCpuVE9OEf6k8nTaYOPS6yseJ
x4TuYwyYP8cenF34jSeuI/r7WchpX/rIJ4Q3bY+/n/VEfwJ3RO/TOo/8ajrZh6ZO48mAxu1Hpjgp
DzVVGlffi3iCW+8QJxzGDbdHNaAqqySe8m5saL2v3EPEcHJhlfgy38xGiFc5WhvBzLzPjg532jed
9eFQ0dXPtJZLhY4YWJImjLIq5ufG3aoPxg2c2UuJNwaFCl7iWw4/jZhTTneaznTGnTq+5YxRGTG7
lsXqi3v7MnCQPWKGfxVfq1SiGU+zvGLxAA7aK5sME4ONyvYMizxJGQC2BtKdN+6wBw5hCReJucze
+3d/E3940zpEKkmzRbdDKZCreJ31VJN1SMJREqS9AolUp5SXkvTugCenDpn006SOeG9NuODm5YRh
2kPJSeDo8XHw4V/oH5fiPm2ebq5MYulXkrxleHUoVT22ZQAoemrY1A6jB8BT1+kGtEwG8jUtwnO3
saVZYP5SDJ7lO1pmMbZlzxh4BP/3TQ303TQ34CLJOFkXiXJewjL3qU3Hu3+/bo8piJ2Mf4YWjej2
mKh1VBhGUIHJY+ASncnvbeMWJpeClJZ79f/C1OHCSjhCuL2evgkbslzVmm/PL/cmiqIUx0ebUpra
A6E5HqqoM78E0Dacg9Bj6mXHQqhuEkVnx4qkO9c14dxksiInF3cGV2lx9rKLZ/XfZVsMKhjZonCu
A2uuACYYX5pvG7w2q6NFJG9HTrHqDOaXc5mafYfiKO9Vx+pWTKpU+qm8yjV8VA7ltzpZOIXlr+/z
EPfv9kRUplschZnQDKpAPCpMwVXS8LTsP54hDqV/f/HaEqugFMmITNR+cHdz9YmCc5mEcUv83KcR
gTIHHLYjy+pYawBJ4S8AhIRW7dA9mGyNpYQyTJ+enziPz9oEOnqqf5rkEMElMbFLjrEsM1bBSf0R
mLZXDuS8DBr4S+AAw+yvGk8+GPBYI6+4a6thZoYG0rnGY8HKLGCWEoDVOSPeOimV4MIwIvqOot28
+oTP1Vr00BjROUJvocMy7IWZnZ3F99xZflnwGehzox5SZCIQ9dra9SfcSjyhQE7LzRAZuYe9cTbv
+N28y0J4OjmEalMoMFpwlKgN2JdYSQ+zvlJvoa+wgwxcfBkpOIIVBoZ7sU1EOH8NAD+eoDOm0ZmM
4HV8vEHDyoN67WlBNa6kOpRlyQRccOwXVkJ9lnPLa2yZfba7Fb3zNoMufYfrIAftMy8WwmoRFxtX
asaHjL7Rtzc7YUdC2gKg0t9q0n1JAca04qAMLlfV/q3vuetjroIklliu34+T1+MDi00G7SSFVTn5
BWsxBI0CwQlOBCtYtuMQo77vn5GfWeB+N+dEouVLm0AR/GQlmUlK9BgxYml1tO4xWKwQWh1+5g5p
glVReXbYRU7dgQ4U5ha2Xqp+NkygrNLNsyLHkULKyE+29hXeEgU+Ak2SZmofKyRyUZ7eXx6bJjCD
VBhbOjEbrFG2SdX/JIXzoVH6xvO/Vv5noFCWLlJW0lASTP+7p2bYs0uSO6M02Nz0V1iNdRuy+jkR
16v64/phgBLkwuIB7WetF8fLkQRJhr3NzVk/FuRrTSOrgcbnB9hT6TFqnj2oQg2S6ZDN2ARbnL2x
b+RYK66n4pdsy1eyNC0eFjWBtGqlrQvBUs5YXKB0QQXptJGlLCbETO49amJiXjIryOrvNyAF0IuS
ldYxYmK7Uu3zDpxULQsGtNDGQaVz7Iwgr5EjvQOok2ZskaKm03XoGQy6LU5AGiI/Wc1MC6CB5WmF
U1TumoPLmhwz+kMdH4TTYhpedLXlanmHBnutb9umfCHnFa9X4J69JlQHCpjWC2Airk4X1mE+N1TG
MsGTo1GuyF0N2Fpxy5auhU/K5rhrDceE0i87BFOzA3xIrFtUEVxUtTKY/yltuZvpEWGDgPLP5eoj
jMuI+ZNyJwcTjIGsLuRopjjZa4mKogqu0U4xw0psk4Cqq8u6sf6XU0NoYnPDGBL/aKH8TO8dq4Yh
l9bWlbzc0wEn346yY7vMwjrvVv+KLi5dFoTqEfss2MbiWA7kZwv+OzLFiLdEB18GE5fiG04frXDj
MWH1801eBY/UlRVk3Y47ZZZA+dJEokqcFUYiwycU8DFQDbsmxyY0N6JAomdPSwoMWdu9LSov6JhT
YbBWIet2loxRUrRROwRfdLFpNWN991YElBKUVkQ1VHG4+mkBnKJmzYXrCoWsxbOJrdh/9zTkXk1g
aLLl/Vg9XigzSUWzLTmxYggrSI5oV5TyWUtEpDCqBHlL9E5eTscWvJtZ/8p1m4m1O9tpmHVPnE5y
T8htYpkkphthR6qFxeR3w9T5A5oB27DpbfpDN9nNiujeQ0zSk+CMCv+9FR25i8OOIO+eGnLttJWt
vxM6eDERwGb8/ok2DQJXPTeQAo4Wi3Acoh4hNUPFnr9HMcKqqlJy/JWMeo4uARXVrIzVasDapu+R
3dwLrsrpsv9a9LsBjxdbBWdqV1QAKgIovkKyYTx6+Pig3uIOYs70Usm6Ki8dscxZWTgJJ/8tINxZ
7NwWtQjnyGur7XVFh/msP0Lgd9lREhSYLAsjszP+wL+x6i2USZAiR/VZa2RSUPY93cTW2D4JyTtr
VjM1ib4wLKt65eFMnG1R51KLetIAo3s8LAK1gMwfNTK7yV9jpze5z0OtVAQgjU0WymQBhtnm1zyX
LAqetvxasJgth1lG9J7NCfNybryhoGyd8ay2hmWYF5gYP+QftgkBQZ0puIz1BI5HXVDeFfYzdKcu
Y5UyfjL0i5xDbE/yjO7W8Yl6pdQ4V/V2o8TYJY0T6N0kdZtRDYMsnvFjP5z++FBFGv/Eeabxz8u7
vse45nQ/es2GZ/D4FyrlhlCh+NBCpIoo9wd4f/gQ0qVzWkS2okbJg76lUmnCzd6dOc4oboKJmGS4
xWv44+X1moRaCeJhUHHt0RzLeKVMmI4ojteroIknhun82Pe4VWfrEzPzVeyuk5GOZkAl/dlc+Y8T
rTtaSuOump+XmdPh7yMXGqQo3ecNLEQcNX1AhnNXXtV338P4VCAErN3KeNr9tcDpp84Lg5KSeINb
g8OhCGDr3Lf5QYvhBSqHjdMbe5jLluIdgb87pKUl8cqTIjYkVVcv2braz/qtak3Yy5R4BzIQmv4k
Ee/VHQku1rBLkXtOL2j0pYB+ZqoYdj+PiYVr7q3YY0BeVjO29MqcsOOeFZCeYCXVFlayqq76kTG4
xDaS69lXBbFsDY08SfJXdWsmLnGumpzgvNbNumBhV8irR6/mgxo2S/OnMno28r0LPW4ZejTWpkVu
/MmHArw3QDIAvvtI9BgYazzW9wDisg2ORSjXgYmEgQW+4zN1SClr+uZV9NQ4U8/QRlP0k/yuzroI
rcMGTfVexKJDOq2sminvQ/j4EIwQ+qT41UBbvDgOnLO2I7Fr9vj45qUdUN7tztAJ/TOV8BVKZQne
fOxj7olpfFaYcHuNdD1fQalIEJ9/T1K7NPRoztz1GJpWuqT8IYg0pXAQWASbZsEgG9e07Qh6c5qj
Okq7PorT+iLI7cpBym37osKol86GwztjFyzr1xsM+0n4kBSJwgsLabm66iURhBxdrGpeDgtF3Jl9
B6w0hfTb9aJfjWSDxCCeyGWTLD6yt/LeQZ72dCLF2Ux7SJfzBzuw6/eXuLfEJIiFw3+xOAhJBPUs
5/Gumd9Eyx110+hgAAvAywrKOr4q3dBvOB8MA7vx4iLNZWM48Cjp1WK4yHufKaLZOcFkd7Mf7BgY
+CyGYREHUOyrkrO5FXNQPELE7G0fKzt6qLLPgeu5ynsqTH8E1O8useJAn3GgC5NvNWtIcnFwD3Oh
uhhqXEKaxWI/WOHwaqyKGGJReFhXSQeDap2WzijyCcmFWSNOhqMt1bR/Ypt7W3CesgmKhe35jicO
ErV46qkIwL2iWjtHGJ5KkqazbPA4ITWAHODp2QG15YjlAzwYkWv8YBxBoMHgp2yplrR8n8AxpsfV
Mz8/0OzvK/amQOL97gtMx3DsEZfsZlLlLaxFrsZrriJ9lOwMeeWX3NEXBAgHUo5BXWyVXBFkzQLQ
vd3kEInlCaeM+zA43ii7W8HUFx6NG6eJunysgGK2qjO6FaV9SN3qt9m4nWDEmaq5cvO1HPr3Xn4p
VIyQ+EHuJLKeRHYowod4HFkBueofbfoeYsounbffFelc1vu3IMyBMla8jOuG+SNMSSuoXsN97ssk
nnwWmYhPfLHftck95iiFD2x1F+GIkxviaZvCUM43zzRWTVzGrEdCOgo2GMYZqbkzk8g+HubN8EYT
l8P8QK/8ESwtgVXW2F5HgiCgXfezAES2fGqk3zSTZ3hLZ2bWXWMWJabOAeovcgil/c1QKY6pcD/Z
uKwBi8tHsnVsf+xDnLpcycuGT72BlnZ5g0ZyKoJyg7+6cSFG0N3BdPlTWo4cYDuhd48zyxQHuQju
lpCwQ9i+AY12OARGf6Sbo/SOJIY1ErAjsxPKlqXZIxdiNYFHlp5ea7Nucr79j5RJzCJisWCoqnJx
ELIGcs57hpq7+BNB4vJw5iPNtOnQ4FEKwGdBe5T8Z/iJFaylIQk/YZUmLndnzAcxI/qS3cB8O44f
LMH0AEttO1vb6LygBqo/Ffl9CHxbgdmgVAHlRYZwulbnwen9OtVUiM7nPgq/7S4B0jdTgo47dyT6
1hlmRdRlGsnqwgWdsc4R+vfmKDltF95CGPPtEL4C9JaSo+0CXMVKCtTHUQw48LgKNn1UowVyKxG4
rZVK9/qtqXpF6+ZiMDOLX3TbpAfWC8H2jqN4kokjxlPOk9X6GBH3lWNgQg2l7127JQCMggosl3R8
Wd7Z8Gmgah9wIWmLq8WnSyMPrZ7ry9RN0XhTaBxB6mzf3Pu+5opeRzjZbCYB6ss9CIIzdzOMyS43
yiOPPRtUpp2jzqkCkBMcoim2xscsm1AQqrMqFep7dLqljR9C0VAUQk/pdzX5PgSbewkQ//tTQ0+5
xWt4Kd+WDvpGPFTIH1MADwcZ1yfdEnbM7mFqYb1pjB75koEH9mnJk5/+fj7h2IFBxjrWWBoxHOKB
PdBWOhEkTfW3w1hdZV8x+ht+jB/g+dRwPcYgmBaQvBvQ7jmbHq8QIqAc/bCPTqwIW3B+BFfqxcSB
8ge+XUjUc7ewqHp4uKvDBIll0EuTwZBOd5IhfEHgC0oaNxEdLtwMiV85PEj1utAgSObHhWUZ/6qA
vi7QzluTTx/vrnhL43gHgxcesgPOZ8pFVLwAXMO2fo1nt+babYA59wEely6pwuRjA/RJsavZMAfu
t4xTZjTV9VgaI5nPsS8dIFFFPcPKG7GS9u1fQ3mSIWU/hZWBS/GgNRsJye+Id7xYTnrp8zrdDnUt
ljTF3TxgQbKvCsJK3hnEHzO5eOQzSQ1+h82ohxA8UBA6Mv2UYm8MteEB/FssWud/y6AhiBn8/Hr4
ctRScs2FvSHHX5DOOlsf4UL62SiVGKqJmqDuu2sFjOv9lG9OWsw+hroU4cY/kOdhITK0Eyhr+zGb
/nD+lYphAep+JgVuh9/zNc137ypJ3hmhut9BznAbpvBcAswWjfZ5W5ymW6vbh8SJ4qENw5bOwow0
ATUJiHJIKpfH32VgVQmUwMq5MijqExp4lxOFT+Yt+mj48r2uiu6tSG62oHkKhGoKnthbRf6ICB93
WtRdWB1g92UambbEBBFmjdoy+35GNPhB0vaSk/QODhVD0sSbJyLpwsju07C11wPAMi1IysorTz5U
7p2jzzURDrKX0dlwmDWgGVasj0xtPLEP1I7FId+6LEy6lYmYf3W8MtJQHajd4arSFTylpVY+NuOA
GQ7Bcwe78tCNHKgCLAOszuXf8TG4fIjJ3flMtcQriTZmQ+YtQZzwEqKxMPcWao+AKUCXB25Fw0+e
9HN50unryc5v5WnYWCYJy8TELeqGkrQNEdUX2buihfOeBfZjaxV+VIHdAC+QARaMjybxQBfVskQN
7T18MF/GwRp4OZwutd3QpN0B6lHN+KIwd+K1hSI3qlMAArc4KOEGSHj8i/LMzmDE6G+HKuNNqzSY
CSzJ2tmgn1MpHtKDthmSq2830pWGyzZmG43AVBFVn/6Vn2/bOw4QE9mwLvQ21OZhtkQ2k6LtjuIt
pxVus4281r90OOFe/mIV5BCJEmo/jgQcEPzF6S5my3HbH++EhH17CpK1Jw3l8GRKnlIgHrM9qNhH
YTC2YxFJWFi5JfZe3Yq+tDCF+SN6HXue/J9f6jFLuAPtyVtyElsNpuQxHfBRmcnBfa89EOTBzMl+
3LfIcPjKDjjeZaj0uezmrBgrAfHlHEiZOHsa1NyxQ3Rk8i1joaPHuI2QY8AQBMTxRRYWXzispvXy
R3Idk11GeGC0BnVNJIjcgT3yTa+c8JZS+JIgFne/WeVgHgulZFuyoW75g0WG91+BOgsyWnq52LLi
ylXakDtS1RymyrDa5SxZxMDktkl5EztOEOpZ6njlugreazmKWm2/ZMeUIx3ZfM0Xk9k7b4/4kynw
FdwcUVczQqhpJXltlRL2ZTCUHAwCpbaPcf2r0fMmZKGYUo/Odd5d2cq3ImAfmie53azois/5QgfS
voko+lLzbWL3Y2vn5eWXWEu6KWUv9NzwGGrJTk4F2A7CIAdSXTHv3LXHqt6YyFq9TpZ+ZV9pfZ6l
LNxxRsTklIN4utrdpC0QEjSUgfHjQQt1R11y5R0tQpVFkudNVOpQVx4U1Xk1/PS5qNdM70m5VCuy
p89AjVUdZcwp9ehFb9DKG+hlBpekj51X4nusENv3X7Ma2C29IbBEVvP6KMi6db9MraNwWUNp37k6
OA8vpK4/QnRLiQs+9p/9633FkB9fv6sF4StA/fYYA4uetr0PUmTZ5XHNqPbFr1anAgumTz4b4q1n
qxV6TMhfofyPSljX8UlHcCS5NvjfJaLOLUyt8JUpfLlkYGJz6jfHudrdj9tmo1Vt6gygQaYK0hJF
lbk98WMIv5FcXNQ0ADCSw+0lfm48LF2BSyELU10CV0aMrdeg/gqUkG9Ur1LtUOhFvNSLoTrzKLQ2
oLP7pB59N1U7oll7+FM2I0E++5ExCWCjIgJeCM0Wr2DEujydXaRvblWiLAg7/SmFoetZdGsWl9i9
mppxpY3cc/IzzPSfp6utwxfQLWnc1NLdDZfxPDGKiKJU5QWHqVtaNmzWM+Zz56DRxTamigim+z+4
B7dhd95DAokh4pyVs7l1st1Z++7GoLpzOE9sXAj8EVX76eBtCW/zk8Ite/ePL+aR/2ZXMcd8gcLU
lrR902x63Cvsw7DG6jPysgJbpPxSMYbQS6txyskQ4grpBQA8IZFKXcCyfD4qHcNjuVT5C9rVbKAs
fcpMAvpMolHAKeUBJOlxipyJrmMjRXgiIL4Q+uTuJuWc9/TRFSPIzP6JkpWe1/jIIj0HLDrPWbNg
SckSnDZqXr0/YMvV4gyBheCmhBkqjdqqGTdJ6Po637IEd4++IjZvRIRN6/I9nfownneKZnrb03Ia
SN3SVU63HvygmVZ+jgblWDP/+6md17hsaZM8gX0i0+oGdIKJGMmbBb/EB48KyyVgaVCwT/5kJ2tw
oPcZ7atShq3jqVoUM5qLY/Tv3THa4stHuGwEWlvgzsrf37a/xdwKLyPCWpsZkDirId6mqbDGryaW
edMS7v4pD/OrBA3R8sFLkL867iQDJdwLe4mQ3IdGQ4kPw7bH3p9duYjlda6VPFIOSmvRS8A4qjKf
eQ9StefYmOft7wW6f38DZpzvCVSF4R3dLnHdhUs72bINqZJXJY4UVW1M5fAhmYmgZJ0SZlX/KkBJ
schARRPWvG+rMEfoxU31TTufqDBILiJNHkaI0N8pBVNigMMtD8rckni/LO67S2To+gwzRBk7p9xU
kCZewOrah60BfADoejCuGy0SrtqEpeUH9sEk8ciCekSVs1dlYi8zJH55JGZp9KWmDOqxZ4A8UWxc
d/IWnEz2BGrhJ2VdYBTTAqLcYei8OTtVKrDMnmaBGN/jSBXUHwtqAL2lCkmxgn38e81qw0HFKd7y
yAnxSZgCKQi73RbK5WGFC0qxkoXi/p0Ky5CRJ888GpOItpOcUBHMAvWZys6c4UEkybZQ4qHSBxlX
WBRYFmrXni9NCgmrYNCmRsXJilTl/Yj68ai1yI2IPPNTbza7zXK9qHwnM5PewppRotaPpouto0HM
pa9QTYnBMGT8MODDa7cK2Npk9VZKHzJWaDMCJ4B/o4yYSYX+h2H+mb2eIdwLrfUpxGAyHU06kMwH
wl2tjUXGKUJHArm2zLe/tnBkXA5H3dahwmGm7OLxfuxxM40NNKm35zjdH6fS1ihi2xPk5tpER66P
GkDQJDYBShcxxpucVtOnWUAytMpHwa6N8oU1SeFp0oVYmzbnX5inH5q5m1IkMK9n9EHk+yy7ki4o
e5ib2tILfZg5eoBEIjxe+VMOd9zYI9IJuSxhNMhppSXcfYNEdGD4TOBEyIxcsnMS31k+Zg5mbZZe
bUosE/I0EcPq+x9UzOQ3Y5zvVIbfFs0fkua2le8531vcTHkfq0CYmwzDo0ATSdqvpo2tpoF4bsvE
MA/wXGjOfZPY6tPqMuUrdJ/GV4sWtD+ldRiYFER5vAOpnl0mrS448PNmKw2OqdZrHPHPe0qKSpgf
knnZDpEimNwgoB5ZlYw9e3b9hhI+Bejz5ugZ69aIwXs7DCyiFJoqCeM4b+8sZy3fROhA0CryFVs0
x4JlwPX3Mip+E85d/HhVYePAx+SPxBA1JHrtkFsCppaLqrC8TiHeqz9fBm3jDf4mmIyIEPyZap6I
FiBGK9dVUUw17rmfqvyp4E4+I5DL1DAzDsMcQ0sxXM5kLtvR52ZGsYutiief/V40UgZjsNWZD3xd
7SxmT2NTeFu1lzWX28NeYHv1Td1486wt4YsQaYDhG/VeQbm+EW9pdRF+PnSvC9hqqDKcohGNFKnP
uxoNEgYFCrIxkla4sNNBimlfbVJLDYiXxIwEDSGNxOIJGyazvpJNkQStgZYEHyYBqZeqjvNqUqUx
a1+WfnCDK6SAtSyCOwYoPwrzCo+d0AEyINAtpQYlN5vxnqn2Oryy34ut8eTYnTdreq3SoABv51Hh
4Xyz82BxvhOWUXHzq9zxJCB7IBZwQqOE6NCVNG8jV8Wtv40mm4A3fGgCmMQoRT8sy+ky1REwB47F
3C+DMcIpo2LHG2YByEHrtDcK4527mCWDwTq5C+fOmmmuxxkAPj9LXa50qL9zAf4aeuzUpdPBb2uY
HLHb7JFN9Popz+0MfPK54j+Pv7Bas+Jt6ffWnkgw0okvsFDcMqHrL2wt87+x0mc2kcxIUPHgpdY5
5W4bg+3u/+HZgp8f6Vins7wnmaPCG5o68RZB59zb+5JW0gS7lY7u74s9QDR1xt2qHtqR/gcrVWdN
xXyV03FY4hR2gvOpiN/SKhGaCecveeKrHo/L0bCzqSCrz3ENh7MtkX4Wq1xow11Ix03XpUrG/EIn
CrQAB2XW3rUoeUdFJnF5LIA43P4014NhLExa5D2O73eoUujUH9AjXclmIjU/LJIB4EBABvQPShHO
+ZliIWNSmG9MFaqB4bBjZ/0vCwkjy2O2notMNducez8Nra+7JOq0BG7vutOaHEVH2wO/+tNd2Yq9
zGL3bcGesFxY9oqE0SoPbTEQE7wf2TZWVFftPOYr+5GorB3KrBsLWkM0uUfXWX2UghXNLgWLRTNP
ezZo0ZMs5VpRgN+PdVPwRl09++Mfy7gaRZ/T5EHKaTtGWYkh3N3nOnpCzjHG382y5/BGEu74KYxs
ZZwMdyC1kmLkHkDkCPKj5QQiZ/5Mu0Az2zXq1023ew3kMyW5SSXLf2SMKaL1VAaIFVsnrlXuOgh4
zVoM3bIuk/xYZBpXvRqkKiUU8qkd7yMIb7P6OtiAwsXcXYILqUgxx7f5Vlnxhel8lbG4A43TNqz3
Qjj92l+RHgdxbom9osUhCb9QT8oylr5eK7yQdxmaRXlxcsGSqKNsH0RI0Ox6/5L5VJMTCmfi+SY6
5iTH+LhfmbTsOgLSfJUcqw/7PldbS3ekbtS/sdlIEN6XDF4uzqtCGi7dGfOUu1a+EIEIIVQT8qvj
sdw5I4YQCyILOhKBA97mdRRvGiv4HCDpJ89I63EStADzFrcxlenxd9RjkeALuXgb5VJv9HsVKHiO
8IF6SuaW20a9pYSFkYVRwdGJJ4AqLaLQMmyZAsxp/3iD/q1TvewS89r8TIe9ZEHZgs8gIJWUjDXO
pI5LJIaoqWDIcxfxC/04d1l7NS56Z4+l37TbpQD0tb10Ymsh3UFUPfJR28BFiklfP4DXHAcOVr/6
3/Y7GaHSXMhUuJXC3ie5rmjU0R5YRQxGnCzmw7dLRvIIUEEfNqaXRWnXf2N/xx5P7AAdvb7j0q7X
M81wLZpHy036xYQpGkg3awOLSPc+ZvnnP/sc1tnmEgJGaBnZF6E+Bhqf/T5LTd84GdVdDoIs1KsS
Q9+J6KHJvuzIWIpT7mBAgSBJiERJU9DvrPTEl8GLOHCZX/vMfVlMdCZ0JaFCv2kYGzikriCY/6Lf
IkrpCFg3BQk0ZYQblW89RYiNMJ2ApU+GvqRye0xLkF35v4SjaNABaFC2cKcR5ZzRNdC0q6Bf3OjU
zZaJbPQRndLBg1GXN7hsKSUBLnRU4ZlgeJdyjQGt1h1t+vO7Wvek6Ock5E2BmAYv9lUk0m8KmiuK
m9KPgnlrVfkpLAYq4GbZUPsgepI/EJsrcIKrAwydFzTy/rJGUGXgB0O4GLGxqX+YJc+lYC07IuC9
qExahuqH9m1lJ2EXOG+eauR48Cf8EL2m3169WZBPVlrxlvt0QIWSqsWTEK95Z1uQDmVzw6VRBZGh
AKMC3Fak5KODQj2VPuAYWOLtxeZsAR9eJ+vxWm5K/GmaZchjTnNk1OfbnVWdiRmN8KudMG7BTTVJ
hVBe1ZuAvTG8g2LUmVn9LuzVbNyZyRVgpj8TV5VDTkW1NKxYsa1/AsIEuMzAfhrOsRpj3BZTeE8O
Mr0FQlH2AuoRouUye+CB8ODF3PMHwvmZBQOCkXMIf3OtjmRyJop8As/wgrbCVZ5FG/5sVcM+ktYz
VcGP7WiDflyyRDpmdpADg7mISony0d6NFTaOcrxqsjGi0K5/ssFXSbNl2mqFK1goWXkAFK5SWkbW
cSlNnyIG5pAUQkAL7i2onSc0e1pVdMyQI0afQvZOuOFDx9RnNgHJXq4xXVzEVE630xTQ5YyKtfyL
nK9fdFNhBasAmznQAYqYi/et5QWLhY7TdxIvzP1rm6eliPS4KJ9r8e5Ujhfdg5Dkq5UXhr6wFL98
TnlAnwnjTVO2Z9Ak5lcO3KD7gapPaMo00HkU1J/AkJK9v6RRtuUcvJ3UVVS5hYNyBKZKEtTvqIiM
jRtT2IyGiH8OupbjfKpgeykThgFUScR5+xzAGxgDwd1fpa7Au/6cLtOqlk57OCF1fovWiA3NeQ6m
nM8EKi5co9iCEj9BOpxGWG2HnNyirD21K3wjJBX/gE7UaPWKHfo9Wb4j/qntB0yiy5vjZV7pNCyQ
1da5XX7RNqaCAsRcDBHy+ArXYQ/QJnbEN3gU919VuglpOTbi0bNDN5SRgc1ib+laQ8/94+9xZ4HG
fcINtkmVCczSy+8qYuUa+j5nrFZ24bdy4kIIgbclgY91XcQ4hFKEW90shpm9fwY2yGK8BcuTTbJ7
1KN1Cz1zvWx2eKIIrBJ3YhmB+QFykdJS0KJnaBQCBBUsf9LshmOu5Zj+hNAB3CKaflofUVHh0zeJ
//+SBF44EHAstnMH1IqqMjxPV9bkth7YKdqIOfh59KtLfwQHYgu2XCQGk9vdsNt5PRyGc5pFTEkP
XCY9/TmqQYiBcRL6GRkDKnDveTMnLJ6NsOeMByYgxsOw8ZfcJoxbwYhNqgG2+b4WZJo7zRXyLcNC
33ynPtSkCiKk9yjsz/64rgD/ElIxsq6eCpoq4ZeF+RWXWFA9rictp03vAusGjh5OctgI2E6cpweB
PvYG9sLt+F7rzWJjx5w2iBfMw22ZZFGGqW013r3gwDJzobzDDj6wBoiRqWMP1IyyVuJ/Sq18s5HJ
RRO+Vj9A6LIcVAshBKUDq0mp7oKS1zBX6J71qbCrKn2H/PG9udCC7MjbyK853ZXhI/zSRzn93yQt
6mkZzUkAJ1dKOrixpmB+MpApqdwxbaOIy3o+IuXKZArGQhITaGYP4brRUpWGVrMY7ddxau3Qetf4
MqWtjo6iUbVlk9pg8pQSqolXMUYOSBBfZKZXNQK71s9FIkfd/K/N5HQWuDBzGp4NUHQScSkRVd8b
LEdXgDroeo6c2cX7Aq98orcvnv350TjktPVziY4jTm2d8BDR9erDgwFsd4GYUdWV4azCR2uRePMS
Z14x6wt2IS683+rbz3w5RsxsKBWI7PTPyN8ABsprWSlghtfCzZNrctLKFptT0yZs3c+B9nByYBHi
5ro1dk13h9XUlb0yuICWUwn0mbTH9Qn9ms6XL0oA1zLz0Tl1aeX9CQSXhNevSvZj2S4E+/XS3r5y
xLs/YpAmvb8of6QtE03GKI5G2LSK+pqvlee2jL0uuIhfhyFKXbUPWXc9tHZtkhct5tOIXHygXJWH
Xp9qe5ynQkklWCuFM51LIQseDUfA6Kosy4Y2owOSgBAB3R9RsIfZPmb3nuCh/6zdnDHCWEwST51y
vjuxHLMPo8ZzlEJYtxjdnnaqPDABhhMcEcPNne6egPtDR4jMDpU8jdLCFgPs8lPaiPr0wsKBIuRf
DkJfaxM9OC9k0KFzzVr6VifjONvE/L8GO3ZufKCSjtBZmSDxlJkT7/UMZwf0tCDLifLu/n3NwmBs
W2HSgYiNNK20HJBFwL3k1b67nYZFKgQWUK3FHKeG3jrKcRaTVYCBoVHEPledvPzMNamKLurBAVYs
3vKvAxuPTk/QUgnQUexFw8bGWIIywYoPJusU8BsSL8szYhoORcAGIqLQXBuxehuLe6opghrrj1HZ
jBlkMRG06SZtjr+7414Gd8JbCLxRSLotHja0trGsq4wynpyuzluVLoHB37H0qt6rB7PSq/uRaG3B
ckvH1iRu/Z6GAucUsNIuW/6p1efcsUtIYw4LWZA9wgYW8IuFQ042A9MZRi7sl9WTl0aOughA79OI
UuSjo39xX852ZPx7A4e1CDo+HyjpZQHwKy44U9ElU3oob98dXSq9tyIHhyTgjVjNwhHthP5cCS8H
t84VDGFfHtc4ABnCXh8HCWQv8kkb8IKlx+Yn+JJHV8pSQ6vopttYxlNwYJA8GC8NdMNQ2sD55PjQ
trg61yjkjP8jOwe4NpLN4P2nLuwkAjryHzTUeBYj5+3EUwLCL1VZ7dH87P+Dl8aTnrtquSfLANKU
YsQTajEaHe9MdXzvz5YQpUV/J4JY2zSqWvRdOYC1dCcqGGLkzP/P1Xp4Px1iZM2MIv9fb6avhcZB
oie0Q1o05/TEeJHTd/+HWNKhg+Qfh8lLdyhR32uGChbx0MErYSSCAM9NoGL3RPSnk7EYzhhUfMyi
ozcND5AgPtWVF0NCG53C75a6Pu6nNEt9yoesJKrUuEI3eip4nxvy3BcJtHY6jbOcUX17pcirwkEA
+dvfkgxFEp6L1Xw8+vBOC/bq/MrXVU8S9Gd0IYCyEz6liMSwz1Fd323tp8XXky0mbQTdB7hauT9Q
R1rFUQO4FNbK8DFRtOA1qS/owwXj6QOixUmfxXXGhdHadHm4EcgOXS+bUpOHD6p0/+yMS89hKmpP
u6ictbsvUCsbxXKKwPhL8G5eP5WBC2flzD9fpFISrJirNQlW6AV9YMoX1jVFQApHjStKxm/O/39n
yQpT1rFNweq00JDj1t6TrlGy+Dh8BnvhtYTLXvFTxggd/IA4uUgV/yEADcUJa/D1z+rRgYXdyCFE
I8RcQCcalIOiHUzyLjOuVW2RarwV6+Cu00yvXcAAJpDaQDTanIeeG5XDJe21CCfJbh1lf1XSbqcN
51VxNg5TgBxuZupIboGMTXG4jsnPYjyXNq2+Lb7Z3DcZ/kdoa858KGj2YvHk32M4INdiA0lAKCV/
/SOupfP9wBe724jGubwF3p0S9YIex7HyELYg/8xbaR6ErdSMAlCJWocjgQRtP1+c/dUWl5MjtUNc
Ke4CGnbzF3Z/HdLDEtrHDkYtst47jPrXWXMmY+LgNUB1eGWILIRvC6NLVzHynWnWh9Hn394C5ajb
ZM72uHyAx9pRTb+VTUdOMhNoAd3vlv/nyLRkafNlMCrMNPuWdMTXx8KP6liI2V04qXzqTPz68Wzg
DoH2t8lWJcZKWl4dufywQdeY240NEHtghDBFUq9ZEWWN/bOJJyae9T+fV63UcalPVq1x1NXg6G7Q
rapbEgV0O6XMs5rNDwKUO56kjZID9MeoncEuFhQGkunK53s4xaQBK8dfB64SWjQ2bfHT/4qTyDQu
kON2IWR0JNRWldM2u0uuyRyJCjawx6Fl7I2xbwY6Cef12ZxAF3ltapDX+wFDOtouWMnsTSuNDuMY
P9LjGiVB5M9WfUm8JZxv3/3LXutCW+M12790dkKwtukhNnhhh76Jr8gDpYUJFt5PPURGm2YKXsVV
GLDPcfzn1wExGEkxEaT4aFT0Uk/d9oJermRVxUvpUj491yGes6kitprhfTFBReDYXEQLOVAzZwPM
CHXibIQYXQhLpnw086p7Q9SETmdPUk3jui6fUSvln7j3sVNBtz/PkrUFNsraR2H+iw0BWBGnxjoM
ar3rXyXOZkZK+9gQCAEYtdRXPff4qyYSPMN8o4LZwjrYLiDNUNW2H/QQn7dyzxIJZFyYef6w2KPd
ZbKP0aNM5ZqxMnEGIgjx8rgdooZ8ymPTvHOOHtQLVSh57Po2pgBKAt4rStsPEXYlZjFD5aL0wMwE
XT3GlsKM1j3YQwOeqyPcxT/IIZxXVsU89WhkvT8Dim/uc7Q4yZHdq/kmz9RBIv1lF6AaCSgm+MYN
VmJVGsk04YIQTH22RMtrH8kZTTQHfUEvJ+9SDADsQ+V6H5H8G8rbfIV9oIud7hy43jeT+Z2ZTr/C
XV5EUXRo1Qewfwg3Eslfv8w4+3S3sdIn8gH9RjygsWErfu+MrUWqH/p866aq2fQyoLONCPLdjKQp
ck55eM+NYiE796qFjeTyeXHrM/QpLDMQNV38qamPsc91ocemlUepXlJqZs9MzQjaUvavI1qEyk59
h3swptYWego3vxPsLeDfjx2vfh7Y3WCIfuNWIqcg9xhvArVly2G8mhcScbSjilAQ4/xaysVBF2Mj
fkvhiOtn/rZQdeN1/KiGlFPwVwOz21uap8V/co+6nhN95W5n1STS8Q/Uoy7KEeZ1TfV8Wj4FbhFr
MPnIEm5CeS6RsU6mcEvey3wrCoBO35KHhqlJAuN5t3v9Y1vz24LcKE07vM+Uzyl7VxKTtRtvZ0c6
cYQxnwD31Wbfwr+p9qLLOICz5lOPJ+ejoaPu2rr0cNqZBvVEyI/V+QwBEf5ei7ZeQrL7HMx80F+y
DXvfIeHszUF+As+HCYXeaAPRKP3o6ni1rQPsslnZ+02edcCQXyUwCQo/zH5UH085dmlS0AdAmOlq
wMZ+LQ8lRTdNJs9OBWAmnSs6082ehEDLotl6/sw7jNHlHsZbdLk8rrgwB8MVVabsd3zun3o7/kov
0d7q+NlTyb0Rn6avShtjhasSKAM93qOSGjZ3auhFMaYzMpTv38+91ynXrkl93WOwAQYxrU3FloIo
q9h1l2HvdT3ufF40MHfHsM9+fzlTWGMDob4AmD9/QykHJpilHH+/gcjNs6sowhIM2MxLkwktotjQ
PPoE56otmz8PEOpVUA7G6NVQYHNNeF/u5/TZRTVwof3NN42gHGSx+Jm+eg8DQxyg8h44AuZxYxPE
wHPRaZr+yg4v5efLNCeaBNjxwcWM2vvXd0hbLS6URXZFuVZ/Gb5BPANTQCF7sHxMHSLdxSZFgCmh
W8sZqXVBVn7HDDry/fiRvjt/ZSNwCZw/wfNmWB86l46RGCn6WJtDxfZ81tqkicNz89oqWU0atf1E
uPyyRMAs+r7brvIRzKLXtyzq74Ip1lj/rh+kNLnE630mc/+a/CImbDcAW6vQfCCy3vJKXUOJkqB/
ExE0ATXMHzaBeSdmaWBgNCnqIG9rfpSMbSZCgwE92srosey+Vs0rz8jWCfBOmitJvDr6BP4epNPn
lL9zj2GNWrWe/1fGT5lbO0tZsokWnWVKAWide679L20W3BbBDGwbRB8z/uODH8UQoUbPGZUao6BO
bk/p4D/h1PDKJo2KzhOKNOQktgJNJNW/ah+gQSNmKr5poz1pFlpR0h2M2MQQ3lZeBdxBY8xJJ4vG
PohVNoIheRsraeZtz8f9BzPdI/F1MfQP5KVeTqE2Il2c7vKJWX8PYvdQUKjUzzKEXB+mAGfAnmxa
eniKu5QciidQJdEcyYQz5yD8dicZ9RJK5y+VGmONz9ZD9lVmdDSCzixNH2SR1Uueyz3w40vIoZ9Y
47HnFh2fKQwLAAvfCId5kRkimwLReYrIucdYp8KgyDMonLDpyCXfAzSXiqchvU38gn3tT4uHOkYm
pTQBwYyqw28zGSiDawz6edRkzBTvzLEKulAjmW5M5Y7LWyHH6ewHPm4gKdBGq1abEqwMODE0W5GY
Ft5IyPVMnHMrb2CPj00G2IbI91cBSxckxyz5jYPszi5PEJFhmkzXkyXW5S6afqUIz1BqlDL7SMUM
GIFt0tuAkAx0d/5Bt5HG31s0j753EKuR/l70euHjBS6P8XrlUM8CNNRu6SWgXPJziA5DI90esUFs
gAsTkJT/RnPvavbgr/60n0pcicCccUrtaWvDnmvY79iviuNucR7UUGrKtTFpQiBV2yxKhwSwA56H
izeAsuDGHVQkrCmpnOQ7nKLdcBvNc5KNt/yCKRYD4beSO2SyKUh9fg/wCztoRep+qCKQfIqQm8VO
jKJTI2AVvwR9deZdLCSunDbyxWg4qQAXXfv1I3//BAdXaKxtCPEJabaC0mtOr2FfYAUx5/OYiPZk
WzNbvlvewzjFapxwXZ0n+Rhz9iuVvpT/G0mfkC6LYQ5FPeMavaIaS7Nbs+zyTiMGJEMxH6CuBT4K
65Fcm3fM1FDKT/v3d+r8K/r93HhC2OmOnboYDF2+53C5UbvHy9sWPPDiB02NGc9RT0M9YCJ4CUs8
GV4wBcJLokdBw7xKhLso7uvL2hXeNPtgvu1iJAygmdc5hwunGS6IOZMj0xvdRd9VzJh0zGqJeDlA
tHEGKJ/yBm7Y+ZOLkciC3fKdlgdyD7FCL62LV9JO/5g+Bww26qw8rxYC6Xndn0P+cMRlvnjOWI9D
A0xGz2nZMpVq70y/tJgxbR4gygoft3PU+AGnqDOnhk2kEgiAxdG7MVI0/qJivrFEdTv3eixW9k74
DQIXz5sZ7aa5eAOOnp4nBG202D3M/K2xkUq3wlZ4nb9wmJtytTybnE7t61LrG+vgBXsBJgAv5W/n
8dFlwCA2TabeZ0N2NZWHYLbJSpQENcEaTT71Hdd7HVQvvoEth2kcvlAPDpqPXY3gF0y12pYCsCnI
SacfYKJYhwYwqHUNWuvNLHOw4s/rr6V6F3qn6Jn/OJNpisWTO2jbawkYpIpZx80Asis17C3L2UnO
8wy2qFZErpidEkx/KJRUt6Fd0sGOq40l0RlgRZggPl2hXPXKSlS9EW2Xpsdt5YM+GH0Ce5YQBCsL
3tCzngNsBjdnKq3A9/MbUYHZ9qsn13WBRwvw4aak2fn1XON1dY3eyZvepLaB09zVc/H59JLdu0ZL
F870CYKzNrao+bHonCgQkKSa0WLFc6lq22NoyR9NSbX+fMAzERbiibmTmvkWY0p4MAsmNhPcvjX/
urFIHeQa07pofQL8fC0g8wGfAgS29LwaV37VWQDj5uvDJI1OUOXNwZYmE0fHVwkS+gplS1f8RaM7
UDdV0i0+vOzHrF0z2LcdHZgUAMeI0vH80cBUFvd8BT3qSkrzhIV1e6JNSKgFANF0j21gYxPFzkAa
L1pXajv/AhFduVMk6hMCrTTCuTN0kraV2ElGaFtRJKQPOcgNrDtoIJUBiIC/noMJeXwWvFhjmbvd
sa2RVINkL3GSRd2MotX0TwIexcJCeQPX70Iy6luLO8z74XPm/iirQT3WhgjAx1YF8bVxz2jvLlRv
AaoUoIyGZNFlVYelhBNpHFAqfZ3DJrJjQEpQ4SOUHh/G4p66bhwBdyCxiHr3fcP055h2I/m4Cc1j
+VRCN4s5qJw5bzgFIHNSTE2j+M/ZNX5RyB6u9pLn7kPCMsMWiKBD4NsBpPymafjRgTforMVSGVta
P50F22IN7qKslSFM4hx+uN6S9b7McLuykQE1nPkkCuTTPiWm0MpzMr71ymE1AJevozMuUZpHjXVn
rOkBO7cBMVK2nr7FH9ieJB0q6lkdy074Cw1Ya1ZP/Sjm3TwS2/9jJU0l33QKnbQG1+bttdvBTld0
dCt108DgNCuAFdgEoedWdhdCidf1nDakoiyLunjtB6x+pT9sRlGFBqN8pkj4fLJrAMdiHb2nUfKI
UJ5gmwnYFU53ng1T7zKCU567IkQYwSUilcQ4V56edhgFcxGRCnVRcVl6I242encpzB/Kc1fguJQU
6oVA9gqpJhcd7LrOz6it/p+oHFqoK/Ywqganp1/2xWljRiD/TxN4jdm1OexFETlwc15W62/TRTUI
5z+E7Ogsk2AP6L8+G0Mcab12cFX6XZ/wQbnPhlfZqeUQ8/BHnNwLXUJSMAcRhobtWF2OrL00IRzE
MeJ7eqPaBUInPd1AawnaQJTTU7RjU1hEqsYFjT57uOQb7iU73hwYp6WqrcaYCLHPbryKwiRwrabc
K2LrEoSJpVUu29lsgRS5YNSDaaFEGjuR+KxquTI/P6M1Og2Rr/YdCf9XRacL7rZjOcd2VCgpecm7
nT6A10Xq7C8/lMrEtfthpUXAJ0nli3l69pdgjETDEv6qJMkev7UNLt+wnFUwtkiNaVhmHHzTbOrM
dNjRCtUPmQDjMVynh0L6eHm6xJsn3GGzYjGhKb8OO2zUjRQ+PY7etxuTt/10IM8T7micfoxUfyDO
9cb7GIBdXE4Sb/fEb0kdzpEDgiknAlwf0zRiDqZatGnpQZM3joCM5CcyEHM33F8PKNQYNI+jyak4
yCe7Ff98BqMKtCoqwie2Q6XqJaUOf7+4YvceiV/Ql4GedlVAFiViloLEe2foIK3YPCopeh44706P
YbP6IJq0AJxwGM7d1X+Pmv8Wasp0BEkPLUwGTPFjgzcZbsF5UMmhSwMhn7VA0zjoNDDjMvLcDdpB
Se95WYXcexWFud7Or/ZJpoymmcGBzeDctZOLB9mYG/sKlayziVmS9zCpaeEiIUlSDgy5lUYGZiPP
2Cz7gVMNrWtld3DngHKe9ioquOf4xoLFvKRqun0ehrpBHh/JvmLi8w4xApgBoowBbPCE9/QXKGqu
o6hhsAB7dBgo37eJS98wjlrLsWSlEh+jSoZBU6X2YtnGbtEOzSlLNxPAAodxzuLYiBMfgSH8FlfY
Eq5/LT1RW/5waJ99RyU9IID6z6QNHyzqLZhe/Z7l0SEfYIkZQX1U+Xz95rprZg+X7rHV86KwlIkO
SQak0mtvj7sX73/Ys2aMfi4RzD6ZebaBdgoxIHbJDOYPrIxUg8ZOb51PMssfIIwao4vqHH1+2GEU
WXJibNewUCdE0gQdwjSYF8HYZJAxR/6AFnXstQebf+OS7in+s9w9nmrTujPMRnPouVUt0dExy+Iw
FgWrYHPVV8xPqnzJgAQhATRHeqSC/d7mSuH7sd6iDNLQuD5THAz1rSrv4hFqYu3lr59o5TcyZPKh
UNdOc43/YksMdnPmCgVO1ONKJyKPm0nGo8SDPbnIpEpvIqpOn6j9uApVULJEIdklAUzyCecTavHT
ekVLXn4C9Zfl5luOa2IdRiLJg3/ZkQcKWWpGrRTxF+6aBuD+pMzehs9faUnZBYldmEaR73z2eDil
iV3ck5Ipu/ptwUpRPPRjloseJsrDFQYXG3m7+Unci9yMLEH5ejC+WpClRcgVPgmPIBW6SKLNzWQv
t9Q/GWKdLAlFpH9EaVMH2XduNQ+eka4tWLxUYTVfVCxRcoRqC6AKgQZz89UDpFob2qRGvwhgGS3/
F9F8Ojqk/OWKz+YIiSZCLhY5iTMWYHUvZRNZRRmA4Sf8VG7HjD9X1yHYfvKFnWZ4N902nyRkJYaS
Cd/4t/+rTztDQMj1d7DnzDAHfzXjH2bIx7Ja22t43g+6kbKkrP7359hraMznAVyKMQvbmIDYpSfA
uiX1LKpxc7snu14ovGUHBCAjKzmDk3QDboFkTOKNCp0ZVzWujV1HrqCxZvXnqjIaavlTJ7feU01B
CmJ09GCtxEMijpYw7nstmmFL0i4upkxeGwFbCB3thk6HZVrJ003IrBwjWM07B3EvGiZ9fci8uUZe
rQmPiSscV+H/EG/0A+z3LV659M4NxJ80ktfFtHsQweOh4G/AArC8WEpo+oXPUiTkb+cDC/hNpKiM
AE3vgn6VQctk81Lzj42JM6Dnz7ozFyFcx8xby7Ht2BVXwkMsNtfvK7X5uE/ajXugz9vKcSecA6iq
aAGTjZ4wOlZoyC3vyYNG+rpnUhmd6oj9kw5NDoBJbfHcrtn7D6nfdpvvWznhjyoPfzl0VsrEWZFm
XKc309k/sL5t51b6iSn7aT5UpDGd8UUHULtVvYuINX0DRNQ9MmpomS8xNxJ5y3QGB7ORAIu96u44
N68uPHy4WAPtAV4W+HRrEFXiY0EsBZx15acGkF9cz+U/tYbnURRPWS6coNUS1Ei9g4/r36diNAdO
v1QRkV0n/kqOv2lZTmsZr0P+nS1L1LgzgzRmyxyxA0hBDJsgarJk7VovC49WOQUN9QCBy0H7mrRj
pfexQA+laPAM0td4aCRECmEfS38SQlv9f/8medkABYT/ynkyXYk6xAkFFpHm46ECgxcYJ/U9BtS4
xJIo9t2IuCA1VIwr4WKYIOXUoDANmyCDQDLP4TaCJtgGXwYAoBPR9lIVNMdrXgHH1l6wz8im+IeJ
JlMsBXoxB1h9ufhZspk8lqYhykpA66cBnRIRRjrxLhUpw2s6TUc3Rtu1i9jPKsvqQzH5s98WdiEy
aEl9A8rMuiLT70R2/Q8DpN0NL4fqa9qGy1OsWLWkJ4jCV4GaciaeWElaXuXEjawULSbO2/Ktm1rk
J608WFgyM5Pzymv0Hzd/8I1d9DQv9WLuWVA+bkVdxBM0uyPHQJxVQYUFGk+SgjjW++kD2M5j9wkR
dQuIvatTxaD8g4XxChjNXeWzh0UnRB/qwjgPCUmLh0Eqxfsj/f0s2raT4oa4y7jsjXqBKPIEZa7v
nJG1vsXzizEq5l2Fa8ggc0KnuUfRT5IujBe2H7OBuS9UMYJaDIdE9fC0xmkrNSZ9HhNXPutGe1A5
6kuKnuIZnPfn1Hre3F//NVqdQ41nTJnvEUgvoJTkBXPzLVZP+J7GUzbWdbrH9MJGmBJHqQAcbvn7
Db5PW5pZvyM7IMv78ajhS7aluV9KAdpOavt/3GHaT9TVABFObF94TfazPYQi7q+qCzw9CsQyqN6f
lEW5ZX87WcgITqggdF+T/yxD6I13UkWUQtTUMU4Sg8BPRockxGcFRQVGPUTvpk0wTjDAb7Ozddnj
zWqJCynKwtace/o2LLYAvRy6lYb5G1idVYWwmo+bZIZjUpNyNv0xQFHxhZilcl0t+FZEKs2ONEAA
uD9ssM6FQV9X6w+ycBCkMukUcKhv1ZjCkT5ijNSJkoJfe7QRgAWVIWUZSLSOH/Y3ZPTDsp3EvZ94
X6B7eAqsqwA8BGUkopezw4/zmPV8pHKhmVroj7QzSoBvAI7swAIxFNM1eZJBphP0Y+WA4txBeGl6
URHT5SFG8rlVJBTuMA/tr60lb2jWzf/mkFasv5ZEUdUjLJZlpNeWs6A2p4Fhh3nlTO77bH2vlHat
ObjGzucVEbG5IvBhD7JHF2gzxOnvH8dGk1mtxlKU55jMz8x1tHoph1SKlIiLaQRmkK3ST9KzOScW
V7IcLWi5b9Gq6aMcBIIVEohTBED/VTEgWKyuz2Wa7Sdn0a9t+V90vJVwLH4ms6cr4K+Att06nq5Q
CkiOK4lP+OTi0Lyfh+850mn011jZ1wAbSHHfppV7T/trcsUbqLIdUjiovVIKGrSgZIbl/0gaNAX/
TAuc2j5HU6NkAkQHCrQACNIa3Ff7ksIsGMW+aYfFFbA9jHWM5+fnKEBb7/DHBLi34wncclxUYJeH
n2IVOXu/xT+BvihQUoECa2nrfcy3ZgPPhlSounPs/+S1aE7BxZNXgqmAdIrLxsU7Os+ehp/BgSyG
49+WbVbn6RzIbrMVILTmCBv3C1u1jJgmkF0GWtqvjp4kk3+zOBwgdUjb0g3jkmHSacErQwN3XMKd
2horE+QTXz59p51+Q2fSsk30jpn7KJeVZNT/HKYzbAny3qzYsjT33KWy4rq7P/AMh9Ew8nKzZ/pZ
DPOlRTRnBj9ZjCVXQRbevOhFT8T0/0a4yzYJnOk8xDGdwtUYQcVKyQpwhju+8CTQH/Nbm0EBPNFe
nOfijOAAfQYWIyLHEp6Kgr0siNjyBHaExOKepWSjC1bVSw7YI24Jwv3t1c+s8lrE/lEBFxyqykNo
xKqpJwIxon2kX3xcjlxgIyF2NtV1rDxH+m0vzH/3PckKw+rh6SEWNLj22YtAeVann9SY9d9YYPhb
Hsa+zQp9e/tzyULrGJuTEDqoUUJUAjjoLf+Qsx6D0uHu6rOq0uI9T57wCqU9jRVEpoyMNVbO4s8H
JnotxYUz7ejgSN8cCbgMOGSZHM2mM2hg/L+vpV6tPj4LmgPRYGtegwTq5KTFvxCvu9VXjBbz3q99
gknWLJ7TrCtcvSrf6c5zr1hkfslhCZy+lDWCE/phOwpq/vwByhcgQqH+ET0cy+hoEgqLCeOtl77/
kgE3IuFPwk3D23LjP4HavBCm2zfJtVrGYj1I83l9Xq5DJPxBQAayNgyQn67FTNxNY9Iv6zAHHm5D
n2ORb5WTob4JdoV1fg1smv4BlVzIkXKOGsqzZOUZEZL0lk2tFvn0kdg+1Vneybym9m7e2mey5Vcc
YiMesZoA5fAXhVtm2/snuTq2SYQaajyw1v51oMOo2XD/nmLUyJRLIiQE4P+6Luw7J4vdqq37FUEd
NxSSDMHKJ8GPGlsjAtLouRlvYxqnQ7bF+mM1wPY6hOFkf6yUcHd5fd3PR33rPdjqKiC74tCpH9os
J1V05H7N4cvzTLRET2Ev8YDJ3VfoKoprqmI0V6WO3YYiQWl1xNkPelOWoslloVqSM/cmxvKYhN8y
Oy0U1TnU3IVdKsbiSu9+lIF+lFl6xiuPfSs/X0yVF0v2xzP3m2jBqqyxSnXbzHFknFfEwPH7TUFC
+nqlukEDOKGBvHwhR2RRwg9I34BSB1MUrBG1zhKkiNxf23QKIE09EQ0Ey3nsAm+oVJv3xmjgTi6N
bH5T+wRktS+HgCGz9UaJ3/1YYFFLJR26wANj6F6gc+YKttniqMtrf+Kck552kiPFKe3HqndRMTCy
Rx6nbx9pihghNpna1/FXf+G4fg6zYY9vzIYvkGCQsvbUXj33p2LmpwTfoYbSmVnISEfP5nB2vV43
wMf66RRWjOf7cJfxpDEuzQ6Cb6GoiwGAs1P86jb1xVo+Du8HB99IBacau0Dn05lddNhtrOLN+ZE7
3ePxpYKUtO5I+24LJHjNlt6v7BmnlAghgHwkjHWo3cjwiVLbEUiE0la23tV7r0GqJM2CD387qahB
+1WdCQebi/KksswYxtKpVUZRfPzYLlBRZ1c03CP0Arc4z0o2lKE+IlNGKNOtpvlKeT2Oefu+hQEL
mKSoSYSvm2cUJxj/ymwB3k2wwiCsQSDpuNx43WEHaNe8RiW7Lq8FCaUtWjNCXpgNfB48US06dJ/T
h8jXCIdkLONvA+1rDFYyPnnvjpwpMW9qiz+V1VbysqM2B/Da1rHi+5t2cbmUdMA1zoGbtfW0BYPs
d9OS0H9POzVavJCnsn5Qc3Y2tOP4vYvoWEDncFPUKt5+u3VEdjiDnGES5RNtwH9TFRgM/0UBnqqA
J6L3t+NXKNiuMVoAeXMUc9A+k6JlDEhHP1g9C6rEaxzDRqAmJtoKQDhyKZrEDJWb4aALnARi7IT2
BBFOL0NeTwB//Y4B+fvBAK2SbpsbsiSGH3c6juabIBB27E5RszKhXSOryrtQkgE83HQsujxqkBI4
P5n1sVXlYVyFYdiyk+5sz5w12sgnl+Je/xnBiUa38xLgVmcwDsrpEdTXk68neINTP+Y5dNId/a8P
7h+p4WvPqG4VQWzZyimTCv7XgqJl9Zhj/ZlvXI89CwW2h52giZgvuRI4MQfFlDgbh2yIi4ukHOGb
NSFKevUDZE6hlsszTVJKADh5VpZd+YDogLYCPqQWWc+pI5hTw4dyKU6nrvorkFusDjFVyOk7PO8Y
U1GXenWo8+6guJFJlGympvcpCn/9dK7CJ2kDfJ3LZNf1Dlp7g0DSwqP4M/DJwK8sSK+Qi0Y0+w0K
M0BpKbLogbr0VWGMy+WRCVp6Pqs3dJuvlKP+LqzxpKMERGzGn88iUCyAbmjKnJqUdWN0+Dt2pp7T
Y2nO4zoXm1lKrq8JyU9t24p/NaXig2b6kaTIPfv2TGieMVrrTqxYIlT6l6YpHko2aQkXoFR/tyJV
ARM31t/6LvapDUCvMmyu3gtE8mdp6uHuVZHQcvRKkjeP+j5VgffOAXCC3fvDK5zFiTdg0DiwTH30
a77BneHCFWJAziLiv2rwSMqyspgYJye2cbwk7JLho4wWwzOfB5B7YNJr5FKbm4q7DjJ2+4kJ3Xd6
vprhK/EZF6N0OhxL8UxRcs77KxWfOZPOhw8Sem+x7aiM9JLRLxVT5TdT6BjxWWXpBxCSh2a+QsqC
/c5WoRXqQTHmknuK9Rh2y75oH8NHvNSXezYZWuWWr07ucx3zXrxZf8iHVya9hkajceFcVIYh/GXf
l2zaKl5arE9mPveGlkqXBf6rWWcd6tpfc6/QmU2t8rMshswZZSe4DeNicbJ5rbao0r1K07f2rSZG
/t3jHjHwUqY+EryeR90vqX0cDT8jJgllqBq3I0DSnFf9yBQErjzD6gb+W7O9/7ZpXLabW2pYtl8Y
xI1dc7lNEkg+aAuBou43GW6ezGDhowt1RL+5F07yOxBZ6YhDI19FNjtb4vlJWVmrxhhn1gOJ8RPv
FVr4FEBs2GtJ2nB13PKa1FUkLjrr/rfC6FwFvCRZ3wTUpsxAqHxatRJNMpUDWjocFyJSr+qeaoFp
gKc4dyYePSSQ4wJXsrW1wZ4g9H3uU1M43ZO//zt6fIYWo/LokM5qWAUmbN9c3N/u/dsMxmVvSTe1
PxBbOuMmHUBhIx3S5PqZVoYZzC1m/PzTz0pOfzjUihWt49wwfsGJCnVQqpfDlmdhLQsEcmqHv4v+
8B7RaNALhVNdtdbzrewv42XpcTv7mhXHEcV9Kn7bRTk/WlvnOYJcH5i+z/Aq7LnoPZFb9x+5Mi8F
x3LtMkxwSGBBKy1thvuCTZknVXAb/uuITQwYZFvLmjhpZSWlIGZBmjWGvANa+7sFapBMbSPGBhy8
OvbYdtvGgishZ2IZhjeQ/7F2ieneMnR+Xz32JLdlHoJnXiiI6CpgSjLfDkvghVh7l8WY4KnSWfYV
91igyUzzgd395HFvmfva2W9Zt7FvIhzYDklaLOsh/UECvegFzkexDJvUwlyDQQt3QATtRK8acQiu
uqNu4n3NsiQsoQ6sVF3HN0Ch9hkBMXAoKYszI8uSRUGTxzS7o0KveCJ8Y/0YCsVXoN0fWGGxOhuE
xr4S4giUFXHQOI/Ty9caEXZBhpO3T856+VUviBkXa30vL8tZhllpkEh6np/iUeAVoKK2642/j/kr
z3jIcHT0ihf4Nus8JihSDEvFyjjsXL03FyLweYA3glYo6kv9Fq6K3zLIkyRnKQr9fUgP6j7cumZM
VM+t/tL+8F1cDw/NGWhKubyU+GJiyROVtmRBFJijLDUP8dLT6Y4cwgOEfM2xcXuBpYk00bBmIUTR
0+yR0MfzWA3NJrANjLczdIBVxsDvay6CvuzT9LEfmDx4ugQPrRMAJHAk2fxkqF9CdPYsmbwYMKuG
EPt1g+Tkfphc8Q9RNPjHTvHyBGsoaQkK3A8CYWiDX4q9dSYFq7ESLFFv/uwoXjgi9yMQ/yskZjDq
ZxyTliPQvzdrdDhVb8s1uixNjg5sS1FX3s/ojgvNhdmUdlKsQc5XTHRJMsAMTAqvqdtHmHXPxgns
QRJxcEX5BMAoGA8R1iT2gOMYcC2VJt4JD9GJUpoOWVG46MRZApvHqDG/FZV0FYdLKg8fZMV7tr50
Oxu8hYcF0vn4pj8taGzUTZa+CtLWZsl5pyNHVHmwVSRerOM7APmbYV33MLLzIAn731yC4QDabgiL
aYCIkb4ABrqwdByX6/5lzwqcR0dZj8bz9OX6gxyAMR3Y+q58JozlvCiLr9fVbi+X6GO5P1Ju8pwt
bNxgf2WI7e8ufE42lA5AYJeMBr1WDK7Yw+laqPjbQHpGwtMRi15vLx+4q33/nmtB9dI/BtuflATf
LE19KfXlfXfE3KEOKRkDHzRpiKt4XPVIzYEe7fa+IgkLqe//NWnxm+3GhVrKKTpX5BGXUuid3d7c
nkayc/Qit8rouK8ZCdW4nwJfj2qe96C+n5SdTDcc2Md34W/UDt+XS//nkthIMt+R0fpV4smyE454
Y+Ds1OaFCnmZL+tmO+KUqMpY0WlysgVDsuJcpL1PAZAA1LJUzXqVPw8/ui3Rwk10L8cxhYohbkEW
OyAVd/RXbt8Jvf1qkh9DUuY0iVN8Vu0HBMffJG6494ZQIdlamFGrKasA19hQI31LUX+FYUs5Kejk
1JblJ/LwplPQIy/DvriA5qZfj78iX6kyLdDrI6fIFiqocBMjHLfWe3iJrMkULo/OHXK7RrxSb9zR
3vbgw9+ZK0a4iyPGdUiY5HCx7M/ewsPI2sHh1nI1W8AF7DVjY1FJnMmuO/QQRXB4cTHzHWbIWUoM
0EOmBbDYS5ciKGYToY715oD3cuy1T9MRJw1LLTvsM4fZG/NZRjp1Dpg3ltGEIH7A4NR//y5sCYd8
LXTKw54Qvm0ykHE2O9xlHcHirw0DvGoABH8RadvQaL8dh89TENGqSpYBkl80hz8gy6htCXgjk5tt
Gp2FMzvqm+IjATvMz4CeS/Yu5NxfURwwLcjiWL2nNtvUxro7CZCJz3b4s4wAz8lXon+fHmLafaHt
dkrL1Utw4Xi/JuhqMlLbj8DS2JGfej2LnEWvlARymHDd/Sr/mC2uMxXHLyNOJPHBcc7g+t878/LX
NLVrLdOlSGGwtlNgXH+XQB25ZGmnMKzjyl6zLjoDSDpXOurkVEu6YaizK8OJ+EVP2oESl32qNERk
iFWNIfKyNlBahvqSqfbT2OdIC20AgBrQSEZpWn5MkFNJDoSHuuTfK4g/f/v0zrQCjbapFhNQt/tt
9flJDPmWgo3DqhF3LrbnRU8Vsmnthvxmov5KnCpXR3YVK9VKOvxpwzVvuCtjb1kBTuF+eTLIXPcp
DEcdydMBEHdlSoKivgL4H9QzHqruSJPN9Hcd51PtuteGTU5e1rzpu1etfy/X+Dq2jDLW3aEJ7DVy
uMDxzwRd7U2LYPvIiBcTwlBgb3gi58o+V0ITTDlfuA88W/9jfdBZVkvKb7y3BFCMFErYkGZFaJVB
Khvi2L8xD3WKU3MUsq4jgAH5JJipfAIS04GoAebphNW+E5SQgO/dJwPYxKAVNVFb14P05so7JNBk
6PD30kfl1pacOj9ZvPY/BnsH9EOcGSJG2rCWE4FlgcyUpkHAbwCEZxsIPbavUQ55RNjNOZplQeOj
ckoOhMLfyKRuCzAp4WJrkrdqpI9ucJR7IIf54e766ODLyVGJULPtvGP8GYVCmhQDGYauOls2WC33
MljClmtoM5SdTgwDX0zy+0g9LXiH7iUuQWzuRjMURdvL0wYzfr9Ky1LHXr6M15OmVGC4qn7G2a9I
IdKUwn+F/S/mUFHQ5eaXFPS7zXNgEaCsymCos0vLMGNhC25IENUyuOko4Mr/Xh19/cIxwjCkC57v
xvkNgOjgJqYklXeO0UVGq6rvln9GEI0QkB2uvDkk2z2YK7NsoJyu7KNYNMWVy7X7uTdBaqCWuxgy
hDQbi6DzggEyE79/ic/+6HRdoACrl81OS/rah2eaxyDpefAQDlghHD3lImo58RNEHaQnKVvw4gAi
/rsd8uvOFIzoYFrrkoQtRRZxFy4qooiviZf/m4ngXVgcP2WM5rnd2InOP9tPKj7EkFzmXgb+RRpQ
uPt7S2IbGqQPXJMQPMyUPOlAZxzppAgmnfMNzVsmAmBHTh9MzgmD4nTTUVSRaqq/gR0pQYDOrOyZ
SxtSJUKVMrRb+gClMLSd6BOqlRrqz75y1GsxTW6bl/ItQCoQm5EA3fe89B2pNwTp8Ade6DiCR+zE
4yOa1uJQfj4ayJSKiT6G9v484Bumb5zCJGB106agJPjroLZ074BTC+RQZq42VAHYAzDU+7fTTNtH
kIASRJR9vGEai3+gb0VhG3yKnDzmKIZgMeviOCnBwWvTTO9TN4fL/scDGIp2EonKgoqD6Vel5Z7k
6UOiSs+zfZraVrvlcQHpd02AfkfgP1F/OKfT6cK3OdzRpQxIIwGeGexMmmI6Jr8P11F59ZQlaj3r
so2EShu/9SWkfuu3uiG1b9j70iHH3pLZDjop/SxSJl51IdwKVrY+yiJveyHUnBzGpviIY0MUQ2Xb
6TV3xdMH57Unui7vz9xkWvyTKs0R1+WIpyt/xk+buxND4V2kc1QawXhYoVmnIu5LuzVFInl9IoFw
HsGZafS1qfGU6H7AOM3bY43ZgoL2NrKltIGM4OynmUXwvz9j0RGC7yZRDMtq8rzeIZZlbkb2XkGf
519HrqdVn1Zp2LtdUkQ+LjRgbZrZPC0RRDhBDlIO7fUW0YQDyJ06DuEqgZl7rXStYPlHuNAGrFYS
Wga0okqw+FFH13hK/cM9RNZNrZs9wDYW6ObjW8msuToGke0zJF/zoYCW+W33VLy9IpBHuHnhvCpM
jfGfCfTJowqDhUWMnuCiTDz2y0v/jDp+QcL669tH5f0sUrZIObLc6TmsYMSDjnTZB1b0ZGRfFai8
Q9D8plVB5NBIABNE8BYQMsIznkpMbxqWKbbeI9gVA9dochUd/nw7/ThgQ3Y8wo+zWtIaViH/AbTI
pd2Zo27nDKwB+NiFlA2k2H/b5q0WN/pHTcewSvG6nZ9kx5KRi3aQvfhRCL12FogOCC/glQXC+yO1
chsLMyXrNE3X/PhVFQAldpiU9ZeR6Y8LLfXF8/nvOTb7vbzYu0nc/cHp4nPjkfOWpnU5EfUnxrrb
JF3z5sbClff3Nz9vXk9XFQNTPMQklzJ3heRWVDwSseM7VwpT1HQ8PFtXqRRp6fSmE0e+tO3LmUNc
U2v4vppz7XtFoSfzkOLkYBYd+nNNwKSXEZTobo2Icy7Ku9SludVVaE7k0UHsYF+3hzuFUIXemqCd
gwWKiik4xm+C3ObUHTwqss6+rmaSMCjuQEL/r5adidLUhYk129xta2hgrvM6cEN08gInp4Kw4GM7
lJ5lUhNAVNDtobr/PIpgU7TDR+bd6LZYUU0/iWWRmRKjwhbFeyThlHf/HO4C5agELJ6AfxS3K+h/
P6UALCo3WHFE6MqP7OzewrtU0teDEnfN3LMp93i951f0ESVApOIo+nRefVhM+kM4gXXBU+3TvSQJ
2ucYMXKUIglXEbWQo2T/lYJmjOOQVU0+bL5DXSdE4UxqbBoadxSS4mmF0Agd7oVdCoCaUvM9OQI4
W1wW9kkrZg6K6/3IpKBi8ABMYgTqwvM/Xgn0HgAs+UY2AOpHhFlOopPMaVmjFL040btM+0/4s7/C
GYsDuEiLJ+Wb/43ZJaLSl5Adwq1zreayt8hH2/HBpqgktLqAFZcEBUf/bio3fqxTIZrhhy922IjR
zFpbaN2i+wXmZfK/v+Dgd7FcYwQvcHDZZDYNAOqpNCX6VFRJ/tQ/au7Wxlq+AAGyLWC1X/5yedhV
dWd9luewUN6dCV7yx85RHPPF3BT9xzqvI1T/TuhjsL0NFD8Mqu8yB0iHJES5fJk/iw5GPt23gGo2
b5THZnyRbLYhmdbI8T3BmYsjx0tlqGqschgkjA==
`pragma protect end_protected
