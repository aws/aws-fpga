`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
EFMp2rswSKsW1KETW9naXrGbFU8b0qB/m4HP1IqtouB8qt31Vk66Q4TqP//o1ca6h5PetQb0eSP3
An8pmbdXh4qAdpBI1Fehj7JF3ggPGTZ+5/kO2GN6dCWWlMR1+Leqj9pW3QmdtJgcGV+C0lv3DOLO
TB+iQaELaeaMqZolHoH4XtiKBsnn0ReXwedoyz1rhhBTPlt3cJfW6UQZrsK3mObg34hV5Wefyb8R
ZLewaxYYxz/kcvJdrzZyduNmR4l+6m9Hv1Pft8+Z27uj9MIN0+BaqbR9pXcInBDmMVZmQWkSoDgh
ZUXIZjr/StJ4GkHKOpaxo6mYRz1bsFCiYeTLyA==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
MrtXBZNxv3PikKaZZ1lqaUSqtIjZWccK01w+zMBpPjHWcYRmqfOXoDbkRYxcSLXnCwVZGAxYRgJ6
EaH/2ti4qxpIhEBOn9LnT8YCEsv2jWqnu390d2kpXdmCN+6KtbiHymgsoK0gfq2hMpRUAXMQkCgN
AM2qhZiR2BZWsh4SYTQ=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
IPTJG4Ei3oPFdFBAzvzHwLKQ7RZtusBmt/LpXqGkaaWkD9I5bpBtltwm4/z+rNF/fGVAyJcBpwO+
U4fFzBlPXdrgaws6au2rjDNPphlp94/pSl4tOb6Q1paVuMUuyFgPWkWXe5z1HGkxN+eJj2Buyt/k
3jB6RBIb7H7WgoKfG2A=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12016)
`pragma protect data_block
ztH3sTUIflI9hQ6yf+ouzACWgnC4hcuZuJdnKOcbmTT5zWlM4W1zR/wvUWBlddp74Yl8IqfLhse1
x0rxHrDZJkkTblfwN4XHN4pgQ2za2wF9WErh3T12SurDwWhfmm8xEAcqJiJ0/wfUltmZ5k47PNWc
h6zccMq4oH8iI9om3BOcXDmz0u3Hu85xBrj+xsrfCxD8MSkajY2nbAts5iWYDrkWJjSkgSII3y+s
GtBRFh03TEZrx/ITy3r6Xt5WuOujdXi05/w6LKfUvdxn3ZOLuNFuCzq9qgdTi6NaF7qFFF0Ghhwg
aAdHFnFpPMGsiyEB64XmKMvT+OQJhAH9wkG0EmP0VfI2n53YGcqg8WHGLml5paJcj+2hGzthX8J0
GxObGwMkg4CBZvzdhPYR9zZENjIuYsj4/0eWSg6cUAwmbTHpc5O2gTO213eyDR7sCrXJSHpy0GbT
aCAcMbhQMf8cNwn2wJDdIQl6sKhXaFmsmqpnIt39E4G/y7QlOGbVFj8BCOahJhzqzfa69rC635Fm
2gguWh+j8KNNGCP/D7+gXpNW6uZLP4286+9a6fZMC6SzyQeMjxYMtA8ShU+HTtzKawKGaoYGq+Qu
hYdJa7N+pNd1b1wpxF5mtwMJLtRdnZbBzjE4DeWWaraVaE5MffNqtJAM6e8KTurhuN0hOSOIYZfX
LvGYlJYwk6tHNq9PnmdV3lJzL3S8TMh3lAUqRQ3TY2vExMy0HTq9hr1/3SDeO+K8dTd5ZvXr+xsI
PUlKWeIVWOltAUk9EeYBsAdw2vD/t3Q0SUQIFI8X897jSPgedHin9eIskpwYskwwZrYqZ+p7iVXj
BnKh20v94LiRXC6rcdETlsez8XnDnU75yEUJ/0kaO1NIu0C8sxlD5eDAoSnzRyk/bVG4rqeh8DHu
f7C3N5XmqmGBnJbG5GJem1IKrfq+LD/0/BgKcewcrxAK1u4PvfE/6isXJo5MFyxa53ZQ0sYvdb+7
NxhzfR8qOTFv+0mB+pUnbECf8afvAN+4dnleYALh7YYDJmPhbz7waVMlRja+75s/K6WbIPh8eqxL
oPdjMCwjQl/hAX+skNnROPK9ArsU6jBZaUNQyMtJCroBtuV8sFLnN0JJFPH/eLjk5/JOKNmfrdJb
Tz87a26iS9vqguZvbkCg/Oa6phEkvRlLB8xP+Ofc017d1MKko+Ot4sTsIGLkxdBtYy4+Jqou2TC9
TBnsCAtJNKQ3T9K5BnA/pTH+NQreBE217gxcUr9+MnUBKT/3OXYjh4O5OIHZjkqy/0LMaVjSnAbr
rI2KnSAd4f2xrJSATZgVi6I8TI9murhCOcV9B/jKvOTxwchAtiulztlwP8oYa8eB1kN+UZ+anMjH
9A/pie/+djnSypgepzwdLb7sMft9O0nfgoTK0YYflumHYxR2R1FL7EN+vC8Ztjt1SpnrjUbDSwoO
mA5uOsHOO8iGN04qg9WZ8UWCifzrP6esPkYgtK/g8xMaG2KXdctTqI6DLa7ALMl8tSoSDUK76uA6
YPgd3IOMgnfMl6MVUL5dvudimADia3Qp6e21BZ5mro+1lVremz0ceye3+lmUq7xGVjkgJGWqka53
RaLAjIiwhJqDMfm+4+lKDlWCj4VLVtzOUzjdUTaQK89Tk3lQ1myWQq4SPgx2REQ913xDjpiiEmUY
BIEce0FVkFwMR93by8Ar+PIj0KMfvW0U0lcKJPPi56MaZK5HicLK0AEF3deql3ahJX+Kkftimk0R
pzLIS0sULZCKcVfs+f+7wVOLd1pkiu79KhkW+oXNEWD87ECcLc35KC2h5aVzWmxlu1vfa7OqHtLN
p0w1YhX4srtDg9Jjmk72NFaDvDefEVsTOpNw0Yh59aQmuWrPn/qtnInk2h+Z3h7IcAGAsVaKGKdK
MOD1NSEY8Chnelwl4Y45PtujRfbYQkrXjX5LeCBeExEg+kJK6H9SGX0jzIduwhdnhCdkkTQpy8jJ
3X7A24gLs5G7z9fuO1iw6Z/xUNFG6qVQF5OzT9z12q5odFM+h5+2mrT0BP727FjZxKRj2NFz6Pre
gQFL7T96Sb8kBxjRWFrQ3WkHkXyKU4ODOEd6Vp34paCJUNKxlxKk/YQ6fTs/0z6zwFvUtIQTK0+P
P7hdHxYYOQnzCoMwV6pJkRowsHlrUlUK69KGyuMY1DWYHc/Zy5yyQxY9muU1GSbbdZxECPezp2Ob
XIx154orhqlQNKMH37zNf/Og+jWk3TfaTqK0ehdGZzs3oBzKIS0K6TkOrgxFal4iCG7EpBrjGUac
K//X26X4nUT8V4WGUXzrQMKakIwySh6dBbftORPTtGEU2GpXKow+KE+xgXtqZ6A3nOPzaQpAQtRW
jLrVZVfWkjO1GSWTdzO9WyTrk5826gncpIYfOTGRm2bpXsbkQdAsIwyFpm1DihpDN8Hek5DAU75n
znvnO+50+20XSzJzouRyuVd67NdVnkWP2Il6Q9u5MgM7xohoym2fwIgR2jRsQxDbi4vt0i/3ZmQy
8izBJxIu8YKyoqMZ0IS7GoPuA/BId5lEde6qUHsnV0EHdw0vjBJWcMZ+OsxgM1V6LT3ILsGBlO9J
DzxdnC2ok4Sy5myUASfI71mJ/nOEHt7zhmwrhuFWPoyQ+O42nMjNm96qOWfmB95yDjtKOiz42neU
LEd8qtkZiKI5eNNjLLGseujMF/mFSsAGO6bWMiprKcklItSK4HEw3pkBAIYyQGITwTSUk9SjGel4
gf9m8P/XXpTicljdd2uvZktAJpnMUcRu2qxJQa146mB6PLvnHSIvqLv61PvBc/3Kj5JiexojZs3w
7zPVNeZCeEcOtZy+XKoY+Z2t+t3p8NUU47pW3WTxSBMraPpf5R1U60LvEcpTj+sQ9Yef0NMMe1zp
U1f7LR8UeWD4E14htOdD7XtzfOum3vDVvyascytVlQrZRCQNquf67hO4RfSOZ9n9DlKYmfAD5cLA
N9QHQ9k5l/B9RUmfkXRRfYVQDE1WJvjI/fDX5rQBUgMc2ThtqTQvm7WJVsf5ZKfCvC5L4bAFC82n
56NNe4Q+N6Z23iFb+xnokXarxNSuwYgFb1xhuj+UJQEl26JkpjQwMIfXixODmxCOdnsdBXJVZDyM
frV7dI/2Tb73G804V4NFqdj5yJBP/3S3d4MHsJvrMSmAAWEWC5pKY0qG5g9KuLm+oRrRr/YGMr0V
lfkJMb2bMk5FGYoh6czuW2X6WdaC4uejyO+ZiQU/F+fFrs9YMjh3NpsPgDVwhtz4E8mq4tAdpUfK
iYX1Ya8VUYpXnq5CRZQicOUfBlwdgwd8Ei08Vu8t3juKUQuRTZtd6kRv8tHdxHCD/70UYlu0boB0
yJUAgJNC+fYUa9ONK95vaE0254v4fkhQ8AXQ1EgievwGX8mYLmMLIX4IdOFPOkMw5eNfiwovU/Ye
SjoI5gC6s2htTtwINzStdo9K4WZYt8o/mAfLQEB51T3vpN7AsrDdWTyG0hihcCg3X/Mgt9nCFq4E
zkdWRowqlTxDDdA2bIkEzKZjhfhJTsziS3x8i5tkrGEIIjVO5gFzXYqC8k/z7dMdMnrMvlIH8+QF
6yZjKDfttL+bsx0qTIxvu/0Tt6wyk/to8VavvcaZ6SeIs/EtYdnTSlRiH6q3POyGpB1anoEHAEXH
X1yoISFj4YsqEZgZaX5iiW26KzzMfCvGP5TNl1+KfnLJzYd68dFLp68GsraIetzvCFQd1SGkDg1/
RGX2BRDAvJTxUpw0sDVlrQRVe65uyqb1NiQ2awBFyYfFsIWwtfh1Uiaxrhv/juXrYlTZYygdaZdt
NYOcyv6X9Le0rctc8zQPr6AVdsfTLqZGAmFn3omDV3lujm4DAbew1sEEY/rT/w6scN6WPzk0CRoE
JkgBJ9zU1ktAbQc9UhCrF+gjBX7usps8ovL6dGB6pRbVInQWCt4Anp5zKDFwGaJSH8eSVnrNlGsl
nnkbXJJab//eoDe4uCJo1M4YUZVZX23X+vA+OOCD8M831t6PkwT334sBRU//GdOcUyO7N/A2ekOs
Mp0YkJlF3gfUc18bmcql/i4A+4LkokQ/QQ7K2DAWGzM+kBLvxufH07JRNCC+09aLF8Zbnm3ta7hm
UHyAKugS5eG5yj2/jG9NfCpRZye6nxAvuodi/06EK+FsnPfTXPJHtnRRjXtCmYS0BjnjqDzi3NaJ
7dt74b3iel9GtJVLzZVkI3x6WfuN5oTv7e/M2zdoD8f0HZd9eLxU0mftSk6S7ZKG4glpnlcQSfVj
mpmfiaeQ15N/3mnerK2Vy/FKJ0FGynAF+ClYe+gCYEiL3VpUXZqHXFJjuVGDMmjZCROGQz3TIeFt
6oHdif3GaCjHJEz8SDGT/460UPFVpCIgZzsKa0eDKfTtfamzRv/JRwSpkqhdRu/DHJ4cSJTgFUBF
UFb7sohZBWaR5g7MAcgflxza4Kmy10skM6XI8AAS3cPPXQ1UsBdz2MSy4Vg/Q7rSbYvrLuwHBAf7
QaofdV/d6GhXhhfyud2fmsrzlEcETYUZ+xLU1Xgt+l/DKSWqihdrzZVP4A4d+gAOBLiepoGCAp9C
QFLNB9HE8lyTJUL6Z0gh6J1lQRuvGvQJBd3ogkMVhnSaT6ftXX+lH0P16nZjE4TnHJJYbaEhElun
W3Pqen7mXBLNzUjp7BFRTMAYpoRH9pdbl4R2SOJXsquYKTQM1Or9p0ayeZpLkZjMWhnkp1+QDeP2
zurJFVg3EuKLiYOQrQ/tV7HeJ7MJudh5+erpSCkAhx0oruaa5M5Si/6IsNeUilH2Ls7kw5z0W08J
nOIFe1d7a11E94+vU8EIEVmag38Gczc22Pf3q7ck1gcCXfq4PXdUQHjh6BPOfqiHSPbURNRcZeDx
lu1ePwqE+wpja/1iiDEqOn0aIhqqZSNx57t1HTKvpXEFGM6q2orL+AbSuNc8VBIqHnU2GYYmn6hu
iG8ZNRo+oy5UCmbz2Z2WtS67EyFPG/j7FSzFb//txWkrayJsbqcG4B0U611Q+Ujd3YV3F5k0iTS9
jMmV5FwsNX1qyxN1IQEPUoiDJUf5GiZKdy0N+pFVzmjhAHFEIgeXGzPeD6eHWQ7BlltZhLLcohml
VYjpiKg2Hz/SndGSBaQL3SbiBhE7R8bFZdUnyKJsWTnHDyVgC0O/VS7C6PkrDJ6cTxeZR0w7x+cl
ncq2sE16sbCn53YbVMRDRWrOL5hRdWII6eRd9ou9KpE1F9KDlbPeQzdUnp93hdLN9nUEq2d3o1G+
hsHOOlJu7whTjQCJT2JSZk09idqm0daHwMdskg6drgXSJpBvOpRXVyFTrfAZ4uNNeHvIgzeAEEbO
xNk2TqcasHFnQP7ztD24RMm9q6Q4k4Byn7F76iDJ8behMKWMzJCMIaGKW/LnjzzdIEZuq/ikRllm
Z2BTY1f/0bBlvcKoYuwWEqxwpAbo3GV6DiMuTv+lI+gmolKUpK6++tlqKG3n+GIXvq/b7Tz15pTz
eiy+0LzfMhZlW4EqZtjd/qa1b9aLBybLNWShKP3GxEQSp4Na0tgEB/XUziqpt5A00Ym2WsSxnFvu
VPKmMr8MjKdkXnDwDuORKVBspPZVwjsL+ol10+11rqI6iDGsBzZa8kq9oxQvPtuX4UO0JfsMWwN6
uwwC0WgxzBLRZ6A9j091cG+foyB9xSHOqoIH36CeJNNqpco3S4m6IXmDxhgD0MnfiuvRbKzhWwQq
AkgFUAcEA7TZYxCsZuzuwaV2x6fZ3P13stxrnZW1Lybxng4ycZKHt8W7PPFAUedPfxyqOQ/P6aIv
1Z+xrUOCLb2LUy3T2MuiQjUrBftEYkqJ2TMoAMytefxJ+r/dxjQlVo6wN/1IWWWi6Mqs2fUavLQj
278piXkeSyZnBpEarl8UwlkyGkXEZMJofHD+/jDie1YgSibRBHG95GXaazcRAm4O4ZT+U1/vS/WA
px/iZ2d3LwavSW0Jus6eLPE36r+XuJT38iYIsQ2VDu3DftTP9y4JJqzdV7GZ/k1WJyS4oi4xBS8Y
Dw/OLiGst7sz7Lt1ShIhl8gLaKNnIxwMm3WRvzBA9MdqGCffaLm9fqtiHADUzEANquXP9lekE9ND
EuBieaHQ8N4pzeqh8srrIMsKQTSUL9P9475vQDyS6UmjSnwaRj7i3YqAltdMd+ztVAF4PXeEOxHD
tpgs2DnLigPU0SEOOu5L22Y6C2v1k61IuBUCI3fPHZhFkuYwzPX6o+hnYAwmhEmGnoFyFf9Q/59L
1boNxQsGlLa/Nxw+gWJn1d9fpT2RqEbEJW5JQRVHwRFHvVOXTJp41ggiQMN/+5PBu/e+52PO7dmK
58GQhMkYgi9DrDTZgqCewj4RxlbnQ8lTrMOrcJPYQhTs078EgWzHqhlqww22KOIV6OvAbq9M+3RU
jJI65Hq6/DHavHHc0G4z3eDmS7FO5iz0ouZZmpGpqhTuRL7RlDSezpAtvgc25cxvWXU++xmxDvou
wTpAZmPV7NLwVvnckGpi76Yo24pN+5a6lcTeQ+CLmPkNH6BWsNhlMdlYNq0Tdeyh0RPqsAaLgAge
MCpq2rZD90I+6ZgP/aP9Vm4GqzC0shwiExpjoxcbDV7eA0QfArbLg3qhbMgKQuCbz+C5XloeZkP0
5rci6/Q66tLgqJkjbqvjZ+EKbbkCY8ThsYvbaTkSP4B0mCwZzne5ChumdQXkbBqLEmj3zc/aLr2w
j0d5q9T0NcnKtvgQjJRWcDVkB4FjYiVfdyEB5QFl8pUOAXYNOYVjSF5BYIdkEQneV2lSrL9c6pNO
CVtPlSRdv/JMb8Cyi0opuz4Ci00YoHSqDDalWidOXF7+ykEe3Zxzgq81Tj7QHAQaIlMaOvbpoa4c
qaHwil9kgj2rs1sC6mpk/heBxg8wlX4gbx0CZOW7Ru0roIH+yHFuUh8lU+jdjNfHf39eIneHDbjo
Z0oGrIUrqXG6YYa23f66Vx5bN28vzezU07fYg801Dr1/TqBAZ9/hI3s87+B/kzA3HjCfw6gzTC9K
pWcBBmPCn/kEKn+tmbZDyEny8U1V1HX49G3sYW+suUC7Grjuc/xdwFnS9sTiW0TW3qUnhBBZqFYH
/fVk/m4upH5ByLyL72rJ6LkcxoffIx+k/VFZKcFNvVAXAi6IHN6kJFgave+Q/OG7k4OvKJdLy5uV
N4bbeHmdiXPceXVLXAGeudTOmkF1rrUFh3CYkUVRLGkYHMTERz4E3k0M5ZVlXi2x5t65n2TP0Kbe
IZ37YqvWkpxK6WwO/YSMhWxSIr3tlwnHB0H7ybOIztSpbZ9FFeKbxoL23CWMT1qyXqiwKixSlcMA
ryFvJmyzkpfx15xoZxrK4Mi6rpp5IEbe267C0rGfc5mrh+fi646efJTa1HdpK+5zTFYDQFa/SNur
cJTvYQUHniRDIZQtijQT5/rhIS7GxHPPQJT7IJzQMfxpOraU5AQt8D2NtbBYIFybPsZIBsQLpXgu
qmd72ws1ECQQOcvXQz5Vv5C+8WAMzUIbj1l/AH34tWUyBG8FVlcJChBEi4Z6sfQAI/maJEJbJX44
x6Q0o0fjuYILrEEMR/GPtyRUEsdmmlxkuylZdeTG+PZ3FF+teE+uRfb3lyrKkdlf67QVUivsgrgU
MIKdr2LG4ZtvrGeI1yNSpNZXsdpOHhdey2WvtfEGA+Efdq5Eeo/1yoz6ZSwZPz3nZnI40pSVJnsc
kDADBwG+hyMHJe3W+4gK71aVTxES92J2RRqrZMhhiOIyZVbHiAzpVjNivlLo7BHOUMdVzpJKXaQD
UxpRk4FKKDVL75EdXFOiR+TFQWB6KqmfOfMEiiwvSl+G6ebIf9/pTtcQwpHe1j1lrlNWqn5BXMui
J0NJqCg5KAEmwVAByc+dtN6HzftI6OZ1O5UwPhldMwozVh3JWyCsAYOVPq03y2NlcqjBY5kZf/4t
5UJ4CamzsmIHVmX6lE6hJEUcKjYs4nIGYZtwOCOE0i6t44nRzssueuOwTBSf6J4M7xDsPhg1S/Bs
JUz5mRD3v6/WODK0l3FSXgB4IgXAV1wwiSCKDg5c4Xpct5EPOBAIXDRKqebYYNxqABml85c+EvGk
iSjFNwUMv/XMxlw9fBu/d8c2vwPpODu9uHIMv3DrasPjEGs5Qhe2lxknMjv/3U5xxim+/zL9ZNb3
iXedV7J2/vpPPuGhjz0cPP9/+0JzDFj3HDcIUwNNb5lvXG8oMWx3Y6xLtlHZX4Sy9KqMK85byiz5
ypON9SuJkEmDGAN9orRjGE2j7isz/LQJ9zSQVWqnHXhXFKJXc6Cf/km8/wHcYPtFjNHDOrtCFTAV
gmLB0Ca3Rwlg2TMNtGJLDUtF+BHq0zenu2Fr/N1Ju/GSHnEVByS9+x3h4G5GJRG2Ep7aYInJ3QkK
O08pPXGSXS7SUItNiwlCD+VSV0Lhb3w2LscJiGpXCVWHhN7jZtWLOuMtv6+DgbWyYeAiCcNyHBfA
a7ljjBjKGONnBAUOisO7+CIBr+bNsB5chi81auwf5kInjSRUfwp477QvKWfjR1XyVAAyYi7DR+HX
D6unyZXrpG/N1If6i5OSw+1/BbXJ/64HMpUp0vgLZgheEZpKm8PWO1A9PE/DkwL2OHbvAc8p8fF8
LM2Yq3Xym+yvESY3tRbVFwNlVlgR1D790YoOyet6UIGe5G92kHK0lx/uctlInuTzsuKxAW76CWpr
oHN0U7tST2xn9Oe/Hp+6K5gerwJO2pWjM7ni5dvkzGfatlAY7YIMpDLH7qDdX3g+nAEVsTBylRiD
kpt5AtIB91o9Yzm5rw57ZEgREioqjrAgQMZt9F4jcLwe6qPAnG5u/tQuiM0OKCAVkAyQa29Try05
RUAB6Lj29I1xcQZ5Xsdyp66ZaT6+XOfi3m9vBJDgg8zTB6BwlFQhB6s7lAmxlhGCMrxlHzMve1jk
BKJAPFlGaWeodVRQJWmfHvSUTEDhbkCPwiDL3IhHhIDJJ1BlIyRoeBssbU4G71ZCazy1haYUlUCA
t17OSMWxVZr2mnzJFwQtnd0TEyzHzyzHtWMHXPS2lPu25eHVkCoXGMXSXlPDtspsTmUadHs6IGlb
tVEij2VMQXnVKG3lQZaKtrSgUAEUGlynUFF7ffWU9w2JbaNkmeoiKdajO5EQL59Ha8t/pmrn7W36
RtcDElMOIB2I/amSBZ761C9suvTjFdVsHYTLj5dcTAZXNclO6RLrcrpQZCk5NStaRER/AX9ZZKXO
rh4fZKlElhJp7ZCh5ExqUGZpBfB1lEUWk6S0Qi649/+S6kti1P2/W+xGMwIKmqqh35Mgtg3iMBiZ
wh7pqJXwOm5kjCH8/J97/PycIBaTMsFbng5Ypq1DMlNBkiOia4qB16LRW/eRAIxrPcGWtbR3kiba
RqRxOHZ7Wb/2b8FDSgUm8Z02DwTU9DZuv059y3ZLXnvWJTj+O7EH6ljDTWIo3MOvc4bJEW4u/Se1
UJaFHZa1gnXDeaMYLyTXrwBAFy1HvHQdm3Ln6G3pK9FB7AnsWtVYIUdxx3SmhikxyQsZXOexXYpo
7agQymMg7K95u7oS1W2zgg2ji0L8+Ma4YHhg2xh8NpW4OaRKqyxOCK5jm6ldWf6FqtxHwi/r/l1E
6n509YLc+PHU9UcQVJHXd3/5avfog5lm3gdDp86WwlYsuHREZgeUZUfMxodQQrLZeq3AwZR2zXdS
F2rD264l0pxCYR53FMKM9urqbGHlgLjZxVvLU+kPi3NfBppUIhU1tQYLXpe/5RMuuVJrfl8DnxwE
lLPZBfD7Pki8GL424zNi858KUBv0SQaKYPBQnj73sVGbOh1zeyZbCamNn7eLpNQGqUsjrKBohZW2
yvq3jjmW3WrQmhZpKCcsxQYD5NlYnRunUWiqT+IN4LRyQkKlr7OBDXXReugaD9vNfYSCZoN1YYUc
LkS8yxnHtXsO4I8bL65BdFyO8beslGhPlC1YY8EmAajIQsuaqvNdaL1ELm7g9MBA0yJuopBfz8SL
7p2a9Q165qqFgJ7H5BJDIPuzwybFzXVqd8MLmtdantycviujZutEm62WhXn5Hskz+j6O8HLNrGG5
3GEB3UGEp7kZNM2sef17QEZzhF5nE0u5xvDytNceV6P5CVepepL40KPo0TOEHyqmbHWXpPRLXX9b
Iuof278ZJJ5duntaVfKatfj5h/AH6q0/KTU6Wdpv6lKsZ9sKUEp6Z5D0GgFFAlAdIZi+lAl7NqY5
kts5JSVIwLFc8qlWTpaCIwnt1X5qE4dGBV6G+R8IIAUlndDamAQ98y56qKBkjqHKDyo/vvCafUtd
T5rKGHOcgJtCljwpYFuhOjxcPdFVLR3iDzf9xiP+W63kZw9Fg+C5zZz21o5iz891o7LhgSDUTSqB
9tp2YQs+fCX5/teCuxDhslk2prb7kV8UMLEI6JBnBhy3Q5+jdkFowXtIlmPDbg3O4foPQ1BaHrqK
0ooUe+Z+fBvgnG4Pwof1/H7YM+vfYMxFGUpFQEEZkG0wU7OKnY4Pa0UHDJReYQnBpS1FxbCbYAGY
OAAkPhxl0NfQWFuOZ9G6dfBuXzEdby6A6ehBvWddRKTN09WtejWlwAlGw/2UAN8gto8bY4Q7ASBe
+vDkG09so5Udoi5V+EoRbGwRNBp/SMcJrm7V0g64DEDvDHdf2UwSKup64fUXBZuG5taLZopPJt8X
xFaYC7+BT1t5DQtiBxif40gmsU6iW8mn8CxY2UPLEVzjLUKkgesfSmiVApi7vSvkVXHka/esBwov
DHguTSm9Ip8ron8FZlFBQb2YZrKBdEL9G9QQ9FbiWteqB71aXS8PTDaZzoFcdyW5dNVvYlPpEHZG
Kk0ynUrQQ60Dmbwfeikyb7B0qTSoqDwqIxpTG98YuKGDv2/mIgkfc2SAAYurktfGUBVXxH5bFKUT
40eJlU6/H12AH/lhDVaoroyWPgZdNmby0fu5LfSr1l0bnSqHrpyX/4MgxUuHgEbpFB/0HrOP31Wv
Wrje4ntzIZ3wpHb0c3dDNfy4hwvnuCuWRObJKrw3Ak6fJ+NgnbcEZlUASrd9Aw0cbpX3oHSax6UF
xY7Odkb6rLUZcFGdUVtKklzpIbUuS3GZOZ+ZfXz4dsx1iAyNIF8gnDBDFqLOlRwmD+5PIPIOlei7
7WEZFb66VwEvE+skOlDH+vTHTqpWQXhHx/BzZ/2zIU36HBGBcwRjCAVHjN10iINKifwvYPp6z76J
Ll841HyR+L5hU2Qckar9LUkqxd39Nt8yikyNR33/izbykM2h6q11kpEsGWRtQRhqapnq4EHSANMU
cm1nOYNdSktg1Hq+73gaqXyb2Nnqd/OPPfB4kHHI617D+iL/2kyfe0jpEalaVWOV4yT0G6MuFD1T
RbewZqsCruOzkDVlo83BoIpkaI87SE6CLluqCGErpg8bXaJcpGciJvLu6oBKX93wJ9RfXZW1nV8x
OySfqP2xT1zwNiMgWY43d1gM2KIQf1gQcerEbMC9AOrvjIzThZj8PcCOs3xGhTcsjnq7fteRaNaW
D3+Ko6qKjKnIEbHCQSvCPtLCEwqze5C6GkLIcIu1Hpb5jL9HYGde2gAimAFMIYQiOHZjhl69/5F4
2I2AOCw4QjgZ9a2bIJ/eaX3Mu/JD2V8iu2sugkvC1NfYIDDivtN/d95yj8G+0pHiobvGYWRpmsp3
EeWCRdCHmAxwFzEhFTa8QCSK5O0yWuk4c9rH+ncz12p8zNOxFFwG2uEBBJKF/vloQ3kLHnCZ0hp8
/cBA2iGCbIObvBVQp7zB/VdWHemJMG9xA4n7/8nqngImi0bdEGjxfyBW+Tcqn3aWebdzf8uI7lSO
TKeCE3rnd2HmTfy0GHG5Gpu+95ZjGuMwz9IkTy4SOgzia1Ea4Oi/ERpWTJWiq0iazAXIvdP4I5oU
DseXsfeUTfz+AiZY6BJJE5WRnzBWEK+S0aNkMj4XBzDEIhtppalUf0N10BKNnEgEKk81KyMq0G2X
v+nfyk0h9q1AU93ippFzatQssx1ey9P6iV04St2zxeM6PsGV6ZqZCyFspr0TtUdsMaBTR3qCV1Wk
x1u1+pjeUKaHVj9lCxrswJYExdpnjMc/lFMmE0kDM8aropDEF4p+g3QeBrRS2B/nHvSI4G3jVE69
mycCewgwcWIFasIYhYttZjOUI2UsJFRhJl8ypM5UvABAOwc4BLXWVI5litpImm6fGqd2AgIkyhtd
BC2kJarykeGuPgRthpxKQB4g6q5k9VRRMDzGM/CygbyMt5V3Qq/wZRwUTU8gfcwAzEGb5DehSpwP
uqQUglbBQbIa38zxizYTdnh3nBDMeK6/Zn9XpKNfR7PzMeh0X87CFNBx+IqHT9MKq1PFNrT6VGcz
P7+W4T9kNNefuICnJq36NhbCmS+3TML6Tx0bZB7Q+2xCklZ6soQhShgV0nmbjG4TcBjOQg1s60yy
gB1lteZCnWtuzw7nfRcniVGi3KBROCobFR3DHaOXjndBglPZO+dysmpwkJExli5MGn+rW/eXhz4w
HlM+FkWP1mrB7aI43onhQTMS7L+tpoRfHc9X48Wa4+3hRNLR/2Vnvd/2872GTNixDE9DNm6b4Dxo
GgGXIqjYSb/c4lO16bQb3iERX9EU25tdGvtQQ3E/B8KKIEa4hsqnKvhEx+Zn8ZvXx1vwtjIXu34c
40oCIMD1gyfH4U4suRdFBiYX/OgfVdK/nBFGx55eFO584bZdRH0Bp7kuMfzpF43pNPLtQD8eQPtV
r9xooRApnpcM2MP84kw/0ytnAgPm95ZdgcW/x9f3ENRLExwhftUyJ82kbiaP3EGi+zLN4FYiReOW
7yvTfJV225ghvCqe0OsedRki+o8iuADLCQqmQVkIlgekPbPxDxszQ6EQsdDK+2VxxhDxsJFP1+lf
nu90H8YTCu0ZytnV0fg0KtUxKu7NsVtmkGUDB4epp85/0Igzy8mDt/5Fjdgoggg+3LhGws81uIO7
ivv0idjcgbYKkSFMOnTEmcug6NWd+ABCySIyHMM/HTl7BdJC0DhE44grAvvKfWAk492qbXp2I4dX
o73tEny9/HV9Hdbb2q8pbuYpE9Jrr4f9VJtkYtiIwBGuxvRqpUPGCx50JCUJodjG4d0e7dE7EIh5
YGZQ3qJ1bcDjDlqpOL1oLdT4jnSJ5dBrpTDWiVegWabch1eusG55y4UkyQErWIzmNYoSmf0F/6C+
0ae8kGAnozJjUPtn4Er4HrGanV40ee0M/IltfcF1LIPbBGU6ZAs+qDRE/6ocMq10PfSFq2a1NmmX
6djh8Z/oLiaR1bKLgcP1cXtiYft2ZYGiqmuucAOoQ8sl0jWVxGaGPrAR8Q2eiWzww6cnABfGrN7i
kTdGF1qXI8JVmnCJ6UPomvldShCjR7kAE/wtjwcZtWiNHBI2R2fH+r+bK3PIwkj+F2l2L+IoPUV2
sdzyehsttIIf8s6LL0dju9AiHzzGv7WJc96ezN9sulHeKqyy0Mz3ZsQ3YtYnspgOP/0vDgxV8Lrl
BJ6h2gXKT7A4/GwzKPa5H+Cj8QdKr8wMmUODqhIsXOjsG62zFRt3ATQyrVcbLxBaQIIv1NnsI9tW
ZyIHiJ8CNxuWkn8l01yllORR8BVbRt/R3oVLxTuf+hA27+Wz2iTIIFuXhfoSqxI5zqhtLBZvbFQ5
q/SfoLP+A7iIMlSBDqfZVBYdu35xLAxmkwpWbpo3OjoVNmKcI2y7cZ4LNAqLBhvevHtE1LWkOFPa
KebtZV3EMjitw0TpfAQFkQSm7l31il2MTl/kH4YRDmmV2iUtpRst/DAnZvKvnTrzpaBkfXZm3y5i
UhvAdn+4EBEC6CA2OdxBXNzjKjO5bdQmfxLeQYLlvC/CTqlYDeglqvn7PgJJIlNN8AmTAx6XpnIQ
lAs4sxXdCktBLoEH6RuPodGWb1B+y2FEtfvy4yuem1Dhhj0Wl/H8KqceCrrl46At5dFRQy2H/PL3
48oDb1vhcjOm9JlLYM+JcMuF8OqGRdo+HhxPvFkNbgJ60HyO9wIR0XH+7VI3p7WRjVHdwdIf99AT
Fu7+4cd1BjncqxFb47+Pw+ZT0i85gyKmNTC57A6KZ/LY0H6aYXuv4BuOJMZhtkyS0Ki53O7CwAqq
DnbnkRod72O1d1G79UE8b7TPZORJSQ4MuMrbtl/ZtkfUDtRX2qUmu3yLuDWX0iVE5XwsBIBPGCzo
j2SyoMhM+WRyvK/OGoTrKAOLiF6fySV71kG065WxsBiaPZdRAOvn9wZsywONdxNlBSEaj+Z9olX0
7hL+//eRCfnu7OPlMEKZ4F76lsBlBHh4wHxhv4NCSQPerft/zjdOK+yw9fAl5ck6HQO0vqKavv94
rLYfhMqSxwkNTYVfr4IZE0i/McY85GYPVfOYyee2rfK2AChE8Kk4Fd+2vxVz712X4/yQuyEYBzSI
fqSPxpG4SVaV33uVIrMXrV0pZxZDeYcRZdCLqfsfibOqurl1lqeyx0NYnMvJihue3PNAArgyAHs3
Te7vnE/ELcWUFF3mxrVCIX4PiWSe7nAGYA0jr4x3fy02b+fTe68EwfOO51iZ+HZgyHjz2/3D8IzO
BGb6RsLmk223CNF/YPnd7XsHMY07YU1Ts5XKbNLTy5APF1y+g3gDUBnsg6sqL7Z9duEyI0MCVkGj
BbjABzvaBxjUXRgKMft+WtL/m9UW8LoLxtMSuxf2ZtQ5pPAcwpDBOoFWS/Z8HbQYRDpzB0+dN5gs
eDGZVRNMPO/fBpKTVDBtQ3yXS0vlgAwJ17Wojgny3ZlnwmOXZx1JOKEzvqsAGpXELrd9rGFCzbTZ
cO58BffeUE2YrY61oYeCxqEcJAoQMxthiO3BQkZ4PZcVWtAIO1rj05Uuu1iYnfSHXr6KLdtWhFn9
GpQUmpAnF82xv0SDuyjg394AJc5H2kgs4AwHxz2GmBuEJjymraY9W02MNy/jD78WBr7GNSkn1ujs
EyPTejEIUUWZMoz32V876ebk/+ggHfrRqNmedhhmGNQTgnzdbQKPaSs1sR1ZB6jAbyiA3xqMUVVI
1WjP0tgXtthhvqZEjrRchliF4Q/c4DVJVlfUUtlI1SZUUkTmy6i0G3w6aUCPQrQAKW7sB/qe8cQR
lGIlwCFuRyPz1kzrsJHGm25h87SfIguupK67wlVHEcV7XcSiy3cBjS9mQFx6+v3nc4U/8udG1eaJ
DlLoLkH3WaV3CSvZ21hmjYK2RBKnwz6VoXjjZsxbO7WmhVgdPXom/XtPB5t7dJvj0vCkkbcV3j1y
/Icg8ZssyeSuTExxh86CTldg0zSjrgkHANMEfJnL1EJHEcetkT1lAuOk3n5aQMwCtYvjxWWtZg0D
8Zt5VZqlxeAg7Kbp64ilqd9FmeA5r4W8SOoHEzCD2GxYDzpzofXUYArcv9BjQ1XvbigurPdCEwsu
gJvRKnIF2hAASa4AaC68+muFBGw1RoXOw3OpzJn8Vw9MYzyMGVIFo4LbLVadNKLDXKx/Rctmjenn
ZoWrSYipV7quolJNgVCl4z4Q/W8vYCqqbmH3WiUKdhlsi0ta+LbO3zHr+kxslc+m7T7ziQ9YNCRr
bN8VcykFwvXaAaBu6XdL8rxwCWHuGs+m58OpgQMadFJ1kCePJT/8eNXGdMd7Qjh4Aj4zztVRkUOh
KwqScB3iuIQc6BpAEHEFYnPQ/bQaKqzMBRAydFH5G1FlLLXvP/7xcnFycf4wqTNqdkZdjxZe/dxT
uOm83e68BRaNf0Yo4rTg5oj6+HRdCwDsdhvnN6g2mNDppt0C07cEOFlLVKAyrGLKAcOu51WEqKO3
Jry9H6k8fWkj6GF/HSjZYb1JBHpNuV0qFZREJ7SqUhcGFE3EdLDXFuMkW6AfkYLM4cB4cx2TanWH
TAFmBIxr1sSTgQGRzAF+i/Sg5Z8jhq8bHGE82rDH9XKkLLDELYNSqbzGCDV5LlmL3J9a4xhXHGtZ
8wSUZ8Z90fCd2rt2W071yapObEfGDHVJ3IQ6leeacRUc1f2o/K70kRH0KIRN4PY9GT1HOtqut/1G
U1bo9AcsX01FgUzimJmCS6qjARPrDa+mlrlKe6D/I7rPIaHyTRrfgjmlAf5pGg==
`pragma protect end_protected
