`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
EzhPzTpW0Sdcwks9WUS4y8ddGIKkTL/sFIAreNzS1rhHDE4mNjl+rSnwB+uHs3+7oB7K47vO8QlX
82ghydQzhdhETzowfqAhPTDpIZoaGSolsHifMLvnyBVSmAFvc6/NlpPlKEtsb6X61naQMsdkZRre
E4kU74R1nuDZ27ho9mmbV+RS9u4vSjv9p7L2cuqwoZb1l7ysFPX17qgy2E+9oyb4XxbSFO4C/y1H
Mqs6anRdRhpblqbiYMtb646gtpN4aux/ExT1+9R4u0gs9HU2yKaBKio8rsPdNQW77G/NTIWDbdGc
y7mXkqZM1dl1BFrdTFjEsn+ORLGXlAw00+sJnA==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
pAm4YAMM3+1onp5zWlhF/4CrOjeFAO7CHTh8pm8OkYtUhF7AtzcEyej/RWg1YDSSdEYbzbLbXK6Z
XQIsuOMcMa5v6PQ4yDKIy5FzzSnp5Gr9cAQ4+ZO5QbqriW1zPkRJ79O0EDctJo/ZS02MuwwtNq/c
bxP87NP7rU7SWqXFevo=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
e2RQNMizX6lgvpiNnbbh2+ryPESruse3QHAiEqbJfYJY3yfZ6Xh7vkKrdlF0M8oTVeVxCiGNmvma
6zMPBSqY7L/Bw7b0SVEahPtk2GR31YlSlQwVRmDHn9vth2Is7otCCyVMjDnmxEAhxixnPixbYS78
9xKGqzFOm4YViLUf/iQ=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 21712)
`pragma protect data_block
96xnBguySp6Opf69B7rzW/cgBagYi2BPp/skOu5jDqLXnnZCEMgoItnrXvgLx067rjE0M9iV9qvX
lwSp0hUxhFAjj0LT149s/dbUV+U23j0rzQqT2bhJL0AjpcPbpHutiFNlKceQOtzUjMmyNodER4kN
XQL/IBXs9fRF0/EUGfVX1Uu2j8WHAsRoU5phhVNlcurMIG00GqGIHskNn7aL8w4Q0M8EvXkVechl
2C+02NO7JwBn+gf1BxYD5OZCgcct9y061UOU1FSuI2Mrdm1DdPG9Qastq0uma3RRQ+R7/7AJpcnj
bsP4rXmnYa7GMpQzUJIEP7Tgj7EfofZSiy07XS3E5z1dP6dQWl0HqrBJME5xH5n0PtNg4ZvT4mMW
91HaM2OWj+pLNrfHp+J2Ow8lzTfDVl97GL70UrfE5Xh0h+1+v85nTjbdzEAedGAxKdz6pg8m7yG+
7lN/AbI183B/K26FaTho8cJ35YN79x6uMu1tw2GAM1it5EUilE59/VbuRQgE+WLvWmpC6aQJJ62J
zzNKRd1RECxVFa1CAH1/lpDZprCa+g8/u8T7XIGrb+huDp7l1spZ/esGynF72i2Amhjv4xMCnfpy
HL6OY6m7WJ8pbKxaFRn4ovMA7oWr7Sz4mChrpnfBeapQ2dl0xGCAi3fqodrRaXZ4m1kXiQu8+4zl
JCiinwFq3auMI6tKFV4uIT+vKRq81Loe8bwrA43XDN75KfDZUzICwwFXaU04ONUt7VNZeXU8a6Da
Ep2Fy9oZPMm/jOHBbn53uQdNef2TaeoXNrxinnkFBkor3vOGhckx0zEwRB+CdgocBU+VbwcmFhI4
zOblNgylnOEf3cqATJQAFfpetER2W5EK3msyWZmA5fGX+tNeDRi1OXxFSUXCxKOIyIh6/1Wv5zp/
mIqFEfUSpImn3oIR8EPMA/WzwWuhD9h2OpHsqp6AixQhxj6sEGkpkN3g9Ad2TAGHxDlxUMnXwgc7
ZqdWMfeFSra3opB5R2I2IxxG+dPqYhUcfvvq4GO9LozfppR3XFQ00Ly0N7RkHNwK8U1r79aG//fh
VSc9ARZVP78Z1yUxnXsQ0eZhrciUNoMTttxrW9jHbJeW6Mos6uhf+o2/BS7rwed8hzjZL0xJrS+6
O5YVVuqFW7I7Hu2KjaKKdOvkfTui9QP+Hmc7uxprkLDx/wqWHyALdDDQJSHeGFYmx4cCMZEUtEgl
ZeX0XsDu7RqM6PKD+skZoqtBW7/MINGr9vu0cV7SLz1ESDv+AKzC1wnzmYEKoFYmORWcXPiemGxS
bGTpxdgjB4XZPkGVPmPisek7hpLG8+F36gzI6Q1GZhdOOE/aO/CZwqiMfyHzOCRdoE9lIKrRL02F
TBRRPovBitpiSw8m8d3HQHv8PJ1BcolWDDmNE4PviaieKYxV5kAxih1Dh3DfgUp9U9Dgl0s/tcPn
39vJvUN8ggEP8+zUIidpP4IO+gDWFUd1okX/HsnUqZACMFZLnMzmL6CymyrP+c8g6mjk6BSv6Krg
ZbZS405MXn78KAQkwakEVbChXBvfoAL+FRCjnzzAs938kJcBbJIM88s8Cr/nAWM1GPG2I8PKITEd
QDECyZHEOmYmyDDUTQ1J/Emuai+kbK07xONqMfA8AMwq5GT/gH8aP26SUTybWUabWQEviJOT5bgI
HWq589hhJE2A3zVZD2G/ekNNrEwqNGi+TCObvaiVqmnKZWUo9y4i5IAeQCfAmh8dfzcAn814xtq/
yk8LuDXMu5c1kRQGR2XcG+4JYv6VXhp9pYHHK0L62rBPQrY02IXzUblTK3Q5C9xr6aZ8igjSoRrx
58asI9foaZB4gYh4ZH5FtW6aQ7vu72XcjGRJNiVPAAcuksGGSmJsVitctZTRua2QtwuAHCEzbE7E
NcmgsjXXKt13DD0VXbXf0WwZekNnx4a8x3QuriCI3vyWogIqokgNRmIP0O0zIAoX76kTNWRQ3mWl
YUpFrX64rYfup6RVLtNpkb5Npq5eFgxGU7Gd3R1gqUqwOZpm+Yt8upI+ZaNXUTE7pEuRnSDe8THW
10UkNuEYaeYBRoW07hwy86lC6L1LMQd9cCsn95cH1ZeAL1PNME19pYudgVrFscpYyyHjL5MYYTt2
suVadX7KelxnkJPEaXzPJbo52AcGG7LYSzkkylAxcK+DXyPebi7diNypd2LrRWLvwLJY8n3PthRH
77bGAfNiBVRwuWLwXj1C7AgHYTKfjw1xyk9gFMH1HISmoD76I0w7PE2zRfNeW7xxj1JDuTEoIT03
k589OPREZWx0VVX/6l4+Lh/rS3lqwFAb0a68b+L0SVAGFYH4usbE35Fr+sCsUqTOYnpdYxmAg/F/
gQn8NP0ahThqcaFBBeqKKWrG/T9mDdv0F7qxQcl5DTT9QLnQWhJNFrsp89gHYPaoEG4KxZsIxrHq
xIVF3vggoI/2E+g77Ee0dvm2rDr6V9CwN8cV69BciF8Rgo7hopCnKmeEkG4zw4GYZbAtqayB+ull
hWpqag13pDidpeHon1MaOko86mC65YlhETo5i9m73vKvphfXH5MPblirO8kc8rHQpT94gcMAD+Ez
6e+gSXYPJvSfHTSiuymRUDdbT3YY3Dsz4gfG2hoEf6rSoaZhrGJlnZ1bGQrHPXnEEP3mvalU6D+3
fj1JW6I/XdLCfHuBeb0lW8LoSHtDanl4TOsT1QTswi7oOquknrTMBKS84iVnc/fcIzWD6xuUhyzW
R7IuJMWsPvQ9aTjyUVBo8aoqtMTxjlbervhM14LpKV1z1Z8u6K/1k5ax3aHvHUT+rae4Bids5FAB
RqqIYZNtIXeQHfK16iNvbsh90L5+kdZJcAapun6ibG/c+K+gyiYQw19hPAGNdnbQ8qTafQutsWY8
Fum3K/1GP06b4/N5t51s+l2MiPISV+mA2x3kvA80dF0pTRZK7Fa3NmNqowEURv/2BN0PXgyLw4fr
OsMMJn8Rae6CN+xNF9j/TGLjFWK5+f5GLGOHVJPdijaVzUnNVftQxCo9/iBY4F23pwrN6ekqWr8h
bnBspDwp5y1AqYpQuN/Ho3Prfyd94iq/yneDZMsuJpVJ9/yKIXlmZX07Wyi+OkNhP00BFFoMdeXa
1w5TfH9xceztVyvKQwyqLrvmwyhcfNdikgeqRMEhconSbZZKmph/NGl0UP/yFGT984+WNtz3GYcW
8OLrlt8KSLySDGn0EYFxXOpqbLMEwznCBs1136ogYqPyVd9vepi+VPR6HkDSLv+a0eBfUcIXJ0QP
4vN6QCpZ3LPVQUTPh4GJoLNdZXd4m0rueKoFiiU7ZCARwxDLmDAzqDyDHCxzLA+Xa1gJ+v+GxTPl
1a2IwzcQWZ+xzsclLwuEtNkTEBBzh6qQF0hUcYCSNny3N2KxiNTRVX+NtTUbzOTcCr4kipfof7wB
YdhDDBgrMBZMRsWP3qR3KuOOUT2gpm5xyvGPApDkAe9N0/yIkZJlEGMu0OAl5rgAaWFivit4I3X+
pWabeW4CXnraic+Hs4iwAov7mF0avwxv2gTVGvKlvc3Bpz9PM8mIFK/NiEiT2s9fcjhIaukuRC30
JO6phQ9qUCybANCPiLuy0Hj4ZDe87mzYtU4/ehgWfOSMkYqVOIC8ZQDB+VAHEO3dOK4aVhHcj87S
/VO1Gr4dWBMf9AYRmX7V10yCKJt5hBhaSxHBQWwLfNh8TpvK5k0qiHsaZnoED7QnoPBGFFOvJpOb
quq70ZZbKYPMTa4N7y7s/5xxJssGzUnqJfZrQsD80FuEsKv7QP1VKN13C+h1TDLd8/aozKhHEh7C
p4RqMga0b5p87ld+gnYm5cdpbyMGBdYKjc76FFkCFWsuSGPAm4TBf3kLFIYmMVqw+67TwTULN0g2
Xs/KjjH5IaJIXgXMPSGtehrf1OzvSJvK/vjtPBQhfHL6so0rhtKND7GPe9czuRf1sWZw1yoVLfKI
E7HVReQyMwiJJKveoVgM1RjW2bgkBgmoYHTSBguh2T5n5ZXoonkbdNX+zDiJKFx/2nUUL2BAoYVd
CfTElc/rc9UiVZiIkqsPRib6DazKxdblZt1yjDbxtLulmrNv4IT9QpOGgfU3dCJ6g1F938kgr2r+
awEmxzAxmS0Rp2ZmVhOFJ5fP0wZnwClCxFoVZHPv1zVfP7ZwnEFP4rYSN3WZKtPsHJtRBVXEsnoy
2ahhcp/JG97mkBE2mJp1wORLND235046U1KS+NlavaNJG4jc0I6Kae2xR2eZupcswEjsOZRSdMoy
ryVwA/fJb6HxE9iofpYfbq9LSTqWzL6RIJv/G+M6iD4WjdKGH1r2C594RHq4DYYsDBVnNr+fqTka
+1EZyhgFnehaiYqKyVacnhiJIyRq28x4AB1TAnRuxY41CWdgqR8gvvx8lRUSJFl2WJzYCcnzBrmJ
rXtgFCfiSH+PbfE/HBYkuUyWYPTnYwlbO1CclzhXkZRqLXbwL84XVM2SDiO5FDwEVtAK605gPZ3X
Uw0vYydUw278Z3ezTzl9Z66AE0x8UZ1N+tjFLBZJR2enGr72lDuZPH5xUHodJsGa9eEyNCjtCWJs
thOFH1SMdAAUjLDzi7fkP4kncnT2P03nJVkaUizwIHB2TQpKdwJhgYF1cudfkh5syEyBiSqIDZGR
maCE8S8ByaSB7vtIx/58RyGCUo7B+GDbgRu+JQe1XBuBeA6y2BEpndyW+RD1MLK8sxlAYV7gmroi
i3LdDFd4rMNkLrjK25BotrmE3CHJfJtnVjdLsigi2sH/ERilx04zRY5503UkF0rneia9AA8yxLdV
ZhN0+K/YRezjFZjvXKGPptfP5sibP9wC5g4PmZkZdnhA0tfMF26GrvID+HgEzDpLyuogGmi0H5ZG
iwiHgOpzNCQRTngLyANuSsgejBKL18EbEptkKtXbLFNNSlNWuwpDrgC/xusInXkkE9+MtvXWtH7B
ynudHYGMb41Q5YIxt4TJbDB44IMQ57lAV2eHTp2o6lIDJQoyxrCoFr7k0DmFDUzhh6KhFoHu85C6
oLJpdmj3gwXEzgYUVVPnr+zrv+ZSFi1GBFTo2R2ZrvkTPv1HDNIlMEg+2hrLtKmh6x3/cNEdmz7M
LUIC1XIQB9r3sc2m7ZtLWSAhoGlxOy/rg0ocawY4+Mi8tuUJb/K00N+YF0xyadUlJVMETdOB7BHn
JMu4A1OAf/auGODDcI1ORgPXtw28AAe3R7MA7Egwm+V7/C8a69qzqsOp9UAdPFWI4yOCBh55DQex
egcCocxsO1aYRyy6kENfUVsg5+0pm9O1oWDsNXQLRNbVcagYhEaTPLvJT6ur7x6losxyIO024xKV
jgCSHRLmFgq5chy8TB4xIx040Ty4yLcuGNznphtL2trdDNAfD7ojFgXBZjANk72ZQYaR0duTyFRf
TSvfgfqelNauuXXxIqstwEHuYce53QimxflPEmVaHa9P4KbKgTVI/dTH/GqOSHVq5LuVZ9M6FNxw
PhCeqovYMrIujPE4vJqyH67XSn719pk0SeJJyQ8BRbFciQZ41sFhc4uDJjBQyO5XMBxyGp/IbsII
zXSdV2MB2JqNvHBVXJQVNisY56FH6ZzVHCe/2rzRJoNtoEFY9m1/KqO3L9wowUFM9nD62fnNQE3N
u/y2VTiabhncaUhmHf4FDhzEOrQSuYQUFW32s6x+XY8f7zeD2C8DADsHPnoBtxxnVwqsUyioxkuH
vgr2asldffcb7q1A96OKSleamLBvffg8jog5x0NuebUymdfuWdWYCseV9pFl0ee9x2GxYB1uW5xz
GRpCyr5Vqeib1lQYSwn9RdFp6mUEXOICPXX7qVWz3YbIyf560l+HHtbnqiie/RSvhYgxzAZCHfKX
mDKj+dzHM9BgSZEaZT1RerWtvjwfs/8JSbMD12YNX2GyPVBOG0zmsytUaibrRfEcDE/yRQmQQGMF
V3a66TLI2Szk47Jqck2htY6OGWBtmP08TJt3h8CqH2qaFhtUTkVU2OvfY3vBh8k5CRTwkSgLiqXu
/9XQrQqnZPC89nDuWr2pGztiQPOmC9p7fr8MMIBGtqr7coTzndnsJUNMUVxJZyhEewky23FzcLZp
xHE+5reiQ5/RvpybusuYvcleaIqT2BaOqM186mo8/nTqt2zb13bjAq56vcFjZ6+AG8xj1RKCV4YJ
5hs5rZrgYuQ2XL5YHHdX6LHEUexbu/TvIGMYPUrNO8dXDLpQEGtOPNNK3RPriQVKQabHu0d3arNn
kBrJRPofQ34d6juHm5k8hYzyQuzz6P4KV2We44c4e9UCzzpkdJfX5YZHi54pWxrkQtWQdOXzI+1A
00vd/bAYAYNA+qyaa4a1vjTEPBZ58JDs4zkxGy31Rrhcz2g2KgZcWX/izOsVilV2NRXkkfw7ns89
De9pYhwIpmQf73kQsWmIG/y27cWYal0sNqzQvg24GcgMbAd/8yjnajfc2x8gs21ev1KVnEZeAiJm
P00bjuBTomxKvQFAyLMPs9SCM5eGstzG7UHAkDpNIy0i5z5y/tXGzFtFqIHdu4ibFLaGHrx7Q0Lm
0SM9cksHV/GNjDwS8Yt4m19tBmiwZE5PAARd8I4JuMnzMHHXiAin7019oBOjYGR2LAdfYgOG27VN
FDNmK5lTB+klbB6C4llB5Lzg3xPicGgnsUuHOi7+pqPlJFaLfebuqry4EwBdDUSxkhbV4hj4O4w4
t/xxX3PW87S6xEo4DbyTEeLfFTgvQK21cTIqKFB3kBsczl2CCrhmnx/q8KESClVCQRfqJwQZfGmz
8PHcTHu7pfnDZwm+d0tSWhtdRhurEltl2aVeuO58S9mchIIb0+Tug4jblA7yWNKDcv2a35gvTgtr
vqEoZa/KhiGTv0MlN9Gp0BzCgW6ZouuUFxv3af2hEYAJCqK2oZhIdYpD3LFXm2U3qy7srDDzzjir
6hdM7A4+Mc3FJ6kUv9p9/D/iJjfpVmEfy7SaFSPYLqp4rSHUTVMCs2mcaVly9Eb5nAU5X2oGRwO9
FTRds8tMljpSgqy4cqi/DEGtMFNhjR0fRS/f8AxJ8aGLb2S8GhvcKwgkuMQfPTMcWNVkQIvHF2xJ
MLljHoNpUvF1RYb2zUQjsA8WaxlG8aZPrgIdGzLOFED+MnN/S6Zg4diOayVvC7y/QbbvM0NIZxpL
0lJFZRLGOSYykLGuPBpLJecejaxRdkMNOFu0MNSn/eZEKKYgyeO1Ttwxyjk/xL54Ttsoub1f2+eI
bE3kj4raV5JmAb1ikRNT5Es0WVhXnFielieDkY9oLFVTxytDylwUFixrmtyFWe98E+lz8JSXb05/
EMt0pLejSF0bOi7Qa1waiTgmUgH311ofj155dSzMF8y7mFaLyaQytDps0X8QI7w+i2lOsq36dDlJ
Vu72MHLVigfKTXAHVBusN1Q/PF/Xt82UUYPNktspqFTg6ZtDiLrEb1AK3lzmZs5tHzTKjt+qDxyj
MsyofhxTGm2erC6ZShIzWpDpau3vgLTN0TwDRHL+XaYpNHYenomoqEg/ysuWauPoUNuLRl1bsqvK
3o2LqYhz8iZlpmImbdtBSIN8P/2GWsiato94mnSmvdyDx2VO/KMxO2Kvz4tixXZzAK2yqt/sOFfS
2YMJz9pTL4uwGjUp8VMMlyxDhJBwuPJ8dF+gvgl8YmuTmEMMCVL0ZVOAZp/kIkojYpm/6kXxGwAI
r0wVWzvijq65dDi3s/xExV78bL8f13XAVQpE0DJFqGo/uoM4IhX8jM4/qMmrp2CxAlsHDvjJJwke
Sm3dZeHNUKPxJljxQ1sfOgc6xk1SNKbvPcxYCxSuuhBHxgnFZ44U0PBDZ1vig59rDS1sxg05+JWE
PCjPIA1qEDa8RI7r6GrhrYVmpHXbLsQaczn+GGtorijIT1M6ywE46/LS7CXpRNLKN/jFbijrlYJM
grJnnbfFW7tzPUPgV0bWAOP+/ZnRQg1LFdBTDUdvl1jXRcRzacD+rLV1BQcUnXp+f1yx6rYpTjSF
BAh0/5hVgap3LrGwVPZBpcVvFYcsVBCgolJpna0CyILVjlBUsOmiqMyuq2gxWyNvYfyqu+9PxQ86
vCCb6q2zEsbbnN9EJA3A4lD2fiDDwpMcPyQvCb5OJtq7TvwZPkl/A0ASRHEXqs8WemeAVSWmFk4f
mLo2SAEMh7DUkPSSwpXJuZylBmJZh0FW4YX0PT42KGq/+UbgphLPE5LFXHS4teJz1vOO3ZeHJxes
X7EOA4Xx9wRT+wPj4esucXNpaHyY2rt5zzk/qDbEKn9xtclyhxCGY+Z+xNjHsPc+/kRe4KdNS54M
7ddQrJuUahxRhfJVk3AM9klrj17qt8/CznRaBJDnB/tjB7OUubFw4CxbjRaVuvhNIxNNtmTHCzPf
7j/p/Q6uM7O7U+hT+fkiCoRTOKL71QKNtatxZ0CwubMgHCUR1kHAmDPqLGq6s52pGH/DUNDxIqkv
L0nTULUT0628piNYbo+lmVgs90K0QRezTakwlM9GE/8+l6MivT0dooZwXEK/98DqozixOnOGhdQr
QHibVZTorT4gOmTfLIhH8n8P+brEAPAbRSMezwu3cI4PHrrKnnecaugQqcZJ8sNVM2hsIbppImsY
H0Ca0TKV8IJODRwuy4vehKY+iS3Moxrd32y+tXAfXnEqRJGLT1NoKgHh9DNeHCr63VxcFn/oU8qt
zEVuUQu1jQvHPtFgJ3sXn4+53TQSr9F2BijaejRfm8LFn5apCOzPVF9eYeXyuf1kWd7OCPy1xAjn
18T4WVaIpdVEMxKiB2aqzqgU8FN+ejz34KYQI/t2B02BgnRmcxbF52YT3CtU7ZV3jtx7kboqBs5q
Fw7B//pAg+PNQgRNTEAcPvbr3o/0prY4q1QjheHxotliJFEhMpa16JuA+l010gzRKFa46hgEB1t2
oAZ+QvO1OFqGO+EQ+k23yKWf6W7dKCw7jwHtl1FH+JgitomW46tPFCbN0cvRndJT0ONMvhbzNPIL
nSqEE5nr3kfJckUTF0WyRXcqdB6GVNk0wWIGzXU/GBzdnqT2O+l3Xfczo34AJPtHFTEXqhG1YzPa
bhunS0/fM+CUwdChdPQOl15klWLZOXLqR85EfpK3vgx1tgrU21Vt2zIlqspFfbXVlKHWBFL4dtTB
zjyZcwEBMxTbrpTB9jb3CmFzILdpqnarqdnD/kjEc5vjRCR2lFr0M0URZw0IXDs2gwoVLYZ+aX1K
ZEnQ/z26zJGA78iWq0+28/sF1pgIzR0ukYDWMA0krpBUQSOkNbd0i9GTyQxe5ZhMQ0htnKAPw70U
IECSmxZrbi/8uh8EMVEItgDAAjPZj6rxT5Qx+lqnF1QG/1otAt9MhF4oXfdvqCgfHbHE6DxJrdZT
++nJoxb7CJW45e0cExE9+BoAKsqIUZMZRPCPs6VPvnSMTahIkO0V0L3i6cnXxUPXPNfnGGwGoCst
rf4KJFvv91r7gxDquC2h9agBRxLbRGr+dz0FemuO7RuWZUfCBAwNjaAYi1PBz9XC2sCABMJNXaLt
LOMiiZQjgpsoYJkX/+4ICzWztMYc0PmoyXjA3hFc2Y0EoMb8IX1pdLTocJPqw3wxpy2gnp5p4cmt
XbC8u8fZkhMMXyUQAEGjhUpSB3G1S9Gbk6uNY61uMDw0ODQx/NFtuCSViek+qZ4P34oMZkYhihDK
1CpL7giT8dLm7hi9Tx/a9jjw7V974qQ/g9777+uct2siPMp5h3aV+jEVloVmOCGAcwyDAMii+b9f
YJ4h6VA+10jMoOqLBt2ybP9RbQiimMr16+mcAJ+0S16Bk87BqHyFI/rPrd5w22UP+YvozZaj9wJh
bOZL/bGcFWar3/r2tYxCep14pgV6PfcimSoRSJ6PqbESXI/VMqxpx3Z/njAG7zDtNacY5dV8i1jG
UgcxIh2Wzd2ItJRbZHxXZYXqoGPHCIihpET7rt/gXXNnvdETu4hj/rXp76ICGWsz8SBNiDVVEYMB
63Gb9giS7BNhb6IPm1uysfk7BS1Lvjof8dN0aI7zVU1Jew/NSXBix497PL3o6+UOhzcwUQRqO11D
iwTXJ3ttmLjtwsSOp0/Rj/3KzS6egtlu8w/V34bptHVrGaRuCsaC3FY9sxLPxrjBsnRUqCyJM3BY
Uv/SegD8I0pLWW5qoohHiOQKWC6n4sQf4HXDh07lpYfgXa6C8ErmA+dZ3nA7BstfBHp2rhQW1UkQ
s54LDmVvdyPmxk3knD0nyQeQuh/2usYZ6PM0iBfAknSfEDtjJTDFXEKcdvlnRam6AbdE8/cXF4HY
mPvE0qpetoTqrD9ymSY2bvWqQz6Afas8QPt44bX2pivXulyGMctM/eeFpA93gV58lTpItDTJyTGr
pdXjcX4hAKTby7iyw+rujPD60evoCvr+iT0/HdpJK5Q6NmkxEsLnkBzgaWrzgUqJZDNMkKeKrQ2c
q8DSSdw6oJoMMUDZdIJrJIN+s2mbMgc0eWV5cogJuXCxc18D8TWz1TnaxhYc6fdffUq5B1gagY2u
lMdEQC1Q4uP4p/WapZN5GPcONtbuzvCPLmD0868Bqvo9RjgMMVjA4rfYVRUPkNdosqw5/Pp0t1ZX
3WEsJzsVxcTCOgbqjN4ajxCDQ/zTFGrmJJWt3BaswwS4OiTxZT5Kfhc/chaCwd00T0UoZH/Kc0al
Gey9XIwP07csyZgKS6mIOAfCX6htONMuyI1WaNEmCWFCpLHkIA3amGgIR6usCL4L8Qk6iB1z7n24
itKB9CeA/4WbSRn/AvELcKpr4PJbzWTeUEQ6qjUawmT5Da0r/GiexmDYQE2jhbnB1dSxIQwHkS40
wQkXPBW0n8lmdt0VfZ63uVNQWNcBTEK4a+hur9W6gSanHacrDyKJvA+Up7m4WckjrQT5yF1RDn7w
yffllCeC/8sb5HauCFaf26r4uzak2ILyRg8VbqlX+23lxKy3L1JFeQFip4fh0xEFpfzooCjvDiqO
nDTs9imfLbG2W8bR3DVlsYt4Dx3S58l3csD+IAmkvC5ZiwwZ+LnUFcLRsvqAKWX4ou3J0f+OYYFp
7WXOCTW6ETdAAD/v556MDltbCrOhqxqxOyizsxAWkrfJhBa1/7tK3rMdxPsJRD97Tpr9M+H5DCEp
oqK8dHfQFYlZA1JEbJ3DMnj8PFnQk5+3eNr+txokqmDPH38r5TtI9NkBL+JDnh7LJ5ZVMUAOr6Yh
QAFsRetWcVVQ98HZ6/hW8VJtGVdcX0eHGEczD4uXGD6vnNK0fxCAtYnuLAztJN/WUINL+KB0n89G
mj7IJc2SbFPnA3UK8sZaY3HZsLcnhAOlfedrymDXQFbPRDjUVN0HJ+c1Gu9gJnZY/mbggwsGwfTw
xOg2+cEI7jD8zS4vb30XDOxCfy/mY7H9PQELrPkBbgckOhfUP7qVPKZejJ9bugjstKOekZSbY2FK
Cj7k/4EAHceN5CYOdT0qok6ipWKiXjaxsPFuyJYKI+m4NBPOEqhBR7IUp7+h8IPwKVORNQwBk8IU
isRXRTgaulGJrGdl98cP4IKFhqbtmOatoE2XBjaZisq7kG6odlGnKNX5b09R2Ry3pg9vaJZdzywN
6c78PibUZavvd5yRNzLFP7sQk6X+TKTarYOtKZ1J5lgB2ip6PPc/KjAJ9/ownGWiAdo9IBFw6maq
LzMnMuywCSCsiCzP/vlRk6vxLtF/0HZS8hBTn6ZWh7auVsQjVMiM2LJBfPfB65TjTvSxHf+hILdQ
/lAe1K8IXq21Ymf98soxmcGEqNbCl9D+owIi7D4i9SuS4STT5nh05FcTppMU9ahFcKrKH1iIeF4w
HSeZLDDy1gVZ4JcuyTKA3/GraVzPOsKrxR+6BOTzioHdNce7wRGwqaTZbZceAe8YCt3VWlvHZONI
PMx6gQtf1t5TVtoN0bt4vBUWKb3xuH0xLSFzjjEGc0ZkLEpnjYU6vDeOxf1VDU5rSKpuYpIsbREj
HMsBMLS19bvR8U9oj0B/lTcLhxTAOsSPOjKDMH9IBNYa+R8GWkcbXyGvTyW2nlUVLNndSbiIDnQo
m16kSSW8kMq30pSvWpl4Y6XKiGrAlephabfF0+qvCeesdXV4iHgCJUVhNdWlj0ekh2On90AlVbXe
W3fhTcGsfQzjfCzLbJEGwhrD81ETSTa0zcLe9+XEOVhMNGzJJs77h7E1nOKGp0W2m2j4idUd+MgU
BpIlvQrIMXqDCncBrbInlHkhDaIg1DakyIGIQ0HVorVFq7Zgz/+dZcNl2+MF/3LkMxxZJvLp5BUJ
ayzwJxuxuEs0YtgQePOsS0n27xgyeWQnaxlFeQbMvnK+Q5212JOxysCkbaZ0etGsusyOJNRzirl5
dA42ygmrboOdZZv1RPuB+7iv2iSyDD8xqwg5zMw827nEAPZFSWteBXE0Nu704y2BNWBronTjYocx
RF5wH9LML9agiMeSCFNeSestZc6Lx9L+kJgw1Dg1+mS236VA+BIz8y3jUfHs0SC/BcbhipwUKHAg
6pPx+YbQtzZz9s9jkZkJLGvNnmVwsVVnXDvvZGk3M4R54KqDStHQlwi38w0bL8Yth5cF5DmyT3Se
Sv+zMtUBJYriXg1QmnXHTfbhmnIyM74cad5kq00XU3M9by3as4rG6R5/EkeWpKrKbB0pM/pkQU8s
fv4J+H7CN2EibUoQxFp+ahhwGnxhiZnxN1WiGVBx9wTtSxB6VOX6VGPHWgyC8myiXWVjy0uahQPU
+2Tq6ybHpjVjheFhOtkO6V7byU34BEDgpggddtFMpXvKgjNQ3ez2vu2BzzSCwXpoeLm+oGMS6oUA
mUmwvpYZpD26lNJMpTeW3s5dCSq324fHJrnqVWL/qyOqnXSAvqw4tFYRIpu0Z3p4tI74bX2/gFdn
aKoEHfINqbOmAdwTnfIJ3YOCt9DE23kIKA+XTkUt3cDgIVLakCnK1EwT6BEoDqtS/iPnKnLkUrET
nY7/qpIiYqEV1/SFCYcYy6+vF/ismv5roA+iG9MAgObyqZSt7fQF4yFAgV2tPqEKKGXXdLHcG3Ws
I4y33wcSbcX+xLDeL9/3//yh/tpEiP/IjQsb0dDK1H8lpaPe2oA5Gz1SJOo/Q06dg5Yjy97wBmrG
L8GiSctwoyX399qZzFGmQBoH13NIoZc1fkFMh6cZAn9n0Q6MVps1bwsP2RS2Ob/wDdXA1WDuGbwG
UCs43uWq3gfo8yQPh/nygNSTUI1DXf6lzNuhI5fkqhDVmlFMwa1r3tppZrDTKF0hqEGAw8Z0qUG8
hstDyvisWVNqcm98s1GTtodO6+VsLRk1Oak/q0umhik5NGRlKaPC8MJrCvYTLjfQ8+CZ2KUqL/Ge
4fIEQqDU/s2yl/21HecbHkgh6bS3dIRde6JNlMlMEh5pvirKP33aD8ix1rV4PLxqmE+/0AMqyocQ
i0zFVtiTOxgmV42n9DcakbAmEW1MWEL26Hp7fxebFTifuq3YZ96rUEZ4ejzMog2cjRskkp/b8GvA
q22XKDCV8QaX/i5ZA9G0ubSFgbtcg21KhPIOoESo7PdOQfkFAZI0tC/oMf4WCtx5Agxp0H/hcHbX
KL65gy6WIoNEy/VDu1Qk6mfWFSt/7j9GfABjjwAeJrqaSuyt1o5olG8prkWYdZQGkfDKa+cgUwDT
4gnzBvSQSAeYmZChpbewbhb+mslPcqPytcNSylRVhWxoXThOPfu7Xenfn4SRtpUVfV0owINgt2yP
hU7rK6sFx7AV6W8FWDnk/4/hqhR4Gvd2S7WUzPHik0LvBROkpcVXogI08ZWrM4/uvSYp4D9X2Q0Q
DVXqi5X4gPuzXXmbWMy/fmBRH/dmwZM1gW4zZypumcDu9767rzfNBHCsDBG4YilTZ8KHTuyO8Bfz
fvTygvtuJ4feH2zsT06mF770Dv2DNUyzcnJ+1Sb/7uG286/kD6GpW1l6jHXVjL5/GYDSFQv7VdHg
UWCLy753prIxESw4AEGAuxZecg1JX46FubtBeY17qlzsKS3+CSQ11vUPKw3t0nIJoqheKSQ5Gvvk
q5RXrnWc0bi77rB/17RfEFzwDd74XxXulQswcIzIstnRvMloeUfxKcYQgep8Vn6JHx9/DoR/nKcE
bwLrz9O0100a9bE+sTpGvrnnDwTl7I84zo4PT6gJvm9Q31pCPnFOi67vwDomJsGSN2t/Kl5SxYBD
jcZdGI+yy4t4ml5ZUVjc3WvD9BF1djQZkkE6lDRooTbC8VlmvsHQd6jhOZmGQYGXzrDmrVO1knzf
BxLW4xITUybUQksWcHqu0E15QT0fM/7DvLb9SFlE9GC86e+SHSGcRx3DtHzH22bt3hFKLtd7+bHi
LBhVOypgJ1D6OxjeDHOC4zmc5D9/RlRfGa6zcpnKCDk9rZJjuFEZM75BlQCviks3lPrBEx4KmILn
rOtr8MZyx/Ebp0gQ/a7lC/xg/eM2kHefoyl8d6IfAox+Amv3fRnGtzQXite1fhBoyQFmMWdikWBO
OI+D/NdNG8pfCIp3FdrnAJFTgj638PTDqT/gViVVUGpJHNrZ8QJxNjwGC4c70kgN/s0fH/uO7WkL
aFGlQ0MybvZRIrLsXerkQrN1Z0MObXemwkS2jsjBw3/kU7e9fCYzuyv+MaevzhDa6qlkHzes7Mvu
teHX5F5PrJtoqR0Xqi7xkD0XwfQMO/BiNd1IZhoqN4Dj5fjvemCTLLqUcaHE+ct8P43CEI1KrfkC
RDfherETZhQJW2o4CxUtPzkoMvJOMtjmb3cczjAMTMvTC+pl3F34pZ3VlgJksJXqQ+kSHGxKUiGR
7ErOW+znfNn2WZQuvVKsL0meyInQHr3Gom6jjnfZN2JH07lrKQwK2LPw2brwVycxKHbohmn20Qj8
QRWi7pbxfB4kwLyd3BXw0PVsWjCYH+qm5g+2VKPjJYwuiKkZLp1YTH6cJhg3BwmPNXjqayY1L7g+
Y1QsxUq6FYNt+pyPLEo+JDC22Lb11RWReVnM5wutWiltwODleqRhpey7jozCHPi5VkRpeVNyrpEu
arEJkd2do5VbJWurS+i3HteEND7GxRewYC/B2JpL/RFgyqBlR8YUlqn1cyI5Eq2yFcS5lOWUhoku
OVk8sLnISqVWo2ITWIetB67fu9oNHB7lcf4+nJyzRgUpsYwY0v53LN5OUU9VLwbQPYRFAihhKNDA
uEGnmpfdAU6WN1xYv3aBFm/dCxN9T9NuurFWmZdv07FhDHZ1lpIqBh15SHZ01ctj/7WYXD/9AQV+
kQ6Eh3SqmjwbDndQOF552lrxlM8Uc2QoYCJX6CQBp/9anmnqKSmlvfAXN/MfNLZpW1sWeGOwVwsX
NiLZG52AzlIhb8TgRY2UyQixIIkNMM1vtzs9ZEQKm11073kxdNbhz3POUMWodup9I559a/56Ra4t
6LMNL9+5jJq32GApafxzLGD31vopd4DyCifbWLQIx3GsQDjToLFcnHWo7gFtPI3HiO9vYUU9DhDi
zLp7SVJQtxwqm96hUgpmRnvKmdeI27oj+aextDjDUXg7hieOVNT1EafKBKSOzvEKOV3dYs1iXnzo
8DfOR6pxxU3KonXLCvJRBTA6xnvJZHydHklCPUAwHhwJclyJRXWTMnIQqTeM21inZk6uh+Rvtcja
T5RrKktFdUf4sGuhIzO/xqXuw5qY8DDMb1qZpP5q6TjjRJYf6uobqqTeu7CTSeBelO73SfJBHvIX
+PItVDMT7WsrWab/rK7CKFw++/2frUU9+UkzW33Myx22tBFwlmZDSKQNxlxrwT+aFfOugRWh65jI
pgQR7/pfsTEYcl/0si7eZbO3m5KHZACoz8ptbGjZdtW9ih8AfOyKuu2dRcaIequmoPCpMZso5iZK
mzC008Z4smSrOTOCfbdrkhyGm7imWwKbiTj176ZTvdDzstkKEJjHts2QrpPJ9uyHrWH/4HYawYcR
9vysE7YobQhCvNGk8DMSxt043wx72Ivm070dTICQn1MH4cdQzOWXvOUVM9idx8oKZzVusTj0Scac
FoLl5L0PviZeZHB1Kq6mPeA0ABYQFOEzvRs9Jo5kpBVEcCHUSps7DRzmhP6kVeQTIWcYVrWuEdfR
YRKDWrWHA6UyumDn01///1ViYoIjCGTmYYkptssl/MmWQBMPLEDav6d9XIs/w1JzYIYw+cyDe6cP
eR9OTKqnh+PNSHQt8ppqelUjvoyCHru/eNWC1p8zdyJQO7QSokw7/osoZt39JW/Kapnrq+yBaCHY
wpR2QRheMA+nZSXkuYwAWNswg4TY0khQ7vBjzJNAaLvMZV/dUzVdBANaUtxhE2WkGyzOsHMgm+h4
f5hG9DTTnBil28sFhILtRWOcw8BAV2yUomcQ0YSMgp2Or/Vk0nGrXNqyWAk6Ivh8e+pOw8oCisU/
j8r34s+F+pxf2+TXhC36zVlrUTJUHOaZ6dLotH5OftrOrTsF/sbwXPDzr9UdrAR5CaixpVlg4aIu
t5pHkTH21RV7fKED3x/S+QZL9sviO87xD3QDx0S9unaJAiLCwSqhU36dHkuXfeZPaf/dBRtTY923
zkmKCY/oJ1CsBLnTvHXynsWXDs0DnzqnckqhPOKyf8KRglBcjTq6ye8LLjBUsr8g5fJifY9k9CCx
FOt1xPeN3+yukqnoyZBzGc6kLMrEMElkmxMUqt/YsdG/4DLiWe1GQrjBq4tBCIrQNu+dFn73iAZJ
zdeohI+WmLWc5WNnTPcaahTpbH64bR4Vf0CdUoR955YSh6uAH1eRmcGwVqYvkth4veW0JZPNWZFR
H3B+/qn4WQufXZ4m+KQOJD8bfw7aC8x1GzYvpZYidcrrzEQmXXk/drFnkr0vEsjSlLN9V6saxCMB
E9x2Gs1oNGZYHkzvhNaIQ6gAAWoXvzL7WSZdvXjMIoi/51vca9Lh4rJRhwKkjfE7AhRgtVoAcuCO
v89dH8x8w4/q5C8zZeyYgA0GsrK3c88lpNjEyKE7mjsIpf776Z8EeyhfCq4/Fo+cXzvw0CVDWfsa
ADWUV6eBNjXqCPC8gUK2/NFH54PYI7yxXBcxk/qxos+HZ6i/r3vQzHOR9zkB5h2yXLq8szqtGxZM
eOJcN1DMXWIEFEy137XjaICLkviKCNvjzenskuOf/apxD+MNzDCncrxKP6JN05gXNHznlwM3bDzJ
w6W64a1IErJQtrwpxHWhjvOsIZTQLB/dzZVoVli24SG5PWE55sL2LHkogSuhaj6M0Dg0I/SkC3Mn
+qVkScw7LGQKkd8nM6/1yH7RTlg3iMiw/ZrNYPKzK/0BfTQjjTvASxwza5J5yWi+iqNcXOvGdQ25
XjI3MCJYyHTSFNVaY2Tp2HOve27POlEhmNJuRhfV0fjLeo7Vap8A8fGDKXYy3n0M2SBEir6cJwaY
5lKtsGP5E1mBGm2/QyUXg/p3LQW+xkzoYDJLQSQMRz4FVPuugcr0QhiqBmYcep0trZc5ysWKG+u6
x7Mx+J/SypnukP1ZBKC9errWvINl3p5zREkCfQxyMk1LYq3/TnGrOS+WOexm62rWsH2l7eNHjHf6
fq4a+tleXIVIQkI4FcvUJoTYnAM2tP8LybTAilHxReV8eJRfbEfLM7gcNiTSbKHcPuQMfliEPkOl
8H+ChZlGcQ9cOgs9/eGlHAmkhuyFObQKJGkEj8Cn1A/PMibM3R2fmiOdxo1J7W3eJnUQkdy+VU9P
yeI0DFK94ZJH7fbK7i4npz0kQdI26DEKztj4AcAJzJI+18XKXrvjd/6hTBJRVoorHq1Nft4MQb6m
iZW0U8B/2VqIGcKfGvSF2n4Or2T3qljy/sIFYH9loQtu9afiuODDjB5dOvBdZAEwAnbbMrqNHhh0
0ok7NG/WlVESILJB/eidJUE1F9uCSd7vw4LMOydcG6a5AnyddfdllLnuGFJqED79T4zel6sCipCb
UrkslT0UEYarYMDdLgvO8r7SMN7jAMluDtLY4mTyjARkgC9dRoO2CCE1ktVWVzfZCvPjuRUZh6l+
sjq9tMrLHaPjZO4Ht+7srOYqsDd05GVYWqRMWnK+ZlBS2gOpTqCG8Y5ksnGnDDIzIc3Zminoy550
5Hy6kOVBnAMpZdgbYq5mqOrPth0V7tjhGnwk4Wn94CIK9+OU0gKfyAIEqQ0CLTDqszF3bFmEDLNH
dPBh/3eHfu/GbMDDk8WkqW9OuL4qk/hJVxTdy42mTaTE9RmhLdf27R1KKDzY8ldjtxKfO3unHadj
4HoTZ/mc7gqiX6GUmUgWxW/2TrjhW7OlsWz9q4KWjDWHpsMnsWqA1o43fg+4DUo2YCywmjp9kuZh
YZYZW7uTr3brqE1UOE3ochyWI6Mb0vnYy4QzUJ+RAOmv13wQYIn/ZVuLECG7G//zQCHfY++K9u3J
KVrVUta+scygdR95xwFB8ZvSqeSd++VNmNpMP/aapA1KRJQfX5BBmzKRx1cbXPRj4m24jviaMHyb
RsowJ2jOgupn1z1jQ+FihO8hJJEOdHyE9fkdiONRl6F6Xek99zCQ30Uyzx6v8ScEFs1ipjinuyAa
jULEEnENL7FsQTQphgNVOVhcQjTqE6RY8I9YbQBwoSq0untC4Vq+P5oU1YxCwIH6UH0jHq85ubY1
8heg/er2QsKhJbHI/Fi/7CDDuZhhXPJqkR95ZMBOh7cyOj/vMA6qpDJPQqgzJpdmjX6c/CuDBZVx
vDEmje78x8Q5JxruLlu3sU9qOKylIaMy1TuQdLsYrV14JyM6aJp0RJ/DVDF5T7XkuTSu2bgpJagH
TDDdi/vI9EJbDs2iz16lKyH8ROZ+NYVEnqzYkkJst00PIpaistqtsuQPnSrI+dUKr/m7pXRYweEv
MZauYZ2D60DmsN5Pn9zc0AfgeMWBuLg7QIkY33bxtfHUxgik2wER+6akaDWxy10MkuO75YwBwDvp
ubz2lrMQbGqcRW5pYL3iHGmtGmGUy42fPERUzrBTJ/PtsZD33686cAE5XDnqawr/Us9NripYPxZo
KjF3qAh13KfExHtktwE195gs2O5OfHATfupCg3LHq3tk122bMMSwNotXWcqJu0BmLm3xpFPwQ0jH
vihFft1+Q95dOLRsoxas+y6JpqMb19nXnxxffHeYnq1IMvjHQCp6bpE2N1bDPJs+WaiTqkBUYChv
JlFX7SB6NwTwQzTilGriidU7wap/d4SNR1PzSddKmIdt4nPwuh5vrr20CoQtRcs4HUTLdfChpRRb
nOxLYDFYc/aQYcwd8s0PcdXSozRRQpfZmpbUuPqrusBUj9CXeKZ2DJRDCFUXwNOf6EuydDQejKg0
c3GOABsPcl575rfhUtkgLv5eI+CY51a3BrgtX7SHepN5ssW6VBbyBbJQgj/Bb/fiEC/biwIdtFlm
3BvfrcvSJa9qfTxXDK8HfJUAEQrsnERLly9nZdsb4aGXCvlpJlZlQG+nGfnt+RYMGyFCUrFxsNua
6VF1s9JgvWbOITBzIncDsSXeMTyGoR/DJhyFGWQ161p9h9P5E7PXgsvGlQ+Ui0mLXLQxM3LsQaQC
XkfmqaD15StEFDJ9PVSygEyZufMU9UfTL3/sk7CJ/O5/4DsEZ6aXzdd3XGqXEoE6lgAdCGilHI0e
6GwtJQBittceLXSMxKB6Phd+y7cSuCMY5PRAbyUuvzhNkxRi+RQhFuGJo8UrHhcDjgvWZjxN8A8b
zqoP6Kn2q1Lfigzqt34cE4+qxiTNn8hFujs5OKeG7IYnRKdcQJ7R1yttDd5x4tJdt5zDZgtc9CX1
8N8dTq8b+Ha88/TBSvWDmYVhtyJVJGLvoHkXkGVN3UrfsKvde/s2iTVXAQYgRHr+Z/Qh99b3Y+t8
q7Ns38j0rgPEDC2sal8AUi+1VPyr2aGTHRHj80IXBqvYL+B/pqSL2KH4wW9clARQBM605JA8oCPX
mX8pZVL1x5PGiJka/rDhGfdDezkHQS7BiWxIawvJ1TI6YN2FRCvR+WOeKDJBxG9mnMwJu2h+8Dj4
RCj5XzRASg3mzn/6oNW/TnSuHIWTTKrxb/enkbVe14o5mEiNbR02N8sL7euCO8mGiQjT21f/UV9I
qyI+6k4KHvAzzWuTKP6i/gajl//33s/RazLgOXBDzBNsf/YFHGDd8/2fk4VdG1g9ojuc2CV6gJQT
Ei4hhzZTgszv3T5/MsSANuUs3cuJ/QBueQ9wKlUsWZ1D3ZKuB7g4sVDLAMMvd+UU4zoMSqKiLpQ0
3Rq+kwZaVcoezplHMx49s2yoQomKEBCi/KhFS5f6/We8CTTZh/khsj7S72Q6a5Y/2CBW8oZXUVj5
7XyGsPya28pl4yHxeDg569pgnG8m/ZuEQSj1mfB9PfopWlxjVECQYI8BFo3VBVnP7u6Ut/pQyFRd
2zMaewJMxw3d5+Hgss7S+A2TdwxHVBtFRAoDSlVSsOMHUGbpLWCnXJ6WoFmAw+H07uai/L5FnXVe
X2262Z8+aXtkQ0gwlq/FZQN4BF2P87aEJXeFlXPl8P16kAXsHy5/ZAknpa8VtNvOoar3bGATZ7qM
ZBAI9r4CcNZTWZRm3A9kvEe+hmNWME1/xuw/sgZCEAmO0/gfqnGM11o5iLpwBOkEp/yG87+lAd6t
A/CkzX0MoWGAsinesLF1JNHRwKqwVmPohmLQX9cnjFHTqCC1cjQG6Q6kMGJxKRvFNhONpZn7jy1S
oJt+ZAXpDvmmXRqYiKPkrSCpzmY60To30GCb0Y+vgSmMep3HTawZYTtbcODhfZdDNlahwYedl+iT
ScvB7xkSqTwMoCtbNV+dMtCgRAvpzUo0u1vwJdO5l9nlK9Be2POwvT+uzYUltFpacuIqQvoCWcem
dZQHTPtAGFYlXHZ1QWa82wCNXzf8UgmG/dmPcA/NxQQZjvIad5wzFuNCmkYmcpDJktzFBSh9VBYV
3M49bqOHIuJ7sBuT6eoniMucudUUw5V+S5gMMdBe1LURObboLKS8++QEzTGfnaGzmHwjwKJ/KiES
uf1SLBfFEfUSW1eI9X27JavimRgp9WipoEfcPyumgRhVxYZKcx2x7vDzn6YmxUzaMg4iC6h+9oeF
J/Vggb6mL/5WMHtzWnjEgC+FWr4Nz5gY5/Xk67fm4Nv6VMY49zonQ64MFo8M3V/Q6cedOQqK9jvT
7k+F2unGtpv4rBV1AdNF3YAwtYYrMVKY5egw6xcfuMygqEwSI57C1Ue37xUlXxB5I5uYnb0ezwbc
hW9lWM9Q4L9qmmXIYP3rPywu+PYy9VkOYaOeKLIL5hDxZpmHmrJ+3GkQ4xx8jhl4uuvNRv+4PRIK
z5rWS3nM21bgkjU4OT7t3Z3nOzr645gjcGwzK2JLDDuN0WnzFxB9b9uijuYQ4ohOmgSOIEyeHMCR
pau33X0Kz3YA8hDjDkAWXedcfXfCrJ3eHYf2uezYyueqH6Ppv5Va6jZYfC30vM0mczO5oea0m4kM
CkpiLXR8PH4DLQyjnnmmegTnhIrJVzL62C+RXISzprnZqaziVqTg1p8Q1KCIW3KHJ4zLIvT4mWZV
T/WUvqX6v4C9CslVh+nRqV99/pOnJ3XtC9Ov8PPcHEAISvUI/2bY6OyzxOnzrt+kaVpY+dUws5EA
FfQSv2m0rKMvGf+/lBkYDz6wzEESumPnNyz4kybOnixsuyL7pllVNj4lGXyDXg9BFDWVsEpWKd36
K3hqN1n3XQuPzPHCHzVn3aKlzk+67wi0vLr2iZkmCWiCjQcGMozv+6a+4J2CvFWqSjVxROsWCbdK
MReURuuZFAlJ8wGW9VbUeMwT7Xs1sPyVleLzf0RXAVqxr3WlrkcQYzSeDGR8Jmwujlmd/L28Ktbz
v9sVUaxEdi4JsSmXTcUsr7LP5lV0Hu+FerZvuTdXAYX7mK24UDx/Zby2H36513UfQAoIAxh7VTN9
qMuhc7E6YIXgSDTq2bIPkyCKKqpkefEw+F5QQUW2TMxzAZZaKf4yN6kdaXDFZo2I7S/eiRUN/f/b
/6mZu/Kk9gh6dmPXqUsfccIIPVp9YjhjKBGxZ2rB0CXBFoCfrXFGsSVRhV3QMz65t/Vlmsg1RciW
3LOjfqRlvM5cfHPLX9RKXYSTAVCcKAm5keOmElke40t8GzkB3LuzmxvNMx83irtzVqUHJP2FcKF8
8buojoPtfj50NK2V2cDkp/jpcDTcJ8slbA0GxbRWmwz5RUnly2cSwr+Z1deIBLUbjmaDWbgJLHTT
EDpcy5y6lY6YAdKU+ipM3e6fPI9e76lCyQ7NylMCz0lvyls+XjKagwvpChMnh3hqh+cRE8apHwOl
J+sP6dVTzhxlsJCz1EA3U+bz8f5G6YXZR8gPtwe7sJ3pLJwBKyknSA5wuZQg2TZMi74LxSS5mrsl
z27Dv7dskr9kb+uq9NXU/INsE9jqAZXV1rqoS7zdjxJ5DdNnUtm1N+YEaRceN0Urid47OeL27T7G
bY2iUbB/JSx/B4jFxzXv5efi/4F+7hCeGebMGfKi8uYGkzftwYFi+W8FBi3mX1aMRrhWHwVjD6a3
79Ilt1Up4MykAsCfQISJbzJkEqWPnCSLBpPwuiQz4bpU+cMbygGrGOMRLwKUP6UFofGEYIWavFL+
LN7Bed/fttpYy4Ulu/0eBs61zhsNP7hCBspTXboaIadb3M9kjtJdKDZzxB4y/WIqvtM1KHRxdJkU
A47lGR/4E6OGz/k44RU1SFVAuFTccFW5cRW1Z3EmHDeKsPe81+MEPmV5MU6NtgkvBJp+iUgLoiGN
t4cjMuMNmKEfgqf0LRDcNScRZcFDU2jQxeVYQcLcrNhCOkww3k18NeJgvR5WVVjmoLMGBjRTNVEM
hxZrOEG2x0RXd8XGGBcExAeh2TISWzMBSV6InEgFdpJ7di8KqhdOWR/jduDMldaghjbnt3snNeJt
bq2Y5+3cTbP+RW/bl/k8OwG7RRvfPnaczKLx4/7VUVcrgpuWp822bhiiLli9iR8cA4QIr8yZFhpD
qtAsFfLQJtWj0nBLD1Bzrl++AGQBN/DrkPomNllChNXDIibzoN7wkijoEZiXDyzOwC9AQ1RIEah7
EH63XLNejaZtSCBG415YKHRqxJyHPxtdIr5UgLazCewWZYVcly0zY9OcCbC1z3wrkE5b+B40jx0i
pxNe/gK5FoTQWilhIw+yax3RWPQl/Y+ns4+zrExz84wBwHOl2dEJfgpsLjOiXkpR0ih4Eifyc72O
VXcE+ErUaClzakmmG1xTSxDhysIpzPk0VdWWhplv0fZqgvqRsrrZrhyX3/yC1gLqPrOVBxaFr8ih
XGq0HyCzRVsS93BiNz2fLvsE14jMUZUX51aH9a/mdUDVix8RdoRrF9Q14TTxrol1X76+2ZPdD74J
aNn+9qi0fO8KBcpPEs9q0r/GNj093LQLcbEQf3J5jUll/tjWS1jazrWvdBlOAwTf727k5XgLCf2S
0Xhgl7kEIhMb0FMu6bu3HtILyFezzMOjeNIq4QWTHi8VrNT5l59fdpki1hk6orb1budJWQoc2Yr1
r8DS89wT/HyEt8NQAZfur1PV7plpBjttGtnC+H2ertm2pDgUYBrExMXibqht7c/FqolNaZZ9x6Kz
+SeXo1eV0wIv50PbZcBE62U2bxlF47r0eTMLIIeOgT933Oqpt4BzCHEJjAhiCKjmkGV53XDa0pk1
f3RTqHjaQTNyVtAkNUMf8uK3bjMBTS81VCdDN2Ljpq+UenbJxH49Ae5/Yq5yrAJCQF8XgBytkFWI
s+a5d5cHSv5RTSRYERZYQotW0ta33VyQW7U4MQUCMzfdMgLW5VpNxiarwCfkuBEZH6+Bf3J57Wh4
DLFwU1IIwa8Lyguml9GKxO0OYBUAn9EJbeZpGhNJ3yyNoBEYrIsykmbJHWDjLNt5XN/lC+lX8Azz
HndlRVsl+m3IImjocwJpmSTaTiI/Lo4ZgdYmGnH2tabEaKh9AKV9HYaaaN3yCvo0AbKzom4mtCvu
OgN5MYQ78XSzm5rIrjCQpPiO+MG9r58QJpjEpOYNo8Drt4fxqnF9YMMJWoSrnavw5pdxJchdq7Ax
Y479C/91YyoyR8psGWzhbGdpe84SjcjmK5zNRzjwNp2dOHHIjYfHUIasK0FEcoiLiCcgx4wiTVmE
MX+wMvMw2h45pSGer7AswHyET2ukq/OcTRDSvkK7EYQu3ntGx2vMNIuQ5ihXGl2f6qOSu89B8YJo
xSE8h6/QsfwE8QPlqRsp5/9WfTlVPcpzzoWdSg6CmOXOQo2g3KLeq21MZUKUxN1GDnPYf3lJEHVs
54oU4ygWGn9uRsvqd/lcCy5bDz43UhmBfTnIY241TPyCKkCSBPuqf5M413nh6Y+RTobKSuYzTnK4
S1++5/FAc8amV8fzgUPefCE0gFpA/hibsV6L/73AogevD90phU60/bCBp/QZcav6c7WZjNxLcMSi
WrqNA30jhHYImz4ODUuvszv1hWUcEIHAPfUojWEzR9roeuvzZCDvBHTwksnDeiUrgpiP8NTy6Fv7
yqbtfwpokxwTURTOxRMMmbd3L3fTdraXxo/5+bmPBiM3K9Sy2pU+XbpXz6+2fKdgzXBcfnTLtgyN
1hRtuV31+MSMSScn/Uwwa9D70cg5hc2XR6jqPZ1God5AeK9If8RP2WEPvuru+jiO2YjKEHa+gnjK
LtUKHkNckOEe/zLw1XRu+Vh30LBd/BsCrFBcviLV4qbRX3nKV8EOLFd08e3X7OQnqHFxeNesxu/M
1JwHC/QgHfA6qYaIRzEcEzKQrtsPDMFYkfgjoJnlBBT4GNOIqZFoeM8u5bqQqgue7DpSwfagTVS6
KxCwBGOfuoegkYc7JOXV9RszT8HTQYSGDOaoLT5b7t2VKpJ9+ywjdEftlaAHwtKqLY7rCzqiQGYg
cH+ujRr3+2LSnakRVsDQX0sOjzqz3DPjfcnI4QKj23OJS2QgBj5sARfW4u12yZ7hBnniLw3/BQHq
0K6eMhk7HBgtUxnF4khAxTY71lWJHMLxX75Xy/A6q+wdOI5i3L7QyMlbD8qPF2+srVBi+e6pvyd+
6rZTItEEYPhWK/s85J5mwTXKx37PgiBQV7Oegg/YhDB/2mSZCdJYi2m6mgB15XbC3FHVXa9VTvId
h80Em/StVrBm0WQd+AgibkGEN4AxE03uc6maIG9S1dxYikoiuqiRLrjoJ6xRp16e3lkzQttEIipf
oa5feCMK4038o1m55CpPFVtZ7Hk3su1u+P+o07EBs+TAbmyvpSsjNf411HR2axdDhZ99BoXmP2jM
63ntzFKhdeNKtrHSiGTsXvRSmPzBoT1NV5Ksex7/8NoWiFMguxm9QP7orAMyZj+lcbhIpVTLawX2
WrXSTAMXKtWQy+hEN8YO51CMZwPaFm+ii4MlX4FDyvJK+k9a7PMpGV0nk5me4ZRPvcDzC8+MR3tL
IncHiNb50JIPcZOkvt/e9aVS5fmmxeXB5CD0l8rHYCxwVrgPlUtyXpmcfY+CjsV6CH5Lz6srvkIi
Shx8id4/nIEyQXdg9IsWMmlyinUpLJrOEGjVtFcYft+a//4SndlvaqxraVPJW1PVkRZ60oxJeSY3
3SC4R9UAeH2M7xRv55/4mdb8TIprhAzNCC3LUo8HyN7IVSxqeNE/NDFzQ2NjPb0Ih+NtlJt8JdhQ
LFvubA1qqNrWHqhprea48XadJ9HWDCDboWkAv/RiTISHofbX6f2/mbXcY7WVm8gyac++60CV29gg
6JWo5ulGcsU/LPWHNUqcRAIol2Dft7T2orsd04LbbrZ5kbBzQazuV3uHu7X3cFNcRo7brVMo6yU3
rbu8IvqIqyAhvYwkp1+T5oSC4QXaSBBGVX2Aibh0sMnDTHpmKgENHJK9tJ9QP7j1mPbgaYhTtpsB
kF1GP12tBVmRKoo8wOoNY3a+7bFzOa9Lin1jxaMDxs0k0nJEReP3n6WD5CnyuUllzTyeDNnGaUuy
b22yp6Bqg7TkPG0HmNt44TtrMUXPybY19+vtpCnNS/6xyPtYjAcGDj8a53Z8oWMIkpdwEYJHnS1w
doWxFJeLp4TdnhI5y/ZKyONAToR2lQh8uS28Lb6hzZOYG7vGQZNswHhs5xLRDxoP+LqeZGNXiXNS
ufEEEyhJBZ96g9IUbBOg5OsMg771l8DEsbJnjTkeBlSRUFtRgKFXB5lylRu4IN6FK8WuTTHYW/X3
i+Gmw4YYruYQ9Jp+bXtZ2qtOSVWrybaqV94yHYjpSuajB4KX5azHMfp2uBLh2+wHWO7/aUYwF8td
W1fiSbDrw/1cVh/WZDmzS9WrMvwuV7B674FiV7cBqK4Ze0iWRfCVP9nzCulWxn0GYsGmoIjqQlyj
QdL9wGP19pnCgAMUEXupBUcmrw+16gGUjEAtrAwNEyBx9mk73+rVbwCG/HKHv8oiKT7/Y+fB2brB
iCWkay2ojdGhhbpVnR0Q6pfmNKU1/EBJLLCj5ZVXF7pi3WVhxGso4j5P4jEFpsA1idGmhRDycuus
R6G+6S2iCK/Sr8Dreov+cIClcyQrQ/N4z68AQyptR++TzQ6CT0SOW3kQzjAN0HEzjxNDJiUAPJrP
teDEz58v0t4PXWlPRlMgKI2rirsxM4qE49hkEgl89mK/RXCJV0ozJrFmyiU9Fr9g0yFzjwjT8PCR
B3XfUu54Sx3/bVthxub/B6MC21bkIqSC3jD5mKLSDkTqhsnLYZKKCtsPQVVkEaCwzahcHNr8oKm1
2C/8Z5naDMRRkkI8USZ59JfGDJJfwzZ1nyGx2ijYvIaUt4WrlljjA/DtyUhvXaviCFBP9yjh8i9q
gi3FHHlWkPRKVIue4X3VbXfufddLOyMFZhvG58Bu+On3OMSBrQNCgw5qAaIbq7QtUxzLcPZsisea
drjej6T8jVJs21JSZM+iur6TBSYroU+IhC6M/8cX/wpGAcoIJqMoiDhg8qHRcSnBxSJlLLkMzjSD
ub5QW274+sqFsaa8U7hqV5KEncU2WrRhfApsd5qkRClcWO3smiPUfMgYfDxAvrLONk9qLfEHXr+L
aRVECnI5+V+EQzUB8LtpBi8WXxbWD35FeyEL7T4dqPuLovVi5+0G0PmvY2cXTcpK+RZKHW64FzXJ
Cd2+qKtd59mOs7qJSpnToG5HWn8HtupA2u6YKfhRXEY8lm5erNclmyAVsXJhi+xO9ZM4oVNNr8m2
ehWq0s5pATZRWhDz+nuH19LnglFLCMHGSljsyQTkVD3ygKzKT//15E3BGfjnHvl48tT3aHzl9nD3
d+uB9xHMfAr3/GbVcAbjzXqK1CkDwgDTCvX6z6J813tYs0CI8gC4Yg5y73iXA/ZM70vzHFBy85iE
c8HKs0XApywWTn/bfxLpRl9cnFYHq9UauZq1DEptprtRWzqi5WhyIdFsw8XjAiHFEmnUlPxrhimB
mQUr2Xfat6u/OXJYyq3TvgEfpXywyKn0tKWd/lR+AxsnMKiTZbuv24GJXwNtBiGdCfhWx7xvCvSE
qvDAQQllWcMlYABZPjPmEQtGGHjts3Xt1zmItJ3/hG66Z72O+7yXXfHZ3b7QlB5va9l1HS6aVD55
QphUCMhAQMO4POezDhkUmrPjHCZW4KNhtwfaJem7KAx51HczDyhl6Hcix0Kcem70dUqnS7WOafYa
BKnt5DOdmODFLz8o5uxnrW/LTRPPjkrB7gBTu61fHiOrZaerlOX6voDO0IJA6GC2JyWR9CYICpEY
JteAaXSaxfiTPMZpZIiey/7YlzAtxDIjPqYy1sE/fE+E/HU/rInlR6R3RLvZ/H0GPUpWR+ci3+uQ
pWI8TiT8OZHBiFlwAuXEKJQOBMoCFWLtIY5fOkurT2XIzxk9A7+PFnIa7HJnVJ1hPN5GHIOGYlhe
UP8HARuen+CTaFRmUn0D16XbaOcjkUmApHKKepmxTwhKPOlS1ynPZPIXl7K/C98Md+E/leCnZbCO
y7uR1301SVn4zxHP01oMvigFbvX3pf4uykmRMZ8aexgH0TO+hwVP2qjBf7Bk3TrBnQqsoAsqxzPx
Nuu8K+cLHtpqG3rHNlqwV4n5JXZqk/wtaO3tMFnzw5HuRsAj4Lo7iDFBdPRIhcSoE0Y3cEd1/xTY
xCvXJnRih51akFStNp2CDTLl1WGs75rMRLaMU+i0nS/Y60q/j7gC8gJT7+rJQU7+6G9ViWmTTPrV
BN3N1+l2rWMXp+WhgM0570n8Z2JZ5Vv+IWTiwazZnSknAkWjQGvbcl0r0cdqmlg0dPlgWd42fOAn
OR8RnBvVzR4kUmPkrcIcpsyq6+5EKXLFB8thffWWJaI4Rw3Lh7vMF7iO6aUjJdE2mxuaS0wPiIl9
c2+gU58Ic33b3GAfFsd7WTaICqdnLCppe+aIE9zUG6p4mCN9U6rdUKvNI4DUPj83XHDJzMmokvmM
0BASxeTRIqZsPl5+W6lohA7ZXGL253hy+Oc5zbBvLVkDmbxC4MnR8tMSeGb+96eSCcwQrjRJ2dA2
hUwh4W1uN2jWj1ITF/++oa/+i/GmTbYETO/mHvccrEpHt1FfhRMHfkBexOMdILvN98xs7fQ1pgoh
hYuvBM+CG1RKwpcW5SHShvsHjugYA2cdtuhWGh3ojAQFBKeTYkQQqlM1vFz4zv3RTp5Ji4oij96p
Bg7MsByRxLgIvx31WCCern1HwbWkpw/k1PKVV84y4ZYe3aaX1AQ896F0D9XWIesnj33ULApVyEVa
VOS+5iNBjk2FVX0/0NBhJNa/lwsK6YOLo3Te6HAhzPyiI1uXaQcdCBAR/p7y5VVYqL1KX+w62QN2
vQZUQc5vPK1+LYezHLCNRqXJM7iMNDrumhFS+fYhStlxMZwFYJrRf9bfb2DjQgu+FywywqC0RzkX
uBlFycpqBGeq4tf6a6LhATejyCq7kUlYatS8FuWcYn9ZZ4LIsC9eB4ufVW2PUCfQtNyr/YBbsZ3F
N81bLPOg+4bgpOo8zRN1liry1xhVwy8P6oGw+UDdgNpTq7x++uU4KSVw11+9FmlK5DEIK4o3W/pt
FRooFVdwCzdV8xv2q8SxZA15l1jvOtpnzwu8zhUWCqlGrzYIaRXp/drYGMC7oM8H9IdZng==
`pragma protect end_protected
