`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
ofUWF7tG2yivB/m/er3bTr2cEb3abjP11CuPUNRb8GCCZn4FiFO/SixJGWxIv1hLtyVEm+MvKrnU
FeTV2v4L1H3psjuL+hBi8eLtKdbs6JqXHX6dTzPZcGxfXdNMF0rgeFGT6XSNDVavPZ2vDnlQPDhw
/eAj6N34+6/9a/op4zWxGikoriszU2MgmO9UTa3pQ6BEDriecfZ5spdoW6pPiuq6eohKngdBcMK3
OPU36ByMe0dmfP4NaJAlGlRUyn/mKa7uCXOVcQVpWsCUVLECwgPrhKcJpyov1HDP6mEMVXMEdHV2
xJZfakm/xjYSHzGGI0oQWY3wSVeSTytpKlC1yA==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
4DvQthXm2r8/7QKc+nPSJhyw7wzCFjnJqdUTsztt2p6VAX5dk6LbiBiZg+goOnX6x1DxHtpIO/Cd
1jRV31Eu8C+sTNii6kMwK69DHZRek/qbIPws4n5B6XJIkg7BV+pW/8dWrgrR2UiYjy11Xyww4xyV
GVuE3IKUetT+tQIukbc=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
GpL+GFpGd+9DxHbgihR/SBz/WLuIbd8i7IdYq9yGEJSnJNhqD2Ogtfxuh32kq7MROA7UK9gw730G
gZOcRQJUBtQf7Lo7+TE88rZBXUJXzOYaCQSTarSD0IrLRa//6boTRphtOLm7FhT1gz9W/sAxazd9
iB7yLMl1TCGihNllEdk=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2720)
`pragma protect data_block
HBx+jNZ71I6qYxI+X0jN4BZei1eOA6vsdvOOnq5y5i+lw0FMyT6BvsKinR2V5w6PEjEymBYJ6ScK
xZ6oXpro14LJg/K14Iv10aAVOXjW7yHYIbOHHifzRtJjmG2BxJb1CoSUd2mAOd3t52FLkbsCKkd2
45weCeXARRoXmmfcPqDgfKUgTYu7xAkllLhQwFXZLd6ZBP/FjDrrGnatWzn5pqKQfUxWtMG/N0QZ
nBmUt7FGjfGNDyJauAcbMIfaYXQEpiwJxwiUcKnxMnQeYbAuaveJb4bj91I9ZsKNAfWUBniYOHSe
gle3OKW9jqberLJzBHfbTiKC8uvThcwo1Bor+VcQvTVHLz2/5YI/3p8BShk0ZAoBR+S1eua0qbgL
88JpxXNUPzEyP3HtnyYueOdHoZ7pHXVgKDvzrYuZlpSZhttBBFI6lK8IFTf2un3NEfWKJutP/DZp
tDp1iBUjUOJn1r+mipep36NdRfsjoS4qeS+Sdt5l4HMIS6CR2a6RHsbyxR8MmVrMh1uAqQ0MmUJ0
ZcCR2pTuZT+LiYRxQtR7QwXTPI/HeYo4y23YZXzfvZqGmJbldW5lQM06doAMuSCrlkK/UsSebZ5p
35kJI7QNfWHKN/CHyd2r4jEnRmdB2eSTg6o6faf0kmraPOgV07rrruUTZlkqdY/q/xNWZ8M0LsSB
vDS/lgJs8fTsExIaTCY0fTqJTolVb5JqBCJXDHYNiyHb0PyRIRV7YMxDxU5M3ZyVNzpNxtr6OXEB
nNUEF8fd9qZNo40tZIDg21l2qTs84+64sh8pOKDsFji7EfSw0HD53lY8IU6IfKWY4ci+DCdZvAtT
cMVcvlCqIsZDnZRwp4dfTEHjERq8c7YXr74565kAHVGA3Jl4x3VKid06Y2gg+MdPJZEorVeAgy96
ySj4gFwcCRVPSnNGq+S9CW5kYgrvKauGk43Zmfd6epdd+xJov9tUB1y4j3FxhUjOkRPCfs0gR1v9
CGgYXki6fQsys0kaEoSpzCNRh6hUk55tpgsJuNW1RIJOkarIQk/ZwATmH3MsFZDsHMUBG+5G4w1O
f2UEaJ0j5X0LzBT749AqDRYLolEJgllSVr5HJGy8eLKnmeWN5yTdrvyUaZPl0NRCoa2dT3diosnz
RyRyhtl3YmZJgL/D9i/EwaBo12lJBtr44fFKCUaoFZVrPogavCik/WfCjiWYR50DkftXhgNraDqO
tbCtPR7WD8QhYSHILE9qujbpAKTIFpLLbHFLEuTQAH9OKhPlGVQOFsnvikBFOVoj6V85dEb9a8YI
LJS5zisc/6KdUZUhMeTx3NRPofugOhvaBZAGgpL+2hKuMME3fzVJt3bX34SHsvDgXWgkHO7bHbj9
VWMpu+qbMQoAqzMToGR5r1/RZSHjXU5NS/o3y618mt6ZNfmxlYUVuMlVxRx3jcmC3FjlaliyjU+P
gfpTT8qHkYsZ9YlLRIBXlt6kLe/r4kNIwfXiKb//fE8mweFzHzLXI08oMDSZJV1i6hP732Vhzv3e
zE9GYzDOBNeO4v3HMy8exfVsm0IHs6HFTF5rfTDzagGxFoKYdA6gQ/umraHg5yLsqxFaNo8PlikX
XAcBOw6AB9YT9kgHEdNBBPAbzGW7G6CLMxpj2T6qN6PfjN5iZ7tuwD1Othi4kjAKzDSZdnbekUD3
n7nR4uu/hkSXYMIygiJZoY50m1Cv4f7b3KMKPZMuk2WSuJMQxvL6idAWBWrhwvrisu3KKXdG3vla
TA602JFffErFCi4UY1PJsjlSblMdOutwAe78TTyc12w4TmqYTOgK7CTPG5AzCc472RiJbuf4sa63
qRi14hvpFAengYsJbt/td48eqsiMbFWeMpY7tWvOqlACQg0x+osBIwbPCApmb+yGae4OF7WzZcZD
Kevqgw+EmBsm24AEofqG30U2FEBaqHtfFEPD4N9UmtWNeK0kx+1RicYPdyZFOgJcUEE/kckUhAFC
ugMv025l2D2aB4JBQLNC0B4B2y2nzy7svsy5XgX7fPaS2AE3hI+T6gNGvhHpYj7tLNFdl3xwM+KQ
EcIqZBbZO6LTsBe2P1UE6n8Pwy70Y/sjBZk5ZWjfoQHr9EwLWtLzvGMJyHR5cACC3Ajq8pXJnP9w
vgPV+ttkwiHmNf/dgQYPl1vc99muQ3H3CKxDG+HOUDgf3Z7ppAE6F28P9G30jdXUTQCVIRlEJ0k/
K34jDVwZ9CxUTcA/nEtNYh0Q/pvUSb9tX6b+mu8esLwxH9nNCjtVzu78GmpFHBNDcFZehVbZxHMH
gNIN8aF+FFfaoq0gSk/bzAM3lkulzwKrGR2tR5fQkQW7tqqTKigtTv2xlSWdae6hP+L5O8SELI0Q
USJphxWleTw+RTWfPBr8VGPOFPu1jqkhcft3J/BUVrKNRY+anUJZ1UPr15QfvwaRwxHayaoIJohS
sfLtGqb1FkhbWyNA8zxSewrvYTV/orNF9VocWFFilDwljoX2VdoW+fQbXBb9hPeVSgjPrCwLSNlX
cmBtV8M+6+RDkBJL1Oxs965VP0TxOnr4jXLAFPN1hqsMTTu7u5GhrLnRWx4p3KkzC9iUmcwqhzdc
p3fC9VXNzgXiwgLIeX+oNaMhQejEhBZSI84trF65zNGWUxZskcScxZTV/Qmgb2Fs6EBW3y5AhZL+
8zigV5GyKp0fsTvyd7hwKEnCEmuGyq/bSWQL0I5dXTOKG7BvkciOzovSYqoCMZnWz4uaU9LzvrxH
GMAOTJkOGnCWtK60vkv324/q9X9VD1s3mSxNlBqiEAKUbv4XRfg5/qrO9aW5OFQ1lAVD4upVwCEu
RWFneuPiPT28wh3z07Tltdv2HcpiIDZ20P+FaNkc2mOlTw5fzulajYkJDMzxE1eVF1pmzcncWluV
zWl94Ty4zJoVH3d1Y0XThyQQpTxt8ROuwJz8jyCzoPRJxmjrkj6XX3dLZamkbge51/P6WaT8aKPT
35iug+bJvVbZU4Hry/HC3k4iOIC9yz2oOtvJCDdezgh5hGjpK2aanREK4iOF4EgNp0zEhi7SkccF
/gqR6k5O/e+t5bzzWAKs7WuOqdVA44jriEW67lEIkhL11C2aaLIFoJ4K5wEZbxhHHcwuGSGzBQ42
Nci8Mgw3cfCknE9yWRXo5IEK1zD1RJV514VMid4AARXV5V6xr2YSF1uPx5bjdnFeWULPYqC8ZQve
3xYhTfAvU70o0zRlfIBysFfj+9Nij5/2Q+NhDZOIDqHGGAphfsVgiJtjsAtTQ0HHgjqf0KKXOej7
EkU1coG8QHZ5RjpK9yHUJN+Kt5youvDP/aVnvkdC0NsWce8NzgSdmEu1AYUqYFT20nwKPIHcmccA
0rsbPFkudpvrSmTSiUvU6G67d4Hvj2AN0VKdWoAOUoWmHijcUY3MehUcIqzG+cHOxlPU5a92LKRP
82hg7P1OEaMpkXrQaePEhvjCWT5aKjcEl94RniJwPR5+0VpEBaFWQX6JByelV42g6gda37zqv9Bs
/LaI5JSxr8n7NENxg0BGZCYC6tIKWzuET4lxjDwk7w1+DCCEiJTPu8/McECk5QziBm0da++sPGHj
2XyFVK1e3nXxVlFLRStJv2+0cp8/XBYyd8/mcWBFmqrUwixp9PTFNlU=
`pragma protect end_protected
