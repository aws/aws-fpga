`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2024.1"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2023_11", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
YdffDp8BrqZg7IZyBAsuNFFIwV6KyzaFI4BXwZNWDun9ZRAcFAnlGXkR92O+tcaoQVVh+x9BX9pW
an9Lw2JUO7InKWe7aTdcbmzAJbJ29Xf8dmHyrgw8wMF69A+cB5jLXrCPYajmikThGJyB8sUtwB47
zMIR9nurHUOOMubaPglXUboiNXt3YZS9Ep6C5rZ+4v+0VRB29vFv8HRY0nc9PQp6Cc3G3WviZD9e
5MR2fj/PpheGIWnGNaJPF6r3ZqWsCHldLEnl44dYmYVNctmR9mon0CFffNXJ9uWN1c0M5mQaxm/i
G4Isztfodh6/IzWlxHq2fs5nZ3NecRoHCInxqA==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
Y9bLC5CWpWtVdboNEUrdYj1DE4fsz/HjyCOtfaUH3RygtZS05v2cAGcjmWDL+LWB0tpfPUXkilbk
srWb95PEDUkz22I0Fj28q1H/NEQA0EHYlvaMQAMIHCHVahjHfaf3swWfNdJVn3MX42SgW2hKTmD7
rJBkkSSqsODGXRrcakE=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
mh227YmSR2QdIlRC2tlEV9S9AYnkoRo3rJZKc7bBStUENq43DUF4inuE879/JR6j9l4YfHPyqmrC
4vUaxnTVBhIamqs64FRNUmo7OxEJAazqh5kBVVlx4/T9cog6zYkhgjBqmCuVC1mfrVftUuxu3lM8
caCHUHXvqsYaK0FkiCY=

`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
YJnSSwtEM5zgEE2mH4V0uf3DhXj52uhvpdnzgM9/78IgPyQfzKFtCFeZrmPbTUeE32PQLr1bYlXU
r4c+t64X9A==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 82016)
`pragma protect data_block
FXtnuG7y0G/NBYKK1rDbKHrzXDND2mdm/tFipk+5ke1EISGVTP1D5knDEq+GgGni6IyzSe9iq/H4
lhDV40+/2vi5VsvpI4QpSnt7Z/8I12Se6pMUjAJ7otj4t4a0KOlBEyT7F6kd09r/no4R0hqB2W3y
5aS+MOaLaT1w+jxX5NAcox1WbSSc6bA0TDHiXLlG159GYzEWkqHwV1U2IIfquJpffOwjPxhVMNpn
uxk7kotJVig/z9g8OFKHWbqV8SaOg0sPQml+sWyuK0cYzOi/DRPZdLNo++Y/+iebHhdxXOLBN1zv
HyeGSqPqe3+HUaNcdNpTBq1XuglgnGSF31mLR4nFNOOUTZ2tw9pPj6RasAZXHrKkymq0fI8AW66n
+iMS5EeYoN3lshW568ls2BfU0Q+8He2YuvZkLxmcVwTcLoPLSa3tHqRTtAy0XL5F5kOSW3Oockmn
jy0nSmrFNBURQ3QuLAMsxx8Z6IM9C+JO0/UClzbQ/AfheUClszHogDk1qdj6UnNLCGt2DPtoBPEP
zMj43+KKFRsXYxDz5pI76hOhqwPaZ0YScbrgFVApCV/BjH0qEBisnVwP0K+K0Jr6S3tFGrjor4nM
25Q5zVGNcPyP1TaNQqkMS9vq824s+9v7EE8smRtVaq7fRDV++pqySXciRJ10tYjreWdhcqmPf/X4
bLyb8XVhkJTHkOXBfweRGTLZMVKJDHX0toF9hFSNol8kTmZQiEy2qd1BUZ5h9qjL25DN138BVlgL
UjUH5WbGrUmUG6+nugHVsmexzzoVTNHnPsHWUCFkx9ZD5Sj7/FxeSPiIZrwERb7JIfDEHxInQiAj
4Xmi0OLdrxzEuAiEt3doLp8ABMzIj4kPk1KTdl8ro1uikyM0SXjq3LeoGvUbzczoOrvvyBVkEVd1
S5kxNQY+3U4TZj83CuHmuceDdAULguB+BEcgjFR6+RrWMTOJvcMNRpJ74JovQWLaCrNYEnnlvZO3
R6+H2JdZJQnz7HCQuZeCe/Q1d3SvFGRyLhuRJJYjs4Uc8VUpV4ggFCAonyQ54FroKcYZiQwXY5Dj
Yw4MKtfKf9mRwjIdqbLcjL9pZ9VdN1JnvfgJQ+Jpt/2vTjceg9HLe5QTctz1qDdOxdl6wedkqu0r
WB/jG7nvbk4Hzkr3k2aHWksrmLssIMhvhHdC8P4SWGBRTUINftLYQ0Fv6B4xJm81DBL4ydF1si1H
oUiGJ4gRvW0M+5KaI1S5m+yCFKemJte96ESdfwWJ0bzquAXGGBs75em84sdCo33k1QELkp2vrm+A
ULQqVcJ8asbVxyWMRk07C+5ECBXCWypHTYzBT5jOkUWXv/BeGV+7v1Iy0A/92jHERbwZE5GOQ7av
0wa+l8Dg4XLLRkk/KVM3kvSOKwI5YRn+qVxfl6xN91hHao8nGVk8G5E+8zG47VkEjLWTpPxM192f
TDzCrjAqwMevK/dTM949BWHo3SUamnEfAjN0XLTNuHoE4HOAWKId0DwwiSyuTfc0Yk5hn2i20OAn
/Ff5Mpytd14n7vQfIyQ/a1lXg1J+1rg8NpCaUpPL185/taIXh9e1UPs9YBr/XI+Tn0+o85OU/qRr
anNDc2stuZ3RzMrn/o9Y4F4JcNsBP7g24x87e+w9X4dPRAyrpQR2tN0pg0SfqzPL8LKBdbEAXG1n
z5k1Y4+i2LCt/9oyjQMy0835m/1McrqrQLTNdm8X53lgENPtXmaZ8unsYILrphTsJnrswlSpJDtU
dYtR1u6ElHKLjqq2iYhInR6UEQMJFZBBvqQMkmJKwfVszuCv4gCZVfcTWJ1NSRDRBgLxH6o1lxWo
X2IhPV6G+kwjtC8Pa8WQwlM9tvM4EvfERqracAQ8LFW7+IpiI6OoBSmJ5qPGFaLhMgmBXUV0UXoO
zyuPB3eB2BNmDWBlsbqr0YXRUQEK1/NoV0bPrbBU8Ra6mPNjvK+MoUXIJwa9nbfZzsCf9iRJrrDe
8z1yBwveDwAejA1h5u6PO1xosmZCJtpjX+27ZhItbpc2EHOYjHGR/NQH1Cmme3k813AabZ0rWD6Z
qUBwzDAMOY/iQPptCPk3ffjpYa4ut5I/UHkgGMx7IOEkiry08SrkLuhKcj9bpvAxahnSzwrbvKjq
DlxQXkNRC3UPYN4Ke3e+5rsUZb2c6OSjpxNax2mElmv+CWEloDmuJ3ZUZa6mmyucnyYTIKR9pG/e
04cZhXAXqETzO4YTsy0WttMQush3aIuR7ttbhuCB6XDw7a133wwgg/F1rezJ5JpBae8tAVv8JaKz
8+aQdkla+suRMQ+M0bo1g+6b46LgPUaoz3pJZTSx7kqV8DLuEXfieBjKuQ6EfHXUP7bvq3qnmPWv
yisLjeIWLTIn+s8Kmj+/ZPTyJvZkUbybBr5SgmTiwzKyU1o7cMAqP2kr9g7ftvrjNRV2dPGDaaRa
BVNIi04F3wzmdN54Xh9TLVKswfRlXWfIv7gJ4fOmtB9wpfgha59UBgzzCFg5PDTvLKUuWOm3OboB
jvYTtL2DrXzE2bubn9MYeW4dsWWQztakA7xHl1IYLMiHFau6xZs3g8WN4T7Vfde3chbvRds7J5C1
4noskkdS+cO3aIQseofrX3rRlunjL69+/syjqZSwFc2LuS5V2w3TCiNtr22n8fBIZkRlSl2ZwQjg
YvOXXrsA5geEIWNcW52gEP3XPCQNyaZM7wtNywF2lWREeLRvT6uwXsefIlCd/AnRPjIR4wnrMrKc
5bW1BvKicMW+ZIsbubHumMurGogFu5N1jF3EBjxOh+KGNDp16/V6/DT3Q687aFFRDA4j6Bdm6Aom
WALluMVprCD/UM+x86gpiNWgqAFcgvlKjGS9WttxZTovrYGfMrHkpr1AXGn7WlehdVm0gBIQHO+y
ThFL/NZ9FgBsaPde1nJ/aQ38sgyKiEv0ISTLlIx8Y12y2K42AM7YEtHNePLKj1ghooIcpfeSDzza
ReRQ2LALmaJNBJJZcX6J9CnVO1eEm3yilpo++xfpG411pR9oJmGKV93B5Hq2kxuJ1nRm05Fm/lDK
Z/xypYKO9Q7FBNlXrCetq35agVnexV+W+xJVBNme68elyp64HID4hmDm6CdEVHkQh9m7r+qCoDU+
Ir1SNWez9M6Ja47W97UHXwgECtdfnzzRjNBmsBsJlFniwag/7utnoT2KlWNC7E9vwUj05Q/ldQE0
tzHd2VESd5AoEW+vkephNHodpRUQZ1gC91eRxSpYlHxi3NPfV1DamoMRNFRH1ERK4SldQWfSU/+n
G4Qr7dHDTTqmhvv3S5x9at9oVcUfUHU1CBxenBt0HfbKUHxlzDrEmEeXgBMEGKx318dzR0p4zd9x
US7ep/VVm44bOPaSn8MibeY2PafCRF60hqOzkyZ4859ISc6EEq6ihXXjvX/jv59GcS8KHWhUY+Lr
4bdoJoJw93RjTHVjjVeLypcSYxYBiyshF176kkkX9f58/3mqLA7XcWM7rEfjsnwAuTh7OQNlYPIV
9EMkSGJBrIeZE6N3hI8W+sWhSALfH1UX/5SY6e9jn8MAQKKnDKfGzk6OZQTPw3rbvZb2dolHzC9L
pRMGlh5CXvftnK6nAgKRhDdlk6igyhnKmk7ys3SKrDTHdltToV8MqnrYTIGzoT3yVgaoqVwJ7Ebr
IOtYmuHd5hZ4GCHj50P4W+rP5peUUZSNoaNmb4ESy40wSNRO268e5VNHcypq5qIuZDeC73fxzWeQ
8Z1Gp+k3+ncPo4qj8Fx/IeS3FIKIhbLgZ7e5KF7cvuF2nTozumOrnVP6FldzSUSPe/hjAnrjpytV
k/AniaKnjJfLSEh5NP/HLF8KvTQZRiaXzZIMvIUp5jo4wFcybEIBxjzRLzw3s1YJWfIMDlCu2keN
aqPKd3CfSEOYh2JsTKU8p5wxe9crB/ogxaov0ZCbAFbS8X3bE+9DV7tXkUbEscx7T/K0SrzaxuOg
ehsxFJtDn6pDTGciDERdl1BRCNbb+gpmoz6Jhl2xBZiUBlN2cfb77ysB1g7vdPcYKNmbbqSxGUHQ
TM52rtSh0G7Wveu7WtN2vV7na/6sOWqWE/ThO5rLCUPampV408FiqwwQsE9hsbQbaYV2I1kFnwA5
gsOy16DX17Kn0iTh9XA85N/9xtzR1a1kVvFya0Fb7MuDAa/gkcpxLXEyNLqJ/sZt3svZJI2RsFEA
4fkpL+Yfpp/AJBE5OpUUJIJiQgznUrjFzYfqvfOPIxTZv1cXzDd0FU5WO+hHmYMf/UFNuhwDDzLV
45ATzDpNunkn3Mrkp1wIsyXyyAE+0WQ5hmHDwQc4x45LlgvcNWwKtZB2K2MGg6wFZ/z4TUFhAj5p
zMNCMJOBxlvFNtVK3HM2lSSOHwS+VpMxwRFuiYr1FN2b/CB6qKhHCG1fQfWLo1L1B1+xcuSieawB
b/u1ZxYUafeJz2RXZ7aFXQ1wXngkUO+u171iZDRRcTw2nYFrlB5YXq+w04a0vj2fgjFXoWKDM5Id
ZlSnKZUGZykB+Tofn7Nhdl6I85m4pZzQgVvF2URXvnnNlHeEaawicgzfVL/VQOYr5WV5t2n2TF5Y
aplleUiX8TCmqKp5WqIEv7t9WWlz4sH4x/2b6n+B5iuHwMT6C8Pg9IaOX8A1quytNBFRA8oCZMGo
iw8pSw3NG93rxZdnwryVYFK2sScf+H8E9ZyAKsR0upXQZId+OFLWyasR5MfjsvvDZOzKaerRpic3
l0nnGk7V4LWBfVuefjEaL2RP65N3aZvIbQ86JQ7mCK8mkeuOg6AfQ5aS7OXHoEf5z1wnkZldWe55
fFGaUbbFQvq6hLlGEjiy4JEm+kW5yuk2XFDlS+95gGbTlVaJnzaWrdpiaiy80SawrzSdvD5xq9rK
IoOLvKhMhk1iDQy522NNWRU+PuaPz1lTH/2gmorLRR4wbWND4LSXkcXCy0Q0QtO4mtNptl/Bmp4+
K7N+HsrD9ktr1tTgNA9evYWGXu45n50I7FBFwXR0ikqnbbaZYSv+2VwykWbmai3qQfJP4QbdC4UG
2JeL3RGyxBWKOly8J/vOoV3quj6Vm3oA6qjyoSLRnoga7BJLhE5Od944hqYqB5DDrTP4+b4IL3AU
AIceqtEStXCTPLOU2XpQkVdGy5xulQKOpf6SpB8LwxBKzXOyT26Cycfs57dO2GmFJFhtD5HgNm7K
m5kLATS4YEt3u9srfNxPYuOulOifqzvKcWx7MF0HIFn2gyww80u/+POEIgH0q+pmOkifC1AeP1i/
RtQflue0lLjmho2ZVXyYXcfMh7ewEBSva5V91PJUCxOdZu8qOr1Jj8mzQ6PZP0rmiTlH3/zBg59b
Y/xl6SWWOPpRB20mCltp4dRASFFINtnbnJoSAMA1XGneHoaiMwhiZnvZyNVkrLRryHGnqvdH/nXJ
5ej3d1Rv4LlKg6gPa4cb15pzYiiPQ1frk2RmO1bdM6ZoLbZ3IvoxTWS6VRyCq84x/KfZrSHIe5Fd
svTG8GiT6YhrIP38eU/Uwp0ghhbWk55pUeV5sqapbEceF0vWh+K0xb3Di2JukpIfCPe3I5Z4Rgr7
rtzCep1hi4EABEhZeLaLGID599ECj/Y9Dz45yX9sk0aP64x+n3R/4+huD06peoYobfaSEt/V3nUx
kOzCTLv9ijhMX/tPPToNgl0hPb3Deqg2KhQlgNgx+8w6lknqzRmH+HNbSPRRUuRwNauV/TF71RKt
B9DbT6/lpl9lpn4vmP744vvK4minbYGLKcYrZ7cPTSUBbcqg3MDO0OmT289bD3aykJnzcHzVsHBw
8tvL2xoUJPSfoMv6Fq2ZiEDZyQOR7g8Sm1vEUP8s7QKzCe4CYArXpYDMgYdSe076o8JMvQ+NJSMb
40r/0C55W9O5dIBErbti5mR83q5I6diG1fEB08eZYGOjfv8xUwipR9zOawcioYiGnbNXzYMWyuBu
2JXzO6tGNqidHK3ILUoinTUh24hCE+5ErY0eFi/XZW/LcE4g7RZNHBcWZ/ijGde2FWroHT8RZGK/
Dy/RlxYS+x0LvF1+A1FewINhE60NL8jGfonowdK3usAAws3QoJxIedTXQsYclLspGtDUENKzKsnJ
fNFM+IKbud63ZOqt5b0WTmzbxEnSmzqCmOb7EpiKYZXyyPnKqYYxguMX2R/LNmeFKe0bawlvE3dt
IHhou0o89wCgBGfxugS0dkdIVh8a/gFdRPJNbkO5yPO3bwtvSWTqPpJmgB/e1tJVkSpHWviySgDo
y8DH9GULuloIJULGWpDUZtd5ECKwXpWNaSDjLeHDaDZfR5Ic0nn3qmTrHsO7CYNr8nvabzw/xBWU
u30ZuEG1s2Pm14ic9hWyoziiart6pog4gfIiCFBb5dIsg1zsRKY2NvR+tLGBtmqr7c4voQb+B6uF
FaVPBVJw3LFx7tXv65DQzWQUSj7rmdLY61UXj3pWGZ32obIO0mtyheZ+8MJYTekJtPS0I2zNbY01
f19tXiv1Yr63cGcnBBbXG2r5mUKlyaZBzD0+sj5aAzOIf8V4hWX/f0QMw3taQJuJMh6Odtyop1Sm
QL54z/vQL8KsnkLpVaQyI1XZjt6Wg1gXFvryEVzptaicxAc2joFqRy1a6ZB5XhOAd8ldWnm97gts
Viwaij60phxVoY2SArGR3th4x3N/XTmZfqLcF+obhu+/PDfl+b0Ursy6HVv/ZZmIxYx0hcC8qzKi
pR8fYv5yEN1paabsdkCHuGquOo2BnwqrZOn/yuyBWA/xAOkY6ysthLKgk3YOwimWVtCHL0cJp+5b
ggSdFF3OGijJ6ZRyye+no9y6ags0QuZgPk4vyqTsCOH+mJBeMfSCbGh+USJzgSYpHmdJDW8b6LQ/
5H8siGGjuW+KQ0iMukfAY15wGSUXxFhraN8Ola0k9dFvbyQG6tOHPH8m5qQYNQZs4SPAGCHPEwmW
xTNHOpCdWBUU8YoeurkTjB5l+wbVLtmd+1HW9BHVLtcYjt97VCa6BEBA87/W3pYB84sLmJhoYNah
74XGJc3e0/LFaxhq5lL9QeSrwgaIcjxddeQDPnLZuPjWbEz04tfF3PcKMNmqSrIir61yTgIEFxRN
UlPjoGWvANVL4P1WlaeIjvYg+RSYkucmpg+S9HddDIlUW4mo93wpAL7eKLl0T0qDHPrrpYYL/K5m
S55hsj63VPo9ymRvjfFuwLZJnj+cyHX5U0f34UcqtY/5+DSzn+ScfgLwlNCDOZpu6275wWcNqUbi
8EPEareEkbDy4prA33ZOQkVqgUUNTuAtci2xZJl0Xm3O43ncxxPzkJaDPFuG6cIC7Af2uvBoqMlG
YbpvyC+cEVSIZN56Z99tHmL4Mlb+bOaYNxTBrf4ZVxtfflB9JlzW+zqmTnvqvgu0W5xuEGSIoYeX
HL16iuxGxSeoz1jQhF+xni0QiuNTqcuKB8ohSpC5XzifcH4OfBJHLU+rLRzWdfPAqyTRJwkZMW4v
2WqCMHynEnWDz9qWFiU9Py88svDfdWENfxaOEwX6Wc4DsY43hTwjWWWX5uMxFBEBOopmRtc48Tjq
/ydGf2tzbvSvRvsHSrR7sQexiqonhRr0odGVLqcMpQJbS47hZEPzjnNrIbKXawcYdxjM/ZHWo2eo
febGKYLqb02Rg+j+VKYLhAmMHQWURtAjm0hAYz/+2WFCuiCp2K926H88cQMK125aNk9SpLjyus3A
qhesXN1dlUjWq9WlnsXTlUMaaeQBumtoPdBKFN6zA/qdsaNIn0+FuL1b81cV64vFnm9yCJFhj6b6
JfLz01w6RmD7nn+kZEA3ml+exN1VqCLSvCu0bSAbLZzKEvIfXYCeK344VUcbfgsm1COVG6ICZVLm
4SoIuUc5IQNSjj1s9kNZWccZt/5uj3AMUbWDFxfKx5MjoHrxIS70XKlVhRX+3zmBVn+l0Mu3re0r
wfbnIM6uQiCBqo9MAx721IBw0rA1vKU+JXRpzYf5VCFu/an6yQybtQzMV5J3qXTWA6mHdCiyVs2o
BlPDZ2MsMIGVkq1YIfLR4VDplhZfOrmQjzGJEx72EAO5uLqqOHsq1bYid3ZoLvlEV+WdriCyrqAW
IzSc+VgFP0tHcEXTzIEwpHBCAyAGQdGWHLls3YPiOj0EuL50hQhm8azth/Pdls1D7MXzNi1yrzJ1
XlAHLjrZp8iWHYOaU5E2h3LqG8eXWsVfTROG2m5qSW1FTpUIzCVS6GMZld75ydcAZADVxFmaqzps
g1+RatSRchQxb3WG2X0NIeckJEHxw1GJ/dbcR9NzUoDhW8k+/VT9OZv665AXVaYo6bDolXnHL089
2LfPPp0SOxkMC4AHsRCnj6TD0zJRKU82UR26ILOyypiPAJB+EWAMaxKW8Xe5eOmkdZbFoyQWOERu
bhS/0XRRFmt31v+657q2Yyu5Wf48vUUo0fDJzEXsUbTEUxNr0X6v+PaFdjzY28vA7XVzdgF7rGlH
HpzrXJaGzHUryYX2JqRON8pauiVDErLsdTH/z+bQ5HMbHE8CEd/ieNUru7hWNWwljKFwL+4gYZ1i
Hr6rRkut3Dy9nM8KZhvy/xRSU7642d5FwIh6TUihlJy3LtV3BaerrKmMlemYGbkA1bFST4ZTWG4g
qkpv4ATUxa76Jfeq6Psghs/LVhitfgAUrbjqGyHNph40dxDAGL+hy1PpNHqWJ8TFWfK9YnRpjNR2
WE8U/UFJ+dNmgbXXZUpku5T+GQTULFxL1BnVSWs/EwbcqVLGdWat66XOluGqlymRof8NZL++CWAC
BeqeNzzm5We/qfY3mffCOcWZoQ0d5Txiuw9vsXjlXQdXXxNoOeb70vL2Pzv2KCwvRERu3aeiHkbF
qJc9dXBxUvJRNvmYMYevpB2mXIzROYMrkb2k8bvGjttyqFhSj1BQ+U/V2EPmO3U1/tLLnK/BEj72
vAsGTV2BNmOjioAAH9pQJgpEvMvllMzTJ2p/fZc5xwQZYBl6odCD7dZBg/vMxWBbY+OQqtTr98/3
1UEvgXbUXT04jAILP1OkuGKflR88gffclLlp1Mu2ui2NIQImhrLbpwaidd08nuszL+kc71R0K3jp
yp3ZQBx4pohO0iI4Hi7lMG4RYTFmBvZbz2+gu9SzGQBkosjis6UHeGODuudHEsdeY2A4hIz7O96M
+yiJ3NBToW5jfKsdPgJwxtQL1b9ksSk9caD53ZahsZbH92UFxfDQmB0sta6aiq3FNc/l+h7yqsMc
eGMA9TxGW6bycCQaPVZT9xEv/bLB2vSccOmmqFecFDvKLbOKML7HVKPkL7lBgb9Y0AgWbqetWDI4
vD2FRCra9T0tkqXI2cEM//wdSvv3583nikQD70dzqfMg9E/njS16Cze1G3R0iQ0Vj6zZup7fAlDg
nsGZngObjbEP36i4yDcM3OmwWSBNCXMzeheVtpCfdLeUhN1D1pPjHGaENzzU6fHqEUYIyjRahu87
RIFh7AfgSnj5hBHw+/7cGRtYFG03ZMphBe0zBpG67WZJGW29s0RZtU2gdK8vPpVMh3+/jHSVnORP
KTC84Acm3fIYvaQGzObT0FMAWdCaey/sA0Cg1zLRV/nsqVB96h1XyBJNmXP18/5X3k2n7/zmyF8L
cbxt+/yp27OED70Spv8Fe67StSvtri0YF2snv38cG65aA77yPr6oQRSyoBPBKXM3QtWpvlvs2Rgq
9nfrWR7gM+vgtkp0s8L+2TDPZSJ5Q2kJGAWCl9ORa3Fo6v1MpOAaOY6pgOBeWxW3jd4x4trAUZQ0
RKLpoUrqVkIfChIoaFp5QgoEJZAAHcOj114oORinWwjFj1ZhgUMG1xt6mh3tBC0luOzBsScd7KVu
NKwzZJT/QrxvsQzauZ8TQTdz0qTeWW+9upv6K8gIhEWf7EhDI1L94jAQ0Z9+vJwHmGlX9BSzm7An
gmCR5PPKI0aR0QtaFygSCg9mpi7kvQKQEBekZNza2e60ZgOCoIkoi12JlkljTM2EsQlKE8cVCFYz
VV89eYsL8nF4/se+m7M2zABytbGRyh4IIoAnwpgYSV/wyydlYL5/6wypXsBNBtmEGFPzt1Rl2haO
6wdGL27nQBKMfORgDhjQYnmmxsYb/go1CeRQqsae8d/esxwo6I/3MpAuDkKkw3w5jk4d0aFxfoR/
jMxQ06W9qwzbcfmPsTPn30RmYrgU+Q3e7kMEC0Qwq9fqTNgBpfB1y1r6aUckVcVTyfHsuobaKY1K
Iv2wPquco4GnE22mMUYCCIgBdYFPrbs5UkwglO98Ln7EIXd+frsCodVjyRsmdcKxThPL1LcULo3o
coZ0tlDnilZiddJDuBL92wh/q1C91Qhys24YNFQhCvcOlVBiHEFGu0f97F9a+KbxEkcdSV+o9y0L
g1s2rWa3elmKtAYrydWDhLbBNnXZprsMsdmECv15xvVSH+p1FMuaMmJI0/tcz0Zawg5Ij0uvpz0K
z/ssbxJaOlL3r6TrrctApE1SsufQ5mp4kerGNNVIejW+iaWSky6P7/hgxT2hntd4qgHS0DrBGhnn
qF7zofk7BvIC+5dsljxWVm4Nz3iJu7tH//9pX60QurbWU3tfx5gdjR35bRWTQbuEi1H6acNzMCSP
92yiNFk3Lfi3Apkw/nsYPPsfBUlsSW0rBjW5vMUcDOQpbCsafe4MiV04pFoE/JDHU1xwP0OZXgRL
tsM2aJeOiKAsoblJcpgP1Sk6cFl9ZszQs/W6DCzeS/p3DMF07IhcsIX3DkSfeeQhd90qUMmCIFVy
r1wGYbjVThxnSpPpo2WxCYXwf0HG8rMnNPIfKjX75vKotJvZYAOHPyB7rPUM0mLGxLTAe5dP00A7
JZGiQ3DDb7lEuCf37XYICNtD00xIUFFnieojTGE1jRlVyb++BiH+rhiRR9gsBRYwQOkgFC3Bik8F
sFgTcGAirK9h8f0WxTr69T1h16QVvtDXOym13WDVm/UksqSrSgp3uSFC2UstDKJdM0V8Z15aoiWP
PE/TDOA96vgXsjH4i47usq1oL2XfXOHXOY54GFlPcVU/BtjpvkNgJKmQ8susrxmj+Pm1teLEX9Wv
FOLvxWN5OauzNk3RTwfwsFsfXiz2UoJuIGCjEgzBFdrPlt/cV4Q9GOBz1JKez1RqdkaS0VEVkXwk
X1gP3qteVS/4AjAVy9vP41lgQljJ9ZvcUkrRI3tVDH/gdHiKkw78my6iRwCadviFprEv/b6n5yqD
6Y7DVi1s8nzKT+ujjLNPwv4NWMD2JYAyCBs3eDomdLI+Xro3ZUeLfQ9ls7NkywUZN8FVnkynrBiG
yOZEU2hXXCMrZDavLZvFz2trsTY4xv5B8y2/hSjx1xsmK8rssoMyNYGKKUVL705hWNVfupomVOLQ
BBDTMdk6B2AeK9c/ukMHDN2BwnM5QSwjWU854+AioKAv6IAH4tppzRmXmN0EGY0BP5yrGA1JJoK9
NKJL3Aiy5n8BQES0V/o0wpZpInNnOsQkc3dFPw8kRybvqjfZ5IQ+Iw0x3sR1J3NMUY21brVMbui/
GPzGfQNORySOK4i5vH9roZy8yBaSvVzUBuA9MBGnafrrphmtg8VRAjDR6Vejqvjf9SsgHbBQj8HR
blS0C6/7salR/soeWFbe/YWb3q85IxH+4tkrDc8rwKGDiiZz+nVPaEqHctVxJjEtIJBCX3Viwfxt
GiMSbpbCfKLvEW1KaYEk59FkREoMNETaX12yXlBCF7gdIgS8Muk24eVBPB584nm9JlIl0TtHceow
KYakoCMzGl+D7+m1UCwviYct7rraMadpT1VsN2jykO2VyUu27w7ii79/bytlIqEOYJhMYOdRwrxB
nfuJp4kFUP1o4cE2tZVpT24B6I5PnHrryFesCyz5kO4dZNNbNejhpj6ZIkVh1Hfbg2N8jOfBm6Jc
WoP5Z9sJwwYZdpg/DlDkQDXDwTV+kUi3lmevmIfbRn6A06CGJt4kfGn2KHfvkY8cqorCb1RpnAhn
KdW+VaobHY003X7n4xkClikIwOJFaoH12qQZnWpWNvqsFXjI4Bc3zX1MkFJw/+ZaIm9ov0KG+1Sv
XMwKGsZR76wRARyabuq/netxqXktrjnlcLQmx21zP79ktlnGgtocqMvsPotlFPd/Vh18SHszcH1W
7bnlT4883G3beGFfNImjjgccdR967AvOtF08s6s51FBXhM8LpGz/2dIayLvZ3on+B5ebO+8+PaCJ
X3A9tWqW8+I3r8h1d4t7AnM1HuDxZkz/MVHVWdruzymL514OY/2mD856oRJ4G2vQmsHbo0wyTS72
krmFCS5hVG7boLguJXQ/TMu8PQqudh/Dlt87VJF9geG0omtqPG7+ptlaoj5RE59Ta57Si6oXl8il
GJcSov8jQetMwUxaN0sREcIkGlIy/u7BdBVwxdXOf7k6xl27unRZo9iLh4wlFJs7Uo6vsuyShz04
oIMz0gLSCGZCo5fbx1iWPMuIfls0mIu1fPvozzGKRX5syKcKRnLHyW1OV0ONcWZlMMevUqlIGVB8
ou0tJajl4TTYj78TyctHPVAM3r5WbemOa072qpGcSpcCdUfBeGSWSgnrmoEk5YJ4yOppXBd3FVhY
8A7kizQDyJZX9FQDHV7K6oVC6eZlfZZpUvjGBhhscDsIqqGEJl7oc4oRRNoaVZjeOGW6c/i0PtQ0
HM4bytlmrhgMmXIo95RwqxdfhMrMnA9SRymxxwDsnE/Ya3BDffUzz2ajpFm06xDjdUs1kvQLR0CN
oDQqdr3kePUiJ+tlb8ZnbJTGTaPvyTq5A/7Iz9ZRK7X1q6y+Egk0GJrorhQDGYI9kjGPQCFo74wz
m4T4W0x/vWjprg1b40tjFRkpbriXwpHV7RH712At3mKabXAfsDwYxLR5plu8PMIOQhnQs6f1SUal
HsVXi1pVi4+4Dg9G+Pv4DsMI+cZY1J4Ryo1aLVjNuMtsFZxCH/IS4aocLQ1FtWmnSthRWlychrXg
XImcYkFFpg11AKyVH5j76+eiDE9IzPWYoZ4hw/T4dzKv9c9vPSTj6+gfjhLGZ02LH9KdU+5y5oHQ
8ZpkGK1BsVTdJuHOWKUV3t9AMMjSb27IvoMwFRo6qduad+SOoKX7AZrAyXU9xHu829eUPxPR4lsP
IwImOFs1CfrxJeDd9jjJivpogpyqCDGV75rG1fC0p9moGBkaQ8KlLkl7tq7ekZnqKXB8p4zQb8/E
DA1d5nGFY2twjKs5cf2Zz8cvArHCr35/0wVZ8I2Ovks5tkOZe/VPGCC86P7tsNOOQDObNN2276mC
jhRbeO7q6kaLtYUQ/d1h7y9ASjwjhNKAHp99ZywElrZAwhIX++nsyG1ufZEVhk3AFqnVBUQqFmnR
IB4OCaM0EwVHcig0dhoVapvRqTCppOVMhY3Zy4Jg9zEn5Og326HRQxNzVkFIbmENLHIkssxFL7Du
g1TWEcS+RV6WfMcDqBu13L4rtPk6ZRAM0TSYTlEMchvPcEayVXaHbvWP3bwTqUeiPc3P6Y3RVwoy
XqGrxJZstmxB6G0oUpIk5lqFsMO8IqLNIYuLw3MALoEdsOY0ckVmO/vZ5YdIFr01PoeJG4RXTTt6
D1acoJrDZx9IGMWUa4pr3cGV7oCVJE3p4QBpc4YUQYMC1M2p1NYghxOg/gf3oxMrIx7fwYorygXf
ctbOkD/qPdSJcr3MFAFMjYlXZSeKoAaCXCL2y6OSlQ9kszavlsFpt6KZ1GLC8rPrFBHfPleer7pH
WlyXvTbnqaQkExRTlWfhXLcRXaYo6AjVbX7HH/n6YSqQtikAAh1yM1YDWNo/IEuLFcFvBickoRtQ
FP0emNxzN7XEq+P5kYUbLFHGcriTA3YEUa2rEDj0B+QDUOXbwPq15XC3JVgUOudnsM704MI9WRWb
dvYExOGZGsZik+jKQOoM1li1PiIFvYo1fSrxfQeg9fjaXkz0Az13FX8JPD5R2HWpF5zXxeevYrEZ
q7yU4+LxncIJgQ0ppnqWLFucwuaKJOvIysP7d1tuTBFzd2ySi7aEbZjz4mnZ9BbpCfpuVPk21Oqw
xVS9V0Tz0HwJgcA3QD2fCUN0jRCgfWmEiKP7nbB+b0ky4M5MRYck7CFSUjDenp78FIxJycfM1PSP
tdNG+vRMTn6SdP6CKzOqIdhPPxI6oipY8EZywo+aFeBRpkGDsTfSm94KU9t51c8Fbn28QJFJM8ee
UXOj/o5Coo1l50gxGipMs7SkGR9hDsM3grQLdFQJJi1izu7ZojGWDCFDmt2Md1udVrvDbGbErE+y
ZNtN/fiQ0uaiojaUHOtiFCifScW2XOWULweK3Ch4Na7V5k+3Sk7/MOdH1U6SAOkIt2aqMSVk22Bo
niV1zaw9BmFskO/6Q52nnGrDmY6BxiEow0Mvb6w6vvcwXkG8tNEdYWijlglk6B2EN4V6b9uxTPCw
KeXhCUTGomtBkiijItxa9gMCtquELty521J4Yi4k52+3Mxf2h92soQ4Bw7w3Zo6Njy3TXs4Tygaf
Jam+Wz30OPmL6Wue7wxnEEJSF0iIVGpm8r5WcNOKCAhNh9jeuXRZ8BosgbjywU4QrtqbtsRDCgFf
Zv6Up/Nphio8Bhfp7XtArTCj51ojP8p/jse5M6qYXPGmMZOSqoLW46LLESK9ra3yFolL2tTIc+H3
Jm6WQiv8ypv2+koWw+M68RDm72SrdwldFihUcTGgh5GgGxE/i1NKfbKCCL373y5Ltdu2pN/zrebQ
kcEkVs8m6Iftu08rIpHTtmJenprNc49+vVu0tJfW7bGjVfLZ3JsIYJh1Uc9L6nV96pkFPd4ylHUh
rqQcXAkAG0DEy43XGLZe1FrF6pcy/blUlD0604/e/6dPI+VbxwMkdcH+wfRKnXrSsMTLI6KhUaBi
u2eIVtWkFzdfkjKBQjB2hkPNq2w6ukfINuNY6EHwvhyuslrBkIRUXdLqDIpy2JgpNMwON3dR0CT6
v38qUq6pKFVKK/mZH6mNK5zmLEREjqUpR/taaCJ8GcBM2ZUEeo1d34BvD2Y8TiscWo0SbqvjTzbX
3xa/RvBaLhdzyzH7+AriY7kx3msb0q0GkWgYZ9Wbtsu1GkWV+xLbjClgnlyHMeA1XebLkWA8ONM0
e5woP3qZmfMCnuQ/VNgy26YjWtqqVGSoOR4b7YvpYE74J2w2v8AtAtYyx7KSZAQKgLzZ1ZLXyxDo
EB7rbYtRDy7El4uQE8M03mjFwvkVecIbTyPSgebTSPw7KnzWu45XpG6G3TkE4XJyDzv1AuriCzxz
onU8ZChcacd5L1uXZoxGwFuLGO+AJnOUsA++SfeHpPB9xMUV6fMyYzrqFrQx0ptoXUokJXvx1Nbc
KSR/ugfx58BoZk4hruQ/PSD47oDl4YUg+hSmn7CFc0czYc+vG3vN4poftfCt7dApymha3RU5tHCv
n6O3258abt0IktirmYNuwyREf7xo2Lg9X2tzLwQVh24l/Qc9tzDIv65zK0E8+A5SfcGPOg6NfJNr
5L+jOGPpbw2tddxfVxBo0TXnCkOkJz7Qx0bBzUNkzSEBFRQyyDeHTdfT3MvX3VTpvfa9oAId1jV8
ZPKHgEZb3dvVoUIPXdBRIApTIt4EnMBMD+2vhOo5k9rNQkTjgg5Cm60bjiWtL/XO1s/Bhs3oNIn+
TsZBmcHYgqOi41IWO6GNu+/LVGWY1sArzPLBcLyGCy6Ise9lpcgzUk0UOQrG7Zqj5Adi5X///EbV
6Xu4xkXb11vU5p0+m9XECN6ZPUhyuI1Lpw4gj7MBIlqe0cpaaIXNCPrfVHXM5b3RNR2o6ETZZBmF
j4Pz82YEXP8Jl+OizGTyCMrOEBsd6OahvXIHKVL3di1LVVKqqJYMNNT9cKFXyHcS++dkkAZdIE6d
Wfa06nuSvgJ5qkidJNPgLKAILMUnk5v3Q97l3Wvt9fVjJ4mfx0QujTWlEUvAUGYROArUD7Ljk+f1
BOd3BChFXrP/KLEX6VOg7bczGJxWAxlt5m1au/xacH6kzGawOKVBn8FQgki5TBAPMTXvVSULpFk4
pJzWHeHl9XAfCzGSQ49JjFcERf1wq+0D7RACxSEuv+K30tpdUM41595QqiBeRdF7RjONuf/MkJFT
lgSHAZMIHJaEBbr6Z4AoSpvAKTxts9UcAXLqal7YNDISmB7BGjDZbtaAOo9rraCn4hNfweuXsPF1
YknP8HsTE1638S+xNoZd9yvxhW+3zOI/M+K9yqz9XVM+KJvTX5pKIud3o0id1AHljAgR4SvSi3ML
OH3Tgo8GRn/9qj+gco7J0I+Jn3fzJo1xwrKYY+ISwPCGfshe2PRkWnPmFAbnec43uONHMNgSL0rC
Ztft0BWKXdbLy49cm/fgn108rkITS0ZrcgXRoQ7XydMJYWwj2nQ5TaPdgAmOViUoXwbmAjUZkHuk
JrO62YAH6EaXtgo7n7+MbzctiV/Jk8rQDN+edup6oSdwuq44bjOotMiPalYzQOIRp6DEfwBP0w8I
Dp5Z6Z2F/tJRD4vUUuzmTagU5PHQb5bYdiBs4GzPoqTldlPqr3vCL4oaR7cy1CehTM7+B6hl65bq
SNW2TzY/GAbmrt9IdsJYpyOMvpvad8HzICXhmWwbciRraWixq2X7RzYV1x9JEAnR1ACeT5T+gq30
lreZ7absibg8+mC4X4IuzrGOt7bmQiP7vm1zyqdgpXZJohOJxTcB2KexJbOoEooxzmQsXSHKBurM
GVvaW/EBiBpCdj9rnGervHm3y+cRjjeGxKSDkWmK1GcdFswy8FvvCeDhvrIB1aWZdH+eArBEIH64
8AZ98Fs3jwVzmeatEGT+RWonqOSLfBOEkvbI01e3uk1JbI6pwOiBL/4gZkill9YQYzLg54vzSrn2
WH/82FUYIOJPLe4WmB8pKxVRj0QZlRKZSMuyNJN2WwRXpUd4nlSJONzDw8Rau11JRr+qFnWXrSXH
Wp5aJAvw5BVH3yb4HpZDdv1zv6Eu7Qckli+DB0FKLA3/G5xG5e2nAoOh0UHgx0kzKuOvueNmlAV5
slL2uQwtwd6G2s6Fh+amJwNY+x73FokGtB9i3m7E0zV7oUc/Ukoohu84pqyI3hNwQh1U7367qLTy
Fz+Pmps8H9CxqpkE7H5aGHgcWYQnkSleWwzVolG8N+5rc6VbKIBfTwsl9tfMFx5kwnDHS/pZ08AS
fMnQY0QLSOo1qQJa838WjXTSdyKHTFLY42jOROnIeECn3Q1DXjtYBTfCzFG36hRQG2GhwxaTJWpL
RrwCt8gGKuq22rboLVeJZ+GgUaG2K/7Z+Xb7rCzzoYmAETqOzO6Iwl8cHLwZ9pLW69eVQ0IsU3Hk
a4I6JSHc2S8Ptm97wQUqPHOI0Jwn76EmdyhP3wXKRoahTBF8W+oBPnY0xaUi/Av6JLF/Vc7YAC6Q
6ro7mpjicKET4kiWBu3T7qxLZ8yp/LwUuIdJdGv1NIL0Cf9wUwxfUkDtlkxdnq4+KyDOd+QOPPYe
+lPKzN7lpu5qAG92sLCfV9BJbsTtm0NEK5NUstcgOYqqIrw5ZphlI2o0AhtS5Ax1Jp7Ze5nQtwe6
21zoP2dxOyR3X+xX3sls/W6Lph7SNsTsrLP6/yRIzHIxi3nmJBHi+RGJtlDeX+X3EJtW0pB940YM
i19zWyKwLA7hUNoHV1JELnoaxVmwdWjUFbCi8bUbPGqx96lq/HYZFKb+C37qHunyfhhIQHqtT5Bx
Kk6r3Ve+wUNuSInJ6CP4RQCKMf0RHUzTwFFb/P+nk7Vj593fMJodN9LyoTeq3ebI8VMki71Li2IA
rtTXsWYO5M2nMq50DLhThqCoeao5gNT33TAKZScuL/wVdlwMZgrD7mgPA5/dY6NVvGAfYXnGZJ9X
Gbmt1mSDKnkmABYjv9XzJ75rdZFwmNE4R6ceT5Rx4JkLRrdZuq23sKR5vCLfLP6r/YG7NDU2eJrI
9ZJHSSPF301hOVVgCGgpLIDLtpiOdeKwLgC5IkQWNHXij9MsriHGEOOiJX5dCG1cZwHxogro0FTn
oS65lRj+DsaMLgjmw6A5cyo/ll07NtXot1mkcTmpD4Avzdc3ucW2znlvJhKXlVzn9PV522BS/jyq
RDrBf/rDT3P5M3HC+Nr7C+kbDc1h7f+msRRc3f1hFl4HbDCRU3up+qkiJ3j4uk4l7KkJibdCfNM2
rd72O302I6CCTJSYOCgbjpPar0qS3j5Qg/HQ2RVlamZ04+HDEXIu86aJLaGCV6u5tj+9vVn7lNiI
GsHVWbPfU2cnmWuPma77BZBtadow8Ow7J3Q3pwW4axZcC//xNXa1r4o/Ppob6qR5b6wDBqDpnLAz
a9Zw4tKacV3cwcFNsdtG0zsH5CKUxyeUnoV+yWuqbEIkC/LGpP3C4mxouvM8kNyDQxPJzVCj/0ib
WrfzuPWED6o0AVgo9racI3jCdAwfwWp0TtNURJaNTwHeIreIPiXFJ6wHz8VFsZPi4VeFaan9XnwK
VygrJpkZpF8gq1AuzIByqHxKYjbDxPwenrhqF3vv6cKf1f0MsZWBmg1LLIdvyaN9S7Rn7RCyfK+e
UlKjBtM6J1EEvAYULvJwIrja9O3JRwIya16Va/CdTmBHAdnb27CiOwvciEl68h3z6ORRAQQROd0c
C3E5iCTpI3qSo+Am/rlCKz2SnNnOnMGhzQAWjYpVsWoBvCT7aZLFn8+NcxYx5yZwxxzvi7J2HTTM
OXxookW8IZoxzysXbOEEKO6oQOFGCtMejUsysFt5gXsiCEilH83xlEn1dNn2gxvYn86rNWyczsK9
B6n1TNzAvnP9AI869GKett+6H7ZK5gCwCwPtTumEtny6UfPx+ZvNm/sdi0NA5ZZDINielbmWnSH6
qeZBxEhO+ibGYBv53tcPaU86nv4g3YojUTY7PwCvpYpZFaXhPQOtaqCKlADaRLLw6QvGUJENi2IS
KGRjVVNrMWTvz5OkBhDvaiEkCXIXVxO1tIsoo0fwZeVO4XVndB3guAevkMi5LHsPiT4iGzeMHhD3
IhYKDEAFJBi/Nhv+6s03uSRVHeZmErWoyvhTrJm/YWgcBCO8pstr+PA0qy2vSWyOio+jckUP+vUT
1kKVs7jRIWI9dDATFJg032wtCw/ZgWSBjwpyeMGSEFEljZkWWFsFD6STJwhTgRKprXYUwdfYdVTF
bZsjFMaV60Ueci08sPZMlzZi8z8ZgXZYSpRR49Bl9mGKhHbV+I0UN3TyMWq8LYxH3alNW+8X0Myl
cTW8we0u1Gp3rtqRbPMZ0OLv3Zopn8Ahpn58GiHn2iD4RBix945XX+G8uXTtX84Uh+Ay9prizfLZ
mD4uP4B0NXlgC5pPiWbfD6oV0dI1QWvydWanM2leqZAE/mENwjHyb2Hc+XUxzaBN6mDXQcihpxNq
7Xdl7KVObzD+guWYUA/uU24gkbdpFH2EQpoeOHpwWxJfL8tQYpHYXvNqEKt7J1fDQzXxcX+tyrwI
AbY167VkhOmoMbF/Vz+8s5UQ0YwhhpCnIRIBuNn1E+KxZ9RhPFqSxCRa/OzXL7C0ygceoN1W5Rtf
AuBT+WKfSEAFMpbMlUqmV6z9ZGuLcWd71CSnBNY3FVImJc2E9nRmt2udObkvYRTx/cgBon4c7XXk
haOaaESe6C2JID2mLlr/D7F4CPVDfQCQAZZMK76D8YeQ16SyXuS2Yisrmom0b5DEz0PFf3JD6m62
SPEwneYvpPkAwhJjAImc6x6i7NS/OeVLXEj4r5C3/nul5VJ2m2PiFplwrXdvsjE/V2gUvniwjXSU
zanenj55lRgZ+NcaWxOYhLKia6FZPoU6gYrZulyfmHXN38HGRiiV5n3Jceq7/5q2pOshNXoJ6ZH9
/QnvHOE1mMueI8LRNZyZWdOAPHlR9zN51ZjG9QZ+FwP+kVVE5nYDzrY26QhqakmfhmzhUNUGki6X
uFs8C8HYyG9CrABMc5C9dVoHe3QEDCGaifEE6lrhKHAi0zYacZepZmQIBcdPB6FnnSZEzqQwQH5O
dZhNdqJt+SZQ210rZqCV19kXqC9DfTirtp4X6vuskKqaPCTiBS9XiC53YjVIlSWoSkQIaJTNyEPN
w93w5/K/W82wMIMu1eL2hZ7epGjOcwU6tX4qt8gJrqfIYjUF79pkSdwE1Y85lITStg7Kly/b8Sum
HHR6SR+V5iJYOfE0aBQzKgQ5a3gCYR6pw8Zfxy9mH7eborjy0fMgcEiMqv2ieU1lWhUbY2WH8zIc
iPmp46b8vKkkknkw0IAAUWY6S+YSBrmdKEkVYF9sbpAKgvZsCOcl1Ki8txklRhUJPJtCROekbjDY
TkRFoRQJjda7Kr49ZiGXm43+26jmZy7WbNkfwcRB0uqR1T9bzmVRDnP/4VfkjekSiaOK3yImjtJ3
NiNQIsx9iCvIwBvpE3oOqyjvyLDZ+erF2JGrk06vy3uCOtoF4GVWvdsSqPMAvGbF5Bc3MEnkIC4q
rQ0RPGNMhAzKGbYzkE6R0SDuoJocnl3pSs5WED3G534gv3GGKIuC1CSW49WZ0pyDOSPvCHDU9u9X
oyOpaDdmVonkujloHb3ZpeSaavR/4DPxROCVx4mZU//F3bVMOFZ2NdC/nUYtfNzzCisdPe10Mkj9
kpkUdff11mihLd/EwMGSpkuoGMo4RKTgDK/BLV+MVp9KcHH71TWRJ6P/vAABdlkgeXEwBBHmExRL
5dG7AR6CuJoHcEQYM6aWDP1hAYrKUqcA7IY2luL+lL/p2Wh8uVysxhnM3JXokSuvxe7jmuJVJYET
wkOciOS/H7CHtifUUu32/sKo7kKz8xLmeg6qBDMEURdrcG3Tx3ql+odSFbu1lEbz32IulL7uQ/tn
HXkjvvwQEsYfNkMZ7lt7aX9SUDNcDqyE97qhDrbdm8z7wByiLqmQN/0nDDg+hc1gr1j3MJzsVAt5
hUcX8u5x/PzmWEXOo1TCr2B7364lM6uFnNgGntpe4WjOMRKvHlf6waH25KfmZX+6BgbYSgfYVCL/
yNpq6v5Moz49unUlWfMHeFwAl7pD+NZU73Cv+0k9AckJuGLp3OBbxlK5O6iP1Wg9fv9f7YBK1F+5
bZpDIwGe7MspZO9McNKmz03DONORidgb0R5VayTF0Na2DcOUCqMxdsB1qeFSqF2pT1gT5OafxsiG
/mFGMDDYz1a0EIAytN6gLbRwlmxOsEhYSUb69x6mpO6Gk7WCHRswkATFGIf3ChmLQfx0q75JMHtP
nYOvFNCQHjqo14lHkLMaXZHU0i8giyuIl/Ks52F0DWZxBnd5hDymplEYYPxRSoXTD4uizPsxiVlL
jYUNXi1MF9uuiL3xzw4NXvS1GwfBaBOFTP0vqPb3EHUDr0qCO0z6N140TcbVZeMSCeEn7PbNmBq+
2WiWhFB6sKMUeM7vP9WD4ZjFJtl4e5dFd8OemcK1rdnqX2sq0UlZpuWAKLXP7TbKHwIHNVptC80H
vjtQsuJbTNPe0l8JeZ8G/7szA16BZahqaBRFFosOMKMQcn+Ehc4TG9peQGi49ki85A9dJz+oGJV8
QZje04ztX+Km1/Ra9uozjHTc6WsvBVc+LCHs8/i59F2XOGBsZ+UKhioSs0U1bSlYTb6yrp0wc9BW
+8ppLVS/DiHOcdP+BUsaNN56wDxq5A8C+M4BJuMReywhhdJAv02rh4xLmosxuBl/JO57e9ppVA0q
fxythK2uWq1kNQv6/ENHVzwO55KuhauJoAuRwyUKjWmMaFte3j1+v1nCuiEJqGRLZDk9t5Q3T9XT
RBNo1+c8eI8Xf3TpH+fQAulEgfL4C2edylSxDWRGmlYnlcqptxz9dBFU0L/KGd1KsMfg54x0X0Sx
SjBwAbDyOkRss/QDtsNinRD8wjZEoreRfXYW0IqYimQ334LH3umxp39xSVOq+YF4VrBivnfwLfRO
wGBz12oJtwX4zJr/BKbxat70K1qHucQX2QIob8VefN9ZlAJLp4ExL4xKDswFD9BbIUkBc75rsE3f
nX0JrMTVThQwqbY0PkV/oto28FuXkwnRJmLfo7wo0mnMVExVfC4bFdrCLrKgbKJ0Epk9kV8KOd/n
vwqiudBtlE3ARrL9mLkz9MuBdYh0DYGKF1bhNhKJ4EbXF0mt0QNtlQ7/R0F5DaBTjOOhNSf81GN4
QkIASCahmpPf/PwlHzGPL9NmeYjGb/KuZVgeUk9/yihv8mV6/gKDOscvcqHJfrZwoXizJWaRq1ni
ZCkvFpW57V+K44JBfoq0T76Mv4Qx4wTcV+Z/asW3rEKMMpL5Lb33UY9OhMV7dNw6Vjh6V323mi41
xfeN1f+WSsUdu/9LLBWzDGJZepQikPC0V8Sp8aeH+p69gKky6aKDPCSjltHM+7vezC5pKOyRTDfW
eN+YvWksQRpGPscuqxnb8VPiFUfnK5eZLtJhoOw6zzxHXkX/ivcZ1UJBe3IZe2b0DfYRwEDUo50B
3ATwqBlcDdg47a/knQLgL/P3Jvpbv4lCBgx2w3AsGD+0eEQQkANevPcFZ77An9WFcRMreKXtAK3C
5zDc/YiOJN9nTZmU6EBYghHZW5jvpjZ+C3FXG0ZNzjrzgsUuSa5+Fv+eFM3G3NB8zBvEYbo+LDvo
WTYBKCSmlVMEWL2Rf9yBf2OgM0+Y4XyKGAaZ9UwQMrrjYpdvlRSpCIbB3BRuVR/ke/MujsbHFges
actMhgjccD+xpJ1yg1ggCI7fd9PT4QCw0CnyXYYWzau3VJ+6PkRDNmycgwHyrn16I68lclPZMnof
XWD3tuivv9QYFOSfrQLAathUjz4Wd7ylV6/PKr476XCm/c0w7Id6oV3ePFfZ2oqZZTibC8xubXSz
bCd5SqcRTstlDCyY0wQ0Jma21lIHnkFDQGikhoWEQHQ7+b8zAFQG5mUOAOOdvWkoba7ZKNUGP3Fr
II7nizTvq+W21hmGOzKqEroEG4C3/CUq6jyvvXXRLcNgk0NPBVSSnKl9rfbdEyGtb/K2VuTKwKho
uMqDlGReBYmL6AcYRr1DPy+VaojGk9TPlw7+hjyagP24JzYU2Z58uSDwE5iJTPKV6FyuSSV0QEFJ
ux5bF9FrLBZcQP1dahwXgNNGsSrSWhOzS0br0UXXpNRGsfr+OedVfOPgd7DuRuRYoUif3xOFzEUn
iX3c3jC6YlPk2pQniGbQsGy/maOXjDLtZPvKBCgRkdHKuX7LDsBrBM05N9Ej96Pwiw/0IpdJIcD4
4TSJKVQWEiKCrPgE52uggGX3aejXCfVqvdhmEpdc5sKLhvZv9OfuAXtw1MnXkUXMiuKdnMGGVmez
L2rM6A/8mTobym5XQDeMbrzQVOtbrlc4vBp0j6gKcsGMUTntuzPcmB8cJiorujphWBQ21oqyBNCA
Vm1V2yrMRAfUCzfVZweFWkCV1sjSe1aJ1M63EV3W3La5q5YOUEXNryvdj17ZMP1kki3sZLzK+7aG
eBddILzzbwa1nWccVZBxIF2+KtBkjbUObi8tRald7HxD/8etey7q74SV1bZQUhFUJ1eUpYcXdo8Y
eoyMzawMn8QcewCut1n3kSFk5nDm0MZ8MV8gOB2GDPVYR0TMFDS8nMOE9U+NNvoqPyXBZhKyhrLK
Gl40Mg1odfsQjGseEZHfYr1f7iSlsCHP7u1tGuGgPMWhcfy2xa3M/2jDZK6i3gYc+wwuR3d54Oqy
yo7XvXiYgYO/gkq2jb2y+IaLQY1FDBWuuE/erBzelFUlYqAXjtSHtVrePaR0YXAOEgNZMkHoaZ+O
P/Pw+RcZzWKPH9ecnRSBSyEHpDf0ajut4ARJT4xV+rjFOloYiQIwHd+isFctqa9BHBrrnjSebPuZ
ziD3uhikRQIWCgXzs3JpJq/slNNjt0piCbr88s+DiJo+kgfYlR4zhQm7APxfCvxKMyhetFTnvGsb
Vt7YogE49VzcIVkf84Qn96tfApeCg4sWXRlSKyho+SV5RFIm7EHOH23n16KuntgytmrQYOASGlAe
JfMou/xWtYkE3DsawSvfQmc/iJzu2dNPCkiyR4zUOsWAuMhI6EOOiFsSl4xRWd6RH9FaLUP0cedz
bA5CUsUT5LkedtK24mZml0DgrI3PZlReDp5qA90rYIsmG38ANkuQI3S+MTtAbIxpW0RPPDVbgP6n
wUaLwI/Zzy5f93/PpyCPw5t7hgfl0Me/SR+Zw1Ko7tXqBFKnHQvzdgLPqK0wXfi1GHSEqRoizsgY
PE3OLxBA+61FpMeMBWr7xHiLbQvivHA/8gGKos2I6Or+PLFTggrRbQKuzOQEcUijAYxJEydFkRG5
LkNBw0rDW+IDIm8AKHJUArBmWXeGV1jzlkLURl2NSnBsZT+6WlA/g58L/IEoYoAXIwWMU7OJk+wN
cRc+xCjHnqBruNzgaaDE1mvAGTzqEo9+/g9U8XVxkK6ZE2bzqmVdmr/hR0artQWBk8Cra5kj3jlb
mzpTxwtUcApDeVmoGC5gEHT2h6caVaPmxGnGDyOYK8/CoKR7eHey1NRETxw0xZ8hEy8OHxfUrJ1/
bWhHpsj1crhT1u9uY04ME3uzNmbhxwbZjTOB1SX4RM90SItjfpOvZea1s3weNiXZcG3NjQt+YDYJ
iQxB72UmWxyDXCTHeLjjFV8+jq8IlG0X9FMQNQINwxqwtj4kbZu/9BOIkqpePZaQQ4hdPkZzvS8e
Bm4pAF9hljxBPFBuvnX7yuUifi+vICPYnKRfZT/yZ3YgnQxvfLl7xe5s/r/9zwPcRfsmdw98XwgK
GZioaZSnYJeSNG1BeMOfDSHpA0ilw1DFU0OWuRCSAi/7s45kMa4C2KMVMdHISFP9pNax//ekBuJC
qFc6yzUn3mfkVNawZ4plSOOk+NEJjGHtUs8JBH4RFZCc6IBxaZ7/TH7gdJsIeR21ONpRKZhyWVd+
j4pN3ohLPU64bcnpsmazJMw8yzEpiN+iRl63gQlJ7Kbmpgo/oiXII6cHZBB50BKKZFTzhLeh/Fxb
qKuFPCJ8mnp/j5H6FAVZQdlb5ZsuMPU0Z2MBMLL5FDuHRXbyBHbcNvsMfkPVy/gs6UUOH7rL7JyN
xY7nzq41BDnNdiNgAOIh7lWLekMVi+ZHW4uUix5g3yfKuqRfN7jNEjDc16SNz/tzMJ0j1NgjDtPe
Chw4zniOXplKFUi1ZmhFzhhQ/agqQ/hnM+WYDXn13c+8cBr5mpxEPvm+/XiWsNZy+zwpybHZJ4U+
iHqyx4Q/H/0Ay0pZ7wOqJ1Srda4OeEdOptAMrAcdNdYJV4NKjLeMGa2Epl6jGtcy1caXDn00dHWx
bHGgo/mug+NgvuSQFQ7QTXTvdrNKdjdmB111hV6LSd5GLZmVuiwVhjg6aRPLpju3fk0W9eUhLJ0h
nmRxknangfUw9I/PElsT9ZgO7tkwcTR2hHfC/bJQk9jp99t3HECb+vv+D2f7R3VDgRvJajg5EF4e
67e/AIisWQLXBS4hfaMC/Mw2hFg97/31FE1nSoekeIBHSE/wHj4JXZ4NEBQq8V0ONAuvaw859xGH
kZ9NGZyVYZKxLbPdkmdoa/O2jCraqJtlYWybHGorsjVPqVLw67zkTqwlkAMXdt9r3CxbozguRM4n
zWsIlpjcghtmo36dQPTpMoS+VgYdIkWJOHhf8gwB/Ezo/IKxSGzdcGJ4xhtrEuGYmHd94/fHbDIe
Q9lbTWGl/GqUFMtl8jU7DKT+R5+hzDqR0bQLX9JpijvQEIO3h/nQzib4mB1eK6p06c6Rp1pd4kSm
spRlIoFH1DXF9BKODFl3Pk/QRphSvJV5ZeOJaADDzLqXh8o9hhabBXh42jq/w9IlZDQAyPwVIUA7
rB/gE659RP+2F15fg1q0U1L8gUEXBlkqIBRVPHsrI/RdD6N2YQvfdsVmZo7l1Sg/UEPUKbn+qXi3
faqltcSjudPwHd42bIUduylP7amHJpVxzCCAoqNKFhBpRw8IZbV0SGK2KAPasArq4IrGu0vXTGO0
B26vD8UVKNqYB20VqpN1uFfboeuLYZwL2tnm8Xm42nLSY/yn9iWvj/eg5IAL8o21Hyi9ZO2+XMhF
9blspz1IARB12c8VzcvsMjAqkkQKcM7Uj4iH2YoeYGeQNfqyj1Nx1AQOeaQNikPl0L1Aykx/WWif
iPFp0BnZIRFAv8TLq/VU+0STmAIACEkoBzuPAEV/ZqhquOAx9VuBhM8Ub/e55Zv4efgHxkfnKkSi
pob0mDPSOL8G39moe/thJ8Bghx3perSc91bcAByygk9yhy/wt9t6OtHPD+k+tqQD35gFKbqRBySQ
V0D7mLi29MoUjm3LhE1bKdAblD9455knxVVG+tnXshyMpLlTcAHWM3GISgv4kjZVwsaeNejyMreR
PZ+vOdgdnicZ9Zncb6ajwQSKM6mM2XgYkRPl7tG49y5Y72PInHqqJgOhXYmEuLYA3Jo8K10nXmgD
ib2SW6fVrFqsgYmXIZ3l0Hl8v/JQNpqvlBw+T1F3UIUM0fz8xGWdMlgfxScriaGEEBghKgjMg4Bs
7+hMJEZr7Jv71fHPMGKPK5mBKZVpSNPDYZG6aHR3T5M4LQJHsA1Qov6ZEBldVjUHHo60TTDEHEey
XGPL/X3YlRxcJmG5/IjEojwIchQnycQ5EsAu0eU8ksxITA8l/HZkEUqduPZ2EBpLKHHgBEX+MAeT
y0VzlXat1ucg46/AsVFw3ezR1GpjhEXhqnhCRcxS+zsLAl5YzZlRE84KGh4WWaAdsgiitf/mXKsA
wW8bfhcZpklKTpKfaud1/VZQsv/Q7alvC2fMHfU0UzCuL3Od1UJaSvT3qSOCilC1lnwlAb6iFZv1
mkCsY0Kt500TPJZhqnjsT/7X25BKyyR74ebhz4hPfYXaVbw+Oi8xFguXA9hTe8o84q8AqqcNETT2
A/C51MgUcd4hFLfiFbeqdc+nKBid8jF5dQ8JUq6RtwrHEcjQesZwh6YuSo1+sEe1ukhTASEr40CM
f9BFB3QbR3WtXIjlB0kHTjlfUiojhUafnZalaPhBB5QCmgRgvbCPZfkWoYpV6ZV/Ibd1V3j4kQRb
7YzPFL0lPOLsq5QneOtsHEEvvRoEPIjnYdPsXk4+uZCxNAN/SrOwN4S32dL127sOSDZN5pR7Vkwx
e/raWn5JIJziXFTCjYV3PjhaXpAOpCIYQSKzzcpi/jj9Enn/MBCld1hgN3XDqPE9qQEz2qKkEplu
qmBZkJZZ0nWXLAheJ5lHWMlTSrpmidyeaEEugN8UGQe6ri+8FbhuQhyrXOwvf8DcyVXz827OrKML
Sri1wtkGF2K92dGFnDOt5EQBlLMwgD7+QYOo+E3iNrKjypLWipH2iN+8zgQ4QdI6VDTNRCKSEA8q
d5ebMfApjjYtoSocrjZHAVQbJYsEDpLuxmE7lD4nkUD+dkwN1n1sdmFvZR7k9oFtadHSlk9LCpZJ
wbobqEqOeavRDBRrSon1epS620rbdI6+iT9qe50d2no+sR0Z1srsOYfmXXMIG9o1MBtnmsNm2fLK
K653UwO1QRZ7xT13OB0RsQvWihgCiGCIlJOktp0aP1tParKNSQkrN75Vwv/PWT0dKsPU1eKPHtWe
liXCCMVj9nfjRpdpxXPG5HwcY7OmqcvCnZQK5Q7a88SWeh/TNsSx4/aap0j0Y5rd+vRfBJk2rsmI
Ppao+LmwyXNxD/ajKA2xflw/5xm2AapDAm5OOrVh4jLAvKXz98oK2q3KSqZ5qYAuG50Xw5hvbGQA
WoAYtSv9MDpFh8djDJVShTkUPKOfHcnE69qrpZGRvobqctCiZvMk8qVHYpX7HeO+wD5Oxsa6iGPN
7JK+EhWogzjzIvwj+1hAbGPD6T/FzCeVp+6FyRsTqCynZxZTBET5h6pkrX5h34nuL1supbWzQn+9
1SeygIMUJqHd5z2rMn3Aty0jOyMwBWaAxanUSsfZPxSTajn5ut0l9JbwZP8uJZThXYBLlmq1k8+G
vtHXuv97LAnXfHO8vti1Avlt3FJBGEJ0k/sq/TSRM2crAp1cAQpZwiKAlukiu8Lricz5HTz3V8XP
v75q4BnYyf3vNOWXFJAQ0g9bUGEuubG4hYGlYuYU7ySrD1MD8Vq+INNdGC7koyIoZ1mmtOj3rV+J
Aah8iXoErSJ2a+Pv0rnu0Bqm1EJnGzFXfSRepg7d+ZMfH1hY7SFQWCmbWc5QFZxiZtB6Z26/xNtx
6Qb+g/1l0uUHYcVfGQnmdDHOeq5rwwqtB56YY/jhkgfZOMEr2WxHrEieuuwRVu3mWxdxKxH7z+5Y
nQUAUed1D1kNl+Qu2DUt1IEhJJwophgnnrI63IyFRTDyQFHn7jqOxbeWZQnF3qqb7YpVLaHu/gjz
4WCW/VLfyxku1Pl4y3W1xxy15uiuTHh4kennFCwLC2FrQm95mAcVwi/LD2n2T1WRRPlFN10C7dEr
5/GJ22OA0yFDsAT2PgsCCGNpfws9r87+cFEXHM0EfID/mIkOVl1gd5Cwhe4LdMgpXO8+3MJI8qUV
pzg2J5BMx2U7RG8CsG+dJUTnJyVK+c/IYsXhEOzksyoI0nDqssFhrtqttgaacCMUoQtN0BWf1z3w
x7AK4Z5skGTSnwBU5Ovn5kjz+uUhZfIuDrBye3zuWOM15ZOTenB0zjFWnoU9XnjB49o+zweLIynJ
6pnq63jQEoFZuSYPwNvw0kPYZyiPoWzUMQ1M+dmJBaEfFE4QChCGS7rpgMYxCI7wT2Ac+3JjrCCv
p7Ru6QYk+bBUnev3F0yMRulCeixmT189zcyT5m94ZoT6uhLXcknv7dJYYDxWC5yQV+59UHu//GRQ
G97rhjmLv+Xw6JSdLh6sXBCg3mQE10xD/xmnQBfokcRMDXXkOYr/6lut0srjEipKI3m+GExLyo+f
ssKgEQSlpNaPZL4H8rTOeVsC0btrvUVy5xOERX8FgW5/SwcJZAygmyLs6FzF8Q6lHVCXjsypLQ8S
d3AbQ1rePliZh2dSdkDulbuV25jnlI6/erQU743HT0H35smxvEPKSpUBE1lZ9XP8HvttD/2CIDPI
0hNAYL01ohkSKRdWoTD43+UyMxP/86tMgylqcu0LvulyeX4iqBFu4xEzl5fMdpWxiQzFb2tDW7cP
YmsP/+u1Odh485drkGnxF86VagwYXzm/BQon3fo+OZM6ob/sY7O63oVeSWlr+Y/T6wLBOVGfrBwO
3WqGibQkAu6Z2bUMxsrfNR7NFxgw+dCl0BfPBx3P77mSZoggpPJNAPDNs5rQm4DiLqdfER8+y382
f3BsK6VHqaLaEnm0+DQL/rlQM+qmuOEOvhBiPmAPp4Qlaw88WBKD0FHG5NrhbgYVWr8GtnCG+/lH
oH6EsuZO0VvRUNVxZxNGpSauVFTIoChWsNI3eDTs45Kc3bI+kSvh1+cjCsx++it6D4kZMqR3eflp
LSQp2mFs6cZYWpTWBUC8onAvb4h4JqTH/biV9e93V+wU+yl9t6ZjWX/yziCZQyehlQ3eMRDQQ/As
RR2CSsQmNGh8+t/V5MT0Z68zBwoJrRkoKJNtMEqDRRWcZMhaK0dmG2bbL7aUVjVbwDj1CFyqQmdU
uGpx/abqckBjBGT6hEDMcKopttbG3wwhJO7tCCunwor654/Bo6wPnoPuJymp6lZAF3ANTck/N5o6
ndui9K6XwfN6UnFXfEj1URt9af+zl40VmRUMyq3a1E9Dp3kGNE+aTXK0C4nFzMyi0Vw8GVvXmR+1
NrKbRY361JEiloY5GYJyXsLv4hz29KEFuxuVrtn5YPym2v27qqsFS/gvWgOKDcH2eOxxRX2J36eQ
RTy2A/jRapj7ixKa6aKTMCH8uTyMhcXJS22F9mFynreFkJYUlyoekTIg/LiKInuENhfoErh+03ew
awwtlvKItTGRUZ8HtM2RAz9lzEa1UMkwUHYbhrdEEuphnlbgtNA+wH5bMv4f2xErLqHBmDeTx4Jk
8shgK2Ta+TosVWHG17lVFlCsvG6EyLnbuP1g3/err6HBVfHYLpl2WRpfGL/9VEYntr69m1RiV3MA
O/6IjxrvItuXRW5ExblsdwIngtjn+MCVcV7Y12ASKPMTB00sE4Os8SBVOcZb+FvktzfdwoR2gyvW
dziE9F3YaKt2vbyzyzJrCGqnmH+8W/NSjnePxrBU6sq+8j+NGnu6o1491KzPXQ5DApn6lkgvzNqD
P0H78ieWqEJDzMxrgPmkciZIpE23ebUAELdPl0JlJkRjjNT8/BhD77pFHNgNQFr61yLgPSe/Lxy2
xPYOENyaogU6GDtbrLInM2mjh/H0FgUeUZfv41wy/PVAwTtR5hI2TjpxjMfG1WZg8fce6n/TpvUA
XNOMLgToMmv2hADfRPLzXpyUGpKuZgkbNmWG9b8jC5Z2f7RQekL/crxfVWHhnRbUYASOPIXQimxc
YyhjWz+tbovm0P/k/hTpShvKa7Rn8XkpL4NT3NX71n8+tfk59MD8PgK0IwHOqsKAOIY0ZC/b6gil
CabYjqlydVprgReypiWpCiZ4I7v0CKxB+IN1wzZ/z7ONSIw/Azf4fpUeJb3+Czp/Xe10CTgZxbrm
CQsk6v/8puiYpFQtzfO9BD7ssWELMGDOG7ec5f7rNViCVOVWc472HF0tS0+tT8TFkL42hPOImmLF
dMFAqKH8B0+9dVbIOTbX1mOJ/Y2f9uk0wOZX7WlOr3wFmmn9w3Cg4nyzUilDttmwa79zESOlWlCp
2H3Oz+jG9bwrJT2ELyKhfy2H5tjHsWsVS6lOAR7LNVjVMn2V0YzHvhZm98vn6ujJr2q+7B0bzsBG
5R85aTjkOhiKlnuCKgxG/CxS/l38NaEbdeiHoxRU8rGv6/7GLXiypnyIbHZLLOW+o8eHA2JBugzL
wnoe/1LC+VrN/pPcslc3ltPqGELOLjPZp/xSin1cdOo4jW2Rw1aNAnUDQqSk3plGAtYGMjEL2pI2
h1g3fTUk+lDPFQ/UZBjReg8dhvSN8GxwpJu4tC4Nb0gZLvBCByAV9sFV5d10ucG6qhMg8noEJjyU
596nYYHGNCI1V0E9MVpvOAlUxmJQkVX3KiUP/BemOR9IvKKtGWAO22F6HujSFXqoMFMUMxzqn1rT
SfFEOlWCYe4/MxHaCo2JnWaH5JktP73nfN9ku1mKly8FaOmeZEFxAtiI9gBgxV71qxo4D5UiZxa6
J8uYRf3htu/i2G9BIVvhwq6jNBSHNOkczkFNkQfXY/LDmCSMVq1bLL5MIg4dFAivz7AA+hFhVbZy
LcO3oNx3vunavBNjUohuWIzlkw6Okr7NNnnRt7pifOG2t0ViavL8iE9UjlTWzyvsiwnTg2y5GdDG
/NphQxlIFzoYcBPLkMUEvdtJSCD1DB+2QZEmuLjd7hB28vRdcSlAvkr5qpsXX9dNp/6lawRDT6wr
QgdU8K30GkVQX5dNQYPHanI4n9HuIIcu9DLX2jNOALZVBqMdCk7mKsU7+ebNxgYCBt9+wTbsJ1g1
VV6jsuwpG4wezA5IRb8QJEsqlFxNvjy9rFiTZzrx2hGeUawv8Nq9mbnix7Ume6r9+6UP1nw45MCP
t6cf7s7PcEXigN5Qyy6fKRE096wxDeg6/66Ra4L2LWts/iILInxS/bvKRt4pBh9VB1CBOsta9+dk
gvNZBA2D1Zq+srSjNwjpFE4Ui22xbaUGDwR5EMOb94aglgwSshb3Myzsdkzc2eSERx0cpQd/ZmRz
ucrJhP9an/ulZtuEsRVS9b8V2IHFIeoyrvUKJ8rEFCNA1L5VElP+HElo7tbqA4KvQfei9MchN+uD
ufsA9z191P6jKIJuNcdjr5nbMjpnGasulriUWSSrKu6dTqqZz5G/QC9Uz3qtC+NLEESzxQ+zML/i
Vr/WbDMbshG5xaO45fqfDMD6rvxVc7C+tSOb7W6ePTmSLJqKPsJgTaiYH4Uh6wO+yrNNwJz6yJJ4
/hG3QbPrANwS1ZWAYW+Hv+2NE4u7L1HKf6E4b+9gAXlj3mOQ+8IVfveWG2Bn7cucbCLndbiDM94N
//S7K17z8aQuftLeR4ivhPAhTBTDiN1Qh2P8KMeRqfUS5/AEbiP/Plp5rhr7+Csrpw3jveyQtLah
xlfH3qUvWOnqtpGlyk/pd3kbDVhFESahd8guidGHRWfr7aI0XMP8k/PGev1SBKJpaaSmdEdpcirA
wQT763xnZoRY21fwXqvHAwwnwb7ZGx3zt14oInh3MQiupVE7/2EgzzuiQ5r/ELHIqiKPEOZBMOM6
twYrBG7hGWCft1gRUPCpbu1YEzzdkl9IiYi4BDMoL2KbI09P2+bGLuLAlhfOX+/UdaLNCwVv9cms
4HYQlxWJG5jDEWNk2mCb56Cn3TmDuNTGfTmw+Is2O6I0V0OMWWci2IdngXbQuoXwaEaguCZJ+biC
clpb4QGUty2FV6EM8eu8s8bpV7ZErBSpgSC2jahAZqRBqep6IdoPg1/+B8FRDN1jbWX7xiYEIZ6W
oLZr5956vogLQ7UKqsxmhw81gvfyd1JnTPN7TpfUWYqLmOGW9zgMUPnIVltZgKjdtHKwHqfJaeG9
mRlFg0v2s8RjVPEOPX6YKCWVuYuV/czAPDkfMtAlxfh0KdSVDe95KnFf9888Nyy9tlONCdhvH9Us
bdZx8g75+8MTPjol+/+iSMN3Hl7nW4Tyf2ootTp1CwFKBAm3CrZZ1K2NG9C5n4SCw4TIVY6BXK1f
wmZ1tM+lUncAMM0UZaCajwFiooWsvQOenz62Ge6BU6MEgwQrtYCLWeJNcONP2EpUB+HU2+C/4YRE
exhtUJiZCnTHY+CANzaqJfNsMvFAAzu72mmtL0Bo3AviJHSZN6OeSmhSHSrWtkObmUodPlxRU9eH
E+5FyNWEn2O5XyBu9mUe6HFewrlUVE66ZRVnpRT1DQLXoeRQok8EjKbi3qTXn2GOQTOED91F40Xs
UhEOKBAOfCEe4NxEzD1pvZUQYHvgNPcA3ny0U5R1IzeXa78aToaXhTD+nqD5uiQ7EoMFhN3k68Cf
WTxCBKS2R1zOD3q5kT6vJSx6gKiSqq6fhkmFaBO9oHxIFAnRmIZWe3Zy6vITA71gfxuAkY6wiaHL
TBSrzgbw5ZUU1lwZ9+mrF4aVW6VRhdbAS3dqG/UOPyckaPZmD1WSd+hCGXq/z6RVHWQQC7xNLwas
WBpJN8F+iEnJE42oDFfdxEZMBGZBsXqxEGQxqQwnyEkvH5q8DPUGFj/LcozgScdGy5wl4m3I/SBQ
4yVX8RPsBW97J/LlH5vBs8kVSZfeHo6MUjDGpPlMB9bKFNSsZwdid8CtGkzPjXWZ1YgpL+a0W/FW
2yUvAqs2IBK/LdD0A3FB67DWaegBJ2aGtkwvc8rkzf+KcN286/epxLmVRwhv1O4pgRQ4VE03KOld
0ealvX455UhIFnk965y0CKg/kbtY7Lt0lfQG3/vuzr2By/jldlccnnPmvqKfkd3ZyWQbF4/1NO5z
4fX+pJNSFoBvzDeumXP/dja5Ed2GmVXNl14XgYzIHkWtwKMsk/Ap1jh9vIDop0s2ubj2qTXZerZI
mZJ3cnGm9k8Jb7ZICrI7zdAIB16UcconwDPjmY1zTIF11UJcYEaG1j4NWeRjQESOvo0VLl//ol58
SEn8sEZvsGJCJxDznN5nHsm2qUFD5yB8P8KbApEt41HfTj6Sh3abRnR+0tbnPRNAcbcqQScId6z6
cnPrTTvYNmBtNcLd0qKbP+t5nv3HAC2ASCnf46YFHGtsNuGeVJKC2tM5opBgqz8t5tjBKZh1/RDD
lUkw4eZ+EfSdoLPh+HJWccObWVn91OgGzZ7lhZxPLU6QTS/IgWianmKP7HimSof+hbePextO1QHo
EC1s/OKuxaM/zFR+aCg3oiJP6mT40qgDxGmg5JwJLBSQmKDn2xN3n4fjb79eszz/zwSF3BYMwJbH
2+n8F9M38tQSvIydwNixm9VZjaqlnzqXj4tUpQzsLHKZxBfow5qIKAlpralQIXbBf8JgBVEs7czk
YGNV9+5Meo+SA4mDZqrDEEMJRjdlRmxuFFSmfAU0xvTA0cw615xrEbXazKVZFKRiObFZSikxRWS2
tvjm3wpkUOmQN3yklM9Tn28gg0GbeA5eOpdgI6L0u45RZpIfBE5p7WFNzYY45IZEl5bOSSqFsXZD
IdUKWlY89BH/+OohIjev3XDvsMz8l0zigvLWGnLtTUzK4F0nTuHkIuLCgb+XH9yWT9ZryS29Ym0p
Dd7kwc35eKZaLeVdJAmjBHa5NNImoRS2j7DLUFbocDQhoH2w+1W0HqeOzhLQJPTNtehK3dnXNOHq
afxHsBf4Q+52tVHdIn+2FNmEas1FXq/B3/CAJi2x7bFrZCJ1hLDxrP7DSCtfxGkRsUrjnbcoRr6o
zIeQJfvaqZ4bJimlxfHzNfSf6k5hEn530Kv33cBT64tLyiq4jgzsiimERHvRdCKyZrtVSCA7RPGV
sgmAgThZmCAyO8hUtbiAjQiYWfLCQuC27h0EBAKGMHuoxEL2z2HZ95JYFBxv9LZcpafOJ7JkPn9K
MY4cugfqUdlynxVinVsDu/dzVYy6R08KF0vr7lgoknRuAr9GlyN/aRnP15lskheXawTt1KJ6j2wo
A63aeSxO6THnFPLKUr68j/Ex9N8JV+DYF4OeRdi9Sbbp2I+kKJbIO28zIXbk3BNqQ4k5wwA9CzkK
QqBsh8Yt42x5XITVpPjvDRtSxrjl13jvXoVf48HsCryDHHKlSO6RPwM2ACZqCf39Q0aPtEGFuXls
934ZsxVeleEfao1ykJtC0/ubeQNGq++34s5N9VZOUvX+qnkmUT+wCsSWRyCJuoWk8iw8oq9Uxt7r
04FTSX6YUsSUM5K0W7cYOM0ubHus1AmQJYV/krvQrOc6TOYPgZyElQoDU93EdSgwDL86Kc17XYgi
TZaWI3bLClMe+IlB3OTXg6Cgc0u4XM7IugZt1NrRpwR+TWwfNzgI5ChgP7xchTbL7dP4qXyyaH4t
I0Ur0ZA395MeMg8iYgJjbsUUUL2uSQt1dM6r26fxA1S12zbARQmAMpWQWO/mO9h1KfRCnpX/dCjs
PLqY/kUcQVcUsrJNfj/Anln0RdWwqVUbE7yYsOWx3M8cPfyDEV04z9XLb7QHswTB8PaNXgxX8mbR
hNbqgd8SASDOVmGrEamaLx26OD/tIbrKoaAKI1K9axev6TRAzFgI90VJd+NDzLXMyac1pCwRoVuN
wcGJIqdIQhoRZ8SdH3NtkpNW+McYIxIX0wQzOPuOS1sJO8z5I8U1Ov5NNky4aK1ZRZHx/fDZ54yj
vmPoZH0Aoq9pqvY5rz5Po7bVraRKzdh6XruJc5IhP+N13E3gNAFDtrJqOQveLdFCGES2yQ1wHryI
MKJAYSqQ5ubEBkojlTr2QrqpLYgmPQngC9WI15F9d4kEhuU27wsDQVVvWay8u9ByjoALMCnqftld
LaczeFWD1Ym7pQz0OqRFtUNtn5rMS3/FuX3hAypA7WTN9EXYAHrcSdwHI0CKGtLP8K4kl8KMxaOa
c2x4e5hgKw/099vVYS04N4OO5WrGUT7D7g9anWgwhF084WOXgzLhL56kxRqS7AqIW37qOmCgjM5E
4xGQ1+lyblQljL0c7+M7FcVdFsPDxVxWTy3Hc3oA2kIKsyNQLaJUavdAQm/I643bgFoNqirMLHcC
oqpw4aUOkn3ehZ66IALMIvppPKF+WPzWclyyQZeZ0C4nwODuz7I2/R+WXTytGTFjVI2LD64BiuOa
4Jt9q87MsYj2nt4LBkVbtU8c3xI9pdgbx4lcQYF5knoq6q8w2CBz7f36tq5j8NsElLEicT32G9ir
XxscDjqdTK4M/2b10/vWstnHxrG3CRC0dLNoXu7HAP4J9uZ21xxLf9eoApYwuRes3keYoQslBjsQ
ecQeQuRFGDEWLEbpOo4fP3PqXw8X6NCZQBdnhez8R2GbLqqF+8F6B5hPKiJcJKyDRCKD3PK57iio
8jWAXFO7kCRpeqWxSsB1QYSECdrstmsR9DwBmteit4u/ptB3N0eQZT+Js2Yv58/qAVgxDN8JL3Ha
ZUTxwU2O6iSqiI2sRrQwBB1nVuncOfdxRb8nEkGV+KediVkRaIyeoDdGT8zPxxNgeQzNlzBHJYWh
TWDH02KgzPBW3wk+Kld1SuzVPJ4UdfwtfbhTKngPzIj6PQVoPTSRIdaXYmoqUgd6KgiKI5SOs9BW
+/nbHGpCHDkce0acziJCfgnmQ7lnX9tGWq3tPBdNOEG2xpN2mKalV/75k67GbRySE1dOoeFCe54Z
TgzvZsQaMnUxm6qG5JmIvI7MfeZWjUVX4QinuZjrP4vYIxbjoWDTGtDGjyHT0mQuVVKTz59JvKnC
pm7FikSBmZsxOxMi7fpomPxoqyHzPw9SklVm950gVBu1PRMuFyqkeZF4nYXgPYv+FHNI6XjeiKlC
JAU+jl2Oz54/8C0uNIW6I6ht94LGDumCDd1MCCRcIRn0pDMjJBDLk/ksqMlzfO05TqUsqo8vES5h
Wfn+MczxIWL1bdD/bp0CC9sOz66lU/r1ZjEdXzrlQqzm/yDJLRV381FwLUIJ2IOlhZRaWyJm9XDC
EztJEG9JWspckNnzRjtwqNJ+gslkWuSQ3Hd+vxE58zrXhTd5a0tAOq2mDFbxz3V8QNqS0XfJmTuP
J0sleW1MJtOoy0NrFs9CiI3atk2N7mKhmSl+wbIWUodAIUQBJNW+s3zxyR+qSJbkD5h838BfPL0u
8swV2S/WpL7zNVQ1rBjrtY0ekxBy1qROj5SgqxTWxO8lX3RSZNdCDqP5oRINheChadHiej6GBu83
st6gxrTckxOSjypT7owUxpM21RWWrkbJ1MOK0O4t/nT4HrtkEkiYibvf1vQoJAVLxs4UQs36peO7
A9kw0noMSBIO3mgd1kyjqB6CNaypZo4RroYEK2yDKHY4EzM2Ag95DXn2aXMMMEoUmW/lrPYzqA4c
VMSZ5JfcVisux+lpz6aoL86a3V3UI8kIUVXsKDfXK4vwG73Vau22bK5yQrQTWGa43zcnaRTLS84l
PPgRvD8fSXgmGygmLhrH+elBZMJmUbHOgWxjzI9pJnUtvLSJi3fglnYpQRm5kP4TteZxfnluDwcp
QX3EBMD8FzdZYyvLThAQD5Z5inv5CUItX8zYtf7AoMuSKc94xmUPSyq5XCyse3aQCmuOOxMTK0oG
BfpM5oJXULl3RRyD7vP1vOnZgqUGVDozmHUeG3NYgC1j99QY7vpjvcyLdasHnkcdBtSpd7shW972
jxvC2A6WYV/8UYORGllIP2i1NBDKVjVm4g3SAZF0gwAas2dbSkvMKAHCCH424ZXE+2/Gke0KbGdX
DgWqMDwQHzCWLq8BHyzrtlo8S8fEBqec2VX6WGcEVzsZ7FN0UcLVrU+ZTdPoZ7RY3w/kcTQwBI+q
FChsG81LFSDxF8wkzMyIo2E9MxNhhjI7jew1e/oEKWyH7lWAWqECcn8Uy99yeuIvvjZHM19ri9VB
hBzSPFDK9P0las3hZeIrsN5RpUgL86PVm9Xs1rPEudOk1R1vrC3M2w0q0A2rQ83AFQeIZT2PmYMp
f6CF0SGjKCTvKe6Tq8T9+fc4209I6YP4QgcBHk7H4s1jNeyL7YszMCJZQCoECW4D7iqscewy81lj
vBourXHySN6vh5PGfVILEwFrxVMp+YT6aanOGOPlzasXv6wgAeJRfQCIrHcE5QZPMj69uZe5sRO7
Rdms1NzZQNvv/JNVJbWOEb0hK69Gd1CNrIoyD4nFAgQXyh1KpQ+ZtBldSqw+wWn1sL2kZwblA2xx
YaK5ygXeTOwpAP8S+CwskIpbY5Jx03ijycNdUsKqCHSvhqlDuieKazK13JoFJHqhcQEYb0nl5jIv
0Kyj7CXXb6ahpM26DZSgltPn2Eg1GgRVjcb8I1Cpw0k6hwsnx84Kxt6Y7/u23ElFX53isShPD2uM
BPNTxn6Q6vAJyHrPHytUt/GRndBLYeqT2MZ0CDz6nTGOi+8209Ub1KiLBtwiLIaAx6W8u32bQMeq
UzhjmZQ1rAQDFWDY8FUzUZ+0gxf+WXtOfP6eUf2SrOb3D6qlnfnZ8Cn1H3hO0Ff9JpXAMHqe8lxr
tjJgeRqd5UwBVeUtmikuardP9h41jOTth/JmSZ7lE1kW/rK5qmSO68PQUrAfwmohawuDWAdUVFQ6
E58Xp3bNxjIGT+1ChvYxTU80UenMrj0O2l4cQNW3WxrqkLeMGT1hKNmlWqMQv10tf1R/T3UVDK/k
ELm5PVPbqg4hP3hMdXOEt2BKqCn7vvS34DFMsYBadvFBs9dWY3jFI3hgnGhsTTfoJV1BILCYVkxI
v9GX3n4R0+r/FPG9ivGBRltS7OVJRoI5UjWc4OlVaPVaPJgc19INzjnQ0o54Z56v0VOhMjBJMFHm
z+LfATUkWezdNxyXuy//8lYPDFx1SuwfzuJdHIyslhmIzxyCTL5FPZvfVvUP6bZlF027Can8OAnj
6wotXWIeb3aQ+FKj3ByNDCYkL/BDac5LBrWUg/q+J/hRNdp1BceMGSeLhNlIf4EpvRlro62fp4J/
Zzz5tF5fIn+BXsfgBvofyWf3RTnNVFNvOT0+1V9jlflyMapSkKXEHYGW+RX1rj/2pnQd6qty5X+k
Fo6oRmmYrsVRJwiFHweF22B251Igy9e6jL4n1+g7hZEExKfrMo457eOBso+w2SqfAKo6GLXYAYOg
V4eu+SUp3wYQUIS6zhPqCOSpp1BBDByik/pbSTujNcmlOCrbZOV+IGy19Xrocrk/25qyVi0xixDB
PCfNognvAC4xQ5d2xCI1PeOo2prSqCnbQClBBsgVfAPtyPUMb43Zwcz2SkzsfnYDQPP1Ia7xpFcZ
tOoU2X65giiCWyCkRov839mQLviBJoPiy5MWx1bOt8x5ykZ699ab2iS7tPNsuz1dgeLV9dJY5SYn
yBplJ/71cIbDSDnU43+HRP2yzuvCX1ZO1w3JkagStVC231WqEFHw1PibDyL1fgovAbURJk0+zpCa
17VfUTHb71b/VWgN9sd6nV6EyhvTxZIxLVkOQtNHZf3Aw9Z0O6FTn2jshwuUnAZ9bjTWqF6eNxa9
4uoUljCgi69CnZVGuOPBEM4IqJ3614AQ89NhIQN+WNMiojSmkbDNdhJwJ8Q9JSHRSmLTx4ETKoIs
x+yKu7K0VhcmYUJeSlpJ4H/nPLeAjgtVa8LjDsz6ErvoB3mdhqaDgfsKLXFzubPIKGdMq6Haox3C
o+JkNXfulanH1yzPVSy4wVF3bpGeX7TE+W3zYPRiig/80m6gZxBelTOj7TihoG1m57e6iPAoOy+s
MbrsHg4gsmi4YsN+QriitDz4zCFerUa4OD4IHqbQZnBHc69FJ/8oIuksSIyGXRIAt1YWzL41jS3b
As8Mvm/oX0K65elSEjkMJF6errRg3n2cdAOX9Z7DyOh6q7OCnZ/6fCaZjrwrrK2zQLL0T2Uo37bb
7ATL4yNjjgglLnILANIeLijSeR8U0XG+m23c0ogcYsbclHwl7ue5vO30RJVLny3w17ew20r0rNJk
L/kuYVUiZmEH6XUyHjS/o1BtD6ExhbugvS4mYLNAs6+7mF7P/Jf8smKCnszlnnyc0YhVmYWTq/j0
caFhUfEFTZIFXehaJB4eBI2nK6nEI5bw58C4f3OGyaYzUVEbWnXDX8U/ip/TVMf/OOvz9OHMiSuH
My6LktItZKIWXdFHFaGLB1+1utbgP6u7MXS14tCDIhaVCB8Iz293BbGVstLDR8InA8sN41Ar7y4u
Fnwg1rCh/iVwhL/9NXUlb+zJB4AxJzneBHc4Fexx7oUZWn1Ww5IM91GA04NytQ7RGn1czuaecNxW
SihctLRxhKA7tGgMiouF/mjBySr+LcqXZECHSstCLA/lLJ5fz/9uS/p/ln7jytN06xR/iUpAuyAR
kyjzECmUOMxG2qQQHyJiJ+t4g1HlLQMapiNRddUbEP/9YK4MlEi3qHJJiFY5OPf6se2vuGKtUcs0
f4WyycieDHx3o5HW1u161z0WBZQWJxxi0CJF1yjsIUroikoYkyhbrjGVC+jcAvACXpvLYpnjyZTQ
C/TQpcd1wVFY32jShhedRqrPuOv0V/s3w8jU4WmrZalWaAzfq1a7hpDGNS9GDldiirt9y2nGpF88
kZNc4BWeb8z04Ov9W7G3TnVWaAmP3InPtwCqVllTJgX3giBJeyjmkgxvJR2FvnK3TKcxfdRa+FPi
s3NNdb0H1WS4fyLjLiDkrrsLHvX+S8ocHJtmjbbu31zQpW1Q8a4YaUG6G/0U0Wy/cPqAtUlyO5Hh
i2bjGinRlSIDFYnvdku1W0ca4sHoXde6g7ufDvmJyjkvv0EwfSNk/uVisW8mRIvQCQFX1UgMeBeA
/A5tHwH/WSN/SLIme16PlkqipjweunvrfOzs3Gib8be8EG1+rk6HeWwf4qYjuG3URpf0GyZKj9zd
CX2wg8Flxz4aLqAW75PlqMMHSpC/G7rZoq3oW3LfDAWfnXuMMMnqzd51kCLdQCQ6zAtJf/oCLscF
p2oZqNbDRfjMwDC11zfGb+jo0nYrL3/sfGsBJI3292pl1aggH8quKt+cW7o7Qvsh24CUu6CVEIFY
8f6r5t/X6Stxksqi7S5XQhABYyhyVplpylP1uboezHlqZ1VQD9nCegAc4W3gQRKKpKtqz6Qbq7pH
R3Msq295ychFt86h93TGD7bIWBTWiOo0+mpBX3kh/C25i7j/2R5vabUcce6hw0PLpRLSN7frd1hD
KLClU0Jflr69OhSWMSxYCdVAaAVerPcyMEGTZ+DSzAmWaMg3qqBNB9Q+06+vDe2OEbZG63o/0IJI
Lx3onVfYhOFmtoKbCbl0WMfs9tFGEkmMZg3uDBG9yvcpAkJBa7+rqdINnPE+CsPfeYh5m9Z4jFeT
61NUmywNtHKWF6lYCLt27sgfVZklflGwsVD+flrAc9h/4npATJfZlyFliX2Df0a04+hgOh8r+yoS
l57vzmXIR8HuJCXpoS2SYkeSl0sw02CfMNcvK9Q+j6JeTQodA5IAL7NFatOrI9Zeu6oS+pLgSKn8
YYNQ2R+wgQAd/SUOp6gdQCtJUEaph4sc2P8hVjSUSNOq1UvVpt6CcN4qClgR0K96dShpkR6wJNv5
4m7MZ7Unzl4yna26OvgA9Xsm4l3TOgSO9nk2KLqHGZFzL4cRoo3Odtd95lnbM8+xEGtD/wiHWyuj
OtD5X4T9o4YLcrQQVZgGac76+kg9rQcoufGQmpBohgfvhR3jEAKi0aj1i8msTT+/teBaIVl1vzx0
JVhEpic2nx/E1Z20am8aixQg/A0r4EfIR0M5Gfeoe2bwQOWd2llVmYxZxC19oit4SjvmANJZeqGQ
OuPtbqjpJPUTj6KVC3c88v081+ZRi0F7fhM6KzBETtlLhiV7/zI26kxEDgBOrrXgN7asnTjb+T1V
KJDLtLP3e6zZJH7vEUiHE9nrOKCUo5hNobbTcq+Ur5WeO1W017yXiWDwXNLEJXF1tDnYvaELlIgM
XaKSDV0i/wTAUBhIGvu5EhqAifdID3dMq1ZCG7Qof3Xjjhi8ayclSO8wgIM4xyDzot37WZl63/Su
S3+JFWFI0YStYws27EyLaHISXDWrkYO3N1Da4kb5mE1s/6tUQahn/dPsveF9tCR7RolJaqt2D8k+
NvP2T/1DoKmQNmmDIDramqFzLtXnhIUehKgQHeIgSEmXm6yVL85OAofuzBqL+mfuVW1qEIP5ummQ
irp6/6HkWR0+6MiPWTqOnM4pWW1yKC0DLnPXpT1t3QX6EQ90IDp7RpkHo9ugFsyHx6SIr/TUSSMD
cRZA7xLoWJAq8AtKwpEcy8R3LAMeWzxKYo/y0AeQ5uBGUh4lAWeRINUXmqEqjxsuVDDx/iQXWCXB
AkOQyuZARhV3TTzaRelqiElarc98kd14/zIRG+Qz6/yCZcaMvtOt6wUV4XhS80rp19bBaLlPlgB3
mJYF/xREVRVBXDqiyxssX6UurqFLuqColdyczwHyJOVYQ5hrbxdTRbItETFB6P+sNtgGTSxbz9TR
Bzf8UfU/UEf916E0LLktcUjTn29h4mN0Qn8b7q4jis+pjpI4RIIQdu7B8Me4/KHXN4iYJt2yhLaO
ofIDTfkxqJUtyJU+bXY+vxe4uQpgNs8KRCblUjA2qzdmr9p1wjbtd7AVg6twYjL9wdz5mxXrcyNR
YOky/UildtM3M1I7WQQiDfTW5JZHDjvOvI32Z7cJ5k/rEDcn3USTS1FHyIlQ2LC3D2i9CFybUAsg
Nq8SZ02XSiDCxEO0PxQT8hKt5NrelkDh6lf4UBXRgBuewOkRsgd4Kjxx6PbR1e8SUxR0TnlOwhOJ
fr+RnV/U1aZL0HvXffPKd/N9DCmcRU2+U9SMvEHf6x3Lr0pG9dB7G2CNP16VXqZc/5Pa685Dg1OL
HI5FGl0G7ZM7qBNu+b86b50t/khap0JPmi3CipusEcUo3E4EiZ9WG2UMoXcc3hIakIyn+Fm5uQhT
TbKXNCY3zz/CmfpXcnyoFgwAQL5t6EHB+1iwrivI2Yf+q3svLMYxcqPNcTvDbJTmiPJhztBRTVtu
NfBiqtJAudZ1IavDSk3L1NfAVswJJyjCxRKqatb9JXxG2rQSSxRVD7TjUHjubAhunFNRcTXkHENQ
rJFXGzhYB+4SMmQyLnn2yEBSEngkOct6woUiag7SRZzE+6S7VgRgVWufvnETfbkstXWdWZOAuFbK
Tk0ih5TZ7nYbKaD8civD9YNBeOIajcZUyapv7EVQIstWzcjtL02YHqYtQQQEFwdb267fZiEvUDlQ
P+QYB5dGu+BdpcQoGe928FNobaTsc+JlN3k+cWK0d+EvAB2an67icl78Zy9uh+AnYPsWfslLJIXK
cKPz483vmRONRnSJGbaKD8SZwCsadwxgxftDVFDcbiAzR8a89+eogOAHXZfLw4FjW122h6ErCoum
lTtc7ysj72yr3Ab4ra1D52/WCauxUC21xuZ+RxGcIE9rPNgs1GU7krTdsguSBLKE4XN6ZfufLPE1
tL1pZr25+TjmiPnWepLZy6RxnpSQx7bOKrBXsis5dAPxIidR9TfNMaT5JtcI9qkBcGv+icl/o2e1
tt/GetbgY1hZ18OoCunhzhatoyr+uE76yXMh/C1qhbSLGocbJoV8AppZnSFFy7SBPeQPeVRy9bSf
516CVSDHvVy8lCVR5Fc8IevlOs+179RVIWp0e5U7tGGeBmUKeiuPH5TVRGXXR9kU3lQ96Ps8pWzr
eHOTRdCQMRl5hjM7efUPMZxVQf4vqe7ZcsXAGOKKNyiDvu8plFhLnWJIhE9fMeiN+mnX1SvhELpm
MFkhOX2EgwyTHDS9haDsZ0IuqQLVmn+vqpktcd/ommiVET/nebp7wXAp0/fqNSeoxyX3FGakTNLC
Q084CtOp1i0rqichGhAM6FhmXHHDKysoAUgr6q1N8sGhGiyGTgfzlmgGTD9kqO0EnatUvs86xx6l
xlQlti3aCcBDnDhPZ4iIm11x2Kc9UTcZ26VtOb3k0iAURrdU0TiSLkV7nHyl3AsfDaPsTqSCfZ5m
slYK4XDlYbiRlp+K0sAlwoIgXcWwHKW6JwwsJFR7RX04wipO4uFk0in91yICreTxKe3HRvAoSM3+
l8VicmEixWSpNE/4rPJRaYDUktI6YVN9htxiAm0Q8LEIaa81mFLLGtj9DpoUh5lnRJ33vC7dbfsM
4iz5oSZuUlcZPl/4rZMIRm5zKEVwYX5HBd6QbUL8W2fSZ+ePrSnyEDHepUP0cZGXXWnWBvuNButm
C+6wUQvPZsiQP0l+Aqd4Yf+NC3qFzJVG2o37QK8zXu+RK+PPnTQUyqYE2sj3TbHh3bbr5KONePpQ
wom1jydlgD+JK+M9c5X3hDE/WvYufqC2VydtccirTtPpwEomzlQzpyfVp7B+SMpx986PDcuhd/JC
N7Gk7lbcPeRpSnd28BjvmalXXcg60+tyZW4AinXU2Ybq4TaLLGTOlZxNsyMLfYQ7yrHK4VE/1TBH
N4yY+b1axWcLP1G5y1FsXSsbC+r47CedWo3d0JlG7CRoCQ7nnXP3XYqkKW/MbP+FPXHldxpTridQ
E/htSU1BvbEKYDROJgdpYOZJhkw1vuaw4JnxR2rifghbhqo+RPPxO3aD7ws7V4vIhrwVanq3d5tS
WXyxV9bRIrj9p/SR2VA/MGzpyl49m9vSYzsivYDFlhd9x+qqBXfTHKXE4bAdMJhP3chOiVFvbKvO
mDS5X8u0U3xtKpscwQW1OxpsbaRR9IaKcpSANfjSM3/rAUajKrOANrUKdpDeiA3y2PvxiJXjNL5b
Z+oqPnNm4FiH6TuHY4lPqDrdogh5RjOCpd+vfhGIj21bsJsMvnQMO9Jfi1pHSI9yJ0Czp43RxGB8
mxBOqzdcrzyo6Be2FtRAebMldukEg2wjRy2rg7zuqZHApuvCF6XUnXILKxgKna7UkjzPwNdmg4GQ
8aa02oAA6FjzQrQOwdfehVhpqFuGfzvfgr+0F0EtKD0ZUYG1V9D1ZKIRxsD+Six3bUYXcRDKkriP
gMcna8HIqVAElI9hxjjaONrIZkpZ9VYqdIMXL9zAVB8Hw77PpD+143/o8q9oy9+Tsgrtm8NjwKsT
ayC0SOGyrJlwlvmfMQuAgCyWQFPNp2yz2v0oxKvSggXzsIL8AnfgcthDia0Nwox7s0B4vPLdJWOc
2niwPRcY/k6cZsJs2bHaDrwXmVpwWMOD/0wrZSr5ELWvUYr4BtPw+1ekyS+6WUjXW7r1nXKVgNDJ
zeXOylEvBa8S8B1FDefqBsQWBqyZD7l5ihiX2rP7U83dyH9OqT7yMsTGtd3lQu4UjWaXEZrhSj1k
k+NcLTQnnQ2W7MAFhHLr9tiYGNEyhqWzf7wyXMSo6S3B68PwQYwzuRtVp4tzkjX5bhcQ/JAJHT9+
UnETV4QXwZLj388nrPOw5O4SmeB4H9NefNiHhSHtpLiapARhJgFg4vL/dFCEZDkW9ll9Jpot1/xn
q+PcGYQEKO9CfccyTw+D0yJXkBAGQq6u+tZyw72JAkKgEvuM9hn7hQkTWNWhKX1EO9C7mxzCPXKx
+GwAZeuSsj3tFXspgzyyhmJ+/eGpXwdZTqHbxV2GBPmhN0XQZ5ejOd+a1prhMMNppcliLAzKd+Ml
9ugUrfPO4HfotKzlx53wgA78E1FvfMhw82HohUIHG9jM2NOEvXahYH6Nazyv/Pyzpw+WO85oSk1a
9PP+gVaRfSa71CCJp9lgEC+6IX3O9Avqdnyf9zILOtbEKhcsEEMzy8kLsKAQk+VMXQ3YMEcVT1de
+vQDM5DgPtjMjoij2XfnRxhouXXwzwZi1YHFAD1SDbST2CE9ZY6HLGgmdHnI+Da0MqS1aajfVso8
jRrSXu+XWXV+iUGz383jApVDmpHzuzmxNPgTbOZUXAiuIRE2KHBJj49CSR6gBosIDuMBpJP7FnVt
Ja69dX/MR1t6kWBR7AoR6ex56L3eswQVu7TQyxJaLLe2y/M/P5a6i9kveMYvJQOx0nCj00sFRTRP
SAegdbjoNmZEL/uFS6zRNcXoVUbOprvgnia9q3lJL6Nm1ksLj0bU0vQpCVHdALgusq1xHRIxTYeQ
BHqyBKtYRinsoxY04mZPWHYVGETzTE+1IMjplQBqEHv0uB1hd+QmXTwZvDKxhn9pFIubsmNNBoSR
6WPnus9Hfwsmgm1J4V1GFYq9Mm8yScik05EsDOm3vhq+lzc0IWh1hPLr3irp28EDhD4eLCxBXKc+
klayTdeTKeBvWYI1+q1gFAdwTfIYuV3rhdb3mqt/9qd0JzUdQWbncLmD8BC2vWdkXgUfugKBGn9/
o61xIrXODtjjpH5TxcLd+CeijYIPVqj0BDCxx7VPlG3IbUBLaOdXZPV76H5tXvoYtnp7tx0RYLiy
iqLtvOaZ2b1sSzP2vdb36wPsplolzENiShQqgV+/7fzernq6FwloBCTC2RLBMWo7HGIY2tthH0oC
6ji3SJEzEmNH8RV4sk475Rg/PkKcbg7aA4uM8zDRwdXzPvA83SV8vIv36/qd/gvn8bESgjAPCJj9
RlnJ+0HLUMCs2r8DHLZ5+pwkWX56pcuhPi3ONsaN5EhhOHthMBNHfaDhVc1xSyztkflYlGbVvaCi
1Oxp1l03KW84FlJXDcwmQhlUfYUE5wu31a4MQ9DouIbI15zQ7kHEu3Ht3CLNR+E19xr5I5Qzgp1O
QJ/61+ykfxH+DAP/cR4WAHTluQiaoHW3JXxKUvtKJvCRtnIpzOJCjajrZDvNj/K2UclbsOu0bC4O
taOa9j7+jag8BpW7wCBlVA9MQV4EH0oAdxmbm3WtiU4U4M3RR2ECCWJ07W53ythwb7WS3bY3GBSV
TWH00D49xWYHgxobdhBTEd2cVPlyV7hJdeTOSTvpdd7dhwPtG8dQcXhILDKkSjcOBGnyUthW7rOD
5VquqUcTQ7TM4p9aA8+4b7A9TIdUoZEDRD7tNsVKuhf0HQdoyUAM7dGzPVZBMvAYtNtyPNCQ4sbf
kCDHpwX30KQ71lwnF9OIRtUKVcRTKMCA1EG+MG/kWwz9ykwZmrfa95px3Gtec29X7mFY52nCUZ64
2mS4N7dUpycvKDJy4fXlkE1znQs1iZTE0hS+LaVTTVuzba94V69Qj3cviNuRaozbJcTb9kRnsAQU
u8/WvxJy2LUamwZmEXvxLuGimJPuvU/bPORvzxqLLb3HFgEqG8WgWTOs0Ho0E0n75YERS2mmk0L6
z5mnnOD9xEmPEfygeUHutwXNBtKf8OkScchiW25IcGvDS3vXb1XoieIuLqhwZfxP6nNVR1+aSX8X
btvpeUVHooeR2NK/QIwqOEBeGjFZXAGnMHJEqoZogJsuBxaqhmE31pvIj8eBHEZLar6PKYZD1xzT
66gaeAXXKP7fV+PXvIN294fJ789/TEQVOopkrFiVNA1/RGmj3/FnILGyDMeU3DFOG8vcAWwmzEAS
lRMLD5rclsUFXWU0Q5DDjV7nFzmrGFD1vvZbB4q1OAnGHipMQok2f5z5kMCPBRH6eFqCv4gxnpl9
0o8fTW9JuhKzFLusa51CZHcZpe8OXpm/pAT3FiczV/vYTBqwI9tiD9qhSd8R+ODTCIHtChbpBwQs
ZfCYRARuKjB1XdWTZjfjaz1YZ69PjQS/dp4JCr2j/879U0lfjIhWBan77YmPQAHxVPWebjMJm7YG
Uyz2lgE7CzJT8mV+US2iDWxzr5Op9tFBK7pFzx8ks3zHv82YOYPlhaYnH+kDDdLg8Hi1TCMLqIwT
/I+K+G1OYNeaaL2k3UwdzFU30k8Ly1mnhfZhNU0COyPv1nmN4Ok7XYUik3muK5TbL1iEYsqAGU7S
x6eW1pwzytZ6Bx1Whk9d6Ztj/izTozmmM7JK4whG5HBt1fztOnXc6+IJTmNx5R/5SZsfZ+mBM630
9r6SnoEl7vKX7bNO0MqKT3GtVmK5l1ffia6STfi6IBsCHk957IvRvjVFhK3JlA0w2XWSMm0bRCSB
3RCmMNyXqwcgNsrmTw7lG5Ekf/Lou3VO5VMMfhYeWr2nHSzh1Qz32UhebauZyJ+6FlGs8Fxdiv2f
5wBN4alWAnHXDMIOAyEYx9rbsKq3TEgeYDFX61SuEmpVcTi9ZWHIBRst9UTRDDyrFN2/xY74Sj84
Sl6FlwbNew9SiuICugmW6EEKNUp/QNERoHqUsBW/nr4KGnF2nR0I0OLeEtNpPhAYcAIi1d+s1CaU
/Y0BTf1AZfgZ8afAJiP6/FwMyDW3Oi3pO/gpBD4Us5U0sCyk0nn9HG+2f31ke/43w4VqNnjziPTa
t+v7Ow1Q0xUlW1FrRFvbJGOtU9UzUMocyNEKNGKkLGqAErzgSA1shAbvigMB/RlmeDcm3tu/WZUP
aOX2tYv5guouOeP4mxzjWfsanidCpJSSg6dOySkzcpuicuV05L+6mdcnUnLGYGrmtAsFUmN7wcLK
i4+pn+A654L3ZmeE40lRoAQ1viXUkt3AkamnDeWNTrsig0gx9H9s5WbYYrBkGjDDl/K5fcV9vlpn
ZjpU86teGhsRYBThGInXD+Humf3LEDkIVT+VCkFkgXVDElL8rg8S8dg9H6Ic6AIvDOAPXuc4SBwW
5x9yarkuQXkyp002IrNP3zdk4//O1qJoO0wXHItNCAyY3sepFB6p06vfkY6kPaFxkS54DjEjiHS/
k6pD4UoqWOxMrpT6WK/ohnGi0LEctJccdOldYQkSB0pah9HNAr19b4oS3tVVg/8RFBOSPrLzXsbG
wdYNQwC9W+LOv+DA/mW4B6+6JpZZ6fLPbs9cKwU/L7L7dziSsvow4S22YbThuVp3sjUrltDLZxhU
BUz8YiMlPYX0UA1RyUkc23zZqYlQaPqgfe1bQ81XG3xY+nnQxBY8jBqO81jmu2oTZG8UhMS3FrKV
dJqn+Twn9P6hgb9XoiE47ilF5v9AC0Z9U+XzJD+Cb29+G8ODUnH81oySExt4GJk7QmCH4HfGvwk5
uiZAqaqRGbqAcpS/D0/zrcOq0EVpBXKe5J/7vnNPASKHKOfBLkCtqbDPAXkUDIkQ9NNy22T4KrNe
/QHmyuXicMo7qGbU6si/Ao0gYBCy05iuP2736GfQjMY/CFWbj58NJLJmTWhoxOKFf/9X1+0jdcoq
WFvihdDBqFWH/Hd5O9n3bAXyRtImFLZBPPFKfjH17OyhdiXyQukSSjR0jq66xh0p8+trJtxfPHig
orexKZbf17lQJAgNiDadVm7bKegjkFjUNRdlhnjcRj9nke18JGNJKuKpQ7BvykoTb0LVy5P3xKmA
Al8nMUUGkFL0A51ZufcInuMUKLvdcP9zoF1O+OXN9Jy/aetHQEzw7MctXWcDKbmoWhYJSmvQQV7b
Rsjtlb0cLvGDsnJB9fxgwSWKLewJ1BD/cgGy7Ub2u4dAwUwsF9WBBsj9z4mXfXx9V9CkA1phrxJb
cJCNPNXYkDr7yVDcZORf/vTU71cgg6nUBLoeV2dQx7BXf87z/c1jlier+Xkt+DFrBY27tbKRMBEa
E6NUtgJ7UyeWJqSM3kcWbh9T51KkVPq0Sks3+7AMUUxa1i2lCo/RJ7DL3OYXvizMK8VYYDQeqY5R
FGIfI82eqW+Zkox/NlWsnUQ4U60p58Nk/bg4DRMMhpdV9jzaJJQMZacfy4RbLB4U6toGGIkwsD8K
k4aB3JiqFCaRAlWOW70XLQA93aFRxbkyMeTJLplanpjKs+ROU4p2gnxFVr5QP98L8lg552DAfhDh
R6mDXVXDZH1EtJ6e9JUS7v50bUEzBcX1UU+dtEnQxaV9iWTtQCnoVrIfw+ShszLP/k8kqWOsM2wQ
8i6VU6lkMxf67RcBaGAGjAa0nDDCzPiKpvs9vsEfJ7+f1Jpq0v54A9S7LGAJqVz7rMSvu9XW2neH
+Jswzq2sqL+RK35AzdLJ/fVzFmMZ81XaPTitD9GBL7DKzFkCOD1nVZj4Aa8HgC35Dkuq24lEGAx4
kDTh6J/1cTSWIQyZV6B7LKSuLiF8R6XKiPX0yNYZnlM2TJtqlTSdwtnrWy2k9LeMRc1939A9WQsA
MsWlx8tZ+jBZ5vGgwtZLQfDJ4HOosuUaJQIRohGbfdSqv51bl077AcswEAMDeQQX4tn8EDXQ7v9L
86LNHdh0H2mjrtsDqzoaDj6JQZL/Y0pF1YwDnooC6GJuQr+wdpWMUMZPnJ37R7WOuTCOhpZbX73j
2R6Cdd6Mn8AlVy3ONVVtU6nz3sK8IEUf6vHy+R9x+xJRsLiz/K831b9F3RaX8EE7wqRMczv1/mlO
5kV+IOBCtU8MZkj7WwIFJT8pIA1WWN9KvNzV+SoE3kHPy3fAMmMVidZqAqS7WbO1uTbbmT/eGnDg
t9hi78u3dwqL6qaLKa8o6wG5xtQU2sYDts+2N0+Ndfw9SJ3ldiFw1rRCpjVwM6oQpPHvriz/vk+I
WedsL6eU2Wiqpr0I/oRnRvjKr2WHRx5QJkkw04Fcw7pWxxeE5LNTCFJaX+8Pyn8hHLCRFP3VMIu0
Y0BGErPlNS42gFiw1tuv/PbNEUvHGWUJSQTu2256g/SiSSPQcauMHpJ8ZigWqdJiDCCSbZE1KtqZ
RjpBLpTbCpAQFUPfjyJaa3AVzFGd5AIJJB+E+eNki/c8l3zp0Lyk2HPCiN4lZwX4RXBua2f6Jbjv
lSk86fHGxFhH3ue+4TaEryG/JLA9ibJ5YkIxnlSOn/zHMLdCW2lxFl3k/UVdYm+U5Sh/zczZlC23
NxSVPNGf/T5i/mQVJmYIh7VhojNZ6maWvpXfkpcQIBGGxwUtzSw6xgK6TfB/36r+q52fKAER37zy
rnN0NkwjFv4YuYct0FthASgHdG23aExRmCl0dsm3j6A/XWEuoXeq5DGZ8HbEMwZXP1+YaihP3ZTV
EKYnlhDHp+nhiMK+Bd0EaFedP/4cBAlSlmddWHlcPcKdfkDBMK2fmOUd30EUl23vLHJjkLmZ3hBk
cpg7guBt+Cvs1Ki7oRPkEpttlbJfakOc6e3eMwvWOugC1V3k6m+N51cMtcoejwpWcAcRBcLuxidU
L89XmlK/jVDhCj+nU3FqJUQVYAk+ScHebtnFu+n6X5H/XE2lx7e9d5sC0w4ZLGq+wvvNV9NjmExb
EDNRrTIG/izWN02WOkJ1XNQLg6zdwuOkhExQ8V1FlouwW89XBYCJMfvCqZX1FEtPcC9pdJ79Lhk6
B2on2QuHCfdYnHWKF00Uk+dBey1q8dRP3/J9vHb3bRgb4am43SxAr3TV4JzAmf/iUovM/28KS0P3
EBdmCJ3C509tr8xVwMnti1MwTmsjBw+Wx+upVr676/ZkDT6D5b3FC+pzgIR/hKThak9bbyKAhW4z
nqSYY+L29uF2hFlYiM0P7lCdzaRkbq92PyBh2HT7icnYJmC+tnPraSO3bJ2jlEJ2i8UPzhvRkyFo
7Dc1h6I7NWeupELcBvUcemflQ9E9URM39pdPOepW5vVYGw9JpZEv4s42YbhURaHzrGllXIOsMEYB
Ru0RgZsO0IniUdRinD61v8LjbLgLz91sHyfcIasOQsUoCEubDMj7LMuO4cpUFFyU+A7m3GRsYBPg
cmZvzxjC88Dw/a8ckZ5LTlAfhe3U6TI6Z+uatBcYkFGZa6yYjxj9AxsqUZi/agFSsuDOAaR0qwRf
G2F3pj8ZWRK9g9peCeZQS8zVSpcTjavR23O9mi7fai4xPNb7GtRTl9O9tgfhYj1q2ifSq3UDRXMc
XR2RJ/57b8nEwdCkQuPTtjgKjONC6s4/UMWILlXFCNivsVB/0gq7oezns5LycRK8/cbYohQAAnm1
CiQisM/QUzbawIFi37xXpgCllVh5dSlh8E6cnCpSxyOn3yRcvUTntpGFPJYcoHL3ILY9fQrGQ59m
NkEQuZvUodtfQmEtniE0GsQjovRfzz7cJ5X+yIBJl1kWLHaLtmA6w7fiDJi4tz1UQD14hERTdeRl
OcEHwUXCianzqhC4Had0DuIgLKOzdNBa8GmwL50JIJirHYV353+v2sj4Wg75ms7+vTVrKG9Qpd24
T16kID1TFr4VPqOTsIn610McU6XqtbmZyzxpLfojiaU6hTlZ45rDoITP8hbt7AvEJp89pkrFwRxt
98G1545XDzzRyOZtFehsV7LzXv9C5lOmputu4s3e3NX5+vTBP3z/U7IqHRJSDp5AqHJvUdJ0s6HZ
uwsgZixfx/7VmTF/HpLS8/o3qGnVwJtalFZNT7zwxEvqscIfgUh6UdLs3Jpa+oOBgpdgoAjFzrD6
aentXur2+D0gBqiobWHDRy3a0ZtOPTRpaBF07+6JPKa5yIDDB8iTRrWSq6+Y1E7nuf2ShDxg0Qu4
7TUnuaDmVPkz24fJvqm/jKLEVHvYX62PTm5/1VEhND2KDQLr47EU8911XkYffEZRVCgEwFStpzI3
TTFbrHPoZQJUURHNu85jJ/wdP2rHAr4gE3nKPg/bfCfCbElidP/Jf8QrPR7ralEB8nVXk7QRX72g
bAIz+jBW+hamCNn0g3VBSshvBNfXJwdBpc5vN3IfioNWEnufU4aWj0iefdoLbGdspqlNJ5iqGiWE
VPCf35Vydsp+FZgy1owkzOwawmrbSW6Ihw/9vuU3EXmPWo0RDEX6QyhXxHKStSFz4WA2dd3Imk5o
s3VXpzgw4tVOSZZTaJ/UKyL5PldfHo9EeLzQNKX9FnDkWg3t8z9EmRtbedZ9vXI+XuA/zGde7HaV
fHpef36nfc8MRk7QR8XYjWQWj+oVFwwpxnCofhHrn9vRz2nwijTyCk5c/dq8SWj1L7JKYgPOc8G5
5DtEysqCQbN09Asu0C9HRaApAbu59CMiRKdhQEkaAbZXxrPTzTVUN6e9X3QdFhMfxO9bs+mMhDS6
b1UuORa6MA4QSukJT1cfMAxSeU9cCw6jdwz/OjN4pW4UiQg5GpHjA3eviuNWspIB4ec11gayVhA2
lfZJL7hfxhoKp+Lc2HFLxOvo/GhG03e+B5Y0YnblTw/RF7bXeuxPPMD5oWC2DhMNNYWi/Hhl0CGD
yB0JH/qQ3r9Y82ASgKWdGMjGR4WxbJ03xi6oBP1XrJ0SrfceekW5jTuVHCWwRSH+Cx1tAWkaQYRX
x0kBfLWrxEyZdqdcN7ftxrCuFplqnZTA3eJfFOFYfbW+i7DxVJy0YfR70D9aRdhpV/Rpfv1+EXVN
h2O32HA5mVLr8wQnTn5b+8m8Y9qaH4o3EDJ6Vqr5zYza1dzfQIMIA7kDpbMqn08A5+9ndklnrQPL
Puix5kGwTqNwri/kenTc1RvuI2iqmonJmsFxoMzULlszCxTFYx1R185NnWOw/JtU63ri716XlNK6
D0P1JpLD0JqglTpnRNC8rVpRhK7gCqDJyJ6Dx/czsGf7me2K7/r9BxUFo9VqGO3WobydobK7pwRB
Q1Y8/wRfb77g0GxNtJjbQvfu+SOb9CkHRuzDbhB23Uxf0go/WITDkbDXr6WCOLUcMOVWJUWT797V
JRklsuxpFu95KfgY+7FIjF/CYnoIDYj7x8zplW9XJjiHmYhpLfN8pdP2iyMNDF6Sdtckf1blqrMS
HekMsLmcMtfjQRYDtoITkN5UiwKXZgwbOnkXs0uMx/nSPP51UirOk/KVGU3otUNuDPZSzo0Js3zh
hg0ZQY7v+C3bxOI+bvdow3Fpca9f1fqlg+JVQzGXtWEiHpyQPSHCjKGD1OsI64sD9LQV8lV5uYVm
wIXA/fCl0KMkGI0XDtzwm1UOkyT+kH5wOkHoC1cqLdO4hHlDSlQ7hheMWeS3BnvqNmumiBDbVAD8
e+f8NZwCFAreebM8ob8CTkANqCO0BNhV+vI4T7DdsaHboQfOYtzze81WqSetwlFaOq9/M8V0HnKI
TEezTnXS2dt0swUXs824Z75He2o04foqPIWmsKVG9qCBUs5IX7L9ZqQCjWpPMxKzZF3ViSnfxscS
PW/d2OyvoQgLBjaiYR3HjiTKHYhVFh3cv8ic6NzdxqOUvC1gKnqfKDxzUxHaHgFPt/5XPczZHLH9
v51kEJshLIDTp5/i5druERwqv8+Efg3tr6LP5B0QOqVb9SHYxrIMaIY15EYF9hfzHL+6JVG7bDbS
4Eh8+CW0EFLn/Y0yVTaVp2eO0KjItkpW4LQ+O7qL5Zuu5Ju0Xepu7K+WqrxxL5XjSj6YTIplbSbP
QbuRJXk5bUregBzSscc782Dv3Qv2wosG9MkVBQtBEorcHZHJHNn/h3X3ICLMoVMcURKAq/p2yEvM
ax1S4jw/DqWBK4ZJ9WBxDzSwiCzk9Z0KnX5dx7iPWDQRrWDsjFy1oP7nBxE79btXHGT6TUxIVJLe
ry+8Do13OxUgbeBPfhrL1+gZ/GTp24jAq6DUnN6pHVCsyxPokFFJQ71dG67UQLCDQalulK4uGaJL
cyzRnd1ZfabshlX8GvZWY9UHbpLXhWJFfyNPfTtSQATQxLJm2IzhEgCxSUmUVaTsV+n4P8tSmP7J
gIjJEfKSnYvami+IpZ6WgsWbC2LSBfSoGck0w05w4rYrRyrSkPmWs/3UKiTXVpraMXHSrj9bcCRo
aEalGApmFc/KxP/v2SKPtRB+S9rc28KRiykmgS7ro9RWnFx/Yr3RIKUqtzr5yNPmjvmPA0Btux6N
uznsBvwbxCkQs/tGTw5Y9ELtAb8QAS5eAdEbBiuxTgNigwL4UL9XBkjU4xWGylMXB0yHSb0MtxPC
4Ya1qyYzyK/RpVw2+hynL2WhOb7KGHC58lNdmCve9xfLorLC9RwP5f305HVnkYIOSGJZIIUQmTqC
lwxyCYDw0wx7jUAppBk8eLFZwgMmcZtr3CcEiPhFe5maFCFFjZ2Rz+jbWMAXWoopF3WklkI0ggqh
RzER8iesxbz560U4iVw8aXefhWqAlRIZTQW8U9Fw0mzJvdREahLtIPmBjPUXJIshpB/Pt/h/9ZBp
sPd5TDScRQGUka6yXikVTufU5zYNI6Wn49VvqZziaS5bdI+rkdrl2PFbfj1JpQNwitQQGUCV/QT/
fKAhzsbqrwnNx16CoL8zn9fAh3oCeWQhoH+eHydFOFbHPgqJZaHNX8C69OD3lAEzwIdLKxtcyP8k
D0fQlOkp5fq3yOh+cC+8z89bkG3GUyLrE5Wq0JOt1tH+T/GRzuK0ixGdG5kRHZ2wf7f7Omu2S6t8
DEMtdVDrdrMyw01bSNXkvxmAfFFIZJpsgHmEV0JiUOH28hIsom8geHgc2/hWPsMmiSvkJ5GNemfm
hrX+nuFjOuutxDMa10FU+yuQx6xxq5q2P965dTIFPXwmgIo7oVGRHfaBZ3yJLlqNu0/4cZrnM+93
CWVYgOoLAxIIAJmBfdk6sxfEQRjHd//o0IGrJClDNsbw0cR2oWQelSVYDFg6pKMKQ+qxyV3UBLFa
FNmxKWYibFDFkUe9VdqqZVY3PkycRRQLD4a0ClmzeTCvS/3diBiLRon7xlwyLCjdQ1P2SReGTekp
em8qPyVKR8fH4b22Syek0C7zK3+Byd7q87N/56yX9HwJ7DJMOzOIgHItmk3uVIH2qJjAYnO3mpTu
WL2WvVBlD5Fs7/yl3znrCS5rQb29jx+vaeY4SQfM3IugOkyBe+UHuvT10kRhdTTm+Qxnmb7ELVx9
MWiEnxxWP8bKGAu+3vZACOzZWzFFeVXQEvcUdH5io+2a6PcbQP086FNZOk+q38jO7sLSH6z8GHkR
XR5db99VLkJAVlJi3f3EfYfh93MMh+PNv4T/SvRr+mBQKPS+ko1R4GiuM5CNRaEqX9D00KDi0KNB
Oc9Rktp8064a9V07D2RLyk5CwuXV7sjt6ShZozNUs7gFT/tqEpd+iODl6AtWRG6CYgPwJt7brKMe
sYIoEm9q6I9rfNK6TydGLjPDPl4Lur0oHTO0VSWHin44aH9etCrhgOW0KuK9iz9Qg4zLavRbCCOm
Yv2js/PXynAfx3xqhHN/vCC2lJx9awnFHWoyvokPJNLG3A2GVZ1Ghkco9pvpvRSHd6G9WMob049k
OzLsNeFw7Kr5BQ+qo+RmwSzwvSDt7tpiNs5OxuiNQeQxUWIA4Pb9j/wxySntzwBwoknLmQJ5mGuF
9hF4dFxu9bqx9UJRSUoWKwBx/FdPx9c8Vwba+VwIZxpPk9dWsbTZlzWGdAWjU3y+GzmWZgYqwrDW
RXq5hrCFOTLjFBSPQ7FOe32mRY5QL1lNT+kZNpUg7f22YiCHhy5yVDI8qpr6Ju0V/gKXMkwov6lh
R8BIuNuW0EFEypTLVKt/TEv68kqBQKfEQt6MNZFYipCJliy0Y3fM+76DVYIYObdNLelsvGl4nXCH
GvrC+YOqBaJ8jsRAWcBu6kLDcUFBK2cNiCrIYOWAvU50TPapOPyNW/gLKKoBzifRuaiG+pHuxIqk
dHaHKH/oOa3NBB7PD9hap7LVPUCdzf++F/L9BVpD/7Oe6Zf85/h5q4wpXBdnRAeKtoa3BFDMqJWs
9mvUFn2zap9Sw0dZx6lMiGTchSoGxctBIKi7gcwca4FYTGgW8HX/2Z7pKxH/Mf2ohvzvHffBpztC
P7C+TyQ2oVhsiyzTGkBVrG0z7ca3WpoDmXQTcpHbEoj+1KLm64d1d9qaBMGHoh9dPXzw3K+ZnibG
sJj8FS0p+x0mic7gGinszU1gMnCdv5c8Lb6OBvA+zOlhFDrtLtVxPTTE10BF7LSLlgYIsmrd+hgx
UQp0g5/p2AdgbS4glZ6Y0kvStj86aEZNuVZE5kqRi5vx13Bt7Sej54eYW4ZxordQBzgzG548d3dm
d7K4OsD7xEYZoiJ8pkmhi+9EHAQ8HaW+FoQReUs8R/QY2T0fbtcaOHJQw8hAkhn9E+Sco/De2bzE
hHCheK9qmKP1wOzZBxc1RRx3rrWYgdkXtLKyfUuZFW7c4+bBoII92AHGvzVfT0gv0bJfIakPsDjQ
v8ghiyXnPWwSojVfBFKdisFz9S9qPYAOp5LsmYLbeshS+5rpoZJe+FWP8ELMZP5mO8yFz9rXoukV
K5djsC6cjNcRybCpzWLEYIan1CIEdy/6BxmH94ekG9Rx8YOk/TtNcJxwpIgOJ6fTgoUmvkmJtxxx
zn8HdOxiYOkSNlARu0QQ3if+cEcvc1Vc402IyU0pSo3eRq06F6gcIj/0oLQ/P2ckE5rzb1a1PZ2i
TNFLl7calUI/svzcLB6eu/cS2f8pTBRhA4oLvuLuIaC1h/KuXV1g7m9yFCCpTlTvWo6rwmcxh0cf
a9gVHT+fDXUNrBi3ukVIKB7HfQ51Qf5DiBkmW9aZrzXiopkgF0237q5NQRKi4FPnuQz3RDyat9En
sLS2JPNNc4R7qcligX7t0MyoYsuhI7QFJsIGoBREcwZNt6BkBOlZEvWXxVm8e7yDM/ZEyqOpr8Hb
iuOWLkMcvhh9JVG1tnaKHJoRlIZ1F3b9dZx0irGE99mRV5/gtGpOSdKNHo3tdPvd4+gAPiheJTCF
hqYMq3vfkoknwhi03+CJ5B+IhFPHWY7Z8f3AGnjhsRiSiMjum+wsWDaTgewBiFMRuwV3SgzNfVYv
D6V+4ylHnXhpt3XLtjR4uRZSB0jdvnqgTKc0CYPrDXBfwgiaXG7DH93XzBFoCl/E+PKsAlCaP+zL
t6YKKT8QyiC7agEIlyjcGl80rY902uO4fxGfr1DJavOhzM7kCqOU28niSXO+Peo51BoBvgrSMAQm
6RP9n/d4a7ZaWb2TCQtSZUh4Wwc5UQxH8SAzeRG4u4HIBXxubnpI1LMOQ7hBEVstehozeQXdztKt
od+QIiceAcEKaKfHHMYyiS68FJ0cKYl9z/i5NW/TplWEPUSAqQXCggIWa4+eMyN4DTm/N3DyGpS6
j7HgGnFexhduXFQRrcGSg3ZpD5RtyxXdtexXFwJLZDF5ZBxuYfZnutdhieHf8q7ZIxApawadiu5a
l/NSy2g8CTqx/rcpfBxTN2Izibzqkx+L+vyLFyT4PN6BuCPN3ygDE3/Zmjmt+F2q4ghiqxDyqdOp
WBGcQ0E+bCbuzl2Pz+wSoBK7Vq4McI2PxDBQ1rFm5vfIvDTHWd+g1ynHi36ZwQfHYWPYJDrCauUA
ABfKSG7CKN9eEzKnF5fbc/gEiePe/CrxNB2WW+Sb5Sg5U+lXf/1RdOEKJOrFc3OTdFnYMEzPCDxs
SuiOpft6RZr9x56zBCsQsDcQjCajiK+BRs/nVkHY7BMAe8DhKwKuKZ5Lno43uw0jjRLfnKU/OnMY
Lwz9w8LL0vnJF6fcI/dya50EbHN9IgGnazGzfLjVGNrrZCTdZuCS2moiptpWawxE7pEEh3uRtMQy
XZMJQdcAbKe9oxZO74r9PwhhBKle31ho4ry4acZNM3CaI6hrwiqj5Z259xoixNrCxAO3/TZ29Rno
HQ+i9UxwQi4Bf8sxJxhO3bhm1ARNsaTyc3vaqIe5Y1KmYqn23LlXmWRaJY+wPcVf9lvsKVvK7DXU
bzpZ7+j5QPwPXelUEm89ZTPbJOFxqE2hSUqMmyZVlUAXFjbRiMlNqpa5HhJKqskad5X6sxcGbYGJ
ZtyH6LzJcOZkZ4pEZuDpD+X2tKY5pawIcab2yKpOyov4HjOAcpJhUiKOt34wqfcqNy96C7v25mW9
/Swfya39Fs1IQlmHzKy3OaIHEhewJvO7qEVA1E1iILC4Xl7S8BcOY2TNqP5q44J7JSa2Ynhj0BRl
8NoEvm879xQtsnrlRTU9mvhICA0mHIg600wUsF9pPIrUiODULR+kddSuV2dHpSO9m+3sWyWDCAuj
ArUtIHhF8xuTdVkm/K0N6DzAl5BUjWvD7Pwk5kRg7OzmcF7s2ZYrqRns/Su+CHpMhQaOHcrFR0ee
RuB8InRjgbMVi7jvXaP4BMCMukgyMIO3sy02ANqX93whTSN02g8OOLyR8vXnDYOtKffk4XTNBO04
KXT2T0/6GqgwotlEmwKRh697aPYPTOcVK1kcW+qoC9EAKWUcNpLowFlix58+/WQXUg/KXmhLbQ7g
tT7kLE2nO80UfoaI/tEldJ17Z+ZEXZs+FH0NtO2gv5bXdNMyOSAQyrxIwx22j81PTKNh34w2U5Tt
2DT+rlewbt72UCAV2Ph+cS6eJM67vGFAIKummJ69mUJz/LtRiGrlHVn/VXjq7hIyIx3RG70KZCnh
ms5j93wVT4/jv2a6HMONFHHbV0ycF/7BJieYVYBIoiei4c7krofaNczd7Glr1jL+KXWSTf487GgT
aGBELD99XSNPYUFYb3TxNcD0ee4N4xDBDZONpGpkzkrOEvNqPFStNjQkUK+gGM4SpqlH3Y4sq8jh
VRIQlUTm04IdW2Fg7+YBD7VT6xzralNCVdHwmayh82WMhrVP2E7CpPlNo8xzq/6ph/+epv1+iWLb
HvIcHL1fMC6/PtyiFaaXAwy5UmUoDvOMhBGtXpXJ9NqXlzpDMCLBfFdWx/Xl0Z02Dw+p0Mkh0/tD
pmpJpV5/XkXHpCVbLc0FK9rRbvxF8Ape4RCxQ0cfEvjp/Os4/Nud1mB61diYxo+/CjLagSbUks94
J1i1joEiOjfmz1ulwk6V7rtN+d/Rqnr/K9HY60VPZ3bLz6XrgCWGV2zsHpMWkzg2nBs2fAkzvg4h
nPyNg4lPDBCGJ32yRNq9b5sHxr0ORgabT8tfm6QkVPXrSJroRrjY/Yy+xktQs3xoZyIqCU+kFK4W
vCj6mKjoobYpRSiJqr1XPMK7e0GShkTg73eYhG6YPPY90h6RnaZjc5vpSqwa4PYr9gBuygADAF7i
u9CJkBBuVHFmRulNQqtbf+pr4tbWFKEKGZteGbjzXc1RpJYw2kKWwbjTDqv7G8S26GFFyVPv6s5U
jy7xghgUZysSR+tU8rb+7GoCzV0tBgN2evvFwEjyEDQ28G6PSXB5qakJ6Lb1if3aEgjKItaWJRMy
4d/bU2eHjmLG4KtXI8G2q+FgY0EPJ+I7mnXnoBVGy7frDU6Rdontu0/oWHOSpPtWQsStGJZ2dFul
r/qwbtCxhNO9iPT4ukzDF4uzom8Tvz2oWffx7DarLfk2AkwdwmzhVI5g4klVuiXyIOTP6QcGp7pj
N1Uf+djxXxUKKeewDuIEIlAlt1lhyeXokAHvI0w9rqc+h6CQ7VByPY7DJJCQ7u6nHx87fDIXq3+c
yenbamTkufLCkJHRbafj6TruCRFp+/a1sjSG38Q2bXobGrikUjFXr42IvKAdhPWQWR9ytJutiCR6
oEkOkCOi4b2xSb8RlrHxgq7v/JEQRylhynbwBChW66zgyfvpayKaurZwlqGofUt9RScznidlNGgY
EfArCwrUC4epJKRUmFAGFzE9rAuRfoRZm6/abSDWkqpDlUQS1iO8eZ6zH+uEJTsbXyiqS+YPuT+F
Qv59SB8BggLDj/FszbbNPnWuzNunYlE1Btb5WKl3/FDNx0Jv4guZqfQgsk9pcKDKqemfp7PUX0RY
o9X90uzJhYqBYvuCjjJuU1laXtm5/n5yUa+HDEu3hOvPwPU/l+Vu95FmdaJUjX6FD4oob4u/N79Y
Xqjn0bvA/scYOmeXC+r+O2FJD5wif6sygFmwejmJs/qgYIU4zBww9O1BzgtMoAMyQxqmRRlDDXgn
3GA2o9611tcF4QDRZsguKXg0b1u5hS/Vpc++6QMEK1fLI6kvUU7kUZ3eh1Agnkm3PL14WJAq91+s
TOhn3VRv7VWua3ikeo/754a0YcAgQQVM3PUt2HiBFpDU2keF3BX3qQcFd/xjEC7+m0U3qbqpU+iw
rSe0vXrZp3zR19qLOogeoFwthEJW95ro83flNENKQK79sNsm2zkeXAfxcC75ptcUfhnA+F6pdTYw
V8WxNazuWzd2jy+yuFfJ0uwbWQ5P1hypmDu14JKemW8b2mGsT700EvLl5RiePiqEpiAKwl8R9rX9
w6NY9yF/r1+NjJ0eG8mmYb7gV8IODmIWZCola/26XhM8M093sRF4Mo4USFbRsFtGwiqUVneQDjXO
7/J5gikAs+ilBfmO297V47rKgvY6T9ShNQvC7rr32utOinjNDhvZqFv+ffwOGo/5eoxiqzDNcnos
+2bc97laEdoZk2r32PYMlui6ijwpEBxyhf9jDUCVD5DD2f44hJrns1tSyR8T0ErH4XjNAa9F8MiW
cPEekrO5qjqur9mdeA4126tNA35pYK7O6qv+ZorLR0bKkvs15LJrYztK7Arrtune6RDXBorG/Br/
9ZNXjIP5eLAE0w0HlwkapWCSU9bPPU4V/YwACspMHI+ArwPjYvibiTucMWer02U0iakbMFg2pf+4
etFds0ToUs0UBMFv3uJHQljTDbVVUbruD9w4DcjflAAPBNuw8Vrsu+YyOgZ+Kn97z3KAiSX13fHy
ik20USFiyaLA+wgs/L9uXOYH1/dxm4IvwRfKPXgLwkOR1JQrOuPICqKSmYcOYUMejYeNeMkMUUHT
8wviqklRDEkLiT3vjD6uGfVgnZl1bRM1Djygt8hf1A6fH1Y7Tgd+UnyJQdB/fnQdv0xhzGvgM8U4
CWLK5LP06Qi02TPk//wkP6lWvHrkDjGWoFQzie5xE/WWBkQItLGOkLpYYYSJKG+a0/IlW9mAaY5S
uvrw7cf24KNaqaAdW1X8BJAS9iR9csao/9tCylUurBGx/7BYcMrMsVnBrMLlHpXFn7aA5T7h3LJ/
xHjqC7JbhxVgt74LQoULdjrceUWkQAIJBoYj6yP/vpNPqUksAVZ1dSoPpoLebFQUnxaohSdn3U+8
9OnL/xSEKFqw6UyNIoLgIvW5WrckHLGwZ1MklTX/ejSCHOXP7Sc1G+sP6ttNOylVJfs9EjRqJJ85
wSsmOHW8H7+UdwpCwDghkCc7/1irWuzbpHQvoHurffju8ccPYei15rvtvSYXA+MDfK3wu5y1cp6x
PvwhECc6iPBt2/tjvgRSKtHUdQC/OFiugPsK+cN3OE8N5+ieCeZAD8WHBom9Ldd71JdQRVtvysdr
C/Or7I5tT4zQyRRok+NBNcgQeQt/biAyIjWy8zWRxHLFI7eQJLxNbAOWkYFmfLhL7WjFGEjPiW03
bmtVXFRRYqPamyKD8LWStoCjgvMlnLmQ7DQqwI1yOq+86qxauKRmcnFOaPfaL0CYYF9+gE9nrZcB
kVeircQVutqILKnGvm6Rhj+GgphAGU8D/jD6pToaS1hwwbiNpsDsxoPE5/kYL16oErRtK+rOc7/u
aiCoJL5YTlk35XuxC3AE9JLPXpqUYntiGuQ6hvRy85MIv7VkC7SDgcKRSHUSr0ltErw2gnq7TK0Y
HwqqkWmUqW/YpRMCehBxlAQA/WwJ2naaUy9ggEGjECUcSOI6tgbYNgmOv+EQVQpJ22OIC359SVd7
+Idb7J3Aw6LeTfhTheR2GNrXEUwdG0jWlidYdM7fTpz2fgqD/RzPaiB/i/aa/smOR/DHMJSRFqay
fuRLh2BcBHiUTAElM4Xidv5Uf8qraCHO/t19XkizNIc28Za9Wn+3tXuCT+OP1vvV71HVSM26U8yZ
a6mkKVNOfqX7gI9aGCma5dsdZD/bB5YyjJFo8F0Uu16CTpbhCqV3LvLYUJc+8SV/Ao0UWGfg4cUF
jU7DjmT0KDUw7BRI8Ar+peDfApnJ9ep9kqobVK6iX8PfIbc5eRFaO5CH2+K9NIScZ3/2R0Hjl860
htnJwL7EhrGc0uTkKQyPXDvOpq7h6pffAB3aObU2nsnQwn9LNcnFi61JUplsUWmG1F2XoM/GMECC
dRB2jB5LxEl+6DBr0rVlp9L7veZQY+36zymXXUAUfjZCMEs70WRwe4yS+9K45iPSAkmOOia1dTyq
bCHSp/Ig9nOdCE2QOxLWyLGCZPyMXBS56uey7n89E3Td62JocGXwingd9SiXeKml6I8NM+Rvx6+a
DaxcD6DuSKoHRSwKukoKYkldAtAQt6H2YO3nTuNcGZxn2ndEZKeZiByurjfbqxilgysONns9l49y
21rtb3u/5T2fnvBUs3E75fqE/5S6tCp0Qiscg46nDd5ZZurclaAxpQp4SqwFq5y9Q/kistmCjXJE
yzxEf/fnB6G5Z/rlz+tW1YygFbdUjezzNt6C5+zMYLdtsCPNfPYqDr8RjAcNNZGKdOgAFkQrJVkR
yV+8pVPdws0b08deMle1Q1P8xoM39LG2fud1Te4f00ZOCHpd5GGuAIn37u3iIvGGH1P2b+sVAHwj
tuSFU29w/iQNhqGnvKWnGQ5ZcT9RvDPGvsSe1RDIqjt4UCFsMGKRay8R6v7uVt0L2nNdHoC+baur
xUDeK6HI0GscqvOeboWkzD9dLb2JrprZ8Q4eSAfULAGsZGnIQ44U8E6cIYwISXBMGYHTJS8Gtfd9
ZQHbz0BQ69BLuN2p76oYht6UScyVGSwSm9JJx2XnkHAPDhATVnSb4TbfMEK9pMtJfTDPoR13CIQ+
78Ck43qDMkImbV7pDHr35HhE+9EEXdWV0UeOY9RKj2S0MkLrjoh+di0vf8ZKYaWjIOjYYmV4CTwp
GzugOqwJYh2JVhdRfO8sKY68CoZQHgvimqtvgPSPvD78D9+wjmrcYM+OztRmcoToLq4Gb4VMU0La
j/beP4/pn36hqLDRzLCEm1yOuvRMmOX8/loWvFuJUa8xLmyT/YVr/mFMJpGMpEZx8Njf2ASloFSE
enHeqBTGYMK4PNv30c0qhsxvaD12Dlas948mMO3gYD1JW77GEnpOzdjo7i0uKObmOcaSBy+QzO2Z
xbHM4LPUVwIgQpfXet0I9WSZvrcJAeR5zrEd/kA3DCuiT/3MAKmxjOa934b+f07sRq1MD3TJ+Jfb
1Fn8n7z4K5gZ5ohXHJSalKpvVEh3kS4AhrXeYqbqICJXuivBZHDnSkrPgRfkp1Vy12JliiVgWiWE
FGDKvHXHImQa0s8VKNPLAGVtKwFntN6OJEliWFgpPVbJljgBUs7uHkdKTD7YOJmvqTu0PnC/4FoO
JqJWNIM+KsxtMWe5NHCl1MSxIxWkF0Ffq0Rxu5y9xOrwYKIfjTrYNeaBueGPEQfk/a+Bfjb1PHze
cO+CGc6kcfePMuQf/k45rxsyV3S3o+3vAy2oVxs3DoLLgA/b7uD2LNQjrnkrBUGpWAbljAkCYph6
zHcyr/ml0Lxvv3LoWacNnoh+hmQifuEKcIRQGnz5Zd2+QYNnNxxeCcfD2cRZmB55OwIbg7N9eR6f
Ohb6J9+fDEdyY+cZuHhITyDGr1M6P1IOXR3BTd8lTK99JEJOom3lpCMKW3Qq+Cj5YtUQvDoY9iC5
qptIgqTXHtrJU6jAcXyfOVebFJMLiGI3DALjixnmM9crovRCPEHpMNe2aYqF4PVSsFJNYlOEu3oh
W/u25B4xiPUI/C6sLv4lrYkZbOy5Fn05fNp+UxRaYoB4MHudyU9PbGjbOB+3ANjIyIuwMjcEeDq+
3XkoCh7ClCizRny4GNg3ooRX6q5hhHfIcbv3kNlkXG88T27KFhLYQ0ZY6ORencJG7qM9P9m8xkrZ
qJ+65zJrkMUN+LZHBTBr3TPi5FJBl+w0qg2kBrBba6YO5ouBEIj+IRUxAlJjoD6PBDhlsUe3QO+9
cb6jtY2ZnNNq1y79F0G8H1awO/e5dy9Xe6EtYP3cvfy4mWqSfsq53/zwzorA6V+hRpGYjeub4fED
NnRicnsGoLsu66HOh9l8p48gJg4hyt8xCktehiUOQzjsFp0RyxSLrVvD6WhNUvVyqO30tS+VUUn6
pzw2L+qn3bj4cjlCXWD6SvXrf+rVR4CBiSBjXFq7lYlz5etclhz7PTIPu/EejVUMn+FuWNaPgNCG
ZWarV1YYiYiZYEVUAsZ+6xKHU3xMCvCuPQvyrCiMQ/4lAdQ8F7RlmHShDXyk1PWdWd8TX18CIxOm
qsat2qtOnXy6zjLcq5oEoNm8UtOyOmMnVxaUEZp/pDSLZKN4YFJeHjTykIxDJ6sWuKkxG4w+AX0u
YA2+58siHpF+8Jg5kzV4cCTb4FURNr6XO1VxJIhVT/jdW5BRgrcycMbN/vW+7gP08CeyOOHvxg4I
pp8hq1y2nrYDEQEw5WWsstLsekFB9rmUTCaU9iZczxwyt+o73L4cRMf+OKZ0Vmhy2ZAhH6vLZV96
Hdyeq9bQmndeGiRXchHJ1fogkQCph+/NPvU+F9G1MB62MZY5KkHze+ra3ATXE+KmKY58NpgG6s//
wJPBSW1WI4s1LCww/lA49Z6SnlRRUmHEXvNp21Z4BzAVMgc5zwenVP84y8GtWWITs+w8lski/JBy
cQiYjKlWTm6cy3gMhZ1nFB/W+tkQf0GL7zXpi5zMRXgVSfTRQ1IhsXPX7euS/MtMgiCynzqlr4aJ
f//HOHypOM1Ff9mfLKRb9QalT9QWiQkPINWf5VXwWLiHlctYkL8ydS3mP7BMZmdjaUNUBtMNzL5R
MADS/eJPE+TOX/ZPhm6fyRkeiYIL2f2dLrZHXNqfe8E2LjNSkDgDFgRHJdsVxCfYzVjAFwzuX4MJ
DUodHhaxJyzvMOC2UK/LXepu1L9bwR0k3gWND9647jb5a3UVVGM2maFSmol2CF1Up1Ry4h+MmNCe
I/F5F2epe5KvOcwP0bUU4BB7bzYDgDzljC8XwAobT0+PEoyfTeu3r4uaKUBJOFqyxrijfBST1JyE
RCy5NSwK2ziyf54auHqeOBgp79/U6XTRNHGsemWuyam8X65fQtx30b2Qg4CgGWynjcKH7Mttr1Nt
9x8/rNILeryhORq9jQPvx4F1fwBTmb/rmuVU2/qVT2edLMvFVJb3C8S7f5lACRvhNLUgJWbyqMl2
USRlU+brhhjxJ16jLYj+fn/e5GqTDGXSpolQY5mH4fZE7Awauq0N7KA10QiJE3oSbdqi2I0Oud0v
xGfPNpPeJPsGHS9nWZ7oTuHizKqWMX4BjtW9uIeFUKIde7iEzq+4w924L8905FzC/8/hazp+HTkU
w4Ub6MOmWMtNynca6akCg/aGX6qV3MBXG+hLeSsBHNP3XGIODEFePEnMksyMlR/tqPwU9Cpwhjni
gYz6YPlcLXpMnwpD2U78vrSOjbNd5FJM1JnU4n+1yNH1+4tfsBqLrQyptYsjPrxQ7l8zdgQACmcN
yWT76ufenUwyNm3KBphdIXMcADuwzP1PJC0jtqMUVl3yD2ueiPpTZyMHeH1sbSwg068agyjhKniw
kD3lNiT/m8B+s8G/nd8xMRbX72H85dCQjPOUoibYzJ98nlTjd2i9kXlTEy/A6FSxziFbRNT3j9Xq
DmrGpJDE8JxOgmfaNu75p/b4uC/G13fj7+FRz5uGInCdUIF6Me6ZLj56R6lOYfIviBOBeJT4OVNq
rIr3kgz/6UgqBzHZvlpPPPvGUGu77sU0x7iJPbgE4VAOcY0OaCyPiReLsOX27qoKKE8YHJ1w6FZe
vjS5R+W0BsXhEuavHR5lbLIaxN/UPD42nUDgXZkXWELam1Tv0y5gbSCNFwXhLgQBaB+7qP2SeguH
3iIRq9/dw5Tc16VHiO+g9hna3kop2rA2Jhgg0qvjNxDtxcCaNcsM06xyASaGaHejzGUQu0PDFfjK
LUwyCZPcqkdEMZfpRwZ9wdBfcaeJYZki4v3BTRmK2HzC/aANgX22dbzjB/6D7gUbrbg1XTf+suwc
mNPO0W7GkSKtdRdW8/HfuuTevBg0SJ3zYBNxq2jaksKmWXOYpo6hn3uDwn3KHnGB5Z08mi38KZRm
GMWetUdJtRR6wqsXAck3+ExNcsiRy4SzhjEjOiJXGrwbvUCZ5EHTfXspGJU+akLf6rjCvnnTNftk
xQXOf2OUE6081uhPpPtQdNaW5SlF9+8uK+7KtEOpts2uxNZdlesb6692t40EtBgp49Q3oFFj7N62
W5TF9BaHSPEAKlVjmMkCLyhMZpuSNbOnDmDZnTeTNaAvtopKmTAi/AgKLLcsxGMqoz739USW5e+7
yQ7Mhk2E/ILWdzt9Oc0l0ADnhJ7QSI6T9GJYsvYgRb3FDQWzgduUbotSddR3wfZfCAUkS64Zs7ua
Jtj09hbE/AG0r7nqFc4pvw3TsGVFMx8bxISsWmzLBW6hPM4z4Ws+paC+Z9mnfI1Up4n9c53UuDUy
8jy8X6ZMFlJzYUeTdf7pNFqlNAR6vWkWXe59qLvLN/fAiq0LFOq/T9yEGqIUFos/gEyXGRkaiVUW
WE/XN+oBfcOzE8WtLVStudp8AtR3GsbOdtVNMX57ArtMHCh4rH99ZOzq0qRxVbGecU86CFYxsjVN
1TkF/s33DhmKbuOgY1PH3BWv4khTKg7ouPZufVKIR8jXj9Sl4rxKaikHGwX4vp+esIXVRMJ++aLv
0CzBoTOSj5p62Ty684ipuDNrUe9+u4Ro52f+URPLKqPm1qEdo5w8oNxHLhcl19KvcLKsLgZI4lRy
adCWXVMC89Tyrg4FwG+RVG33nsMy5mUCMlmR7SrrjYL8TnQJR63shrNY30ddEY2Kzy1hQB1FdU3L
eG4EL6vruhqdfOcAp9z0/9SlHaCkTYd9oNGeEkEj62n+N/khd7d/gPYO7Kn5FoPFJ8Gx+mA7jxgB
HHrTFQhA0jsVrnJUC7RF1XHn9tdn7Qb2P9MwYRRK4/tMs4oNx8n0Sptp4ydlGlaeu/mwaL8NJugL
L8EBnsM6lKxtUg+8YUq6ZAQlQR/yVREQ2ag6S1M10djqo39QCu0x/Q5Sfd/epsFToKecZZEK4wRU
9crc2Gn1rdn0cirWsXWK8hEdBNFV7YEqoXaDvXMYOxjdhbrGLbxaH+QiLoqbUj/ZOuzQyfzjZ1tV
GGfWM8KIkXgjB1AMcZi9tHTzgDTKphF0zpMOFPW9cwmPr8qVWWlNPMmz9kabvouhxEWnL8tOF7Ob
EdENTJ6yBymDjAFGql9aoSiH/IiY1kPQplNLQuE7SCbgNLahHlAt9DMbgxgv7Kh/11MKisG74hdc
yy9dl/1wQktp8tt005jR9CTEd0MJDQIi2MuHijFrmAfmLNh3KC+yR4r45xvBbCEQtjfzTQiKrHor
FSR7cUDWhLb5xlxh1Rmyy2e4hGLIUpKtBzzYXAWHqXTEHWwJ4VhrkVPedB99Sl5MGfrTTL+mwgRa
0Mx+TJOE3Fm+wvQPzG6Q14dm8WEMGk2uuHzCL4PHdPe6FZal8ajahu64jxFuZyUnRxFwuiol91OY
wx8ISNrOYeTRl2iY3//S+W9iPQGM08m7ydG5+bK/dqg0A9qpBI5KhozHgF4oPKyXv4i2JxrZ1hR7
qdGRYR4VkDzne+pjt/+ezM6vSe8IxBiPsbq/yxo9p2yFHTeoUxprNgxRlxNnM23rJhjQ/K5RzbQl
YvIzB4JeH/yrb50VVhwybJWzj9UaJtW/VTkKWiIv35L8Gy80ZnOrc/tNfOs5ocbqaujwXIr/hpHe
MsuaxHbCpkTGBel8Fa6FRepGAzyEUPjZndToA2M5G9vhbOht87Tm+HYCANk6ASa+3UzCHwS0KWzj
6H7zu8VqCHretDkWddyVlE66ddm/xhJx53WYcR+iT+jIYbEnsNwR6PNQSuYQYJuiXuryKR6h6Nc9
b5xNvplso1XNGeLeh47IxXaYxE4OE4yUCciJn5bDyFM316moSf5FN3zbOe6lOlcydnwEE4g1ui9G
rjQLmxSXdH0Mhkswm3QlXsk0/tuyx8iwI5ktEWdbq0gRzlY7cf0THYgBg7UMLKYbw612SoRqBwJu
nUj/GYMDr4Z58jQp9goKI+sK+dTW3zFK9Spg3D4zIN6EIx8uXm2aaOrRQ5yKUvIgbwfeuVgHt3IU
wTZZ9ju1RX1ZCzBRRZr8ZJjhBq+2AhF1Zf1D0VZt9uK+O9z1nc4f/gfLrjexHbCWUCOdPVfxFc4M
hKRskTgd1GfUCuXAlTswmmwYIQhYXAnLcP0uj/Qu7NPEP+RSGgFfncZ2/GTARdsyhrH9WGdSRnpY
SJpKxcPYp8Dj5ZW32inaWepLKWHSNeIFW40blkcUrL5RKm5fYV6LwiHQwsvW2GEU/r9JD0Nul2pY
o3V0WCpzgNB9VYIk6ZPprUFtSsWL2ElMdYsWUeBNMlNqQn5SRtV6ZEmnoDw0oNzAFMVDkQE8gX1w
ob83MgLkJb8ZgIRViStnGDFG+oeqo8zg1P1pVXUaTRfh4RJ44MvOOLjrpSER1QJICu6knFGCqymc
w/ZNYN8NY+/4gp0mooItAFrrpvK6SXeYfdvWRitvngLCJcCv+RcQMhXC+gZ5f4PlEIuplP6zngxs
Ge2E7Zl+0prZ6j/R6DqoQTP1AgDvfclvSVB6fXnBs/T3xg3iFM1edItyA5B8ZwuNHLipxieYyG/A
6ARM9ZT00WbzZpJx12FvoY+KnYba4GoDD8/b5QAKVtDAnRdVPq/jhHVktTyy2mTsENLRIrxSIZCB
rxNEofGXqHY6HWncImxJq/Zxo4WamXBYvGEA2YW+BqGuqjuuc9mqHB6xqaxBve/tblKlxJfwOexY
WHflvGf8xsiS9Kdi+z2Mqe+2bnNVEmnLcDKZL454NbkQ/XfHmnyYv/vlhHBGJZYVXbnNVif7eBlf
JsO81k9Kl7XPokUVO4pIeJs3FOEx0vjKHTj8PpEpsT9TKyZ6tSObEyZQihsBII74aFTR3C8oySKD
6C44s4xsSz9WAU0euFfJKLMf6VNVFKM/QbCXp4o74uimO4i43L5GlxBS3EDotr7f6MS9utyBj6Bz
CxMh9q5t1PblJagrFcZvkVhKu6rpbzIoac0NIIoU06eQ5bn9ZB63kRzo72fT/kZQoofYi/B9fJIj
xJr3KsGi0Xr1u9vrAwd4H62FywLgqgqaEG0OQMOr8Ewau7I3Qn1F+eXZD11Sm00TOPtDsEh02cv5
GooQXUDYwuIlSLJ5x/2gw557mvH39ulQnVSWse/hCXKe3hA79erui4fdLyR6yX8UIAa86jiEzDCN
adOokF7SEpoDbpEoVwV0w6JVwkqpUb3KtLwjmr1aTv2CMgp4P3c/w4g+pLlmzVdj1x58m2LNGFeD
/VYUD5cZALIWSE9hO90KC5oitQXbze5zH9RS7m8wH+6fdxCY+YgYS9jIO3tE8YNk3KkdeQOsFbUb
09Gmn0Ye4NqbXBd2lPbQReEflJpNhE2cw+ZuPJAWCc2sn6YMkwlotb59YUokEUjIqErBliXAnBot
RMJTiB42Gmj/oJLBqLl2jov5Ng6ThvHkxG5k1pfRItoQiYCd2pkYNA/stlueUV9XTpBL1UTW/siJ
WSrzn9UcMv3VSlnxDZ/87gb2Dr0/8gbIuDW4tISgHCaxJblnpn8lpJzofUcp87F3fr3tlDGiCqdK
APdi4IKWT+dEkXu2PUeK2m+Kxq051Yl3ykhRZ6wfbTBOoj4VFPmJSbA+5in3LqjGuf3U5p/0i2dL
OGTpsDZ3qFprWpN2Kabwzb0TyXw3NKeN/IPoPysKUvZic5gFMSqxZQ3TQJwiXWLEeoXeYOIA1xI7
rfojg2hZL6IdTaO1sChRNKXReiig9WrFshBydlfWUeCbL8UXlGsTK5sMX1nTpCIXF7tXh2WpqzFH
aBz+zBEKSTQ5e2IjNKF6QyF/V1vGNOOHflQjyKTU7gRu8xt72J5gnWcYoVZYeF7B/fZirKrjm5QZ
tM99ICNJeFOz6QifhjtoqicPhxkiWJIqaBRmog+gLtGDbBhYcLF2VRvKE5UObg2K4TlGvSHVsFzu
WbJREVvI2v/Q3Qn8lLXRAh+BbcWiN74zNh24IeJFV3+QEREyF6PlPbb4a3IHfSLbDDAXZ2K0qAuh
psxAnND9fGf5JbFPkd9TyDsNFfgU4otliVgoJpX6/4o/ZlVXaF/OcPzuNrrPgVHrsn0UM8KLAogx
Ns0denFou92rFb38ufLGT/zYy/qF5+ViCVkclShWQH10GzOeAHnrWBt0Eun+ZM5/0t7dSx3RM5xj
C+vfReLjHOfo6l34rndTm0ePVDW82dKRjf6/ZtzvseLPqRxeOWGAyuS5BXPXJa0DwbcLf5D+Gj8b
L+GPLqDiBZohgw/5GVkMTQtc9ORnkh11ATUfWF/+k7N0GKVR2i79j+rr3jezvX4uI1n3CmUXjbu7
OOdZS8OntyFrc7RgovIWRsi1tqvo+oSVZZgroRVVi3wk5uwBdhHlDjHUxlmtm2pOcVvTqiN1Wm7G
udBQIKhER7L4wetJtRwQCZls7kFZ9bgAYifUXD3w1Y6E8+8HsmZitfU0UBR3mVt6zB0kp270eFEk
JDiuSuh39fjTSFNvyU4HxO4C2tQdt3/b48QpKrRJTzXvZOLHC0jSU+0lNht89eZe+UXwdLsl0gl9
CLft6xkv3+VXWDrxTPxyHYZRraQw3wDWLgvy9Jvbv+Y6d+/l2Fuhze/MTD4iWA3KajQ7CCmvf0W3
HnpfjQqHLV/n9tHLZgRZ/1r+AhpcqjTE+YoHGE2abreirc5NXkxOV7SEnp5KT83xuIXN+ZSzVJiC
6K/NMp9P2Dxbgo/mApAor/zPiR+emA7kNTEe5g+DASdmMSVTFjxQhs3W0YLbeRB34zQ42fQsWA00
z2TWMH2Gpn7t/UfhHDU4ZIrR3fPiMvwdUsa7wMxs66MpP5mkKlZTDWCXvVUNXgWW8TGuhjiWlQnq
9GyL1yQmg3/X0lf2oWWZiDE3dkgGNVKrFzG77aSC/29Ezij8jGeTMYjyis8mNy5MqJw01Nhry3VQ
zOYqgsKhmKxWSUhSjAQ56fbZ8fK2GGnegvPCi3Akrlt8jYgNZPOYIYG7ADhLVQr1NP8n9J+m7mxu
e35cWW1f+9elHT8qnGXQl91L359aZwCswhwC7EFC4RzX228HTYn0Dcj7XXtFz22nDQCcwzwJAaUs
deMR3PojqxGmeKap6DqX5OCdtPUvvV2R9Ck0spXGQDSEFQyiYa33Wgdz0mDQd6u+57ZpZJEYoc7m
YK7KsNWdmULrXClaYzjGblLm53LKehceduChfjUxbwQdU/iRqpdrTAq/NBIXiTi9X/37nzYT7mLu
pD6FnAzhyd2DSKxol4HKmI0iLt2DNjRSfLn8rcipfIfGiooGqsqg+pn2wasS3lo6albXmSIDKfGb
Fxe6PvMPtcu6pPo+bqGVlCu4ezQgOGkKFRm3cu8MungJlujxrzp4kOku2RZYeLbFOoUHsfRnnj8q
gRBGlloC/31I9x4j6WljLsu8uRCkK4Y5gONd+W0x+c2jfcdbUfTZz0SADi2XOQ38Proc5/zHCVD2
PZo1HZ8YAML/mhW5kPLjJx3EF7KChYGDyGTSvtmKG4RxI4UppNInAT1ZmKt2pBorh9V5b4JLpm1s
E2lyvubGm/A4AlhqB5lJC7D/AUbF3koQL4++ux10fOTNL/Jtm4xlSih9sGhydSI5jJbyWo4iUFrl
2tyz+SzYOXy7oFrBqhMKKnpsgjM9aTfhqRG6EHMjgBGt+qeCa/iMzdj/7TXJ9eWzF2n4q4C9AOgv
JzpsVmSuvpqJvwaanjjk8ZmiMX88ADt3XkaupS4ccurF3yWUeOTuhIFJFfmWkNQOEL05DsTktI4F
qNlCSNkfZWAdVFz+RnG/Buignjaux2WjfcjrsoG1c4bMiL/3aXHngAbbGdLkUDyYJv9WELeKgdPq
t+WfkI0FNO/MUiyo6QnMjlqZaRTrMsytgUWztGyHeV+nLHrDFpn06+aMqVYWtQmva37zzgZoI8Fk
jbv5uclIuVA1vnsDkbnixdsDsIq3VbsqfGJTPxfp+eBunrM9Lf+YzCM6pvL3qnz2nWhfzh5XTC8i
M0t3LU8sxzbvaOv/WRMWCKftnsvLt0WD1HiJ5vo8GTKnRhrvX7RyEyAm6K/U+pVMMcJUmEAveRuW
ENUCC+tqH/rLKEQIk3felFJdmto5PAXDVUqwvbM4udrrM3qhvqibuZu4ZOYntlS7ShvmbJWhqTSJ
QRi7+6TrKRKlqryooszdVNJXNXyp4V/0Ycw2UHhNPW7JeYmNn7l+aGuhipSZGCkf4oPEjgG+Gsi4
TIzsvCMm/weQirUCcoAXamSDUVLF/7BOYDDmfqeb+PA23/AnNUkEP4uJx/SHh4RZtV/BzWoD/EhO
d7ogb/q+uKSna28d0b2aScxXCLMyjIX2it16AHPvypkul6OZlZ0kXPggH8i2Yyg+KoWJarfiX9D/
wTld6dOmRkgKMdQRqColdq7OOR1tQzfd3h43gpu+nzqMAhXtqco1z1TCt3NC8foA3keBm16RZRWb
G/A0uTUVTUPXOD7+r6u5Em+htOiiiOz4zO1P8vEZXVqsQN+FxVGxS2j6xM8Rb0abCtZfw6Li2XF/
3oTzjica515trGEUfCl9PLQ5YVvvLSKNtj1TS5o/HqMe111KgllZep0rhcuN+ABRsTwYISGLxwgp
vK8nSxu99YSYZTome4sdDAH9oomlr/DvysstyfvWurIc7rQKfSfgPZFX/MqMNyzz4ApUUb+MKruQ
Y9G3R/RGvDEjqJMK7o7gu0paL1y5tsKOvUfmcgVNa/09HZfCzug+R8MsI08L6n8MAnN3Yjz/djFI
7114wmDDk+AzkGMcdcV+U+nrxNPn3n48dtQTK+W/D+jWgdZ1xNZE8fJQIw0HejDjBU8Dw1rz89ZH
4PtcOH5yfTlPV1VjZzC5Hlmbsotv1SLWs5peYb24GNpr6DiQv3+yDZRvCSU4UcFxRJQtyMgR0hdE
XlXWbkLjD+wyvEmZds44R3NFv02eof3z6uEPCdSPGiRqMRBvMR9U2oq3bv/7S97rftDPQ7XXf56A
uRrBI7ZXlnvsM60/9kMkYpbWPxgSADd52oGHRJ+a5BhoDKNBbaE1xxgwbpMw6ZXBiad835hinwt9
9PlhT4W2ItkgvoAIEIqah6Wya6r6FNT3IxXe7Kr2ni7fKkzqZLnmnVBOrMVAC/Y97Tg1eah/Mk0v
1FgdV8+vBmqOrevgb/7eluhhHcWSs3zYREzDXeJx+IdcZZ03TdjOtsRHi6JRvB+AwJfzEC79d2hW
xtOi+ZsGJpoi/6dnW9BLhlF7JXWxTmGiLuEKMfJeVru4Cpjnd41JewYmhOfe2vfUoPQeUUl2q4fd
9tvMQGB+opjKfNY2AeyNaQdOXiSxveDdyFocItx5+zKUg/DYZ5Ik860uPjTuHFpKk932JapZowXG
iNRMiVt+xmN4XNqAm83D2S7loAAqpdTB7K7jPrdHU/oT8y0FlX+n5TilDClgoFFcQsvqX5Ty25gU
VyPHji0+LpUq9ESrrErY5NTm4F7YeTK/Kkk6JCqBlg951Ql+9m7khBCVnRYs7wRfq9uQeP5t536i
1vDw8WilPf2DO1Nq3mw1t4MRjadkzv8JyH6uwbLYDtO+7LzXqGRrKPdZNPn4ddbtQOo2k7njsP1s
bvnUOzLi7+XzyLuf++5X1x7iFK57/79AZe/5p7ycAqa8zFXtfTKj/4f3w81EFooG97wQtenbwm61
qDdrPc3o/R9U/R6KOVCNnIsGK9Mrzi+mSimu1g6Cc8/v3KHfH3MxJCVLHvK2OgPyrQci3cmGBzOc
xYS3e8A7qhyevuetszToKjNk5c7X1piPu91/POp5VD47tIWAr6R6A4e5/2K5OQ2B3OOCQH0xmKT+
XPPRJzG3UwT8nYEJCv0NlpIjH1RhJeZ1xad7CdQ1h0iSxhFd0naUWCLe8A1df40ljfIWHiimIZiF
wfkvW6Gvvn6ON5tYkjNOr+pRnmFIAlBJ+U4dYsSWRLI+NADU84lwBMzfWAIzA5PSG6fWSTlzDkNa
F7pj17xvDYbbjiyFva51CdDtlQN4TK6kquuFg8AKBo8eSA+vJBbSlkmvP1I6sSH4ITDvRod+1cBF
G0tdP7dgMK+oXekTqkkrWXx0bMVNEV1DsK7sJ8nKeeO8kXw4hH5t3X+9wjQIc0CdU62aVNe5A5KD
jsxPIqz4nbQLoDF4S804KuyMs1Y5OdPCmx9miRJy51t2feSaNW8HWpaj3OqavQ1IMry0I9DKmnwJ
rGlr2xTRQiLmkPQlYacaWMMbyvg57dv2tvRXHe9bDPW+4LA34/bmTNvRTFcArjQy0Cx1M+FEqfVI
ShJEkymdowGakYy7yn4QHq4uMoR9TCxch9vBC/ZUb66CYzA2+N4OE8Od7LZ5xAq6c/VmCvKcklLa
BZnZcQPb89bTBlAOtLbpZGSYN9ZGYJm1rSMg+m8OYF1nagbe/NRdi+tqmsYp17lyxLBxPZPPW7xc
DkDdwMxIpaFyQEApWqMS9TOrH94lkZMqOZSNQIa79pnxYRju5whN1SynUzcmkcfeHgN1PdT+AXvc
GuYHBb35CidGxpcGhKlxkWbshSg5qA1H2yqoDdR89OLBOcUS9kM3AR5JI0s7JkDJJsz+OdTlRYDh
/p5a8hd7IpJTPfXNlAzKSpzEBIqZKoYBW7dhmYC65FpYtH+2OxY7lHKLVcntMb8qvddvlYWEMF7j
oBAzdy4strwbxuZPnJkn7b8b9G8sIC8YYOeygdaNSvZaYWejRTnWPk32mmBGA40xK9dJy/jvUPAZ
glM65T47Ax2osS+ekQR3ZHdJx43lyd72j5ObqQ0YFoiNw+xY9iNYjQsPFtsEDGo1TxM4VwBud1qo
4Od7uoWjzA7hiDBKFSzcvf3Pdt71zFHD+rhoSyr+vW3gCqJ7JD4iyx6Wt0WJx0je6leXCSIDspoq
kz/g05gqFBiLsbEI0iNdyibLixv3fvY6s/mAa891l0vqJGWJh3SVrgLTSbHGwlP/V/UxXSxVgwEs
TrCcjKtFXJpNxjrsNJjHxXhemyPAZO9h70y1BNHPWFMq676Iv9Y429MTrrnv47yx7eMmW2v2CNJ0
sl/VbdRj8kYya8zlxQcY81wesFJKJoYQrxp8o5I7kquGFjqgRIQPukm9KQuEjPPaHF6/whduUGhv
/mz1lhjCqLxT5y2Vzd/CaPZLdw7hwOr4x5zru6iw+YOxtQr8B59LpDV1KmM2nRXets1j5p4n4mW+
PO4IlOeT6d0gpPzvjfahD8tbt5Mbfvg8vVYvetmuDEeT6W4ZFg6L4VJupIjmribCRGtTiTV+VrPY
N2sglLvIGFUsax589IFkhLOUF3/Ji5JyaS6GeMDMkw5h4mZdEOYZxOw+BcpLcWjfd+QhIiZNeKPm
6NfiPRSCCJRENiSyJ3MxHXf4Sq1KY218fjH6oiyg60mqzTkC443FRWStJysfCgvsn1XBszfZPSok
HXBlmaVzN0bnHcOcA5S+bEb6dM0L5P34xczm/VENuE7V9BPPybBkCb6I3blxc2hJfN/K2VjZPPIu
riXwAM3D2x7eRi0AzTmdFXWlOs4ZrW8rrRq+Tq2wWCf9xklozmgtNbdBex/Ffdv9rCO96eyTJC1m
yodmuTdfYWoIxysiCT2sLrSSh2fLjJ3Dq9gmsy7OjfSfhfOHULXMNvQXX+wt9B4WIXYNbgBSdZ5a
cQRaVNEYwmA0KCGwEtGu9QM2CoD0Gcgx82GW77YfD4iEcuUXXbQXI7eZLt48oz/4XraLmILFoNue
SEanf8FE11EZyitsBe/Bz6T0EHYXXzZDIa6Gx88h4At+V7pZP1+IrTRoEC0x7gCOaNHCpFNjzyoC
nsVB1j91tVTZnkUF18nlGanzUjy9MnXbA8gbv/3eqE7D9H71bGjbn6smXQy2ZytqxhH+dyyBet6z
zoBscWRGWovPdUENObZ0OkzTiH2HwnNtv2YoqzrgIFkbbcXEVwwQo/ITi3xRQO9unx9jFJ0V4sWy
P+xrpkhweeqwCVscaHfJhi0G7RPCrLkdziSszYCySB07Sc1/qeBNmsObaSPq7ykvw880H7PgERyj
yesKEA0QTnfydv5jV/GZWeemtZ0yoILgukpo/D2WkXCLFloQOcH/fBQvaEgx98ItSh/yi+PonVw6
rfCBb/1aIAZBI+kl9ka8ggwz31qb1yoRrDcVo+b8cJ8zwWZ0wPSI6Q7lIsDeRPYaq6KJoBG0bE4/
Ee70puxp5AJCkZ/NOleq4lFXmWgFHj96C/7d7uIonKzbvRJyPF6UCRRdzRcaMlXBiuF3LhNMoQ8E
5lTJribT4ASzGP3U4ljG5LIPFQCjMsgGKWI3X40q4k+m1T85nWyTev1dUgKspiwWoo0kxAm/Necz
InXkbLFMIJFlK0ow1NaoZOlKQNZK6wbEgVo6P7a5VBwXAcnUN6E4IUfqLhkz/Yf6i9M+iJ5SddL5
YoIO3Kwb2AYnSfmDstlt0YJ5I3s7o9gUeBTyg7bLH9wzBOx3mhzRy7KxwMSy+nxYydAW4mUQfL0K
U2g3DXFCnQKve77J4zQMoWnnJmivZt+qaa6A3s2tO/zG4W5FGfBgCfH35HzJXPvfV1p0wsOJcTWI
335nAZfPx1te4A9OcuZNQKTuPTVfDfKz170Lz1ZB8ojEiSUBTGvCQYokr629RHEzHXs+GxAQ9JS8
PQMp7h7U5ILDbUUiKodKNkyUzgJpNrsbvaIXlLIJwajX9bIQEOnwO0hTDOcLuILzsQwa/i0lpiwt
lH6OpuGIFMuQDT7monDtn63XYqcX0NoO1fcrnDZtPAlI+scJYU1yYgUV9auGXU/jN0SR/OJQYuu5
S6xTCa/sGDIPl7sig6v0kXa28iHMJldDd2zHo6LzN1+k30TUlpcqjoYLRo7Kt0dSVoPEuryMScdV
QzAusqQfFpUyX1Rl/ipFVz87m/3a2PRGA/rZrt+D/gu0DRgO5MhtMa8oFgxGECTts449kYJd48rJ
KNCTgrBiKv63zSz73dvf/9LzhNjv6aoms9fN/Ux/W8zTtzNYEARjSoA1pMIivPlA5iY/ykJbjMV7
BVaSPFA5l3s1IYnrz8CX1U2XIqvUlH8hQ/s9Pw0+9MyHnQKl+Y1841e9eEbOS5gNt7vupgHXxkBZ
wckcPXvIpk83kqIlgZTGayiekCQlWXvuRWNPjGrSPBE9TBO7drEwGTdzf94455WeADGTQyi8rWnM
XqBr5NmvcWeMdm9HynRW6NpZ6UOnWUTYIzeHIUttDq9hU25LGnjZjlk7rrDYAWxgz3lGXgHb2LoU
/Bu6iNm5hG/ZABBTYI8qZo4mA+r7Kxo01j9lu/hePHhE5FgvRcK3GoZkGP4PL/XV+tPofwJFwlHO
VNgpvorhi//tN4goke7QWwM338CLxp4nixZHM7TxjUFDa82ZwbHzMWG0K2WKCX1BbDsnB675mP/2
0T8y9+xZzOhmML5BZ6Zf9NVV5bK+Q7AZxovOF60DipwZmyhLZScGJECUku6Tz9DBKBmXEGeyiKXz
JUHvxLA7xecsnPbxLUsFzFSYE8chI89sJoKhWv9EijZncKNJ0kfbtj+jMy9F72XBkO7EESmpzMDS
CkKssUJ72agTIJ4swmfOcKUPyi3RCKUH8PIkBhWRj4xnsMZJ5SgIayNNsWGPufrjEzJOck1IYzj/
xt8+heGHqSd9mONA6g1yxs7slZIIPcu02miqoOLkKcP0hbf7TX0fslzqemiQKrU2AOOA3E8YE2za
2QTqdhX1FFIF5F6BFwSINKk9EcmFvbLDa6YoD+jv42HixUOxrl8BttEPYuOXnHkzKPdjUQ8/28Yg
cfF/+5P3Eoz5mIgOlFR92HacezMY15g5VeOlsKdV89phyuevs0NlFzM7kLnT5AESjM/0xoJ3imbY
rMpoa+WxTZk9PJjFo/zAkkMiTYr96f7Nl1FNywZjj7KffT2S/fKdBQEXrVPIpkeuKxO69g92zBPW
FJ7tryu0522dTLyqG1AjXmFu6bwzUp8RZEZKLpyb28oVxSZQeDVtTAmVS8O5RU6aj2HHIurc4lNK
3IoAczKtX6P9WRdwenXJF9OJWCBhQ7eZKj94VPUTQnQ4A7ULr8bhAYzL+RFOswaV9wpAXWEuI6xl
D8ImKUEq9YDE0IWyST418DO+3S2USEf6VFvLC1Z+KD8Bm4ZUVNDw2tlAsnUOdHZW2Jt3UjqNH1sZ
AlDZZ2sDoRtVcLJIBwUSYiLAyc6tiQGPSI35s+ifK6Np39prXeTWfjt+poaKbHPjLIUYAnOd/hK7
arVU3UGOBLomRVh3redzo9ui4ImtHZui78/7hPdrRYqSUOs7tzrF2qrNZCP1SV6SGAZ4HhOsUXLZ
Smj9aMbg/W4GQB9Bbn3Hn/SYWkTdeSfkFfrZk7fh1fj+OPYTtKW01SDKIaB+kjhijCja030I4W5N
dJJC0spF9RCgpN6owkXrhVAECu6cCt8kDlStercW4T7CVg7y82EJAj3v5Hro4M/Ym1QmJREp4jbR
N70yAgTCHYC4BJcdAPYWBM7wybgduTno6ARldN6QZf56QHCR8XCVLIzPHab9UaynHJgx+33A4FLS
xPdGEIbBcsAvw5icYa6Mzl63XK2py3xazw1+sWSufuBBWPh/zR29fKaR5ewW55kPPH1s5n83dYu7
OJZqofvB947H3RrAlNxZEkb53D6j5xZd+Wzl1Q7ssufPYVnqtFowVvNFgSZrxSIg6ZhdPiu7Mj/c
5zCYwjCxhVclMS4eZVFXNL6MNhRbEsuwS+H7NUvJCKH+ycPagJYgNZRCaVxHeOmJb7HFMtLaS58w
TfYo1ZfTIHZRw2EcVYO147OhuiFWK0avLABDexT7p2AWm7b8IvnqOoEnCeGyaA3ooBY1VuDy3OSx
OrmkWl8SaR2W+fzajAxDwpz9NeZxlDVxC2XI02/gM5zyxxe/wDW/5x43ymXxCcbqxqy5jbsY7BWz
+tQCAE1AplzMz5xhkX1Bn8/t/t0T+FDjZsdt6yCru6c+mi3ov7UI5oXuSX69BPWM2RXZZGuzYgGm
n40Lhbi66Ei4Ayi78zIaGg13EhexdDj/2y0rqhIdCRVBZtS3OZ3ltyUohUeITE1RiknnzOo0EXfk
6574a5MYmVvfQNY6fu2Ava5H4OorRfm86YH6ch3IZpcEuje7k2SoDjAMcwiQtFeaiomiR5asyWmy
e/EK0dvZpoYFeI+o28wyhRLGvcGHIFpeZAA08eNblqBcTEtzKLFapy0pxykLKxBz7OOd76OeSUSS
k91o3MIxsaEG3u9i/Y6KgGK5b5e11VVgVyFl3Xo8P3X4I8a5UtgDsCaRUp56YUTquqFTnvNq1xJv
yve/+mt7QboJqNjx5lKFmxlgvrul+mPXS8lmWuWX1oLlasYwaGp2Elvg5nB7iLS5AVGKNeOI2A8P
lLX6w5eR4n7Qd2gLa++DtFkUS1v+UC1HPnaMfbRa07FeZg3IoaRtNQW+juFt2qvDw3oBnef4rQQy
WenFioVQ8LtULRwUQCLTgYnMVnSUEZS4R7reWpyC+ZginTJAb4MFIt2Yn0vYcFj9XpWD9Rt5E5Hg
dDfhn7PHn8swbF+c77ALMGaonDePRebKQFLr5RXCzpXyrOAydj8F3moTU4qpCBsyxo+brbtayp9J
o/HtBW6UVdGmegQx5ZuTgI6cPstcp22rfPirsdk1IHPsU2asjPxVWsvdi6OsLXDQKh9Dr+cOh9bU
OK/ividd9hw5KTYvcs1/v7X01UISDLFz+F/5qJBSEI1MefVFlttd9KUt+p/Pk7FQLhT+2E5MgIAQ
Egxjz/WXiUwRicUL55WcSQGlnvq6JGePl9QoXsTdH8wljw4qXx31/52VCNNMtTrSKEEPsCs6y/DD
7QneYzSL408yChDPKs+U+2p2wdam2tSa0Xkw7Wu8K+R5UCzEI6EFUvFZn43v+YndSJRRS+Lcjjx2
1a6+Inf4II7IP5E+vkL/9bkCcBwCik8EZsdhd03bfQyX5INOTKbqA//NEByf/iYzLh5/JHDUepD7
/TLzORB92/Kzg3nn3xqxq+USdIm73E885ZUtAnI+dkuFQ/7lrUogsjuFS2qIdxxBYgJgDmxcIwHt
cV+//Mw/w8kFWZ1Im299ERxoDrLdHygnxtVZAX5/qqZT0m9++oPZniSSAKHsz6EAg6CtQp7duuCR
u1Cph/+a/DH8Grle2jWbbGlVDvNqf5pcAPWmblsHEyRXtLpJr8f5UqSWsz5wHaHHCi98ckHJvvV1
T7l+sTFa+kRmXUPHqnR9i38av5TQJsMU+wt88BmdFLqKkMXCk2e4+3L5TS9da3ZDf7bRPHMwTPai
HLWREPZHEfWfzOGhaJEBNSCOA5sTZECu1eEPF0sKC/l6c3c8rBIMbMy4Xfh+1DMkca5FQVr0SJBF
ekamauOBIr/rm/kdYyC/B1ytKYsVpuoVGDoJkWL8RFyVQnDhFHrwpQlUCO4N5VMQv9OY8FdDXe5b
dtUEDvF7cPlgcvyehHjpXO5ppn9uQ4vjPf+KAA6iYsoAuXeT1CKHLQCbz+/KLjaU0ZsL3eNZTHeF
NhjnWL6q5o1Xm+I7g7nEkV7AJqeNdZrN8RmTyJIp4yqHxC7DQGX1NHRMgzyS3URrOjGHvOkZD96Y
TF2Q4OAl8o40yu/pzoij0Vv0J2ko8So6gYjRbynHI9UrvOLzqU8CQxJ2PuAZ0R4S+Ji704ycSVOt
H9qFrFAL0Z9XQrp903Bbr9yw6l5d4lsg3iQio+ffVIfahNBeJPD3cznZ/ZjPXeP8z4IAPj4i78PL
r9fdOhhox82jRtt979hZHW2P7ffJ+8vNSiI6FqzdT98/MbO6OyLwRpTnJjiTJNVtkTXEj7vhNbXr
KIvz8XbULqsj7gBemotEjLVxc2i+By99GnHYSrKCED20pxBWjWCkmxlVCStKL8gJ1TxGeybmelcN
YzRWdKitrQY717auM6icTQj8I4m4g/dIW82A++K+JERJtKKxQcNNIvHCCXV0VRjuT34U/mPZEKvL
VNDpp84ku9K23cM7YNuNATuijyd3NJDIGK5C7zoWSNrFeDzkZqROvsSBkCkuMjqc3HEv6VzsuQ+N
u9di7W6HVQmYavyFJ8rpAqd2nQ4Tdojl7/UUX6HrlLbYByuZ/GonBvw+khWgz3Ts/uQApvy+efFx
Ill/2TdDJqXlA2bBis8I+FtkPVussknfEg7rrSz0ZUC3TOzbfo88ju/ZUtyO0EC+SFfedsiyJ8gk
ifaMHHbMkkUYApqYy8GdnKyV3Be0MZxnXeutc5vI0HnptPbGf1aBRVH06NAS5mb2Ik6zeK4a9//e
mv3HmjOkK6aOGsySw0vCqPPYEuTTT8WBj7uvkkPNKbixJWdbcnF/kMbGdYAnxpdNb3ZCzoRLsxVE
T2WsBKDGPrRjb7ghbUj6bDOYyi1f5eoeUp1OUD0pA6ApraUZI395U+KwliYMtEOXdtz1NK13j76g
FgsGWzwoqURZ8EaJqrpOl+c80ZnjoNYV2tAEMcT04ocht/eIdDyk6ZHMmk9wZqIFtB1QQw5/PMFz
xH2wceTtEW7BLt2oLXGGUwK/VofqZPSxfpAYaWjEj1poacV7v7KzwcRHKdHjqQH1u2x01Pck0qBv
30lhg/417AnzmayfCm6SBFZ3R69AJtuwQA21vJgXkuAV9YbNXHCqzqoxYtxBXjZu+HwWc3ELF0Bt
/x7asIM9U2B+hEmipPhJBhmroGTGAJsBZtiCvoW41OW6ABpilUEhYu1eGsBk4DfkH6wZWLYf68ck
iV5CQlztFTbNXEr3vka23zQjJUE78umPhyYswvmaaTIvEbf5YhJpMfXv/JiTr3iNO3NM4LcxzIdW
eaAg8TQJ2A/wSr6xvj0MVeBhUIxiV0J/+2vPSbMPN11FyVII6YsZbDCTY9HI8xABUdEjyM/nX4rc
r61UnDR5U0aERmhpdp4zTmTpQ8xn88+RvCxrqKz/LFMLuKaOQFZpAQcUVTO0ghLk4E689xnjWLAN
Vq9zwQrky1cIpvXlugtZjv5AmT3JNrH8SClhCUQ03IVjd4yTFTbCl0tLEX7CHeLwqyuUAnDm4gWS
hYLOLueOGhU7poRzwrwKizd9P9IfHyQvd1PivkmUR1orjWSz0oM0w1ylMOTJhstQpUT9gDO0ah0y
1/A1R1JwTcLr304NW3EmJCoaHuAuFrjwCzFQk1dQF+zcLDUl3dGARGfT/oiq0ex/7IjO9usdiOcJ
6jzy+GWdV2NMQcaGVM44zrIz6ImQdrZp/LvR/GxIJ5wamRzGjgkNQDw7yCbVIw3Iakg3bVCVTdhf
j7Wtmgl4dmPKcOpvaOT7bhPfL0ylI588Z5F7h1LeFv94zwze8iUNTRtJm5iTjG88biqs9TDx+dE4
XjfSzvX5NiSGAOLVvIA7+xkFfmlmsdmZPCmoBZor0WJRMzuDGysPyBBt4GxtQxqtmfGslgg/+Jo7
+7HHx2gthEWXpXHoSpYMi0AssqSzx+830W63GFXiaTx3CPHwWUJxoidEVkov7OwLjDTJdlq98ljh
ri710ixw7GciXZlJrN+6jRLCOSjp8BtGEyihA/BzX6PJEddhcnxTjna6G9TiT1X/RWVENL5/tl7T
1kZc7Yx4DHqO/B4kCaeGgl+T4agMo35x8PWuh5f6ntnOk++nDUDdWfSSXd0y6owJWI93kf2fwL2f
oh7XlURFwizGGCXr+z4rTnXOJmdGKGo3QUAfh72zK1o/C5mNooktbcxBkUsqIxm/Ji68QlNZuEuC
R/kgb2rClJcog4okM40sNq8JJqsOnIeSv21LTo3yRw2HVF26HJ8cZJiFd/rPklB0ORGpdv0MmpjO
mXThYlYNI+3FkV2i+VBLC0o9tKsvHK2f0K4klDu05UssndAxqwJAOyu0CmrB/dbA0p17n+NjYMIm
rP6TixpFfkPrNufzbSvqSDvnWdiPlOETiRCddWii7WOuFar4L5J6SegnwPO/DKWzgMzTeVzBsnc1
tpOYfFjIzm8Uv4I2EKMXKlVByD56SYZGyB3XPu+qcsKZyMwLUASQ3nZVe5ETHCzqi6jfVPUqHAvz
cfXXKfiF9bL5MPZfj+qMGTBWtZvdBYDnsE178ZSpP3imU4Awvcq1jnrHZZcWn50kP/oj4n26/adX
SAb5hI2GvfM7t7OzQDRVniaM3wYfkt+gW14Ck5Vl0YegRHE3qMeCErZ3UuWRkKA0+RJfi2laQQAO
ujHsrkoVwEm4gwEa0pcAVQhB2xESlXFvYW+XnhEWIIJffCyBlHPFl76/v2dNKSo/fELsrXLSyIRW
Hlzj7TT4meQejP4JkvltBp6pM90TjcW7zANDKaTZDw3XgRWu9TIqWBH9UnZr0yNbA3KpojwJvm91
uj28G2fyP6MMm+NvHXwKNTIaKdjw7flwtvXjWfq5nEkDIXuVgEY78UXcaC4trFu6Vw07Wv4lp19Z
VO9jVz2x2emWDDZ6Ehh6/U68xlQjCP+e552o/ghSUmxumJ+iZpNNQsQ24oL9w/2AJkZY7m9E38Ex
ot43RN2mQGx8kCkAIE73gkMPx4WSiMN+j52e4qtRQmWHnoxy0p6xG3ekczISMRuOftnFrrbBPKBc
5uaSlg7mouUd3iqYPDarK8pPPgeMMmqaw32Nl7XymhXvo/v1rBcDsTdILPm8mpWYdy8b8yLc074Z
xUWbsLUDo8CcZKFqDIKx1LSt6wOSEjKJ+vcWVQim7DwKll8R/64dDSPmwAMgkKOI14xs3jZhblkE
BwdNefCQclJ+7q2zc42iJXG9xb2qWcsbj+LpsafPSeeHT6GIlRfpoPGIdonWIW0AswtsctiSqkQN
eCZqqqjhp/8e4k4DgXPigPEGv3f/XrTZE2Ic5W8Fs/UCxL0ZrW3HkfuNIXdn3LFjFJddIPOefV4Z
C1ne1CKfyZyZP4tcn+VXk2D53CAiUZrrCHjPa9KNXnPMRACySZmbIHiUrhph8YdswSkf9Yd2rIsN
8v9Ud8T03TsZenbNZAglw8T6/cGhmwOPS97vbsCFHzCZadQ4x38mBI//pAOL1iztsXgw8sUWa/nO
S+9pEN+jGERGFC7rIDxYUhPfiUGovulN/2NOMzfC4G0GxWH42FuPZHZaSU5BK7gZ89jCh0vGSooL
AuH84CvR5JccS2LqVRzNYBKtDlAzxb0W/YjoJlV3d0/XWrRcBp8JBjm6nR5EXtpujbvYxD4xzAht
rKPzcZGrGRIVleMIIdwhyKKZW1gvy1xUl39M0sDGEuUOV0J9nstAKyzW+Qn41xLeIdcPt5mlWRRQ
ChPbteu5LjRWodxZmtuP1cW7gqj8k+D4+MYchAFpxVfwgtLR7vy4nAhYZcVT226uajgBIux/DDIC
ZsmBufCvoVLwSR+ypk5dReQVapl7q3WRXoDtCgh/KiF6q0WHqzQdxLmnDU4UYLbmVUBZVNp7E7bE
CxGR3KqkTt6WGCGNuD98bCj3COHJnxicE/2DWtrd7lRzXrPrhANiQAuZ9kdM9pgxdEsfKvnjBXvc
Y16KX6CnK4xhsfgbwmT8flail8CApmISHQOt2NBvUa136EU6pgnQV54LanRJHYWmA58KAtAwhS/N
BhxVAyUuvewWldOta79ZcR80zt3Rr7bpyg9kj0i5LqShz1zw1J6X0FlbROKjfBXl/6mhyPBwzLb3
pnCpxz+hiDDlZhW7n96ZQh6+gRnsWHLQTCSZqt9RX/ekmCE2EggErGax54WOI+GQ/sDnf0ScqF+l
r/s8SllH4uOV6rWPsEjPJ79UkLrOd6xcN7XrcXjl48h8Kot+hC/NaaPjIlIlL9G047UcuWL1nqcn
arLAZ6pPuQLP1/pXr+K+NIBWHSS8HGSWuDUwtEAsTDUmM7CzzObQEoLq6JGy00BZdLEZZHM7J2xm
MbIiqzopvvs22MIwRq0fHsBLgy9lad8xol4c/P306wFgNVxHN50xDUyf1iyyCbu1syvsVMvngzBX
NVozSDkr3ihXXQ3RYUOZ0dtimgMlgK4KcWFHL5SvsQbVVPqkixB0W65zcI+fG9UQXuhFEGStqNEh
y269nnUPQfzJGiyouYyqN6idh04bhaGl9JEkhM8OCc0LlGSZ7lZxLDjrzMEgdUR+Eibt7lmius7U
3u7Rwol3z+EcFAEja8kp3ZDyXu/RuNilOd41gHP/8TS03LZzPkpqIMwxwPGFOuRYP7syOce91mCT
gIEhOw6LMQJtSAjA/MaGFklNPq9B4hFNpkmOErTypVlW1B/xl5EOdw7VcHwHRkg6mO9y57gsHbC5
TjGalap4s6R13TQwt79UUoF4g1ga6XQjBhqGvfLynxywZF4UpLXaKqrJ5piO08K6JcTh7R7boL2a
Aw7oGYyAqeRMS20OYV1UUZoSn/DtPuq8vpEMdxV5YAs68BwJ+D4wwcd1lQBC5VTHocADXOmJ888b
IdzkgqFhUhfLCKWvidy+7/c94wUr0Vy2dcpwlkmMvJmoUuCi+Yvw9dn2p1wDjDeVOtLVkWo78iuu
OPMusYq8nJLJR8UoWsBlK7yiOH5lJ/DWKqovIkaqzu6l8Y3LPvIFsiI+D1db/bwIEAsf0QZvOW5k
tCWVz3VFOpE5iwiarHGtDXZau3qqf7tj6QU7vBKYArFGEiSGAGa/bp7dKw1trOaS43Tg1+kTNOKb
M3GI1KPhWaTsob931t3Q7p72ibuIHNYxF/YY/CenAM15hgYVV4G4gh6Y0puWjI6vI9Hja3YWa0N5
t6u+aazY9nZEaCiVG0Pp4gHkVHcGDQh/UW9suIW+FugqNPyg58YjUcuY6O+Gz10qnfOZ/DK/MkTf
azesyRRoHQAriZx/EdDcwmIaRZERlY8LijFA6CzlIkxgZrwNQKNedYNt3vz5SUsgYrFOPienLIHr
w+Lnk/wJKgEK/40KsM7vpPstoKPAE5e94nBTmNiKaGLdXhbOBrr+cmDcZid99QizCdHlL0oeR/WI
1w0NaTycOqPO7+AmdK/PSxQqGp5kTGJoa1ABFIkiNh1OnHRdNXZIcdNrnNwcQk/718hahfC4u4LR
+FfUD3QWM5T9XYYgQuM2i+YLVpji5dPlz70kL5dp7kox8KST/Ol2XF+zASZ9k4gAlFNaEzJijwlo
d0K/xL5LhXqGioHKdvEhEyIM6itDthKMTpWyvbNkzxjfqpQZKmaeWyyRiyHXUBVNMlirVoKtS/Re
Za/qoZtSySzz3l/Dr4CdepGsF8qU+L9JBhztUMfKE8KKW+qprhCeSlbtzh3MUINshydU5wX9YMHl
vf+JZdeHF1cKYpigPJ/wpFTctbIJqY9Dv5AvF6zKZGparTU3wFasow7namF9rijYYJ2xwrw4Uyl9
YIkQA8yy0d3Om+jLvisHmHWunzEBIWQ0nJnIHaxyEwuiFH6E4/8K6X4HJTQZOjqyqQ2WNQRa7wsc
9RzdLHk8QHh+Jpg++ZusXoXeMc2n+RuVReh1C+TtgLYZvurqxtYvJRG06Eg6DJGcNWysUeR8RjAZ
jx2J0vFhtRsvdjPArVlVU2qKyMUj7x7Zeg1LIrBFvH0vboLKutrSPJxJOB9KJ1vg+B3+xFgPd69L
2L7GNSwB8bEccdUYb9MyQSz2K8jKwZ36z6FFHjsY9KFQfRhIeha5T7m8blOR9YN+3GeK+lgr/VyY
awe9LXnchYQpxSfnll/9+PFggoFu1oZWgduWoLajqHy3jCL301ROg936A4E8dB5W0yJXSsA/W5B+
UiQlzSc2vyUmSPbcf99Pe41+UPxbc7C5+zC76x8Sg18aF08JcIs8cD3v+6oZK6gFlbhDozMAsxeE
Z9w+1vsMHl5FYwuwvJWSHzOoD2kSgL6FoF/vLA9n/03swuPg3wNRbJc49ztePXGal929DEs6n+bc
ojVzlrKZkmisEhtjKzLjfbI2FhpEfE6hhjzgy35rqWuVgGpOu607o9cAxPa6S2NcCUMx9zC/0LRC
goh+k0LrRRMORIt24pnw9PP2AYG0qr0JjA5VqjGNjCuBtLCXJzsHZ8q6WmpfVVFdYeG1M1YTSBEK
Acb2e7O1bWqj57oZ3ssirgbp3Eulb16ogsJjbJ6KcIi4teJ02ow5HdN1p8GMorS6pRYJ43GQO6WJ
UNAARaeCcVACUwKtB9YEzhvtvvZkM02s8lBgJMfRoXayhEgrazt+575P9L7/1PpHKD3VacveUffz
/dWV9mJqSLVjAkrde479T7tj0xEAnI1+s4jdqt+PSjSQMYlnXSkKU6XfywkHswXScBA+L9KepPSp
r4R+WKkEwel5/uneZkyXeDaJ4I/aXXINf/50HFTSYZB4svBzSlxUow2NK1j+q4ngWAd0/H67+ggh
/6T0zwsgtxiTwQroPwEq3zHjDp3bgcirwMvZt5ir723PXRCkQoBGCJFV/122hAljuwtHJ6iZNOQE
iK8F7T7oMcLhwUidTw0o38ElqRF93LUhMaCZGDs0JfdeuM5uepTrG7s2o7NSUKDZklBJActcDRH8
M79Z/eIE1sTCCp8EQeMalqOuTNuVKwxTiad7iaRlpku04WAC+neQZGM7OeLApsJ1yIAqHTjNDs23
X8hlO84ITHX9t36EyRt8kJLrZssArmsHQGTgsJS5DgDo1HBe3HIMcW8mZNjH5uXyw0w1AKUsZOEc
SiqdoJXiQ0KnjnRq+In484xAahNthHV3QEpYZ99r4jyy1ngnNOTJ++o1E05bO03p0k8Q6xnfYqfq
kyCUMLTjkJ7bw/Hr2N2af+bz14sAbeiSRA7D0/4naCUoKGUlwAz+sJ0R6FsvJEJm9SOy/OvDutco
osmFtfrPo/CjSw1wqEnLMMq8VP4mC0SD+GP+6w923b4slQRQHH4Yey18Gy2lysIkb7vqFyPVdOd+
JcaEquOX6JWE6kSVhGqfKj5xIill9o7Sm+IKL1XX2iuDKg1LlmNAJQiGw/DQnSzztKRfw1nWEeEx
dUQysIq+Vs0SSGtbCyDugV/bfDoH5Ia+DszwmYrf3PGRC4W8n8S9pY0pr3ExipzFJPIB53fspwH0
n9ZKGKoPmholMHdqVAo4ma3epWu4WY1AkSQD7iiFrIXi6HU99Gy/1YqICWkqnmgQu3FKfe7HDZrF
42nVp7GLX8Fzhv+kY3Rp7EnCfp7VzT99xQoxPQ2tEOLxuQw2skdSc3djdVmGWWJaoIZ5PuEyC50p
Wr+XPbbQEKijX0Bzoz7WyVQ9pmh1aAreqpJdAAAnFfHElYzm+Pq7yDzig1OLWYLCn3HeokGSHRkf
atQGehJ3KeazOdWk5CvqXFalM7wUS1OfppOAQwRnSiXb2qTl/pJN5DKyNH0xQPMukgMOVpzQvmql
KxO9Nz1mWxzsSixHI6DgN1xMTFEGK6jBnTOAJI5EAQaQUxy81lFoH7SB05m2fM96tZd+moxPB/eR
OkT3IhsRqMsxr6J4uhq3pcDHKlypR/WqO1i1Ec19UWkzy5JaefpAbD24kd/b2XxQ2C+9xSScqLS8
IwyCi02YhkWGnU0jpp1NaTZTBJijGWiihv3XNbls835ZrngfBbAmBFD+hCYt0Et5TibE6BKt/HJS
PNIpCXDmM0BKU8Ya4G2QtjeKAIlowozcKa4z7lzYuO9GwPXdqdjaWGmXuS3YqIk7swQSx5MhsukR
fkJI5HGuSnj2Kww/++nmuYnrIZLuhfem8Er9Yx83JUr2eJrhrJEwGdUOlV7swLcNc1rbky0wVrq5
RYVzHvIiuiFq/r6XfQKxXoVZrhtti/Xk6BaaNgdtdHGLwxOETPRwA099GiFB+ofv3vFnzR0uRraC
D3pN3HRt5RxzwNuiUm+y2j07XhGrUCiemKm+/Dy7t8lkDZxxm7MkaOOczwaqNOdcKh3GJ11j/N61
gl0YDwevGg3JfLy9EqHnjZiL9H0lBsSCXzFi2XVgqr/qwWAd1S8BXDYivpuplUbtgrqXwjwe1fFS
ReAFm41JcZqhNFGGjeDZtCEmnPwcSjEQ70rPOH4Fhw23BZDGy4Zg5R11LKm9EPrnTVUoj23kDD1l
M3ehhwjP4nUC3/e+VvIrsmEEQcR7EUaNiHB0geT+E594NX7XSA/rL4go8ZVsNsjvlaN5yL0Tn3Rq
V2cnMQISECx3ysY9F4sakb8OeeN+Hb49OJokIbZWSbOX58ictmQPDF1y70bLGO1TVxYlrJeYGYwJ
K2J3jzxAXuB8KCR4C5zJvKfonQJr3eeTZLAZvR60OWYlcg9lOehdJHHFZf86Sm62RcCeuTz+uDwB
hBMjdNBlvJHhy9qyeXu3ogB9dS9TMOK9k/9g+fXt5SxYwveyB6QGgpGPWfAD9zf9/yrQfN0WVU8H
3ZIL1uUgT1mF2Q/oDx8vaz33jWcngs0g+n+kY/O9MiA+Yv5WH/RW2SnGOqWlPcUrUQAn5S1bnXvE
bbmAovi5hWikmp8h1PSZuNIt6rcuW0M5Z3eIIhsEysAZCTK6w0mR1gn7GRdx6fQXurdmMbKVbJSK
dRyq9VY17ZeX8YXGDAKeh7ivv2NsFs0jMkg/cTcgrPxQftm/bUnKPU3gvj6Xk6mI3myEg55i1hGV
lEJ4XmejOk0UzaEqgQmTVercv/ZDqZyVL75+ZStwCvTxV5Gf/mjuFTds9uXNQK4TVu4CDOpazdbN
aCz7pJONcqTqmvEDealliAWRvkAWEtsYjVWD0cqPbQ4wK2dRq4jdCbgATWiwryflmpYB6BLcA96b
8RmZ9WZ8CXH7CGfIhGgwg0iXUIMYRo/xOGHlHlHCRNr0SExe7pWR3CoLptEORmKuSsNg4NvtcKZ1
AOTQzos7xHQMOE91Q4lZwZqn8muTrZJw0cLoFl6ZXrmFt463DAJmk4flZpPNHGBJnFpOJ32iYTc0
pqlfFhvnYSEgWGFscfjRy58SN1JKapjEZ+JaK48Kjl0scoa10yth356EwWA09rciNMJwxU1ycRc6
l38wEMhYcKfu454ZHuDJW6Z4OPayk43IW0iQ8U2VhFU/Uueyho9IVJIG8G9DacuGZlzSv4+vEUgd
7oxmpcRwajuPfJBvMFsWMhbXlKXZeIw2D7ENtG0NodjN2ONTm4yVWvpp6G/p5VeLzvU6OmuI3tvR
ET29267jOQL47ykd8Hp9zfYTO96BrTSfv6wn67djPV4azwHoCiQJrNeeipZUjWqq3wkH+kHrSKzn
KPxoHdWdpD9edZeu79VAd+XrIg6Ugd8YcE7/2ntMnVPkO1Hcz3RS5ikYAcuHVr0xGhDVC6FAPZSX
H+ql5d3wj7dhxG5q5BPMXXPruv/UEgqTmQkyn7IepQgKqYeMmSMgD/cCLjEpxGgjgZAk52eHW+jN
DGH0Z3rsUA7FZePTSOuQvXE6+zMsfxiElvbMTnUoWTacpQlkWNQOTaZ1+FDEJU2EcZJstUEk3MIr
0ybfHjdgaSm77SJAFsHlMYVudtGJlHQjqjwVY/MHjg63kyPQ2MLIYF/4bfrkQdD/gygUIh+FqMbQ
xZ9rUjxK7/b868/L14kSvxzmp7txeQUYr7PcP5c7rZPcqwxKM9/bvFImxSLILeClaYc856Xn2Q/C
U2p65rk9xsJPLIky5bO9gursMk1yJqfp2Q03WmfmzX6zheQLIAoeJisYvZSfRxPxD+lezjal+Pkc
YRwJJ0qYWoxJdtq/yjTR3VmsTfJluVbd60nGFj8b2zCq0EoGM90hEWeoi928fTh5n79v/nF8pQey
SDODkOCXgz8hOiKyYkVZJksp2ZQGP3U6Qu/Hv9r069xtpH2Q3FslXmYqYglsL6iBNUh4suSVWdUi
7/JuaIoE7C0XWTjgebDk4nqZC56NwwxlnvDSaSaqWKW5P+XNAYpxPi4sm3BDrNkYyobVupC+j3r/
vsn/BHMCzI01+yudJgRA393qBI2DZhocKxBXB/4VEQMgjpBgrAU1oJ+5H+7TmsEi2yX67lMGDTOr
ZSdLCjRYtPuW2MfqgbG3Ey2AIXsfVgMRIVC9IvQ437OvMrLnzF1JJSmsxnk8N6vMHgexV94BkxQ9
Nd9SiDZRwDT+/L8UenHUwy8iqmWZjkHmV64moM46VplKzGHP94JGosVv2NCI6nST/VODGp5mVNFA
r/LsYS3Dae4VSwZQOjGhnjhhE1lCKQn08m/T3+l3o/PHvyVs3AfyZ8m31nHJOZHo3xHuuGPF90Fe
w/d/NyQmEL9RlMveoFxXVM17pF0ZgLadaFXrTnSTyVYKaiQpxI+m1T4hKYmw1Ij+bW1Z9AnqpUZV
NzusmOdd82sh3C+SLDrTkuIREpXdXL2jGumBTTbdOEYxL0FcHBHuDyGp/37fvlS2A5c4Hv0aLuYG
yGT5zg3Bk4qU/fgNDEKbBAx9yTRjPQb/IKWXnX7/PN4BfjUj77w2ZOpwWaErYHSfklmFOX05C5ha
t5p6/pPsheA407dMBWj+07AupWYnhqwvdyrJB1aelhhRSIL/34bEyhvnS5qWlhBB8Gbj0Nq8gIhd
ufQSRJxG0PIXMnnoQY9aN+1pBLLImjOk0WD/uxUS6BMxQeZWHytOZ8RWIo/tqrA3bJKCTjRTH7mU
6xaBnnC9KhO/iIw/Kaw9gYKvexnKa+ldIxmJx2H2QYrK0cVgal4AuHfRJkiJ7f1Eo8uF18TYaHMm
aS2YBA18uTzhz1F1H5UuSP2j+RXyR00yy9ZXBsfBJWRWGiV1kNKN+nhczU90c2SuV0Oi2gV8qdxl
IrlwXseEW9Rcjx2fistgzVb+1vCZRfARx2q0tx8jSKmzVC2QbZpc9C6dhBYDQRr9ZJ8ON1g/pVy7
OuuZZAh8MOdpXOHaQb46zxqyaL8rsNCif3XbuxAmOqD9WMeqfHx+gtCQiGh+PHEv4eBtq8G7Gz9A
HSaeyO1JwVTtHUL43+3CX1CVhHMGkvBIqVelra0hOOVzD9S+JmYgVWcvh1lw0RiMIgeeK9VzfEOp
lw9ItB1fTcSrQpeu9P+/jNXEC2eins+21ZzRiwkFekrATkhtL3d3ILIfFXKbzJGrOVYY0bn5VIVC
vMblklB9/p2XTagrFeNQmbaF+oeWsUzRD1IMv3ji4qxQPJ4uCPKy1gOeI62mgZfKcZjYa/wIDnGF
LwAmYeQWNl4179AtrPG98kvK9yEhpxeoFTys7mML8aHegVnUCZeI7MkvkwWDTYyiHyThjHAySGcG
WjleEypg1jRTm7c0epJKG6KatiBaJP6u4b9vajAZ7fTYbtpHMQDjp6sZoiSMQimG0KxPmjJYcEEb
eHhiK7uSGsK5J4WiX4Cl3/sst5SjeG4miTjVSiEHOlMY1N/EcWim77OpV/yBtgvpyGd2QDIZuoWq
tJx8XA0RHKjPS+AisCGiR6Z7spYMs/3vrC0x8a1dJuJK0nyx/s8FCxpcYsSMxyST/A90ZFR5cH4T
WkZtDGWmvD/jjqHMjJYZW/0dyVIOXt9fxhZA7rIpwmdh8nuAxof/jcQVBgVrqg2HABxtziG1JDXj
ngOb0FsskDXzQohBsbaSPlIK48jWFSK1xAeQNdllf5zb66zNYmNmOKrdJawvotLDQlkalxzmFFzg
6fbKab1i2ZqeksF1DUKSAdQytJKt8anBhySrcDqTgpjtzWeDibHRh+v3+ZJXxGWMgthtc/2pPHQM
u7mZoJKu4RztmtYnEmMK+75VJ4wiYw56s1NXIB9HzLn/0friIwynUtk8h//cYJjQfTJWlnylPXEr
ZlpX+A2J3wvYcvmX9qyiT98yItRQzy+AjywS5RgSKEI20ApY0+GB4AOK3cTfHAVbFL27Yv5GjaE9
+ZukQCqm1PZmM5idqHWM6UcDv8vlUW17LHOcMWALVS5fthVU4OlVYu/+luWtAK31D+VSU8aPa3fA
oITd8wuK5vxs11QzDc5VZKchu6T54EDsMjrDNDguxwtKqaMNWEucz51rsRsuEzLHOJd4cpN1XC+q
ZcG7OLgYv9wBXKdmCSDbCVxZEJUX6tI6e1ZEbCoi16KtZlkK9h18HoFt/8GPKGX1hQEQRaVcnVbj
pX4mZw1xBQ/o+C/4AUYXmp5Is3KUyKVdfPgfsW6GheomL9W5EsZyeak3DanzMvGJRV93wDt5JiAS
wsq0PcF3X7RG+ziCjN1TnRr7koOk4M2XGZoOO8NKP8x0HeWvuPIQ8XvGZwxPt15TmUeJGDTn6YfG
R06VhhFHSl8pIhQiwdb7QABBNITC7WLYT2AyVNE8IzDO56/DmDXmFYOksSo8EG9a4veem4jkBSs/
XgoVBXbLeVCb3MP7z9VgJmPQJcrOxXy0xyqtbdpczTBJvAFu5ReWq6l6kWvnM6au6QgjYySHAkdC
WcdBNXov3/A2wZtZ388w43abwrPHDFq27wJ2CahBNyKAUjY+G8YXMH9ZKrnkk+O9w2jw6oU1z12X
2DLIhqykZhX5EpLoF+kskqnyToNkBl0wfCeDNOXXQY8JRdYbq5nqEkI+E7Mk2TYQKCJ0p/yKE7ji
vMYrnv/hrWlDIw6LI29tBQJG8+rrmo1PkQM9bVvqqiPMeORZWhd80d7YZfEZ1o1miW0lWul6zQ9I
5j71O8tboFk92L7Ibe6TKBpo/aX1wNdDl1JKkxBCm9ncy8V3p4ysIroRMw3WfFWpyOrdZqxH8XnY
ItM+OHJECzqV6m6S7/9OXUoLL4N92hj1/SRRF6emQZ5HCxvBfDYJ5nqLQBjd7TKDFA3lME4vv7J+
LcJ3vl6faNCexwfYS6WB5z5u225KePQJxRQKGpN8FyQYTdxQUUsR344E+mRg7PnZILmZa3/mjnnu
MmwXJslE+TG5RMVzxK1wA74oGF3TX9kLdFD2ZwI4EdAL20S/pThCroV8fuS2BdIHEP/muhnxEFke
yo4NFTvpYbo7JRTiuWdXYRkASNpALkB9KQNYcbbtV6Q5dJhVOgsYokCgLUUjDsZmAMSCBQP39oAp
AAd9TgFGq5ANDLlb3wLdH/ZhLAuzlBS3IidxVLth9NZ1m3mardZpvyo9rjOY/InvGBnowHUCdGxG
v+ESI+2nCabewvs53vcJM8FYU6YjI8o/80Y9f0dSV7MuQkDhmfA6uTcTJvfONikni+1VYD03Tmow
rO5qyqFA62EOnMb9HEJw81tvqjDc4L6OcL1FptxjrJThHP6yhXP1GzwiX4tjzIxwkoE7WAxbSl1y
/Am0qsG54o1f6m+jl6nbONBY2GLcV8K15872ruIvK0db5ZK1UMu/3Lwup/gvpN3Xj/+WyJXe8rSh
3qdjRioKZkciKuFKSKsftxucFKxD9sYC8hquxDbuniIBGUpOb8vxPC10plxtvsEFF6Pl3Jf7bzV9
AVlR00EsZ/+yiEmG+24UhAhAt+xPHS7wuoiEj3pjvba8kKdh8gIf7GYoUzg7UIganmI40azaHafo
4o0b/1q+Piw+kXzgVMUpJU+/gOGwiKsUEfIWgKf8WFVFq8TqVhJviIKBAQXk2c+ub2RRInSc0shr
dsG3qiNdJ2BZebSX1fzPnzwSXY1W7mD4JKha9S9eizScmOCzb+29qk20AsOL2C7xMv7+7NFyRmfX
RmTWNVolHQqew+G+J/nGT75psfA1rBIUVai3wsCIiIcUaFaFz635PoC3EkFQ0OaH6DZ86g5jibVX
XHisyC5k5niYQ6ILI4KaFoNxWRByT9+QEyEO7MFIbO6WpzuitAmNnDnACgqg2H22XpgOWZPMEq3G
GlpWTga0KY7lPOwRqzQzPhTp8su6jVPUpkq9QuLZjVsYb7GtJ2wcZCEKZ4/9tbOvFl7N2fIMMYR/
dNpmLf3qXPSdx/Tds+I1v7BPK2IePZ/mUNlZEcREatQMJWtHy+1wRH/iCpRXAwrXSBvboiPwlg++
iWuUy11E2PtYubZJYMZQGwXEcBlH6rlnypD1Ro/jicy/EyiBQcFQ8j3CThebRrvcdmZ02pJVDiR2
gXz/8Lo2CTTGPAU+xRRzmd9xcIjq1A13rvkIOgcS5p+JLjQnlZQ5brkle1xZorTYOOTcMVunvyrV
FefgCGX+ZngGaJSdDHIMjZI1W8PoCc5KEyT/Du/CNhgGEqmOumOwfB2X/Srw1idOH8Q/YKoQr/zn
z5nNUZXfZg1WoMK9VaeMDGnoCN2JssGKQMoGHzbiMtthKzUGhzJfCIrpN1MRG/MHf51s59YDZbcT
7V3VkofnFnVDBjZ4UjHPGAEhy1Nnq5sDn6E07tMt1uigeiegN5XIpjYszb40sLQAsDcPESFnX4hE
LdTiUzFMjWVMVQhr3kaKr99rFtin8VF3a/nnmrfvkE34kDzmmgLV23HRZn3ziYFR0mq0ByNjQtsd
0RYYl6+ZDUdT/LcPunpwFmnRCyT+WhTXdCK+mJHAvjylCBsqqxvM/sPEKX2UDMMJz+Fa2Vj4EPz+
uQDhizy2snH/HDP8OgccqyL56PJdB6c7zLZPTFEnEFRjsUmei9pSoAt9QHSPKCY/h3MMvtDa/DpZ
wCiCAfxDlYTuvI893zqNGKJH+zIZNLqW5yevk6yuyQ0JY9KGTCCNLmKhpoKtosEJBdyMQf3HJdGZ
ka5XCZOoqUmXl2dq8WwkB7yej0pv3kmPBKnpVBdLdpJ1T/HxUM9fPdV08ax/TrEF7PrPQJp2fF1H
FkIoynvQ9GM+sHcoNow3KSurkRIXGSvKRVjaWC+zObt0G/VJEwED0QSWjfZMXwB7b8Qg6IStoBrD
IOCNpv/8A6fSmjEu8QykI7KsYdNsGOH1j28t69vLz3YKWOChxWEEFLk81Qq3aY/I/JiUtMzn/OIj
6oAw6cbgIhvihYpR2nhVj9q6Pjd0+XoHsqkYhAY2p3w2ce/vsj7Y0SOQb3S3b/uqPPhFDyU9fPcX
ZOVIHYdaHEnK7hhyC+9LJ6lw9Br9gwyZycgohyLzIt3eNxifT+LvqkNvAP4QPplA0CtuZLsWzBRO
KYsvInRT8UgmkDAJKO/mv3jftp4KOLQJ+LhxYuUGgraPvDS2H2v8BDvXHYsxYg6/NB5tvUUvMkFv
td6Zil05je4BYPRrJLny5A40IFSAU1AYGxcqMYYwH908I8KLzX4uPnIWUEEzjEqOXrkmfb3UZg00
UcR788yISG+uta+3/Et0GMGCXNInYi4KVEGy8CsNTVkZMUTzrwpYHyKHph7Ajtwyc+JiQp32PKkW
rH8TeW/qmzdg0wt0jfnU1rVf7uy8rZuMio0GbQIM9H+84lSk9n1HC2sYZqs7XfGM+5lYbzx+ZKAP
paYHIIFKcN0sdti5B4QWf5URqvDfwO7yJ4IAuiJKCOya7aNjl3SOvUOfVUlDQkjRUWZWlHnBVdtN
W09eeeyJiDGs30bYtGXuTwbn2PSmG6LgXq0yrrOHlLrddIK9wI5hcZGTBm8WsfPZtoc+ElF5wGNX
cqAi7iNfZTswgDhqN7hIBGtwAuwz9BlzfEB4nJgMl0uI1R9LsBDkpPk3BZzxrL+a85jCLqXz5U+o
dYfBkAPvNyDpZtgwHid3smxkUklMSZ8+wnp299xWhK09p06iUrFbb/vNOCZuH6pYa/R4hh7N3Oxk
rpjyQwlqucxLBgcMokiUz3On2pSG4n7g3F8d5kdl3ophVIRjDdmkpQS53aAcJDnFewZ910ip8L50
kzx/kk2jLMKTMUhzvePB5/X0+ELtAgTnWsh6Mg82yUKYoY+yfNtcwFFS3LYsJr62nmFSvH6i+zvG
E2P38Tz+836YZh8da53jif1XZe4RUocTVOycvcwyQ9mSFaVzsAezjgglpSVb2b71k/wObNFGKusk
CLhMYh8L7NqdZDe1ey2YnMN4ylhwDB54yys8RwrB15L6CkVmhAdE6FqOXMaZMkPjGdY1a0j9MBTo
mXHwOKPvRYqcVbfQCqTWtUFdvhD4YRRkCarWQOb6EYyT98GzBaaDhLOejy1UO8l4wQciSjq9Cq64
0DQeHjEjB8YuXwFDB6XHYazmkPc/S7KeYFp9UXrGekyTSt2ePSgQ2aeAAmHzHGifpMLPm7iuppNO
IQgJGLE3gvsknQDRhGXB2o4IjqTclh+G05xqv9g/jRkSNfphIbm0h7VhY7wW6x1I7iEcORkfVMrM
FCPT7Cnvw8wXzow9wOaOpKVdHHXCCYVXXph6vu2roD9VbcLx0MWGERFQOcLyun+A8ZFkWFt7WWhz
OXjDJaqt9UoGyvETSjWGanV6BwjuFDHl7elnCA0lVBijkbIsUCWhYX/HUOcYn8TKt+p5mSMZJPDH
TA4zU6Br2fL+4kAMNLnRYlhly+ql1s11ZRf5cGV5vgbxe8nr/EFS7lS4L+cPBjS4Bfuujhu/ANla
QUouowqRj69Fx6cGu8g3bJ4dyeCYabMPxztV4RcXDRFMyMgwRxT7D9aaCS69k5ySi9no1hQZU6tv
wgyAqI7dcLyCGfe5lNLJJkBkNBORZBwKajgON93OtrLgpycUs8yd/P7mdqyOep4gCvCbmWXMltgB
thre/HLFaY7Dc0kAnAIqKjLEawTPVlm9/ieikemfhQfEARAxuqOwSCVqT8pFTvwtXsIcm8xdalM3
Q4K6Ibw8WklMYgGFxuRhbV7fIoSFK1eLX29yL8C+3ZU7GTAi8ajgg3lvZjYNLCn0IJ7ry9GOoVND
OZkQWH2dUtIlA39Yx5wHpXiaoQQx+0aZpXsIE25tGZeOM9o2Pzx/ofAvQPGqlUmR+CXUFwlB9/TJ
L6gRgNl7qdB4XBfKszbyaLGER+R5TDvUzDjuy3mpSMK36OafFPQdBvvGH45rUnJTvtwpe+c3X0G9
gVJsvvASOzia523NBzBQmh5tLg9Fs8urDoAbKfHNE6+j/4N2IQ1zp7SQvn+eCt0moJfmMgpOADt+
wDe6WK5ZJNWSKgEv5aAPsZPkt1AGD7b34I/LTcWnj1qKsiM9HEG0FpUxAiQiOldfWWbD1KQzuXIT
i3ARq5pjkrQVQGiJtjLniUEBoFYyx824yFAeMbBhB8er1NuPBEf4h58Y9o/W+WE6P/Ak5+V9lPOO
fNjUQYF167+O0LPHSWueMeiX8YVvYiFDfY6fFaMz+W9QGJTN5+lhrDyI2BcHjOk7rsL6iH5aIZq7
8UlnCsdqBUlnhX7aev4VRQyet/JP61cn5bMjCgG2HSjdW2E5ijjG/Emb8p0G6WDi1q7Jdk2uc54n
D6c4UX08WMrjbRn0cwuaG7hHg3WXiVrTeSH7Vewxk5VxrD5nOsuIGltKZVRDkZEifbR2EJ4xwT5u
KH+1lerCw+HeNq/kJmzB1SCYon5HPDOA0+27QZTcy8WtL/UTQAzceHk9QzsD7Sw3jkqOcotlSC2P
8KZd6yYBprHcE8vzrLC3gAGLn3DosuVsM7+4edAqwX/oR2zdvdOunZxGCC6sZAcKimoh4Z2QA6ZD
+l3Ck9s0/pE41Xk1xIUpz2LwFpJm12ogE4tBTfT/l7NgYLBpAx5lP1RFAXrN+U1UMmZ9ZOClr86O
U0pfk+JQRDkfua8c3JyGXTa7oldp6auVDapbOorxKxZYIhux7Lcl4joZI3EZ0l0Ib49S8OOSpiSD
Jr73rz2fOXWX2qwxBbSHkrd+QtYNwwgDqGGaDPxofPb9Crvg5GlFWC+e9DcxW0nNiyWRnfY8tQPv
UZk0mDPYdx+I7ipCrRHKWLp29G6p+NunY7F/c22egv+nlQQ1sr+FY3lYhO/29D4d7vhlIM10RPxQ
1vGX8zl91U81Gxa3MIW2JeQjNnZZgO8q30T1JSkHwiM1Fpjt4F2kKhAio+QlwjclddhC2lNrijQV
t0wrSDvGWZkx+/AonlMa6F7udis4eBETTcf6trrOMyJTtotsMRbKAjs60lQtxuD6T7x01IcRRhWE
Z5G2OPlHmbgyNG6wwW3MsNZExkAlr3/T1e0LyBMjexkAlByxcZbI3tLmUbT+qK3m+VWtSjwtOGIT
PP7M+fzlASCKGQqM3OuC8yXyS91nv1KGQldAbwN0EY1Ich8DYRtPck5W1pdm0RahogEMFD79sMzK
PMsuWVsuRx2WCTG8/yN2RWUffLZU8marwN8OzHlvHf46Cffqo+j7R+iq1DeemYhNz2wTrNF3ij6+
FYpybJdPN0gKYbBYHMMLBgNDvwA0qdNN0iuVNiy0pyF1YeBIfpsZUuWhvcAS0fNH54CJjgTNoC2R
Jp8uQWPmkN/4QQSAdNeCgIImsLYHU8oMN6eer8RCaFoZDpaAzYWcYeiA10ELBCkK8b5Fuh5Cb7/L
R9BR+eqrkEUz8ads3zyAPTDT1I6gt5dAQHfo3DInOOUvH04MwAyWw3Le4In6NmQa/XsHbuYrAkeH
7HL+KMa3wS18VhafI25HwFxaGempu3oBqSMyUwpOcUoPvC4Duekd0Qd2RsBaiRU882gO7fKfopkv
XQUpAfVWrk2OzNpKi6yMh/22xCjTjYVdGJrVYxqHUNOA9naY7QQU6CJhkjAb6RrBCeSpk52yewmw
b5K/aXRxbUqt01bKGM705XJX8J7BHTvHMylgBdcClDIvQmgUpKA9W+LEaLGduaDj3X6KruE2TqOg
LcMY9rfi9I0pqyCqkmqgmfZ2uW626NvBE8DZPORUwTwUezVko4hz0yj4xUK9z/NNOVxlY4njJHos
KFCmHrT5p4aBgevdAmtX54iuD9l+5JkFdhfmRjBmJYn+31NS2Rcov4+qY7CjYAxOdGtKmwcc6aXK
TsBPGuOos7MEjn9MHwlwL9Ygvv9nbLhzO/dH74Nhtb3ODpmTKuZ887bH0k3wO8SF8ht065k1xZ/1
dV650+Riia/6sPnZn+blu4yMakCpm/xAkhx+j2X1sYQJ7VeF0T4CbSP65yfTcZitUqgjKr7XuoRc
X838NBrCtvQsJKlTf1Ho+lPb7PePbuwzkH9GMYyxP/9dmwKdzP60csn4knK2Kv+Su4VcqAZdSjD3
YQz+oqfkin6Wh6Pqi9MXH7CnHQIA3uy5f0HA++QYY5x524ALeA+ovPfXjujaV3LOvtrqtf2nRtBM
PDhZSywoIZ4zjS9nTjht09ekfureIRD0XMR8DUr1A3U8PvUqNxpbatT71fSsG7NICIwMD0vfkMM9
KSWl+CcHMpjSTsszwScAcuU9zpa/QuCW42ah25ITt84IjuZ053shXvJAv2pcG8Z5gjLiEFM5oTx/
ROzmSt6jLnvUE9XwdZaq+jEVHFrL9siY+X8MJbjsqUjh47KR5xAohoXfsz9pWhqLh3c/sdrakEd8
GR7Z1KKM6pwSFH+sbhyoT8fX5TsFQnceNT3hmsSWLxiPdIENhojTxEpmISxK7LHMME1KSmFzT5C5
JI+zJPQk2kebPad7txXGShbblQiS3u/1ztVEYuSaAuvkGorjBVvgv4cbnWN15c/8U3q7q0PaM6XQ
af3QR2tz1gBUmHDVJeR5+uFtjZEtJypWcOkDJCbOxdb7LVPtrme4Hxygnj/taM9kPwIDHHaiYzvH
jTSoDXYQWKTGxSNplWMk9Mrrv8Bletah0HCW7q6JKidgTxof/Ps9LwGWzwQD49RwBGIFDDZr2dh/
EWXj1/nCd1q+USkNS2sS/WlSWJPoS0062D6XKAlnAzxaiYLFFi85aVk5Tyb49zkj98kJzIw1Q2wx
hFXXl2rqcFethmf1BxYZEE+t94vt8dxBbyL0n+v1PNYw1/h3BdpP1Ap0/KAPwjQFbcMaJOxOU7I6
hkbHu6GKiUix3x2QJzCXjQMoeBPtY4MSLnKM++gbUxxzR9oKtl+UJMjitkx9RYfuZbwPe2mehcDW
bwzhjTlW2PRKn4+hyIoj8UNN+OSGt8e4io5T6kH+FvQW2wbxOXE4wRjifckZ+kozZ1jvFzJHLM1o
c05EjeoyCSxMu1DMBq5l6rUTix8/u4AvRNSpJ2qzCxzIbRPJeUeoWmipIAqugEuh5YrR+ZXUlGLp
k/mk6ZlreL/vT6ub49l0QQalvUDOqNatlK/iIjvZ9gHEDuFBwxhMtyEUQmxWGTMOkmCMzfGTa7td
oV7lDxMiNg5YuzxxOLdMiG4rG8L/yFRBSoHk0PjNRstmT5VI7RBb8l+mVF1F0U1GhkufCo7sVE2U
9ATPkJSB4yeuJAK2B1iOzM+AgPqk4st49ZxNM0YldzLsAiAD8//Esx2mMDhKTIIf8kMCltjxLyvq
f1JJL2Bo2B0benacZOtJYF2TMKONXJvZLxi0N7lGGsrYC217taCuwtcNSXvFas9dFhIFP0JhqSPy
fAHy37x22MyBICw0F/Ogt4Sp4u9i0UWuPs86/eWy8kN4xz6v0ZAqZJkW6iGmItA5V6eMsa2aJFJQ
64ImNjzDq7w+Jf7+ejUS9jPlnpJXHAXmqKFSDrx740tRH8Ajh1tnLtQJy2JIXdyHbbO6iqzFf+Cj
r/ANPuyXF4LsgBBp6xYcshyYNDkV910+F9ZUZ7t/Krn1nW/RAcg6yDsSb9bOCIFM65/C7YD4o0zY
i4zonBqqv9LjAl/gEnb0DUIdAcne05m5I1K0kJq2Kzn4MbzgTVVivPwtcFOPlELZXSySpY5mxJh6
dSIvfRDEwATng0KB9JKATq3u3baQkCcKUsRh4pwA+VVcMGnpKlNz4SNA3RT7gFoWwDReF80LEjoQ
0TMes3sHI3vSgHdCj3Pg5pfNHWdpqT0vjswcsHHE1YqW6DtqaA3FeNFGh3U0tuN8c1eX/LCvcVry
XVuq8N7shtKgctG57t28w+Q/Qw4emSVt8a91LxBFiGdL7u+gjkcc68R3kOrBRz4edVbgS9cP6bAV
DvcBuOILBOuoq8088D+G5QZXNRusgdhIZ17ew4+9r0xJLM32LpWLHcn0R2weFZwM2R0me/nr4NAO
9+Q35RLHtBg7RnxudCr59RyPL1hNGGIotk/x1OfmNUJIlsci3REazykZQbOKtYiMpDu/NOdVcDwd
7cbf88YYvt2y+/vpX4CaKSQ1WYHnw0UErNboS1pN/4ECOF60eq8dYaAvWL+MvQAt6pCtQwK2ufLd
ucEOQSLw2c4cXZ/jEsqyH/+m64Swpb4vdck24ciKUkZAiyIHodMgblncOIf2K4kGQQ5vylBivOZu
dEwky+ecr7WeIdnQtZZgGCAUFswI5ZlE/LzVAtWIfchDsKZWPZIU3HvYXto7m85B5OLDm9GopedN
jwL88lSuas5QwyGDQjoY2e1k56uda9o3PtJFY0CvU59aAEdLeQeVj5cC0o9qfjaqNAHKbu+khWaW
2eFC2+rg8EpnnUKeg/oLTPZEODqDm9e6SAp0vqhuOvuawRDY8/2Mxps0yf9YhbRHl6zBUIWo0OnN
xerr+BzCjaQr6B+JyVzjFG1k4rh9DdJVnwrVTHPG3Uwv0unO2My9Xn2QS+kbWZAMzrWoylBRHk0b
LczU4SLT01ja3/E8qS3rmn8X/+zzNKg9OiqvWiK7C7uiYSNPxP8imAq8lWboJwWgVsz0TtmWUP4N
ItJec/+SGKZk75yupAQIKQ1IuniugM+7HiiQZJP6nqD2UtJk3vHPLo6D0Kl+TszbGCQcjVLuOGfj
xSn2ESxOLTkaVg7jfJO6vVQqy6E1Nu+h58fyCj6mukjomNqEF/6YcoksnSC8Io80QwXDiFVV0iNh
jLIUP3GqcPjS2o1dF/WRbWOGCtQnBR9Nst89jeGxh7OU8lbR3SFVb1LDX2v0TXvsXf4VIPLm/kv7
FqrOVgHptj1vwI7egRaPb4/PDSTQXqOgPpWkqx7A7mhlNg5A9g45Z8X+8WJ3/Wgxrv42t2tyK92b
d/3F7IX2F1dXDTxkticR4KHswAyGuGOAxSsfPcDrWvfbq4DlIyng1szg7EXn9jO+/Kr5EIjbTuZN
MLnGZ/lE7u3dQhsOvwPN9bL39O77uDnhD9i2I+PGbtRJdcnUdSPl3+6AWG8zob+PDtnmN8YI+boT
XT1jmW4OnHv59tq9SW0I3GcNLnKavjMO69YsziWHS4BUJNv8xSzFnr95Pcg+I8Tib+4Nz8f22q8q
XOw0XtdYX86QP3TgbGjpP0+s1OfcEOssBMynvRmjlkfEQyRVPK+m1YT2URa/uhNShWNPtyW3iikW
xN7g0ysxsgX9n/jbAF7KBQrMwD8s8cCfRXv/RT0LhGqHmF94u7SJ5iGpYJMkEyNnYb8Nd9Y2q7XR
RdavCTuof0S9vzf+E870FrahHhU7NtzIpYHO7RzGdvrNV8BWSJoMfSuccxUYG8pqgpwl3DY+x+Ha
NI198ggVqCe/4bwTwtf2PSHA1S4OhVcdYLExM9EeFT6sZ05S9srYJj4XnNHhX0SD7ptn1LWLyKk1
EFXro+G/j4HwpQpO13fQyNix/j6J3fZvXxCX8g3NejwoBXOl3dt4kY7vp/po0xx2Bi09qnk1yyMn
aGJ5LyJ5PaM5k1idyCQqHZgqUbqdaSCftXurK0EwGKTAhO8Z8Lo2WLvWuZqtFXmpzVE7exOrlYOr
HGPfA8O0AT4IqR9OXhJ0gDkb3Iooxrh8ecn5n3jh1k0THOCAMm8Cvg/QM7tdY/xLs2FDZ3FO53jc
eYp3DrnsQ3zbk4vnPp6QJZqFbQxyhOEYVwkLZwg2RUvcNmOUf9e36AiG+/XeAKeMp2P2k+jfPKZn
5lTu8IUaDy+aMpY669EhVCjevCQfNJ9MXgZrVwGBunKqDISnmgEuP1fx52Cjh9pHRiXdu3TbT2fX
s8CU7K3sd8ix1/tkhQ7D5596Fo5YhcSg1gmX/FSX8bXpUuHn/wHPpc/MCdzUErOPTRb7/TTaGOdn
sx1+X3oK75RNH9Xf5zsUqWEKWPDU97zX3ynbU/xJWTBnpbc08B8HktMB3bSAwNVNmtm42t0gqOpU
MXg8at9ncjwdRBZAvJ3sKyVASgC887+coA73kLovVpR/e01D6ABNqoaVu34N7z2NpxX+Zs2GJEYQ
ok6N+QxRrkqCuTg9StF8kzYher9rMp4ovav60Yd8XfuWYJc+YIEFAD1M8GJqbb4s/NQnxaVw4j5S
WltfsR+msza7WS7nGekl6IunbEbZ5jz/1hkS5vTM20xwtZI1S6QrkllJwmNWGt5tuqSdWHCJjQyt
eIbqMpfmwaGWRQhzy1Ki/wASoD52WZEGh6MTI1zKgZ+h7BJp4MFuLeT/dMHGPX1896sVW9aYfVGu
ibpkUEYclI5symTqFZlPnKACRFt/fNaSOin/Q5AIYo6Q1ldIwU7JcjO7jCPyRbsPkCasJMogJZgQ
q9gvDxGGkeyj6j/Qgw2AtJxfhBcW5Sbc6mjj2necBTiLn03p+4GEEeZ8RuxYWn5HhTmRfkCQvHQO
6VQFeVwT78oryycn2grG0a8SLZg3tfn7Da3gDYRyD41uOebohXZbvDqKgjoJYTwYlLbChygHOWY3
SiDzHDpFUpwvrKNknncUgr71jKkmrmmSw+jfLWBcBMCMvlp3jGFsU+eiVch0+8LvCnn6RAK1Tmot
lF5k6+Qp0rVcIZSumqFWa7OABkI62onTJWYcdsPK7VWuosObSUHhg05CAYj9tFqnn209mJY4EfQg
zpSBQbMYqc6THoLwK5CxEguQAa7rqlANQRtjQYoyhFhPp1N3NcDdYeSgb6yZDbL5dPBe4nG6dVHo
2/KFAxLX5r/MpK8Mc6lf259uoYhnVKrVpQUCdlWNgqL/LVF9qlDxHzoCmyA7LiBPh6NeeNMPUeCS
IEZnkmrc/v6UJ1xarKaQ/WDuLuLpHH+TiyDb8CpEZixVonOPi//KZHEljpP0hvg1BRAdcnO/46dh
AZ4MtjWA8ayriyNi/cj+ZMYvBRmsRjI2I0UDeEJvPdIYF4XPN/+40e2xjLEcFy8uUMFxW6/MEPMl
LCe7k/sOnmbdOzFI02dsQXhcOp06+zZW2Ufhjva1iNfgcMkFRYR4tLXfGOPHaGetSDr1mtGR1di8
ndyGgdk1ft6oJc8nQvpI2MsNEdvcTIz+7E8d2s73n7gY8G/He94M4NBOyMVwkcXBARNkazUR6l25
lt8fRX1sH1wm5/DODU4rK7K/t76V74ZKD+uTbO/LA8wGZlAKiq6LpBcEeHIp6zSP99fdJM6oUiNV
QRjaAehxXWyUzj6NWT7r/bFjux7ZzIN7ym7B1ZEYk5kVer0N4L13MJ203plaAGiDQZ+a0Msrz9pr
NK+mPKfs2EAY+MKmZ3RqS5OsBNVkRHCykbXN1/2VsxuVlC3e+RK8EGJWZZwaWCDbZDPjCpo2T+9/
jcNMBnFOnEq1AjQMrivxWQ7c8ZuqbCaFip8l7OW3d1ne93ZV46ZVmz071vG8VN46EWv3my0sbIB4
4qhCzm31lbPdrOxvWGC9OY5ZGM/nohatV7yw01DfMZPpHNp2R3XW31Nm1J2dNK+p+YbOd+I2V0iX
kwKc/K8nBL2neO86gTLs/jsrjgeEB6jOLnpcTnmJOJDCFO9olOY4yAxN3ldRRbuhQaZlg+jNZgM/
TrJqlsLliZFFGxNwOyKmzxz87CqRvC4+hzpAwgCiSjmOqRGa9jl+DXwMaHJSRxFme+md+lW2ykyT
CL+v12z5Qc1rGnwxluhOnq+B14N0aIv9c236MmzbgUTgfqGzoOJwguZzRH4tEugs1WprEraMcgQe
DVXWTNShyu916MOJOAFgLQHd3XlNsZSenKJcTn7Fb6KxSAWhRrhQs0uEbdDY/58EXWX+9WoJDvZ3
Sa8sTKab34N2rExEne124aB8MIJoa16WcIWfVuIZ33ViHaTXH6XhqxvdzTtnklIaae2Xc4B8VDgE
j2SWynPdSKNP/SA0wz1dSHAsdb9aNUqGKZLvTWqU6/p7rhi371UZHsY7a4oLW/iLyokbceOOzjEp
/E+J4ASWaQ5xyYb9sJzKdj7Y7hpyYAqyAGYV/QJBfB6+4E859GMmQeOXXKw52nB9pSXH1iS8ARnE
iOUEamebGH+P1bo599sXijL+vbRu1Rn5/Y9ARsKi5tqC/hGGi0OGUS3NLOpJ3gaDnGCAL0RGrIHa
qFnrKD2kaIhqybEXgnIoQB/mtbwKVQCnH4fvYCrPH9a0i8s/7Gz12dTi5BZNK4TXVw2BWHkN0W06
OCgdUO//qlNeoxFXb3De4/Z4hruV0DHwAJa6d6npPRyVu2sB+j22GHeXwPX66EWLYxr+13VN4UxP
VosKpfoknt2H0m/EMxPXtIFHyKTAKPpBULS+zes/OkqsODc8iuOYcCIjLbUvx8Pct48Qu532GtqM
EwD8YbC2TY1fVRsy7GuA81uzmXkUqOg11DmbngWIWfn5MKyPoLgAqsoHAPjYdWUfkFjKbSeokcN1
7iDJcwsgvuKcdxECr89lc29eXHe5VDmtCG2gEkC5MRcGl4mtXOStKsIm1J/PyrRi5a1TUAfByht2
asta7aqe8bRmqXcQt38lFVEeK0LyPwOf+KzoXZXh9BwYbWrPAn7PU/VzypTu9wKlLERLINFJsx8W
sDQ8x1PIkmRK4jUoDqWFFgtw1GEJccwV5o5O8Oce4xnn3BPYkru1LvR9JFYXHdlycc4+BWU+IRh+
8N3iZ195lnFwHZf121UssAOEXZ6HqPZngSI4pQHdvA/DavlWcDh0P7ghwIpVEqhp+JESTC7ulbQT
XzeoY7H0wRhrR5IDZczRn6g+SWQokelhP7wq4gmlT1YtS/VyIYylEFjEJVyMS3NSVHit5KqQcxZo
ytuxBf/KvVMdMbYVv3BwMAxcoAU+rHNknTjcR/0jousE2vk34+WcAUuErRTGAchO/PYNUm/agMWa
1FTMGXUhqMh0Hs/khdxsBxJ9l4YGgZfPfUh4aS2AB/aScOHwFZLX22N1xsMriH06tIoOA4EvFlj8
cVf0sQ16pmGCJoYe11R6/gZtoZdRqg+YNHoFbjTxgx1jgbWI1QW5RgBnG8Byuo233cFkl0yLoCez
flgnfrRAuYwrxoDJKzSzMgDwExtbKyTUbufu/B78/jfmFU7tgqhX+vwQHgiqcrF2MK43eQf3bU8W
c9B05Detd1yB0GI2cEG4y0vsa8pbhta8DvFY8BjzQkhMBItVDmU+YBnwEbjGDOr5kTJNbtvJmaZX
ss4IQWqDV5BjBuira9lfHWXxyFBmsprrxIKh8DNrrs+HetmXeLYVP22qjnHxj19WJo0ktkavDVl3
IHenTx/qDvmvfLyLyvooxZg2aQVL3wlQ6kkhvKtsmSbkzjyKdTfynIsNoOMdaJ7uJDxSFvpp9pti
y7QYtM7xIVEDpaX/2JeqqqZwrMnt4q0XEIoCw8+pOY9Rg6gdbLXWNBx+Lsxk1mStk34wIsunQnb7
0PWeg7kJ/nOr81WJbHV5jKpgp0cgK0DKZZnlvtoEgKtb1WbWiSrUG3pzcrcc2CY7H+gMSUMJut1a
ln5SWQ2XY3/eoP4DiK4bawkFVl1xK3Sfe0YIY3WXqw+RthR7I2ghdVp2SvKu/uml7WGcyi9DWy7R
yaLUgI7KVpXv22V7LZhU+vfX5mkyz8jwu9I2QdIyDAfP3PcdwnJRtXX+ur9/MjvwNa1EC65mvE8J
qQPJ7AOUfqQ7BwBYvLraCJMNfLDt7B2sI1HVarvERYNGu0Nyv9xSbQtdHh2BfrXGs8kaXa3/xWRQ
crLQMCTH3ArvTVnqSXIJDuAhBNclqyKIwblaRj7YT6Ui6zfYBMPNuT2myfZEBPfLK/KA2oowQ5bb
E4Ku4LRA7XjJrxLandPspK2h5qNhrgGf6sFUwwmARDHrksUMrf86GPq1Sv2QqMLyflSZjLvz/RdW
E9uFGon9/MsH1kAAMB5llIOR4DeoPRTpob28DWrrjrd4GNHynAQr5rAntx1FgsF2xmo7PgdKJNVb
fXr+LEeellSBgDmAiWXhhTVUO0lSu63SfdYA1NZyapHRBbDZkB+v+QzEs3ayCUvWW76Lqjwaf/VO
I8h3T3U9gmwH3xOQ5CeU9N/pJmUbhmAA6h+PVJ/XIU9pGcCgjSjIGr5ZSXjAzDBLoshEiCmYKVGI
0UWCU737rSOnB42VTzBCXFGvKIxoY/rJ6OuMdxgFt21UwcDs2CY5Slqrq6kuQ4ubHssmKuw8nG7O
JwiFIyFIZ/1IiYZJ3DXklOujvn5UQgEmLOeTeaKTe/WvvORrctdIrHwnNhKyGnTI9bWAl4zbUgqV
mzwh6cSBQ63DOhFZxImxlKG6vtZi9/G9natFAXEJN3o8DCsBF/ZCNwYz1CzGg5vgJuD7vmk0CbwP
+J4HDB5J323GPQa8xp2tE3s2fcbvJeElV8gx97J70pmah3S+JBh6wtwhtWOVMrV6qgzCjnzo4RhC
KvmSet2uXwnXey7CskPrDG1LWFPS/kqom7mwM83XemtUDEIXH7OtZNRfTx5xRjl9xdp35EADtOBR
6bjOJ2PWiBuc2Ir9s6yxcKHPluEhR0BPFbZxNk2O1JFPz7Pd/73/z6ci4j9siljBhtjZBdA/YMNl
usd0BWj1kUW7LMaBjxzWJe3pNJ7zzw21+4ntb5ZeGScZR66XJq5WtF7GQnGri8qnth46HKqG4Kxr
NvSdqhINy4KKM0lqJ06YdYZ0oifve9l7inhTFkwREh0MD9LziKH/MbVeOv7NslPAGlGZSUS99VZW
IjJ8AY6YReNusEZNcS0vwztoGKVBi2Ha1Jsyi+7otZ63fTtITIyvqc4mEKjWew2HRhiG09ki8ebP
zkc3ByjFxLnNiIU23RIf+baox6ejlpmMDVnlJ7WQBt/02HQeU0WfvDge8KJB7D6xo3Qa4OpgYFwQ
whVYPPBMbria8LvglvPmP11L9BgyM7NshPvg+DoQTTx2lYphyA9Cj2tMwJd/KISgeqshSJQnX90G
cD1PJNWf4DDewv+WNV3NHyOkrO3TA7xRtnRh2Ineh6V5FrklMmIX0AwXZhrOOxApzgRld5LLNoOD
y5zxDmXuCTvn1DgLCWw84RFhOmqVudRL2287DB42rm7XjjeD0chL6lnapGvM2Ck8c+Cxr3u/E1QY
3NPlOUW9Fu/cnIGpHXLK2I4ctwXVArAgoH1yCUJHrL0rNZzx5szGgPwzpIrPHhviY8rs0spJ/yhi
qx1QaK321xCIpf0dPHiTq2/veMbkdlQI7nhNouBIztjbC+x9eJub0VjKXDL5L+Gmrqbg+jrTfo6K
58Z9RD1e+votanHSEgyxnuTTs6hKSRDThEfr/p39KU96gssCofhtX0cCXG/QkiryWYcfkSibeHqX
Uz6GK1rW4vWWg6a3XjDyGMQsjcq5q0MNB8k2gCC+JN+2lj1LCAqc6nq6uaYcqDYrQL0wsICf3CIZ
ULqvuADVfRUZu5nC0VKQzkdsOepuWnxbi8IIchAHLC/6t1EY/A+IRkLmlNC37LI+t0YwAVN4Om7E
QVlJxRA3drrjq8+SnsH363diGXaRnawLqJcMt1iA2OpgsyUDsG1iCwqqUmSCwfmSMozwK6ahpUPe
H2LQPcHmYgfLLO3NWW4t1TLpGyeWY/RHmZQu+M3luQlVu32qNn88ruU/j8vx/mn13oMn5M4V19Yu
ua1x2oAhq40QNBcc7ijIFe/4X6Q71Tp4N5fKRDwdVGkfyl7UDi2YcTCX5Nl9Vq8qxgqTi1TiXNt7
Qc/Q+h3efPnQgINk6lkbfVpTDmBXaJLnc+tKIK7Nlarpk/KvG3GAX76eYN+KrXiTmbM=
`pragma protect end_protected
