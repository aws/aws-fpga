`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
aNdoLETZdauyAtxVNlGfdtSO9ITFa7UEdvkm7ZC9QnSghNwQwvwrGBiL0RciKPLDbIWJgwJ0RnhX
mrGqBgWM2RlGpdr6HPIM4eh1/LSqLJihdBAXUA7icsw9kK9BordoGGF3MgmdTeI/oKRXIEstrk3O
PVpvayUToqaN+HLEF/9LTXzVSP82GP+AP/vVu6b+0iBvKnenaAmQfr9vNeT0JSKrvy2gxPvgAeZu
gh07odcrVydk4IvJZS/fnZ7agaSoP8ORKx4FawgrT/V/G/XjZN+Nq0UZ71AL0d76m1wE1dO5s9JP
Z4b14hnpGdN7wD5xfBiifZcE8SErLmd4SPzigw==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
NiEVwxA7UUX1Qou/iq4SJ4pZlfNxbKf9rqn2dFxi26HTn61WFY8llMcqJCwnKhg0NsA9VSDjzoJb
7WjqsMRwpT3xQL5omIOW8GXn0/IT8hw6Pff3vikFc2kD1J5NcBlyy37xwayzi/TNd77naZRKtHTT
fLLLPC222dp8kS32U8s=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
RDc07/IFiCO43R20ZpSDAqv7WmkiIz/UCHy36X+r8jkvcjGT89VUO2zYtxE9A9/E3HADQv5ztpl+
30JhKl1/0vAFO2FdFXnHJVu3IXAChR78YO7hJgUUdTHCMSCjR1Go2C6qjlLZrcyVKVlcze1+7Ex8
eUnAceGmoyE7YKufAso=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1600)
`pragma protect data_block
I/fRiieho+rUQkUf3gN+XUx4Q6Qx9oCniBM9MINQS6OodSsbEtfR2dFQ16jN52oHANSFt4udHAO4
xMfVJDIiP7W76gbCaHlFPbEjmnRR06wq0IVMDtp1bsBDN7H4sOYZOBxOb6kbEol5DYHm/fEx0GTg
72IEuh5QZQ+v/WnvBoVqtonaMGqWcrBVoZ/asEKN1vM30SJa0+4Ikx8L0oLOfsI3/L3NHGiRRfNA
Kd4foZH++41VPzsyQCA9z5PT8hbbVSq1cAKn2oVamnuTxiP9xDg33iv9crBQUzRx82s6MBDOanhg
SQgKgwvQ2D6a8q6MU0gqTFrlPFsdVxp3QH8ZBpeoyZsAkrL7ofK6ruIloLQRoGsceWdgC4IqMP2z
bFkvPvN3bRTl5ijr8Os0xY+OKn8P44aPbzKbcrFz1r+d4pP0jOYRH0z/Ek/UINJMst8es35k0KE5
Xc9EmpNT4jRIG2NB1059JrsvpZ7JcRmxqTIIypiAod5RTHfB4wpr9RmgWCe/WkxjFLWedUMjdyKz
ArVDD/j5VO3hERGtECNCeZZV8u116kAt5IhlIqeLO8+FPGiOVl5Alp2uWxaOC336cYP89ztOqB14
XqvQGi8NycVxw1VfCWHbgbgDXvCYcgQ1NHK3rtQcJUG1u108LOGUpaSSEi8fO6jBYomw/FBJsVp9
T9irTx78DLj+mI6BnuFcpVM/jyQu1xI1RONvJtGyv8HWw1tqbu0yGbQvADfl0lj48KzLeayknQ5H
R5H79npl7cJ5r0kkHItUzAlzhzGckcD1SMe/NuaryZjZV3H8cTzzg7gyXfmjsY64+ytA1/z6z5q8
/zsCJy5xYaeJ2/+aWlYHGob49pSiQdf28dDulPsxlIHl7aMy0Nr0vxjdsg32bHyPci2NigLIsmJj
pQbKSePCbfhR13dJ0U3BCL2WB1AT/Y56xyH8Psnq8UklwVbPYGZJvSFL8XaTwYk+tT/zJBM2QKJv
v6U2Bl1sGSu/qe8OT64ONBeWmkFq7QAA524LsT0rAsKc/Bfln4TXLnmVdqs/tBTQ+aAVnRC6Eoz9
nuUNBHdRoV8MvT0C7U2p0zU681wPw0D1ebgRWxFRRe6NYS5o92nhyQ1ZF308xbQacD/CGasnJJdg
w3hJhq7LzaZtP5sM6JngG2yTRRx2Gx3a6p7nHLsCIQQVFoZ2fuSBR9jDVKMJzvcxmFqcMITioFua
N8JrQm8DCcOWXUdozThdbZQ8GuPiwFDVw6FXwm41wLQBxZ/sG39rvodcTYnrh47y7p/4+pxc+18V
m9+AHaE9bLZzA28AEPJxRRnGjf3OKo62f0h1APcuGHRJUu+Od0ToYgx1U0zm6x3fGo4PEay8KO6j
TUdf2389arEdD9PZQ4iLT3p4yQaUuPeA4iKupbluzTsUaTSAmdR7wnMyssu6Js2aD4DG5pTVVeTG
5hiCEqm0eFH0DyRKMgS03pNDOpRNSN2Q8wQqatLoDeQaMu6esmbt554rn76kM/7W03ZogaJ8ualk
Y5thiYeU93lbcP/aQK/5JGKKV6eChgaJ8pSt9987w8UJwEMNXZC89zGY/ViIMRkOfXDrOuc5WsVl
COj2Ed7Ya+FSxpoFa3XNPpqrkYMn3GveuVpqFlYFjxBsRt33sxjOviIevjVRBwcfkDEEbP3u4kOb
tN0oxuRlo2+0p4p6ZvkhS75i9OMr7VCCK2PvX0EAhxfYJQ2/eXkmCa+C9RtsP1oBe84PKi9Yb68z
bDrZRvX8Cy/emlFIKz0H3rKM15bSUWguOF/Ci90dhkBCne5JISMm79yWAWk6i1v92HM4DpZL8x+p
Hj2cdM8EwqO1QnZNuofGsgCe5/nZQ/lvlGeyEozWp6YPMHxM1/i9K/peZhPnsiWRq5v+F4oIREBw
763Lej+lJBUP9/UkG4wAcXiVXTBndVU7zSOf+UxnUi9rxMhUj8QCXqvj6SRwTjOdM9vL8o+imt9v
Wxad67JZAsTldUdgb6M48bMjqZRBgwWA2tPD9P1wyUtOrVnltnczEAXK4QstN5fCPt9VI0Pzm5MZ
6+yovr5V8Gc8GgBZTHN0KVY5seI/Csqs31daDD/9/cxR+XkvsG/rwpbVUrb3Isr/l6A3cf55owGK
iA+KlQ==
`pragma protect end_protected
