`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
F2ysZjYUPgrh5WFE5W9zoQm6Z9YDqltdP+nF1wjJoE0ZMfUkeSFL3vCSZ7T46E5nyutVYIk+mu5x
MAzKX85scsQeaB1JZFRO0ABMUyDtoVDSL9ClGBJngACO5o6WDyyYIMylxG+uVsBtULEnZ7dsrK2Z
+9EJO50R7bJj3THlFXEaGaG2u3M0cyDfHXItxkIi0ySYNrKeyl9i25fZ5dCkBT1HbkcCEpULvcI9
U3BPzw7EENe2+KCd4Ue0psS0tXrz+OOSFNcYQJBnDk2AO72N3S2ceaOkGpm5cncCMOdVt+XYRt6k
cf4N3lNrUp5JhxCkwgsqKvJICiCfhBZn2nwgiw==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
3cqwOO9qJXatrM0dtFn7XsdWg6vqWZTCLCrwECkWfT+3v/A0fAiyHH7XwsUWlD7jCvEfGcbvvQlJ
Nrh8R1IghkABx023QHZroOhLJQiENDHrRSbOB1G2XZKOXkmkdrP2ii5vQs1C730FXQZhBBZRL7j9
GVQXXNH+8J6dqiwy+fQ=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
IE2HcSlJ5xe82wMLef+PLL//us2bZ7jLoUnDNGwT5aPAPl549nf7v+uk/DSliIQkLR0K9uHgAZh/
HkAeRiDpcfSn0WTccFUDuQpTtvg1Y7FcSGSzVEh77iaRP/tMePfdizvIBNhKoHFd+r8hZRjW+XGi
3XMD5TJy/NrAv7F+MZw=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3504)
`pragma protect data_block
jWrpa8CB6/ywgIG2VnFYXZVyiAy7/2Bb9eZwDW/CPVXfWH5CkXbJWi5diQZoChaGj6agr1/vbmf1
YZ1nxoUwy/HXHc9JXdma71wnfANwfgq9LieSlqS3mG6K4VJn64ezirUIfgYz9LAeHzqI+AYUy8Fd
q7ftmGFLicIPun0od7so6qFAGK5XchgoM9dhpyX2EMDxrrtSPIbhFdAY6KXVpsXl5tm/WPk+CE2X
MKeOSG9MXZV+/GwotC7IKwrqXXEu6lEn0ieM0o9RyPVPHnjWjOk8IBMOaKHa5EVFGQaJlUf/JMND
ZhVrQuJ1zx8x1UPTZCX/siFnDIARMuDZ8FjFzvd9hnX/70sI4MzJcKgSYsCvY+A+ERVlHr8gJENC
h0nsaHtpy8Vl5O71hkYvye2c+QVFZCQBIcyhBlcE5oFSb31ddczX1zEoiXA8YrUHPL0Ij9KfIXLv
+P64bydddxUpPvzAMkjsA1lALc9dNP0U5FtffqOT/zFTrTlqDzzfGGT3PBheligK9xyL0mKU0m4h
fBNto6377OiB/AAw3u8SbPILCMbkDhVzbrZ4+zRhm6sVbMoAPqAKLbPbO2giCetCZOCaLwFClFam
aBFa1HmCPX9QAG/0n7If4381bxFQTzOjeMsfxQu4X1voO37Ozx35d8EaKhwb9mI/zIbbYdTKb3rL
il0b9j6pFIxGttv9kUyxspSEIaEyGbUi8JIRuD7puMOGIYtfDFMyeiVhFwrpa0R9twba3hEqV+yb
cHseKTC78gd2AGzpIltxHXHuQk/8th7wrAdLB57wDTi398/sTrK0E3E2Y+uFjkaiv76Fe0ddbhCZ
oBdeklKNag6xoTcSVrsafBTazPMOwPVLBJIZzCGXhPEKivGnb2K/qxhkdOKPiElJv1wr7yvAvRyu
RPo8SaCM91Yrr8Jv1h3iiVlANXkHnaPuriS6JCYu6Wu+EcKlXorGbGQaff2C7kX7ZQLN6abklA9g
BOzzPlQf1SbiVLfUTeu1am2v6f2syw+U4HGtgsa4QtlL/PyLltYZ6gBzsEK7/n50I8OT+1oZxiCX
TQTmEaCT9kIw3BuKcDI9sxqZSEjoli/1ynQywty7I9G8ewcFQHqBmjKut0+Smjix+l/Svd9V+Zf4
xIozabG6YqS026gYQTep0gVpgZVgH0Um8SUHqy7AgzlRNwRiQlecDgvpxEF57f8zBt/dvdqEkuuz
8BLGceyif3aPw79nM1DhWLVKA40QZhF2ZCPuW2GeGhhIRPWC6Ouxz9voXW4kTSz24jqaFsJ9q8BH
qnDJSBzEBI9FfMAaSXw3oGACReJ9XARyVftb3GzszZFG1vet9QubeJuiP1YLkUMKfb38IXUUdl/o
0KvgmtAJlH9ZOu7F9vGSEykGsJEbkBH0l81VNlQurqkyp6v1cWjLFjowempLmWm9UbAGpP4DoHnq
cThuZoXsTlTlLWtPsLTSY06uRjtjJzlJGb/RYH0K+pxawWysk3uZrvfXNknwb6qrl9kxYg5llzvA
LSzlLwoxoEcPSzX9MUZD5RQfYgnaKpZy8qhfI7w73ukl6MvBURIg1Bp+pmrkwPxs87VfUWEIPif6
6gmbARpHO5k1byfaeDIN15JQF0ZvMpIghTlAIh/ApHsJC4dt2muGQYda4cBO7Dy6GRK/IwNCUDvn
4Y6xFwJ4FrzStbohFJuVjxzyCBcrDb6BkJ33fHJDkoISyp/F4+2R69ZiI0iE8mJ8BjRFjFFQDBFT
IQrgAmlUPkUXLA8iL6PDwVDWChKYIyE41IZhN0kjgF2YjMIL5Yp5QhyR7EdDqlrilnP1BwXhDfxL
Xn0e3OpgFfFQRUXTnHJjD/AClRZWLMLHbji85fitR+mUgxSpzsRcAZwCGj1eSIQHCUlrjkOYfPx5
VtsbJfQZMIgb8S3hOVYiYtDyhNr7GmVi8iXm4yNb6fvK7YgrZozK+8pXpQC+LENdGTHPvKd0mfSK
Pud8NnMwcI2GqmIaCE+3mamAIE2p3KMS7M7bWwuRE90oEBnIP3jBHcVVB9DRA9kXnZSh3RDkM+l5
6EwwKQg3BrPpf3xHQPQMavbw9/vJjOUJ6ATyXdfueT4MO3D5BIBqNptjUBBUzThZ+SwGWgtyVLI/
v4YIK26Q+cWkgvOxoZzHiohI/+4rV6FoRm6QsjsqSoxuzXjpvwson7krQJ+o9HUiEF7QvACVK9ag
HH87cDP4pDgbziXtm7uDTOopLyFQ/lpFUxnprn75XzlKQIiDR5/QYcAqK2qywaMZEL+bNLrkoFdQ
YfKK0F/6SXMEiBBnfb6Jz2+QVTPEo531pdnCy3+P7wJhGTE8WtzAaI/czf5C6PJQSCJv7epJA+Ud
uJz2rxYaU0dMGAZifHNNDURRtGWlaUNHXf3rewBVsdOcn7Ny9cuowNBG8A8LszVkCkTcFQxXtPQP
9tsT567JXemp1dO94obuEUpUppiO9e02t7VUu46bQ/HCrth55xLF7/hpJTPfbGT+5aO4xkZY3DIG
dp+Zt2JW2j8+uiqiR54aBFJyc2eYaT21vmv7q+8bpApwXXmPijm/6R4Xnw8ahbbRLA0Fw1/PATVp
jjoawSTyKHJlQ18s/dztxYhVciNoLLYy6TJFCJba0Mx4PtgBj77HcApmbaNSpA0d5+YS4GD7VHHr
aMD5k7N2eUaATZpa+GARfBouCOoUzzGPHLJFA/H7aUHPssZ47uJcdc+LotxLYvc5FBGlNpDM1GUH
0ZEoJkntheSbRSvQ0VlppRrRyLetuj/Rg8x9Dd7LNd2xOFIEk1NufGAW4lLIJR8G/7Pgd8q6YxX9
xtZ9DBXgSWUn04LXkf/RmGyNsXyv39iv9cvZ0pcsZuSE0htZGGLScXT3FezbksoyxZqyTWDQxfe4
lHUITP3ctlzVvC46ogm8eKgv+aJES4PkT7M9ifom8DqSfiahO884Hba6z5By2h2iXKVxHAfwOvPV
0qwXRm4d0VmBtLtJGDuOzypYtwKPQ7WGKX96D2LwYY6zyErghBBpmBKCwjFSeOxi8GPnBrC7Gq/h
86Em1MeRY2aDA4fS8nL5h6O66LH+QDREveEn7349b6LVo/UWWnlVMTOjJs0cDiV+S12mIX/tg5KV
PqURX/Kq479i6uwVH0zJOrymrNYoBgsVdTSDkWJam13l1BljVX7K8QN4pW9W6Zl2YNd2s41H9rKs
Ye0slHJgnlRnl2sIwZRtNLfXP4CNC4UVmgTBTEvLP5g+nZVxYASMQJb/txklS2VULfsAi50oImxd
jF8Oo3UrIM4a6B7oOy4uv57L1U1QRTQ/0aAi8oDRovXpuh1+gCIIGLU1/Dw9p58MfDoT75gkB9R1
svCDfe9oBK8NthpHQLykK3GU9vywrfWsEJ+Fu1SbBE32ew/Ny11OkIYitn1dx5np0JbjkXIJHncQ
K9mEvAAoD5CxmQdXxcJjABiMRQNLxi6u/7+Pb4+mcRSpyIgQ7yuO4tLKcfV41OWY+MhUAWaL9G+H
e/TfQfhPf2xBXb/vqBk6gHDP0vfHDDjLa0YjfxHkDvplugwePWDjHwnJjBKs38VFOnvwU++RDjzj
tSOxMNpZxCT6y/ggdbhylfizVLVpsapYdVZWTQFpk3cWEmUf8/vlGsFPcwpXsVasilm9J9R1vsXp
hTXZrJx/GIxXF8EYfqg7FTe4fE0taUyLTb3XqP7IpgO8Ug/VT3jgXHQz80DRdZ0LUvYoSgT/sLoG
tA1eM6uUff6AY0jud22K2jRm9L7nsT7Ufga+NhbMGuzBJ0GZK7BSlEt/V95jW1SPIudHp0Qw8YEX
QSyXcQmE1/9hUA9IZL/lz35Dc7vR+gSJ81PO9w8rK5Cs9itWJQfIrPFVXfdT4JEcF69pZ9bD1Zfc
JqEHZU5YDlmeI0YRy9noRe1VI0lfMvW8jv8hnFjkmM6VQHdMxiF/vBxpLfyEsj6l2tcYmnhrhKM+
FeceHqjLod3NPlslViTBujXNydVCkLCLWRh6Blb6o7KhQywgSARNH6KA20yr932vcW8OTJalNpI7
bXeAnrfDIBNxYWcFCxOgwN3gF3bXgBczyiw7T/tVPtRRWr7IXSl5aBHkHuOfKTlW8CpTYgcPPuQt
A3mY7Iy0adqLzDMx/RNQTVlFsqinjzZLDKJT3KWUkl/6u44EiH3wPfNV9phALZX1xBkV9pxLGpOR
JYIE82uMAPJ8xSYqnWrQNMWN49lzlyaIEnCccg4Op/j9w14xoqQfaGxaSQMdrT9PlDXyiQu/OyB5
pMfjd0Ixr50Id7LLRmkW5PZYzAJFNAGixdgZtN12/FzysfgSIqcHKVpXTTMrwnVH+rgxLBtr+14W
2yPfFIQObcR3UvysXuJ/h18NcvC6JJePciG0T3kEC6KQV8HHDfGnMNkqIrXgDWbjWxIEWyPy1PyJ
CllXXpx1v/3N7ymPnMp5xJ/LvdZXq/av6bKQN8FiyqtGPyCSQuz1tr7V5Qz22g+pm5CyNnJpq72G
NF4+Tn2ZlE3mB7GjgLepOrVFt4xRZYTe2HAvPb/Co3tmk/aTXg+rZnS31Vx6M7SmS/Wt0pmr3vNE
4TEbaQt0P53MPTxxsTJHZCCVqaRyM2ULKRTlc7ylSgXPBekc9ZFbN1V1wunQFHpAM8ArCf0ugMyN
+t1gbVViZ66pffdqa+VD9CJyd8ANHDPnRye8
`pragma protect end_protected
