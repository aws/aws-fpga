// Amazon FPGA Hardware Development Kit
//
// Copyright 2016 Amazon.com, Inc. or its affiliates. All Rights Reserved.
//
// Licensed under the Amazon Software License (the "License"). You may not use
// this file except in compliance with the License. A copy of the License is
// located at
//
//    http://aws.amazon.com/asl/
//
// or in the "license" file accompanying this file. This file is distributed on
// an "AS IS" BASIS, WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, express or
// implied. See the License for the specific language governing permissions and
// limitations under the License.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
JXm3RR2QGcKrb+XkrSOwXn7WPMk2C5zxWGbXkMFu/SGK0LOeqwWQ7h0SLX9w8ysXyrMQVdu74pr7
gW7NoQzqHgwe6Nbo8IheC89zmv1dpXyBaZKoVLHDYM5bYU0RprcddpTgiVXkiskuL6mG05kScKNb
fExeuzuoqq5qgAnde3AgJ+LHZoX0+dgahtG+VCeON26mGjZngf5wWxKd6hXrzPo9Ucq6EbwzSqsm
bM3n1QZEGzzIdl/TBGneakxAhnzf1Qtxk+yUsowFVfrM29rbvHc9H2SpWh+cGiDccNQNvEatYjQ1
ry1RnK2UtrLeUKUW4qsaPm0YXZ4y2C38KnjYQw==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
msZELicotuG+ebFkySzXcUE6xmTemgEwBKW9rb70jvlajTwsu48/zyiaqQJabO8hlOtLy692Ol9P
em9ndbgdlXizTehpptVspNQ0UELV6orJl5xEnwxyjxe+S88P+Aj3AtgsgY/iPi8irdlELnyg22yc
tKn9NAb9JSHM3OKgdYM=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
k+tEd42evZ0l91l+CNoo0+Fps5+yCzgU1WefKo07be9Xe4W08toQCAvxMNYFPakRdzXgjJCNPTab
hGaaiqaJv1MrZduwFkwNoaQx0tZ0/Z9WKvZgvkmhHQtvszoHlV/Ydjmog2wrPTenjyy2B5M2ajWn
wDN+dVaE1biGI5N4jCM=

`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
PnA9kL3co6mXzyzjIQhJcHbK8zRRF1ZhzafTkZA+5YgbEWcyC7nz/zG41IBJLGLsd8V7OSL0P/6/
zgpapwP5bg==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3136)
`pragma protect data_block
aQI5/7xfwFGjueggeppi3ZfbtyHOicIpoXMO0ZmFfXvhsM+HnYyYXc+95yffeXg/uBCRCtToPUks
Acm5Bud/h35md7ReC/tyO2k49eqaavV+x2Pw38cgfuwCjQVtrGpR+5zfSvILsUFnTyWIVHo4mH8r
4vQsjRGZ6oHZT04wIe4z4nfCCJkmeA4QL/iB31UZo/i8yPrI2CVrPbA7BAWJqIEhdSU0a+alxH6Q
NHSAWl3xGvKHOUt7I+XaYdTOxNIWVRtAkrXmHOLGcR9iBDlxXwN0Ile4qtmTuBKyH41sLHDtTOQP
sq1/US8D018T+uAAMXqVe1PEdepLh8bL2t42WXD0TOFt9agJZRmUTg92cx4rM8mYnu0a/LY8qJGC
pRwcIbHCZw1JvGe2LHNZu4fWws1gIiFIVBUAKx5WCbH5QXITVBsdSKWk8q2HzsEvRBqvCvUDavqV
pDTI6WXLoBGqcrrcfpXSAr60wwfTwPM654gqHniNcmFiMj3bjBGl+VNQLLct/GMgxJ7uZ3VcXlnT
DvoRGbYdLPdylwmxqfjMiE6TnQsuWaKcEKP4VPtUp5kcgRKTy2cmDwifPb3fwNoxNqeKF2s8cCvX
O+eV4P1f/ipeBUZnpqWpFNBmu9aE3EM0s7EPBUpY1U25FMRS04D2469iu2EXUE6/ndxQsR9gPq+u
Ejyd4r7ZH6NiXPLNylRfXapg5yXzaf5h1v/WQskZ7gv77+h4XHuk6Zli/ZUwdszH4HY2MCG7mH3J
tQvP3nV11om45l+cwZ/t7nBThULvEkyO7m8x+G/7AF9WgAxNbk7rvmCiZi+8ctrbV+1ap4acFIQP
p6dyg8vbFp5wEUh+CwM15RJVI9KBB+5zUpzh9ISw1iNkwr5c+3A9a9ZAoPIEFbXGwtAkWOmeGMda
Pp8xUZsJwUq3lz4eaBytBqKHx2OWYFRyg4sUv42hzcWuzZCT9isZoxUmE+fDaSrqN1AH4FA33/3C
gPn1UoMgJEEqn/n1QY2Sgjf/Op1f8Ze7OZ4vyGcjuGgPDsE/4R45wOP6Ja5KkxxDecUTZRJxSSnh
ywdWVbvoiZ00+xpB+obPxQcMs4t5xO5ppFt+UxK1IQOAeCBeN+Pp8SIQkcpDG8GwU7Kg2cu0F8K2
+EvlNYFHgYK0aIJTFRj1u9COpQf8Ym3fwRpJBqKqo22F70G6DbBAfUZmhu3Tey+ZiU/3TWxUHJcu
mKVzT5uuOw8VGbr91Nbie+FnBrqJ+yqSKI3vj/s+gK0RxYbM891pH9vzXdk/jWxqYDw894yriVJP
3QsqW2V56/jd33JpD78bPjforTNpPDrkp5S5wvAH8VS4BMPm4CmVn+75zDpbSuxt4cER3lyAqVee
A9iA9TNUQTc33I8zxf3zpOU2L7cXZpfUJBXjzYIok72Cf6BGOhZYEIlLRYXFuxGlvc0oWE1kwgVl
wUPtFwnmwOVzJ+QJA5SIGDLDezbYC7JMsixoZPznxw11XJq33jO/kJt/snQM15VEc0iG+W3l41bX
bztICkAppJ4oM6wjTiktA4KeuR9M08BpzfENuGRAv9GrO5iG+TDbSJd7GW+2u5HoBY2dFGD0/4/C
thp37kOOJElA6bNig7FqhApGmNfBU06fKtlQWGErUZmhm5qQpGyu/KEMdD22YHEJ6nQDTeMLQ+ME
EY8Cr0s8Z4rVL4YKqEIiKQHjfq36jPw8n5GAZjkoVb7O9tnslNZ/Y07DJ5jaRgcd7dABE7GlXtD3
I5OqpK0Vxz2Sz+35TS5HGR4QhNfmQoRT3j4Yngo1Eh69qCEz/2dp4UMIt55ruIQp4uumfH0jshxx
q7iw9h6TkhXaGvgIPbRPCg7GB3Cb2tYt3H91oUnSWIqWDXiVOkh3xKgRPAAYOTsfpBSp5Bjk9Dtu
t2YAn4KmyUSWJUvo+laAdUWMaqJd3otB0xkjTT8vy8bawjpsBuSBdFOa72f841J/KEfzZ8H/685B
WsiItgRpJVqug9MRa0fQzJOuOmJ/JP+sgNNz2S0Dp4uc3/6Y2YegVqyk6loICs77d2ilFiJGjxdw
gwznxjkeM1C6Mer6s5lb3GTztyTnZh8d6KfoG6IotmyiYR7FqyXOtYs1s1mGuFR5G1o9+W8NCw7h
ESQ5LtGAZ0Cfi98aiwNg/NYM7nFy4qaaqEXn3fSOSXzj9KgS+sn+prL3iW8M/lyCm7ECvsxzLjZI
4Xjo/AZILZgnbotbC9krREvQRJWoj/laclGXGP2u3rXE8idhjozLLET5nWpHT2EC3UFUBD2+afFX
4quPO6CM9lsLoyboQfgAfxR+G8FkChj96kHmTl8WZ2TLwqmHKRlNNyqKWje5NdldkyBIpXdw8alx
CHCzOITZlO2LtRTdzYJQrDVyOjRS/tnN9LDv0hQrSH4xqxYeLH4FGIKuZaK/rBHtQU+Bh68INYs5
WF7Vsh0cYESMf9XwLxmF37joiJ5Xvj+bDakXMGSmzNNXmKv/fwwFtlaobpacPftJTWlcCm5a5gtI
b/NMyj5xEUbmqLDdmHu70ezdkBRVQpianbdg35GdpWGRD6O0T3LCiovtAB8TraDw/35Djj4aWiPF
UFpWkiz+BH/BWEKbj0TzPKKla0ELTX8pKmUQST4+oBufDtdUvSFbTL1gPAGG8eVJO95k+zNBVUB+
kigyUkkjFDGv+1R36HBSYt0hxrQE7OaVBLt/mCYJ2YhTxnnmWkLptg/Qmpi+MXfKNZzPba5EEC+m
v4ztOFNic/1QttDGbdSA1S2EYOU5UcRRYmGP9WlFY8q/SC5RVPXtBcusGJpJ6fawXf5UtVvtGlm+
bU0llZxaOqu9QRRzPBNdy/j6VVRFZEK9RWvDOogxBKnpNfuHuIgGgDAo6NuK7mCnIZVpvFOvSFtD
1ZgBGRBDJmov9Axtw59p8+fevewanStGFjGC3RplYNCP1hO2bahXr1LYt6gRKtCdhAtzlrY0S3Ms
01eDn8C0T0meoafIVbT8Z8T5hz8ikevC0ef20OhNvtffPqTLHHORmVe1B4Li4Xo1HcenwHPm2JAw
6WpMjWV9K7TD8TH9rHj/d+Wcxhnx74y8IVTSaw0jze9p9+JzcTVZd+Ksyn8cnSRXfT8xLlfnZwyC
1RfNAgu+sgsn+TuvOhnB1BpdYP5TiaaQe/Z4XXSfRZtzOeIzMs2ZDM2ogLtsCqam11Z0ZpuOHsb5
5ZVt9ImqazT+sjU4dKg7Kp5kaod0jXnMP0xDyAycx2P1iAfq+pM1tpn01hqY3b9tmqsQerLYj1Yf
aMsBa6crxgWciuVntW/ma0OwmQaeBb7ufGbZNZhs0x9Xmmpfv6QLp0JfXsxYDVihbHKQzASM39g1
tIR/rSv16bO9B4kvIOUWckPPngmAquXw49xh+zhMJHmVuPujwiEoHA4jiHxSYQ4ziNGYMTH6W4fl
1WRQxFClopU1IqR18iYbk7j2vAw+HL6Jm2Xp5Js4+7ciai8uvKJ/9ju1q5P+1Uf25d/3rjLNkKqk
yy5DSv1hib9H7Jx8/9pYPO4lIgvMXb2f/au2u1nhWnMc/f2krcy58wnc107BapPEXZ62vSZFZoHw
oNziwkPTD3zx7t6tnMfALNf6TrJ0r5KT8CUJq7xP49O60oEPFMWbggIAfnvBJfuMl4kKZ07+yTL/
FaZBti2fjjCQCzxYOBDLLw4nsZEiswhHyvWvEnMpzyolmQSHH0ocBD4Xg7wfQWbT5UuFT9txZyw8
KrKzsHuRjxUxNLHfXxE0YAwFbXxNqYxU4sZvvq4WTLHzXtdfQzFZB0zicsvsMQzwCDBCOvE9YaMC
uxy91Lu0GQz9MIL3eaZzNeG8PXk8PAQQP04WbG+DCs+oyKEVnos+gz3yQuH3OmmBiWTmZidbhYs1
FF8yum7Yhm15VBbfnUi9AxsT5n1Q/4+MXUBhetCp3sZFj9w1dv3WjxTunYiPkykAs5/7SN7b4g+m
BQFLV1ZMjwCSHe1dMh872AsO23DsZN5ZMGnTpAVK0MUfEVXoMsxSaXx+VrsI++I8F2i9qyLS7Ncj
W2C3mZLCH77leiTeVJK4vBXEGnbLaxx+3BGn80yWxwBcjqA9TmPIhS999ZAYNmB9Z5a9pjPjNwGR
Gi0d4A4kzSeU7y8c0kxSuNhYCw3PaIVRWjvhDtO5nw2xjhc/Z4rBzowpsjSeAhJ6hcETT3NkO1zk
wA==
`pragma protect end_protected
