`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect begin_commonblock
`pragma protect control error_handling="delegated"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa", key_block
wb9tUZ+LDBSPiO/X16f3W+rCATIQvnk0Dd4QVrALehlEiyhzvKvr899ko5izEj1XYeCXiU6XYdpB
UsszEelQ3ayVkecBwqsuzcVBdA3MHmAiGjqmbZxjh7YMnAb0N1R1fISPvyi7bYfJCi7o53rdd/JB
+h/gncPKh4ee65+fx4uKtqjydvC9keLPGxSQ97I/WM6FfgJEyf2jnxHO8+Ltp9Sey1VN8zkjMLLm
HxeldqRoPbdQC1JdFfGl4+POOg22SXKsvStiQEvt5Hn8BnNfy/duc6ZuaH5XIBwnym1LehAWF24m
fkIaQYDEVSB4Kblt9gWiunb4V4hT/atSqy3+Zg==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect end_toolblock="Hs6IMtsaZvlEMdKTiqfb1x/B296JzHLkTmC9B6NO2us="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4272)
`pragma protect data_block
PepbZanmV3uYRyuU9S+q7sUUVjjkC+EsOfP03AzXE1IoS2VWVifGfj6uLQy5DqKyNbIWN4chFyAZ
iL7iJg71aT26ID91+1wR8mcq8P4tnBxq2JYZ87VjNOhDLYp1p0GNn/nLpKxmbul68FVwgWeZtdWr
ahzuTUDRh487EvXaQuhH9qB2IR4V38A8wmGCb9HhyoRRQWAz/CeA0IZbiua84NvYtiSuTZ/IZuu7
Z+3gKlfSg3eszB71aZsVqv1JiCqKP48N8KF2ULe48yTakhJFovqkwq8fc8IvC9DYyCgBc2haIHmP
zWbOiKPDbw+mVe0nzWVc+RZR1hZ89EcZcHt2klSFS4OD2LzzLTJ9Z4MPOeF8wE4IWj8LeItK8wRo
uZ/R6pqk8ChmQ0k5+0VgpRl1Yenx5NK989DqMiSq0RC3a06dFVJzpeYDu6/zesFbKQ7NAcZLZew1
+iCWPbVWyCcQLKQekTH41yovLg2m6LNrJBV+D3BvreJkbcIEF8irmuRDeS19V9NcUFLcjZJakIxB
ZMoq0KBuEc8UBNj7g28bzvhM4uu90Sul42YBnaSbX52UdDmUGqGlOI8VWwWG/IUygWSaHFDeNhNv
RGGGLTHdoncT9Ayertv+gMaDsw0HMwpCJc745RZxExkgzDUvUnJVwKcYaaxyGnQhUu7T0sMbXD4e
s197HaDcv7wL7NpTDlBs5hjcJw+BadDZdqhplCvOiPxMM+kWSVLh5g84bvUTNyIfFiQY6QUfoSKW
coSr20KLhaJd2QnxYZv2YhRdg0QVONcAqISHqwEekNuGqoWLki7drQJEOPRewJRrwd9QTwM/A9Z/
SXfrXoCg7iBWiYp/URWmR0PKc/e8snzmMZhuhQHjmW300IEzSNwB0gI6lcrMWXYW7f9iCzFrAI9N
Qol/IFnW0lBnWaG2fNsq7uSDXB96wnS9LrV7He7KwR6+05utM75oTH212tMUmBeWB7DY2LDV8hPi
I5z8EaN2jJ8gFFkI7IwZ40t5P4xb/dX/TgObcDk4egyorziB+MRcOkiuDQb1+bkuWYBBvdHsl5T4
j8S46cJN0avfoytUnmk36ivuhn5aERa2/PexqfmVk7bb2HseRs9Fr1URSEOHJB2exjJA7xS40yyF
FiX1k9fVvb/Cl2oaQhm34RzJov+S2ls1SD/K+CWvLen/Vm94V2PklZa4gE58NSONK01NsmyP+A6B
uVDTR+NYDrbW6Iwx03a40YdvQ8xavhNe3rU0XYArR8GgG1QuBAuxdTAYWrMUb0NtiBDCYPM38XZ7
qkfiGGfjCWknAH8Sqnn3iXiT17Z0GTa6HXR9JS+fW3VyWWEBdn5ljOuS/fqsqS45nV4YCJ2rCk72
2vX6eWLKfQJUE5s/Du5gNvVfVBTWxgc6XRMK6/gOguyyXR9U5+9anItS+0ST1FMFl/vclVPh8rIl
kHJezHU8tZyXzV57yGUpGbo3ct6N5c4LvGNxIUmYBOguSmHjJSPOrRVg1DBjYcalGIwWZkOia34P
QWKfrm4aq1PbMEDWssZ24ycrftqNwhSAfxY7LM8gSEPmf5HMzbezcPYjRGaiB72UVKulz9fVtS1L
Olw3iKqUXL0WgDDjiAjvQBAGPMz6Hqe/TopdqX2Bi1h6ZiClM6+UqdjrdL4H2TcjqKS0OR7ahMOl
D50ZuA9uDxFolzjmCujYabI1RI5xlYPZ1D5BpRueYfnFokL+I5jxikew2S0BtZgKpdDqLUy8a+TL
CccfgZvh+rLbq6BJmGBsIyv9+wC2a6G8n3xLyW397b+vA80fqEDvb+Uwi7qc/aK3Trj45PpmfjQW
IP7FNW6HAGJ8bycNxrCp+zZbCehJMbVMYo/qxp/w4qKrj6FwKl7MDofqb/+ob128F+o6gtqxlFbq
6wt6UJmMI4ZkiOdIpfitdu2OPwbyn5zeIxOVVb1gsYJbPhJuFY6Q0X3+00ZohIUFt09F3lDy9cJo
PaGn3Yu9dz9C3MnkCv1BJTqN/yyyC6HXOLjLnHEVSOsnUNmQbpV8zwoMMPdtXRPhJHyKxwbY0RDt
/5ortiejp1SAwn8OzQ0F+NCMMc9IxXVdOD0BB/3kCdEp6h0pxaL+WEkEe28cARqHNsx53or2Ehaz
hp1zLA2anzrYF8i6yJ/MehpJep2YQ8iZyyuQKgNaGXe8DVuYqRw0FdZKpUdR9rO9FdVArBKZesi5
4Lcr0KnEpWv1vK4ke3oNDxHu9LN+JyLsmEYOzb8ScmMhvXb+bbLRMlbkKsWYgC1PLvua1KWbmyRW
bvN37pudg6JnYz6ga83R14P6i/7ABnK56KUgIuox5lbaqE3t5saD32x79/W6nXt+232UHsMNC71N
4zKkGoy0b57gXSFI2h0uiUIyE7ajWKKHHwn2J6Mzo4ysuEwe7Vj+4FCgcguPdUf2J2jd5Af9TGJr
kndmdhdQxb+ohKiAhqr2IDUJwwsOvU7/eBpb82QBRKqISpSy4b41htbXCIEVylb0IX9Wm2RZc5tK
kzBBM2nkUzrNn0JdfTgZQl+5hL0fIrELYy5+8LO8Qfi6D7GQ2QKrCJSXm38bsbSxVDXrysiUY9dn
4X5kUvsPjFOUR4zvvIb2uPgxqHyQ9mdBfoEFlNq0FJXjWi5OmzDsOBceP9ofa7RqeSsfsWo+fXIv
xLoPMixl0lIEw7ccOhfcP0/o6LHSeMybX+Xgva5iq68m3WLecL/yKa8x99F4CHKI/hNUpKvW3ZCV
3uOceHRtdJEjzwWJhewdV6kfaMbFfUFbLaQf7CiG3mJY5B6PjZzush1ED3gkQZyFDrm0hxlyc+8o
Vl6gaoOkopkiWoW5Ge5G8wHS66mgocvRMTSvXt+XnAUI9/sB7aO7ey299+urM2oK5tdaodnJqNJd
2/suXaiZaSC3ElBFkVjYQK9FYz0gOBrX2GGW1yg+BtQVmkUVtdnug7kcFjfzMRNbuShqBx/hCb1X
ZN63xqU0+cBxp/fngkDd4iW+uVmdO5Gfa4lT4iXM/ja7gd1KB+wiJiv8EeZLrDpyCzeLN1g1rOx+
ulK5sUWRSm4kH8eolVivC4DtZrEzrPX8tpiTwLS678BvKojb0GEHbdIrjCCwPeoTX+iq0FTh6YGZ
nPAc8Q1P0e+dlSMR/8ckR4T6KrlAlbXYytfsL1iwl3opfA3aBXtL522wdt/feQgSbIX4ABb55/is
aXIVL/TcLA6uKSHGL/HiRA9HyGMiAU7y/SzHM46wtqi7MVkk6UjPUvIuRxBamoF7xxHXCR5GjMxb
uRatuWWahJa+4UAQAZJ0yhPg3w/n4//RjLkuS7PiV1XK+6ibhAq+yLLvibg3bdz5Gp9oSnMCA/LY
D07owdSun4bJaf1S7QfQPJ4slfnV5gfVeOFLo8+eCtrWaTYvO1aAlHptwagBk9XqxcYegqQylSxF
NfoGoAJ5inpSQ+CjEA07igY8Inxx9VRaHAXejOwNKr2Ye4Q2bIihl9o5HwSD2vwBOuLXzPX9/U+Q
36oJVIfMbAGhv09nZVE7oJPsskiJw13E5pbyxVsUdr5giNBymzdoFHkcphzGh7wgBq3RTjcw6Wz+
f9xab5xsBj4n0bvkiXWQuYxHtPS/hh+sQadcsg6+0opMFhXeas1+08uDh+i9XuwiAxxmHd3UM7DH
Tm6WbXUXdmc9ZhuTgCeb1DducuZD8zMF1BlyLPVluzgR/Vtrmg0Z6XNqnA8RIwOhxUenrROsDRnq
VGc+fOsclbyglaUBNDt7PyJ/2sOZtJvHZI6SRq2NNIukkP+/od1ApT/9W7TAU41tvpje53t1eA+v
VnS3ySUOMLku9QL/rwZRcXu0LXd6ZyLis2mY0oegCU45bZA6wmxzHifQTBODQtOH/i8T/fkJDkpL
ZgXb4WI0b1+yYElg0at3bKDlsgT61J1F+UlQMRScGPQJuoQaNEs9Q5m/leJGVh5j4sc/qgrbvZlC
xM+4xkqSp4/WrZILNfZ06MikOFOAu9PxRCyZtLbd9KAU4Yn7VA+nrB8fdq6rvwlnTLVl1pLBX2EH
2AtvaJJT7QR9JlciEjLRVNvY+ef4fXapMlsILfTRlInQvtjAjZFegGr+tvQ+Xuu3JkouE0h4FexV
7wSLLIU5kelLhBd3hJoIESWhMoC78LSTwa5DTANvNTVF3zORXeBQfOatwGiB0pcsXQDadN3/bFcL
r/paJjR1I+8mmp4aTlbuuNTiKFhOKqlW2S74yWbwd90vGKOtelcvPRs1cTMNzLiD21EB9dbuVkgL
yGMxX8u0fJhzN+stSyBnj+n81e1t5a2WPqZsJTnGai9nk7nzT2ZcR9rP8iMR0a3o+4QHbfSUZx+k
W11ggXb+s1ERro20Qbze/eAVCoEVCfxJsrxKirIMTxT2oOpk5VEiPt7XA4Wi/VefyozCFwFTh5IC
0+ZOcfX0RJodVWcZfYEL5EaebOHUhvdOiv5qGmYTn3u2qlK13z4jcrcLz6B2GWlXb52n4XOfsJvf
69Sr2Evllm3ERFiskj0eNvpi5JWL1Gyyn0x8Fiu1Y+sTs+UxN5k/996l7WKbVPubjrlgSFlu+9DX
7uX788seDtGjrptEQqzFztcU7goQozuFLSywOd1bk9AMwgbf5E6tA7CAa30aDd/5w/zBYo/NBIgA
fPh4+EL0x+1Fo1tyXaYQmr69a/FjrmzAWnGRJQ9ZlZbCWdIrOGNK2Tk/wl9G89EdYuXk/U0YV4Jp
W+ezLjhNDp41F7MyFMZBKXoQl8bf3fBC+HyKahxBIsnCEwpzTLGE3HMdzCpUhoMh4DDtpKFu4k/k
I3hLcAWQw1qx3rDtAZDIItSG7PJZui25e8rgcSSZIh2bOYUVzwRov+cBmuey2DX2V+2LzU8e/UdA
pdeNN4Iki3xuXxneTljVESX3UiLwFOGbm+e9QBkLeXteFL4z2HGWf4m2Oc/lc9pVQaJdaCnKibMp
4R8HiSqyCGPAdQNbJxqxdQIiZ3EFqPeTperzpPXM/5Vse+wkxeEoRFzJlvAoKVaQtrwvISgzFk9g
ZG75/g7SgE6027QXtoL91iYMs7WJy41g5eINwoC9kwHv/7MP3iNl9A5ehxiqHPffmQsnAoNnbWz6
RgjHqiGDSwonJb/zY1n18wiDDzetdwBbym0YQP+kBiLLB0g08ZJzXHdmXiLX+rmHKvA5J8Snmwb+
0EkKWJAyx6hsyxu1yp8jWMDI1zI/mJ/QUsA//SFiGDxJSZrNzyEMygoOLz8pdxDN6DPgtd3kv1il
jU3KwH28RCVMlOuad+9phjOcMiEDBQVKjxbvHSG41zuwSBGrEAY+MXLKUQwD4Ldh/P9uW+cds06M
n5f8DencE4uq+iYmOUUhK3rp9EFhu4u1M0UnuXklHr16SlaLk4CNoizlDmidh8m9m2RoIaU3CWh2
CEQPAQZRzGqoUB6iZpC/YdQm0I+utnE9mWnjh+kXVHBX8qqcna/YU2urex72ZyHBVXQq8F+n1e08
IpnnD/LksULSrON5QjXAqYpt5AK6MCnt0SYg/hlk5xjXt34SkYipBTRluHpqUDkp7bIA9byko+z3
DBWY+gYReSm49e4DYh/vVoWFvPV3oy3QyNeTqONuGF37Azl3LRL/vvROtF8TH1XuXShDKr9JzNUc
n9gCRKIvx14nE+D/XXo8gBRJdJKhbYcxKlpcC/aPMJ2fm5JOoChdb4mwxnFLRbVIZSSLewGP
`pragma protect end_protected
