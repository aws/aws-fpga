// =============================================================================
// Copyright 2016 Amazon.com, Inc. or its affiliates.
// All Rights Reserved Worldwide.
// Amazon Confidential information
// Restricted NDA Material
// =============================================================================

//--------------------------------------------------------------------------------
// Stats interface registers
//Register MAP
// 0x00 - GPIO 0 - read/write scratchpad
// 0x04 - GPIO 1 - read/write scratchpad
// 0x08 - DDR is ready status (bit 0)
// 0x0c - DDR reset (bit 0).  Set to drive reset to the DDR core.
// 0x10 - AXI Address - AXI Address for accessing DDR core (refer to Xilinx DDR specification - pg150)
// 0x14 - AXI Data - AXI Data access for accessing DDR core.  Read or write this register
//                   to read or write the Xilinx DDR controller registers.
// 0x20 - Write Words Low - Stats, number of words written (512-bit words).  Write to clear.  note is 64-bit counter
// 0x24 - Write Words High - Note can write either register to clear entire 64-bits
// 0x28 - Read Words Low - Stats, number of read words writen (512-bit words).  Write to clear
// 0x2c - Read Words High
// 0x30 - Self Refresh Request
// 0x34 - Self Refresh Ack (read only)
// 0x38 - Restore/Skip
//          0 - Restore
//          1 - Skip Mem Init
//          2 - Restore Complete
// 0x3c - DBG Out
// 0x4c - XSDB Select
// 0x50 - XSDB Addr
// 0x54 - XSDB Data 
//
// Interrupt Status0 - bit0: AXI-Lite interrupt from DDR core (refer to Xilinx DDR specification - pg150)


//--------------------------------------------------------------------------------

module sh_ddr #( parameter DDR_A_PRESENT = 1,
                 parameter DDR_B_PRESENT = 1,
                 parameter DDR_D_PRESENT = 1)
   (

   //---------------------------
   // Main clock/reset
   //---------------------------
   input clk,
   input rst_n,

   input stat_clk,                           //Stats interface clock
   input stat_rst_n,

   //--------------------------
   // DDR Physical Interface
   //--------------------------

// ------------------- DDR4 x72 RDIMM 2100 Interface A ----------------------------------
    input                CLK_300M_DIMM0_DP,
    input                CLK_300M_DIMM0_DN,
    output logic         M_A_ACT_N,
    output logic[16:0]   M_A_MA,
    output logic[1:0]    M_A_BA,
    output logic[1:0]    M_A_BG,
    output logic[0:0]    M_A_CKE,
    output logic[0:0]    M_A_ODT,
    output logic[0:0]    M_A_CS_N,
    output logic[0:0]    M_A_CLK_DN,
    output logic[0:0]    M_A_CLK_DP,
    output logic         RST_DIMM_A_N,
    output logic         M_A_PAR,
    inout  [63:0]        M_A_DQ,
    inout  [7:0]         M_A_ECC,
    inout  [17:0]        M_A_DQS_DP,
    inout  [17:0]        M_A_DQS_DN,
    output logic cl_RST_DIMM_A_N,

// ------------------- DDR4 x72 RDIMM 2100 Interface B ----------------------------------
    input                CLK_300M_DIMM1_DP,
    input                CLK_300M_DIMM1_DN,
    output logic         M_B_ACT_N,
    output logic[16:0]   M_B_MA,
    output logic[1:0]    M_B_BA,
    output logic[1:0]    M_B_BG,
    output logic[0:0]    M_B_CKE,
    output logic[0:0]    M_B_ODT,
    output logic[0:0]    M_B_CS_N,
    output logic[0:0]    M_B_CLK_DN,
    output logic[0:0]    M_B_CLK_DP,
    output logic         RST_DIMM_B_N,
    output logic         M_B_PAR,
    inout  [63:0]        M_B_DQ,
    inout  [7:0]         M_B_ECC,
    inout  [17:0]        M_B_DQS_DP,
    inout  [17:0]        M_B_DQS_DN,
    output logic cl_RST_DIMM_B_N,

// ------------------- DDR4 x72 RDIMM 2100 Interface D ----------------------------------
    input                CLK_300M_DIMM3_DP,
    input                CLK_300M_DIMM3_DN,
    output logic         M_D_ACT_N,
    output logic[16:0]   M_D_MA,
    output logic[1:0]    M_D_BA,
    output logic[1:0]    M_D_BG,
    output logic[0:0]    M_D_CKE,
    output logic[0:0]    M_D_ODT,
    output logic[0:0]    M_D_CS_N,
    output logic[0:0]    M_D_CLK_DN,
    output logic[0:0]    M_D_CLK_DP,
    output logic         RST_DIMM_D_N,
    output logic         M_D_PAR,
    inout  [63:0]        M_D_DQ,
    inout  [7:0]         M_D_ECC,
    inout  [17:0]        M_D_DQS_DP,
    inout  [17:0]        M_D_DQS_DN,
    output logic cl_RST_DIMM_D_N,


   //------------------------------------------------------
   // DDR-4 Interface from CL (AXI-4)
   //------------------------------------------------------
   input[15:0] cl_sh_ddr_awid[2:0],
   input[63:0] cl_sh_ddr_awaddr[2:0],
   input[7:0] cl_sh_ddr_awlen[2:0],
   //input[10:0] cl_sh_ddr_awuser[2:0],
   input cl_sh_ddr_awvalid[2:0],
   output logic[2:0] sh_cl_ddr_awready,

   input[15:0] cl_sh_ddr_wid[2:0],
   input[511:0] cl_sh_ddr_wdata[2:0],
   input[63:0] cl_sh_ddr_wstrb[2:0],
   input[2:0] cl_sh_ddr_wlast,
   input[2:0] cl_sh_ddr_wvalid,
   output logic[2:0] sh_cl_ddr_wready,

   output logic[15:0] sh_cl_ddr_bid[2:0],
   output logic[1:0] sh_cl_ddr_bresp[2:0],
   output logic[2:0] sh_cl_ddr_bvalid,
   input[2:0] cl_sh_ddr_bready,

   input[15:0] cl_sh_ddr_arid[2:0],
   input[63:0] cl_sh_ddr_araddr[2:0],
   input[7:0] cl_sh_ddr_arlen[2:0],
   //input[10:0] cl_sh_ddr_aruser[2:0],
   input[2:0] cl_sh_ddr_arvalid,
   output logic[2:0] sh_cl_ddr_arready,

   output logic[15:0] sh_cl_ddr_rid[2:0],
   output logic[511:0] sh_cl_ddr_rdata[2:0],
   output logic[1:0] sh_cl_ddr_rresp[2:0],
   output logic[2:0] sh_cl_ddr_rlast,
   output logic[2:0] sh_cl_ddr_rvalid,
   input[2:0] cl_sh_ddr_rready,

   output logic[2:0] sh_cl_ddr_is_ready,

   input[7:0] sh_ddr_stat_addr[2:0],
   input[2:0] sh_ddr_stat_wr,
   input[2:0] sh_ddr_stat_rd,
   input[31:0] sh_ddr_stat_wdata[2:0],

   output logic[2:0] ddr_sh_stat_ack,
   output logic[31:0] ddr_sh_stat_rdata[2:0],
   output logic[7:0] ddr_sh_stat_int[2:0]
   );


`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
YSNdkTQqe+SEc6Va5IruJ63EC+GQVQX0lDML2B77ereOBv/wgj6l7IKU5UXHmbtW9BmEuXesoeHz
Bdxak9QgkmvulqJX4FbcNIa2gZyeyUvTHTF+AsCkr43j2kI7AMCJ+kC8FulNDASxGgazkodFGegs
9nZzl8hRJDTVreVsWAe+AUksX2SPJ+1TG4EV+em/VNkR+BX7XTp1Op64zqLPV9uESzH+MwjCeDlE
R8M3dvubeHarAIs0OqMPUHnpT9hcafmfCzN8U8PFlqcNAsMPMZxqaMX6FE63WaOYaF4jVWPf74Lb
BoFS86lcOjrp0tOjcVtOVZvtyIdmAFWq+gS7AQ==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
mpKz8OyBufSMt2JfPeJYJawE+QjNe5PmkJHEgqDnYwhEaw3PPRatvCyV0/1NTUZUHVtYW7pZzBme
yi+xRBdeyG54C05lP3HCnVCN+3+ZJLdkffvn0ZU86UlHY9krzLEFfXEzKgFjsZto5mlsM1enO28y
LMkBpXRAj9aAiUvrj4A=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
YRKfHB1JQ5FFB2m6JdNJ1LjDAE3DaVMHCoBVWW0dUKl+40PA68LA4vs/1uFwHGQDYk0eipypFbIP
JmvuO0OoTMhOsugoZ0Y5R3eyAd9Nr7GQk3oK/Rcj+T2h1q/Y8SJMJVGtZodiTf/a2+KbijKT66wN
0Z7KZ+QFYhEtklHJumw=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 46320)
`pragma protect data_block
ygObws0xuBx8sWZ9+mVOL5PSbjVQxbUCsLVJliSnXtBOlBwP3Srq/MN553WalwLhQuLOhazC7sbn
ZSJGSJIQCbnL/6v2fHKg422I/s8TGPVRweDXoMRCHv4PBv2aesWCRVdONDzo1RBH8b7pmz+Tx1Md
BoD5E5J3KYTAz/sT8MDdrEP6gC36SC52Giq0ghUZVhiGGc2E0Bti0Hl1xaK5rlnPXAnwWz2N1uXb
0rAx57HZ/rJcszqdG1A47/USgCDIA0B3MIYURV4Qu8sPJ6X5zk7oFeix/WdpelAL4RLnNR12jPMe
VDPzbq9CpwQX7IfHCp0B5PNyBJdOSs/Vd3a7lWMKYF81xo4YkWGLj434Q61Z3VGNShxfkBFdgQhd
qwWW3qdGjtcfaXDDz78JxA6rrMrGASAOiaQJr3n9YGP1TVZoR0OTA6txoHYbTPih3hXquRuBmT0H
WfydsizRnrAIMp40+QVBjMhIHm05Q6Wec9/ENi0SsDmELuaIEkW4I57Nj6co/LZ+BR8udr4DpBdP
5Kd8O8O8b7yWBD1X3E7kmKNQfyU6A67esdW2UdMagQGsHMf0T7Cpc/bdqxELfkPoImiYrvLMbTHJ
aMFX6/IwBbTXIwD1QlKbn5o9ihLzSAtfZxAvn3+oZqvII3+zCudmi5v04PPNSOObm5nM4keHJpdA
nOUXD0llLATBgfoWPl9O3SWC4oyyt95+NO33OMhTNdKBb8aRZlyxnVrnyXKjQPIiNELOHzTWDiWQ
T07/LtZr8/bsx+D+RIng3VCNel55ecsnNapKlVQdBEFNUOvNTFK/yQrlefIZIvcXlS6+ATBxho0f
zjVs6pr9RiEtPViAZjBta1DSHGHeC1Z43Bu3ctgbyv72/vp+cS2u56q9LccGfNCrvJ5dgVB5tw9j
j8yizpP50a6txfCQ069mXSlFqmcV6zekFf6hlZDd50w8kUvQDCqwYUzk40rL38yd6OSHNzDaD5RT
5/CW0tIw6kHiIF6YmZ1Mi9EraKM3KqHMASYgqBJorXGIFJnEuS7bi8Ap65Y6ZEwkgwWQ0/7pz5Wx
yfrc/JZdCafL7B2pQRcjYoqAcA9GqOlbs0F+s3U/9O7CR4DZz6DT4Aq354Wyh7opSLLoDt78qrPh
M0mkjMI1UYgMB368LHlIyozTUGRRHKFY3sP/iGZdDIBsErOr+G8jRFSYNUvXf1ZhcvzqhCf37hQQ
RJu19PL4ABwW2hjb/vcqulzTOxkXm3i5LzFtYUPUMoBcBAk2GnwYNnhNet7Ov/WtwFxpA+ax+8FQ
rvupegT8nBrAOPh0c22rnPdzYZtrFH5g8qpb8G3FgIxnSo34mtMLCrR8erKwdSZgpMvfbkbtQMuO
i33bOHYZUaNUeKDYV3MAPaMaGi4INBfvEy/OnY7TgTVjxo5udNb2no9vSJX25RMPSwNaCVOg0lhQ
rlIHxB+W3tD9lxcSaXTUUALQhUIrSu2GiZzgIHAI57lK6v7rRFy6bazgXIy+wNhgGI/IpnTdx+RL
cV4rsQAZ5bwfhGsLyAajzRpVsv+c/M298Wkh3hE0Fkhk1WEXypRDZ3i+qvGr1Fs59Lq53D2i/KIF
WLZ04m66pXV3+2nuIdbggsq6ITMtHsDJIrrd1PczQumGZsW640MxhSZtGUB8CAeVvUtppBy0dV9k
WwcJu6PZ5jw1zlXoaRIaVcSY+/lTEzBpvgkKostIJ9/Y0GnZutpq0vKJ6x8rMLaocuj55D9h0JVx
D1x86cMWQb0u0/dQlx3xtlxU04x9Q1GoHe/IYLbzZXLhZvrX7qEzegyvfHT+XhcFLG9N0k4Jyigr
M5ASsmlxT7BSNaBmbrrtwfud0vYL/uXoEcjALdCQ9jPURY+cTtYW4n1fn7HBZBaowbngZPM3+mu1
A9RpfqTRPBifJ0YNCTB67o6TKvsDv1r0ArOQfw382WiwwL0MCGhCCXzQbHwUnc82iLbPk7rkB+uq
1j0ZtOUhmC+KDIHtLfrOgu1nz3IWhClzB6eeZifK/lXIt8uPdRR1aySiId/WG8kSG+z99R7lqmoY
ljUeD+eJi1I1Eb+MQm5uXGBq7pWxUd7f9Qu4IgrC1C7A+sZ05QsPP3W+dup4UixyaxX73ynkJyR5
pGVCaFuDaUAxp0GBIHeisxI+3yoHjnJEw92K8LplXAvCRagRhUQ9kgC5I5HfCCN2/p/ahA/N/P4f
u/xO/ABKPyjxgqiX2wdtJfzohRIkKcUnQV/kebGWEH1D/idY3hRbmRWdJTm3kXUthXt9OpGSlNY0
4Xh5szGApjY3onWEimpGRVwD9pBdo0PULURcmusRCLUHN/cVg2ydOHcd/jR8/8DY29L55eEy5ckP
uklT9hRC4I0SGnMOoWjz4XNjqc4G+zm4vyhvaS3oDLGw/bQLxzXe/5Ad+cyB9U/MRWcXCCaEjPWQ
R7a8b22xtnjyuURVno+F0jkh2ntLqN1OMKny+W7KQ6JWIw8REjT3+QsbwYGdM0NqDpyo+IW0zrxD
jEu0AASZjtOqwMfefPCwc5Vjs8sKb/hgo0tqFDm+RJPa7ksC/7PSG9I6+5Zh2+93Lpk7qlg9iucO
NjJ3gZA4LF+M5MM6sYsoKVdA7DSILMz+j7FtIXZbX2qwMtsZIA0dx7nT76hESuYZKOtgnZ6i1R2a
EumqlwyLfcAEocX9cmm6Lm0iF8BdQu0UDqHAPCiIhcjWx7m9kYA72oyzQli4S5w7rNthfC+/g+UP
qraYd23phhYekqKS3VLGEDBZq0g5Pl/s7PJbfXiT3y88xBHnpzcrNHgp3bTOKLy6iNZOuNNwhvvH
bgJH8JLBeUZQE+kNLwmt68ocbh++cX/r6flnLJp4RCq9M/BWYjgAJv+MOxOu+fjWKdFNb5fQuHyu
Dmwv5hEKc2tDg5xTJ2lr8GGYIvfqRpGVZ3zUlZOIVkxH4yavN16a/tpWPFJJDQmb9T2rbsefg1F8
P5d5B8QDQ6AKoaB9PTSMNfwqj4lCkUao+H8NVnifSZHtWPaDLUavaFNw5wQtYaulFSyQxQ7LOZOb
cRo4wmMno4wbfONUAm3fhOh+9B4rnVq6tK/LUmvxIR4uYuezoEUq0tqeNQQVNuGVQpSQivDAQKRc
/jVrTa0xF/ueGhWB6QK3gfxZZd8j9dtVwZ5UJbyDyCmY0minkoITHfTIT96wfOSnkuc2u3LNdpS0
kGE3DxVvgCn6Curh1Wb0Oqco8/3F+e8a6k9Gcs2W6KsQ2TOwiFFfHlFZ1Xk+yYvRqw0g8EYZZLUj
d7ZqXpx1BAHxroHXvv5sps56Jad+48ZLNlJBoxP51oSXrycB/Oif+S0LSg2H+R8LWmyy1vWXvgRS
1FQwwa/TzfPgrnv2tjzTopfQoys9L3inMD4owmjMWaukkqR5o+MXb/v/0nAUSOzXXhhIlCAHJ3LY
ZLlUsN7tuKRngJYhlVUc5oU18lVYEZQ7OcIPzoeb9MfauB3hvEmv5bVAByhaZ8Hvh3XO3NeoHcgc
6+H2XEXuIV2wvwLwH4EjmihtMdxVfMTCq+QQkjmUehPq6AFZGxkN3aboJmEl2o5E8bKCVRvZ+4Zx
vUYFUW9CCBPpIIDe9q0pNKt5KsQWEg96JcC158zsQce8OxtCMucJU0d1Q/Olu/7J5SOQ4kthXxXV
GVR+GkEYuI+neSEZIM15OTsODjMh+zC8a4z7VfbBdSA6Yt2sYNe3Gc+6cvjE4wDRti1IPpVSC0sK
1Opw9vQSfECSLDvZByo0yGmy6YsIKqoZqtq9I0NwVqB9JQrNj8DaJTBuM9BwWW7bQZLz1S2COpRO
NSam89AhA0QQIct9WGi5L+jvDM9Ot5E+SVW8nTCWDQdUincZNlWyFgaLism5eep8aJxwLtU/Wjzi
/Z/lvBahYri25IJ0vnxNfjWPt/dZRfRYvDjG41uluEgj+qPHDDH8mo8LN/iJimjndPnHUJLekNty
F+X7XQezY5eHBkUHpeaEQ6aXTjh15X2N4hz7YwOQvGBGnWG2OIXFReUWGpUQ67cNhfpcoFpXdLXh
wtlklXszDspBd9qJO8LHOzsacgeq87a31BPzNmXYglNvmkA0Wk2MaTxp8KVD8spdhc4BCsRRB9qY
N8F/3J5AI1XB6DrU6D5c9IJqpkeBGC1vHZDAZrvX1iFx1ynd/WBJLNOUeHmO6UFAZTIJEZ1i7n63
FVObHFlPHVq7JhcaCy5oRwOvOMOosq3uUwLwqi8LtxdXBYUqOPfD7rI3teiLxs7LrLCyGKRHDJwj
bfLbr6aYWRnYTQvQeoKdA7jAKcZzPtW277TjpClB0jx9TXvdhsRbWpchVY2zen0WtoS6NTQMMvYc
FgFjevzRNHIkAYD0CU+TXdowiylmJ2FtwZcsgIODQxNxdOrTAehj92Xp09dbzWl4BrWP6MOPETcn
xVbYhxuGgliqbF1SM79w/GGi3UhPeFJbqc+m9apoTS3+hdg8lO1M1ixkiXr0LBByJnCbH8bCA/Kd
RVw6a8R3KJHKL4Dr1H24qH1x93aZjlZjv1kvTsyC8nMQwM9ndwqRIkEipOCJAb4snZc9LaZnf+Hw
aj5w9Jv43I3NRTDZvckXUTEe7RuesJxUgnXJ5A37P4bGrDPBlC3vkBqbp6a0Q7RGp0N1ihqi1iHU
OCm5zSvusl5HkSksYcV+Ndt5zcnT6O5ZK0hrjcFVYv/aQ5DF3V5SOxR8BW9hEOD3ZIf9/bCuNGfF
HZbWF7NWIK6pa+YMHzDZWFsIREKecaYbEp8oCzDfaVgqt9EuHWD9TFIGkgtvN3yTByrjLHVF/jAH
+AoZk05iUKJ0zOMwpgNGEtrCwu/oIgWs07AAkPT4wz1+Cble/IkKwI+qhyEMD9rq4gheTGoELuZ/
5BlsbTBXqRxNZbT67yEBSR1zRqBwLNwfm8A/gQoQAGtcLxuNxi1FoqbU+uHTOC5/kQ7MHrcszvK7
sC8TekxtJ4ItskrLo69G03Ij4bZlZNH5582GmJkEpf9s5NKOuO7LcRgTAv+Jypurt5Pjid3gPBxC
PAK0VxYygKlcGwWi6v0/VmkigT8y9fXux5Si332SQ7egzFrGgDYvZ3xHvVBYikzPVNOVWb+o5I4Y
nUONZSJoBB5Gh/xzTVzUGAmFZ0gXNb+iFoNkguT/DFq2r43VQPz2wreD+Qt3OXWthJxHDHBYC9+V
Q7Fx0LBKar8CpjyZbhj+FdmG86wtuwYI8ue16GVAgtULHX3RxtoUWxFaAAASooduX/axaL8T7M7O
RJqtbncoD6g17U8o+lf54TbOCCe4zasvelben7iP+tHRuw4Ws07wSntCiaR78X6wM7YqYeRCNwaD
vX/4mFLPGh8IzUSjRYwI8EL577kaqnx2wMRjf6vosv+lQxxreVSafRTUMHHDJuzYllmQVNcRbhAr
eNYt7f0A+8psJGg773w+v5W7nkZOXNDfUsMBx6PD0hB1kMxRpxcFST2j5HA8FkNMZQHFJhP455b2
UUlGSJoluqc67OTLQ+4jJAIsRJpwKDo49mn0REhh1Eivrx7n6D3q8aqsSjNsd7ynL3UopHJmAPRQ
ZOt8wKfmQaJrtSy9ZolDPJB7X1Dj0Gkv9W3DszT5XMfipUhbtNn5p7+P7oZqwIbKpgBN8frpRM+A
mNVwA04gtSWNYXuMNS0YQDsSlSbROu5BxVuAiM8ouU1P0FReuG41hrPLq1205DfBwbDIpTO7G3I9
iUzFi4/6/DBxKwz5GnitqhQNWqgWnHWlc56KvWiNpzZAgO8/2cvqGsqnsDENbQzvH9UHU1/PNN2C
N2CA/Sq2aeabCII6mNtTn/GOZ5W9F/XA4pyQ9G85acF76Y9IDqWbEr4Ie+BJ1wEUI0utcSkyia16
wHMJtoPUgx1eoDPQyiZtLot7vdXEO/6LlxAqVqs8klfHmQrd/KHlc9NEtO0STA/lx39mOWgDesNk
M1UE7CowfHZ1na1seio5EthR/7l2EYy01+g1P/I0qkFlVZMr7VMTLo3jj0PA35VoPF6Zkvo70BRq
iuhcQJDR/aefv1XHIkTJuYpv/irdZ3kkWTXW2qvsaW79VMWwMtYtkqGhGZAqCstUx3i9S2qUymHp
pSmuEx6wN+Rp73l489igWADPHgulXllsB+i3FVMuoUYaJxKDYcrw5TRRgpaMiWZsOFeaVAgSI8o8
EVycMJ9lWBOepOhgWqM66QsePuBmxANdOufy0ds2F9HH7O4orzgwwlFF6MXjLUGGMl5MXqx0+wQz
hMkwkre/mad9+5GGdZzhHQ7Ogfc6Mye6YcEM/PzsgVVWbdgTfL9Ex5JuyqtmhWOd/BGktdJP5V5B
5Lh5tkojl3NpYTrMtwCrggdUl7DVMtYTiDZgZvD9ZtpFW2Ryjdm4QXUfyxPc9irdRH9zYdw/Kwhs
nsk6Q9/Mzq/pXDZQqCNk9AZB3pDamEgq0Tm5ON1oZ1foVnNYV5WeoPVG77mFTKbODFCTn1qNV5qb
KnjAYo2CI59NGn8t8/LwgELKd19TpEhCwIQ4TCI2YXDvAP4uInAXW9SUxMaScXM1I9YlqiVcPXFM
CN+FVV5tgi2y4uqqMolLYSx/+wLkJ11Khz4sNwUROz/fSEUJZbfFNUT5P73R5iCceffv11b5M3FN
MGb/bN1bAzsQLocGu96ubLMgJd/mxdAqvsQXUoPl3z/CMLyedipv/0IP0aRDnI/287u7Mowp4wnA
ilxUsPSd02zQp5ytfXFF9L1n+EURqKJd0WzbNt0c3hUXcH9jthsbdXJ3ICkG3Hxk4sisTiaXu6UA
Y+j7rFdRSS6hlYOFT42LD5w0UEVuEGscKGaScTMwxw6lC6sekbnYoNPfEtetRGvUUDVKJzUICkPN
ErVEBG+4CbdMvsqmuWY2FTRCJztvTXqyJgJ6G/htnOy3xxwgeV2eyVndbyyD+it64dkLlJHWKJpr
3Ew9YDbigA3mZD7KkuP14EH4IUdNX7ZMTyTFshc/uXFmGQ+OuuKmkVAp3+QwF4lzJ9qy6SWI+GVT
ZBoFFcCB+p+KTOeZtVfgnKgmNqUU8zf/SVCB3yv6XUZDb8IRzeB/syUDwjV1HTgaBtxNxrLZN7Hp
fAeHw/tp8KH13DXJ7At7hQXtIJhXbeIPtYqOVh+iKvdCU0cglKm+lY+coCpKHFJp0fqTiRYY+/I1
dkcpo2Io2hPQkGf+XO/CHZ/taOZ92qTskTNBgWgN9WZbxU6YajiAw+fRC30JgqnIHrarQn/x2juI
823JcPyC5bbEDFiUwMpFMf5JCtH2mc1MepEhkPXjH8DrGwRue0Xp389C59xSVEO5ekywW9/9R3u4
cEtJ9YQQAnri/zvWYnmQWv14w3Xkmn6+uMVTRXU9kU/RDGJaCuzOFvH62tonTOL38Dn0wvC7BobP
nwPxcYk7r/q+OkuZpgffyOcCzuftLBS3qJj4JvzCLFt7pNBZnQw9ngnYoM8wNuNS/o6O6rYqe1CK
NU1hly6M86SumIgCaK8WmpvkA3MZRaCuWMIZvFlpGriUJUXvW3EsuXQu/dpp/YMPD1gf0akNhZOs
7httYM8TLHT7m5Q34uGh6DrBSlV6Xq6S0gqfZXS/H5+lJeVJZo4iM6O/t7SS1aLBoEyrXde7pjiY
9qc3dSzshEAX/kwI8L1FeRqczlTA67xxo4elKaYyOhuysBMBPY8xIFdg4rMBxB9QPqa6g1yTnfKk
OEM2RpmAM5/PftVzlf3DXkWIFE38/vw5yVxXi7u8WSQnQiz3cAYTGg+5tD7bYfZfevSjwHbgXyFi
6S8yDERmzDd0w3qR2VlvHAkSBZNQ5qOX98Fq6kMHW8d0j1AKiONK4NepQL7fzlj2Gphux7/u0qhG
/UIFujMyiCtCYflcRyz41DXdDR50rQUbV3EkaoahLlE9dU74bIBxay2mH4AJtcFMX7rjtyEv7YjN
SD/NnN9QmNcJlQscjLTDnRd/0riAJrkgiwhwTO/w6zqhCQaQYw/vJt31iUQYGswxkk+sJ3k85VMq
YasReuEQmgSsljpoifV4Ocb30VNeg+PZoB6W4a7amgpgEP/Yk7+1Q4cM9nhjNaZLgwawTxF7cGzb
u1Ld6C7dncQ1xM/xlyqWtn7z9DYIaqf1Koyh/G/hffxuaf6JaFmOVOwe1hpTY2lGgK0yVZMrGJQw
AVm7q8oONjWqk57ExkHlc/6WLIvrbukMndYrT6RJBCBzQ6nkigaz3x51qy67k/MYalyT2FVk+/SY
/+BwH/XbNKTS6eE/pNbQFZ5LhMvdgodZz2MaNcdyshAI20P4d7rQ8x640ZFsJNqjAaDpmWjTfksO
qDn+diPl5NtOc+SOJy48EnMwd9H1Db0ZdvsS3Ol889WpyaE6sv9BZy5ht+rb8LMUbfhsJpjW4ZTe
7hUB1sZUv7IqFSBRLym4RKl1M2p9PF0mSiPTpZDBD7taq31iJUycIVI6ZuTW+WCd6OSkuMyWyHbQ
gNK807oxbpA+JqIQr8jiGY7ag5euuLH2/Qq1wIIUeVSIEk7nu8aNRRTeq3PfP8YPqBAorb62+zQM
9xHDqzbEXoiZcJpxFkbkO74K17Iu7goiCohqUFYilQD8cD4xE0abSiWXCsxJWip/YRVW2kLgM5oe
nYZwdajnDyvPYkn9Iiluidn0mCj/87tOSvIeykgiHh2TVJuHnU3gJXACxmwuaFRWS8N+Hvuot+BF
BaKB/RvgYqQyv9FjkfYGP9punJbjBh7dr+aWTdNgP74SoSHaN0qh7oHV3AGaQgV4/gdXBk1sfIln
4uk2sA2NnGXFsgAMGeJo0GtUHXkz1ueOFfCEZtw3HN1JjxIJckr8cTFyfPmcba1ibviy3NvPuKz3
W6tq9P/38UMGKjFpgDmV38a73Fr0uRP/lJM9NktafdbOpQqf/MSd6CsqmZWOtFz8oUvkRqUj6kL6
ZuekIPciR2ax+O6kNbzb7CqwMYisYpfbg8eF0fG/1M+aPaMqC9FGkunpAx6QGMkEOP6mOqQUDXCH
HDMYcGH50zXUes1P9oXm7houU6tmq5Ik+ujt8B5HYwQfnjRKr8KRseigJmSyB16e7HRoCejXsmhU
oK3IGrgytBNz76zIAgePlxGcSKJuLxuO5cR8lTJUxi/G/IAbpmJwvMc/y1C3MxaYvI4xnMacfhRN
oUG4v1GN2kwAxI2ve0yi/TP3qZqns6MqI8Ir9c1DqgNdPWzxHcMBRV0gtuyVgfUQkBgrCHIiXrST
MgaHvTQKfcWI7HsakRV35P8fBXTvVT0so/ecgZUUfy5ikyHJZk5DToKXMhLESzNGlxNdHU9xbq9c
cb1Jhe4RjE8QAK/KriPvONWqOvnWpsjLnm6tc8xEQHbR297GppUtBpxE5jypkC2EeBhRQHAQ3C3p
vjAkDJD6RGHUhfKzXcwwQRus4WVZkqc/ck4LNeJdYsnFRT6GhdzvliRi3jZNKm07wzh0QSE087AO
QgNJ/E9YqVVHfa7KaYPJKVYTRqNd9YYAUI9Q/zAp5BkrvIhSRYU9U61Zk8IZc0T8MNBhNzAvgFL9
DdbsAJZuVgBFX57oxsh3NTnCyIv+bxATFbkXEEYVavJshv51NnLGrMg5hqfsVPdirnyMrPk2Ax7P
tpjdjjnZDaTkxO6HnzcbRCP9UxkV3zUp3u0dDs66StGHT3LgXcLfL+4+kclnDOlnQ9UMTDKGCDIe
OxZhb3eh/k7GYxsar3XWGqUQWFnNesxtCvbEcljXePY0ibPxncNM3LjAacOp2tnBhYFoEsRiYUDl
TkPRIsPIKrDookqEWC1k1mmn4ubQO7MFIkr64USn8l0Mupz6KVA7n8G0lQQfihOt7rOvrTPwgxUf
UYjwG0H4YXq3I9b9lTbvow9aYBSl+hrnD5R/3ai8t6/Smex3qfDERBkjIPJy9QK9+faENhvqNJpQ
RMV8v5/qcoHDV7RuzRVVedX26pyK1U0fX1YK8r6SSHbmo52ahw7RHhTunEDDgidGSvF1oAih7zzm
sIMBB6wj0jTEu3pkWrf2WTFbP8Wkw9WhcjVd2np1+8zORWWHtL+GWIZ8K69BYChisAw6QrzxDZfZ
PrRv0p6kf+9hHYgMDUdncyt0iGtAFqUo/3XVGIoiHrWwT3RRwJTvio37IlScpC4jILqpaU4DKyOU
Oz+z1YS8BffOYfXlKIn4cBcGEHPlNYPJUwlBry9OgZ26UkLxvFs9NBnNFaQ5IIQoNpT9iOIVAj5L
s/JXXZezeoLfvKttCeltRwXzpQVkNwR+fQfm4CRAM1VcOOkiLOhNiYt9Ys+G5r1ht0YTwik/RlXc
RYO9QVed9ebvXkVuGpNxUnyLp2gbolSimrh4S2r8xdtua/5ZA+TNvF7chCIh16tpYbbNif9axDUf
qmn9YiNEkxNqGVbAzyOCSGrrbNyaSbxtQBNnPkq2/yh1M04Wyns6KPHzUUw3Jy5yGtTxIeZoPZd8
8lw/0421ezL9I2jEZ3d+TBsYgcQ2vAipUOFZD7mQuScics/+VrbCF1PfciNIEtS7JO8asJXIqbYw
UrfnakpJDyXhFrU3/GB5yR8KJWhtbaFOgLR9XbqfSeNkwWKdSU7Fp0pHYzsaIUWlLDUjt13kTs1a
BW5gCgZVmuJX50dYKnmJkR5K8qzBAXsfDuMDGgWH7czRl4TdGPVPvx9uUeKwfn3l5q1kEfd7WLTj
Deer1WD0CVUK1H9IExzjoGEq7bQtm4hjvHl0phvbF27S9hJ1xV3Z3HHtQVxmy6nxJ+3uGOnDAdDj
p500useWCH69lbPY7U/fEFsPf97Q95Boe4hjL0hghvfU0pzD//o9vn/9vRTawDSO0miyIf1WeGIq
nSWM1F9EtOMCJtOa0gus5hEWOmyT1ISsXUkhIi8VuXN60sIFpzqScTUsumyAIhEzPyorJLNvEGng
lbNRcfrhfE3NnHQ77gJZieF94b2KZQk+Ht70p2ZRoA1llVys2ihZcytWJD8ByASGi6eNfrZ+Wyx8
v5Mz3ZTsymDAuEciCG6PE3vH0+1FgFKzDP38sgyAIvT0zszpsqFWUlwM3AkYkUMlJwyJqyo90uPm
/dafCgUjBbdqIfUYC6qoxWqj3dpJXEln6erXzoJJlds/wIupTOFZ6wxQy7v5vXoPcD+RRnrRdclV
h9vpsqgFTfAfFgA0Vl7B4Ax8n//dhqyL54Vy4f5EqaJNXRtLayhe4pUyu4kuf0FntleLdk4tz6Ga
ER2xWTrxfeUNz6kVbfg5KRA6rsbKiP4SC0vP0doOVjDUEeoVODRyqf/vzFZL+VeAhdRoXugKmoO0
shs7slZkcAp4hDbg5CyQPcbG8jt9wrBPbLRVFtWN5UDvGC9pIAN2h1tLvsCV7yYn6MfeRhRJPGG1
y+DNcjcf4MTS6xmy/SGmJbY1ujQMC036ouFTiaIpmkiMUIYqd8CXjpp9DOjgDBuRfroLVk6ymkem
DswLY+GYWVTh7ASyScLGa4g7sURGyphvMDOMF8XguMqMxJTp5vGCOzk7Fr6TLFXT6S/NdAi/1yVZ
ISx1lWRykjRGwwvgXW1X/hLMIbpZauOJ+dFXKTqNAQcspio0NWze59W/P49+NRvLFHQJxIlpLRCH
V6Tmve01r4edO5LtABiHesBPoh2435zDqH3PMk89YZpX/CcDZ3HA0BBSWD/Q4JPgfZMLQKh81Zdi
CoBM5md+IcCNTuCQb60ftU2AZy/qgNrOWx30gpSSKCT3dH4sWXCP11ZsF0enp3hcrDMEULT3+b67
bvimc6fqxbOJ/b47i/qgoVxuFB+1GxAKEVMR6x5DLmkkBg03Ks3IqasR0UKa1YmR3oFzVUH0Hb0J
s1pmBpSuW6W91bsocnSK6d/F5fcl3G35IBZ+MrAgCFuPx9rjIR5uyZ+B1pU3BaUni6RuX4MrYsYn
KNCv6rOnnJNqaC+uvEJ/MCEsesnfAqcxmbIPsoc9gbzLxzNjhouCh34jIHkoLvJDb5YVojik0Efo
t3c/HZ7lWqbCKYVOJzc7w2BOIcSgFawzSXqWdAb8JkoD7FI8CTfMpTeRbb+H9QUjHUSKbyogbAyO
56WKyNx2F5oxV3fk5MSZooMtEoqrDUuVXHrTaX0mNkUPWZEtHREIBBUDUx6YVF6Gc63cbGEbiVQo
q7+W3VIpZUgrucEpHkrRkYChfueMdanJ3afK1JN60Hk4/TgQAFVBdy8jC+FlNPPJtiOPtFBuQggu
1yLkJz0Q8h9ONMQDlBc0cp8ccCVWdpQKUY3BUwErBhL+t/QD1vFnr+eWOu7b/gKeI1rKQIEKsNJq
DBfiZejynD9MjjlmvbMqYTSHX5L0+hxAiA8UhPMRqNDByRVwi5wWGD2IBGGc1rl9lvqp2VtUV3OH
5Ijm+S037qfGRQsY0fJiPJyvWFpFh9E9g3Y5XhI3vm4hcsavyFAR/PP//xDSfmntLwrISh8dWBYh
bQej5zUv+RFIg5wmhGd8D5564OPPwDY+YKdhpCUG/9vr9etA6LhlA+2V6nt9x+AD2uptrRlJaUsV
6GtLa78YoDybPpWQjhdquaBhXmdUd3ufCNuCLf5oe4QDzfL5wH7pfDlSG2eFohO6X34QvPREcYdy
D4B7mIASmipNBNLBgyG56y2S0TY4kYWYtElUSEY/yl6ePJgghN7Z5YiMI+Z/pEcy2EEmsRTl96u3
/tRa5ajAMuh3C/3SXOL9TBhhuEaZIuyuDVj32kWul6SIJQiuE3sjIHyJKSGWpaDXW3J/YS7XcR6b
g/bGUkPH+P77a/B8QMstTVtSjkWIziXQzapf78Lik/sIU8/re4Ytw1FGJt3UETM6K5aILtWH4mMi
OOhce83d6uVt66WoqXpFu0XN7kJK/x2uBTaoz5KXUL+U5YY9ABNP8m0L3Gr8kekBqB1SI9NMWWcd
fG3AZVtT3y9fWTAXsGu9lOeJdpTM/1KkDPJT6YXxVpZESN8in6GlrXRHyJnQNk8QW3bBLwCskrRv
aCqfkoJxx7SV/ZBniB+7t6S/e7Fr24tyAxf/yAAls2drAcE49g0q6C28KCG/+zPtTwdRtJn3hI5K
wcVox9hxSWTg/KcTFBb3Gdkmk5o66jijCPj1GrH73hb2mqYTzNgI+0YBeDux8Acr8unv9IUfm/Qd
gBVMcnLjkae7y/f/1QIetTyUtHfJ9Hwg4+MUphT2T3Ce//LVMguHFWq3CS64QAMwqTku31MuDJcp
IzbmYGZDNgKD7V+fJniTF3YeV+OhNeOTB+w9ripszcSwDOm+dGubs/YPe6NbN0eg3086tsgyqcJI
hBLSmS2lcZkowsxFDUjzAd33MVrrwDLmGDJVtyJRttWfi5/yxpEEzQXgAg++x6jMkB0xihtYsToU
a/2y1135b1Zo/FGn1fRAnOmdgRVAxYBtdFX52V0Vp7Ymh5Y7rzx7/0SwnNMAEE1K82bpfpIIi+iy
tf56YmDtz4pkGMQpP0Z8oY0vs1xhlPSokLL/Sm/r8sKjHJMHtNEcGVbmdfAzWHYyf6NxoGjd1M1h
xzzU5V51vrrqulnOShqxkEdd9UOZ3a8aa8r8xIWUeUMROPwUEgqiHKl/IIQ/bg3+g9BpqQqX2GNu
pE1y3DfPuBdzdrri+FsYeSzRZEiXd4AiJecFG+YQ6jBkMmnqTD53T2Q6lWvG0qHiIdwsJpB7IQBd
llFEbaAeConNXpSWHFgFnJ0h6zgYa1hx0kagFdqZJmUxWfpe2r5XtZO2eFfTkdx0e5IrReoWnfLT
189+92l7EmabH9/xxa3Mfv3vLb5eVxxU8DfiRrJv4BC1ye1hA5nU4W2Jt27SV1/70/94/P3I5825
+3h5wf9M0rvhzmO6dV053qMyV5qIGqAqSMfD0mtYi10zUwJ4LBpqrynTGCsn1+D1rU2zSBdq1a1C
+wTzT5JqKXXx5qixN9KqEwQBWsKhQsIOp0pRxk4XLXxFnHQpT/donMJzbHgVXfY9k7XEh92sQUiP
0HyBkyMbEKpx/lM3UOJJh8ZE2xgIl17GdBdd9lec7kY9hKnECBOJxptNuUv86rsc9tBIHo95syb7
941ac406oGUO8RE1EyLH6r1mYrWT/CPvLF/6GYakyQOdAODlJbzhGVwxH5m9r8BqmmrsYpFazaVN
GMC6GvzcRXkHv2o2KaqIYxLkwswBCqku/DKJtKXsN+xCpdnmTx+nDBn+nUzYNAJryBTszuC4uHwo
aOBIkGMGMDBKDw1XqBDJPoirYeg9BIBNdZfZHrSOKxj70FcjVvGGohflbK8K7hKkuRE4DyyDZh/n
fWbpUojzmWqKsNwGz3dauyyb/Xg+V9tkYKTlVUZfjdbFN540lBO7FeV1iZ2loehpYAxswsScUmDR
WUAv4VYp966nocNd9HIskwbi5IylwgMl/n2Ygn4JQQF0Co2jCcxLnPnPfrGORHqSuz9FQ9qOIrcF
vzXoXbQfdhSI4glxTmJEkmqLnzqhq7JUpZQkgoTMu37QgqdjrORk5dn+K2o8y8PkeMk7Fk2C4KHU
PxYuz3Mz7QzpouAIfwABJkE0CaRWMvCRtcbIwNJ/CGL1LKz3zU8orwL2VYdayXgS+YopQithryW9
j2pqa17rRZSP27Xh9lOb/yZIgKwQYKEvHnW6Ycr6zl6igvpoAL8K/BkBC4+d+jzDGvCA92eHhHxU
k/yMyRfO4ZNYYeV3n1fe2SbnhxZcico7NzD4ooxzyu3R4TCcTZIvjOi07K82WeENtXDolKTx+BuY
ZpuDNR452zqaaIqmTq9cenDG5oohMyFDs+tWEnYi1X+qkXRYbh7rLcUq9nO70fCxyxfK2d4KX3vX
7UHNRQAf5f3cpc1cDdms5FhZge2z/7uqUsgN8pqEesGYH4c6CU6OpXsiTkbTHtaeCi+tYUthmI5Z
VNO8QLG1HZWm/4rkxUYheoocwV/jOeTABeDCFydfDLyTPf/lNBMaH7VZ7XbqKPtNiYsmvv4pFlE+
xLwkSh2vvLPSLHbs1wN1beIxzBSm88XRLiku/qp+01CYlQYXSYQeT8sNyTduxUIXWjnLHE4/ZTjc
iBhsjZVbgLda99eLkVMbLBFIvOxQLtx9zZ4P7T++MsPCkYxC2dnhCWDsQMjtO/XgkJNMAHQ3GgD6
6F51WvTwu/TB89knAVlDkG8teA9CCT9E6nWofoBtVkEisqkBubz7KmwE7fm9MZt3EKN5ghkXpP+h
QA/khQMOZ+aK7WV7VI8+s53FJWk8RfVi+iAInOlzsULFtp1+GRvw9ZmbajC0w4EhPE7MiZU75AEO
bNZRUiAG790jlYjsfFieeSOe2Qa6kx+7VsggX2tb3pzZa0krS99VRM10nTo0Oa+mNfuiOGwIsUxd
MI3tx+Gx/jJvn3Ga6rECQbacKmVdnHhqhqfHA0lnN2SN646ApPXhM+gVMelzOdAzXnByTcHlNY/a
MgsSiUfMjUSHSi10J6w5RVkIDMJ30gyDUGlqBiqc1KVD+690D6gl/vIo3jMQ23uTBQ+/mHRGkpnH
K8gh9w71P/bbNiZSn6hvugPtIkIVkGBkTx5RMYMIfkfEhkljmEugoPLuZ5m/WU++ZzAJ0b56SHh8
7VfF+XyuQ6X6pLH7Nz4StAfup8H1ycNQA3plCJalKonUSMyIHSWo4l73fQkQ7pDFufR9X7e2mDq3
K2IDCAtPdpbhmvEHmNxPYPRKbXm/PHxZXfofXxIATKgesdzMq/nOehaidK6VNdfi/xcQbQJQ/Kgy
qGK4ofvLRFafmcoWay3vEN33B3fe5JVdtRCLuDqaHDB+WeUrwMs0mIJ/tqMmitn3z7EHnW6obB5A
u9Z51InT/KrorTgS7QaorCOeZrUlJrVyHb5lqhawlCYYIY++qPw6Ar24Ik7sO7yxrqwPBTu1cwab
JozxAtSo6pQUXEhJIxPwxv1v54bzQdGgIytVTB03PJ5bpu626Gr5tZGUNUpSSmMNNxrQvn34Ht46
2qtDCMXVDX2DZc00Xe/QpXrdfD8twWlTXezgRnYTfTRb/wMGnKjIDcsk19EDEEMhpIDCkxkXCyix
FOTgAMsdc/aK2WnV0uiKqXnFWFEoxNTfnAQEPWbNVFZWOm1eu8aE7/OAtwi8SMzqh6URcrcPzZJf
2NZbnNk3oGtzL20gX4BQasuea1pHH2MeCjbo22P8W9GO6h9x/gYJ60s1UhCt19hoSMhTVaw/rypq
Aa3ug3FFdriomelC3aFtTw8I76tbnRKXzoyH/83DEqIfBbAtkVzws5I9CIse1MBpApF8dmKzppK7
Y6b9DNVwDsggHVJu1WRDrCh16wIME62Bl/b5ufrcddcSCcobswJtY1CaNA9d2ZQwPm1ghTyUZYuA
Kbk4j2f+1D8We2h0is52xSjk/G7ELMLhnsjxy6ODDT4VQHV054zTfMvHbMHlyJO50fzazyXGwfh/
wE/LjJDT1/SDelfus3N3glUu/3LrQG+8jMjUKUUMFYzr6LXKMutAFVgdjYdp9ntvcKkAzOzv32/F
RzBWgtg7zdDuOnRWvceaJsVFgHwVWHVvKmvF1oGBjbAphKnWTUEJBUQzalne1UbBoqkx6JyNGASo
IetNbx9HHhvElfLBT/5R6z0dSmJFr/7gEDY55xw3n+5odI5+G6XQiWcUeybOTTXTHWICMKft8Efr
aoKfxVTldHaKE+9vSwjtnTMlhkg9cxLdsXljDOQym2khm4hDVOBu5VIc7nPOWpNrAOVm+TDtU3cv
k4N2A58xes9SLZZnx7y+qLv9KiBw2S/R8jjqDnW2bBmP20q6N+Z8/hSu89JJGcQPHdHCSohXVdVz
XV/YL456jfp3xOm9FSfl5AzI66DeGCN3lY5R9fAEfXmgbaUMw13UvdTkXdVo3Wtzy31BZDCv0GW1
/dQV343p6omGSid3dcam2j6Xv2xLmqiN4XxJLZ3ZjZ0/XOElhJIgITu+m0UQTJJ6FvuSegX5cCTg
27g1pComz/uXPG/DvtGn6rPFlroXVfNqkpXGirWrY4ZIVCn8zDLL2T26hrwTghTNU8McM1u3itx2
zEfNm5V3n1i3C7TSLrotbZBBJVtejXyUtudaf9DRpdVMbIbhpHbEzla0hglyjHlX8i6rWypuGiSv
C2SExEzXl4TZhKwNampdDysptj5/ajq8oSb6uY1Ifv0kG2F2Dkof/uYZ33//AR6RL35P4kfCD3wm
pVE2L+Czp1QIs0goutXOk0xeZZXbPyxzup0np0o4TjrIgL9p6up1569d0x+QtRIIjsp7VR1dFq9q
QkgZuMwXtc8bY3XPG8zoD/rKcQuqEJA2CSJ8JOyv3haiXBilmPvWeh5pJ8kd7/LlApWmm7fmskpC
Szla+9KyZWdiiMOJ3yhmp4vGOT1qSTvprv0ZWR/HRPlfi+4IiFs4IuUH3OZwGKNCuOlmsEGPT6rS
lGo04JIwP64j8kyFmmPeXu0ajxmyvAGNAuL6s+OcFd7nKy6a6MvHtlabxhbY9qo+wuVaRPS1D749
K/gRkmbhbGUJKcSzbggJeFrqmOyi0Hv7nWp/AR82uXcJjP4K4KnDwtM0SZrIEXrdJNLYZUR2qhD5
RM05h/bl/kH7SzbIV0V16qQo9b60Nc+NNqRrSt9aKMxkhyxbTL6QPeXdttLtEHHeS+UlThnZinTQ
lMwfa5b4l6njQwOjGOHJJnfKX7o1ERsRdTO6J3E1Pv7J30ooyft+1A6QunBMrA9UV8Ar/dqVyC99
XykOVOnBFeouhMOp62lC0/3b9B2UughSvUp1YmP0FKMpsAQBwE2pagLMzm9opNQ4trjRgx9YHX5Q
xEdYkwo3sdWLPgAsPIeJgjUOAN2wWtL0Zy+khHgc2q9LA0E1StE/cjDb1KFg5AZqojUxu59EQcM/
BnW5oHj6A6cYPOg0bVxuptjwBQkFqkccplde5ZaW4IfLGXZK2xxlC7WkjuqOlBV79KUx8jDsnuzE
O90+wGXv5oJVvv388UUrStkx8nZGigi+MSFen3xilBaBjT7j/R1XZiML5RylLpSTqxqQf5GRQNjD
FhbKetwwatpS/OIqfxwhN2eoLaykX4Tk+KEAVifHYg3QkXxw3puPVHham/AseP3cloRQnyQhSQyu
IH8Jd2VPmr5VeXWjzgy4Bca5SD151BiICvNmQ86s+N4QlyzFjgnYVc24kmJCKysC/Kfqp9bsqNMU
aS6+B+fTBMMBtQ6EJncYNNlm+HRKjViE2Yf8CW8q6dDu6C0Dbzk2UbcwEImzbOtAwDaBXa4ose9l
MJIWXwBhTNREwZtxhVC6RhsdLL1gD6JxA6fv34OL2F/h0cMS/6Bz8W3AQ8BJMwsIdBDpQyZkXdSV
ifqinN8WJuRSmNajJpNHmB5sc70U7o3AgZVwravmXekE6xtXAJaXhzcvMDlS7vZXogU+YxoxkRmd
XnLfLbALhITlLsOxwdzdwybcaoUcgaUFQAtaNpmA7ZSKAR91qBAX26PVKmH/bGMa3k2Bo2Lwh6zi
O818Ja32lIbCbaBrWMLZocby+TOb4huFcH0jSq41k5yTAHbcmbVwV0kQMSlb4pMfrbQTORlt/k0c
XXivBiCtPkiJ9JIw5VXuixtjwAmBbtzQ3EZ7lIaQzsbewy9IPNoYI4Gnxd2RhxpoJh4mXSi6QgGc
dyD3LeCuYbD8KA7wLEzYbavOgPTysvAyatHmwTxhVJjwVOpJomwcybG93LFd/xTqmdVvzUrrRg/8
0TRUdXaqzOsSUaIFBp2gD85VR1roh28CFe92QYRgJtxhrOWu7tBKegCqLaErLtR6xe5Y3cIyI3Wr
IVUXrWyAb27v5rVlccN6cbM22A7Gz/jMR/t+0NugHuJyYgPQdZckV9jUG7jZ2J209U2PiFKAU3IZ
+nYMemUEYOKle5anTJVSZoQ7pvtg2vt9hyBhs67gp0U9q9nJPUzv7RmAt0Yo/GQUcxog8jnuCkt2
9NHCVDMEaQjouy62DvHPEASEm09vIMTPUny/p2k4nnhElgHbyluv8TemjFdQWA7BtrHVmGYyKgbC
A0CMBEBlvwGpXzxEGp5+QkHjp7dNwdeh/vzF0PiFg+Vk7FU6YxOABpGKDysjZ5KaaDm+4U3+t7sS
eFO/PtyTKQvuvYscPWavnB9p5jKyyHsa7eZSYQFa3ap3wVWw7bu0y7P4/NGlpBZnTrIjvLhaffc8
cg+aAbC5DtNCSetJJn/gpAiOEWvnaaInLt/3OXW/L2cdAQsnSHxFVhmQKoNLEq7L+UXt4OKkyTnX
Rdh/IurDNEfvbEzuzOAchWOJc1jdpDvUz24TfpPLDhend7oGwoP3RRRmEi6ECs3xlICtuys0gFLS
nqLZyNyQLCDgvk7IAm3GoDiuBEqvDKcW9azhYNbiUih1vbPf9mg7ckJ4y4iHgaRvxPyyhuhPHuUi
ZbUSdvdhc/+TiENpJChpAL2Zf2u953G7d3o4qVKA4ifbB0SZDELBcoqJoBpeBEGPN15DUnAnHO3n
5oFmub+OONO5UGnmyn/zR73E8V3mboTxKn8eYl+Hd17CCqzLGYoritTLn4dzTnYVwyAxKo2Rc1BH
vKDadP4m03LCEGVOZJ+M/OngZNQ9LG86ryTQgOyuluzernhFpiYwKdG2AVw08++5rWcRLZq/YrO8
D4nDl58PtA8v8H2u9IQncP3TO3nfdIwGYXwykYRQknx6u3GS2fun8Cx67F1NjkxPhosOiUC6iX0m
j3+M+uEQwABTBg0TpT3nTLCBdgdvYKxVku5/g2YmTgq5OBnc190H7BteWQ6Fq/XUHQzQOLAPFzJf
LrmX2zICm8Kv1FLmKbT/KhRciJVUJkQ21CmPCaFUiv9do2SOKoyipDLaQFY3mnpwnERLBPiCsaXQ
RTA9i6hhmFyAsTrAaPQDXMhlQlPeygJY2ab2txQqDCwIKSLMg8TbJt4Or6sU/K9hx6S+B32pvZlz
cvE6VmR1wGj67DPjXTvehipPx+IdNe0y7nyPEdLLXXO1eN7gSpUeK1nT0XXtqjcvt8rAVgLMGoCM
4OtvEprY51yRwBzsTfASO4LpvctL9dsVqELk/cl92BLQEkivc3CXVjMn9kdgWMoju1Xhgo3SULRm
zxZRrxvGV7rwTndmXm3uoZtVbWfVRhOoW/8g/fFtbAeDbmrxIOWPRoN7yqWcQ+tToDIYCM+SI+rJ
Af986//OY/Fx7vjRXsoki9RnLh8kjxOYuHU5Xxni8REDQ/0a/cWqjqwk8pIV5roUaN7cwd+gBAZU
S0njrDqxxZuhZ44lKBgE4JxOwAa4uadNjDW2CBPIbPl99SSWzbvQ6BXvkDE58w34qEhdS5lzbOZ2
/cqS+MDDoTl7PNOzC2hueM+pXhi0rFj/XmVMg/eel+TXldGNva68sI2zgnSwdr+u95inDtGMXyX4
dLrrMehBmAvd5AwYsOBAmpnkCSSs1CGFUSuDy93sLNV+M8hmA76ooqyB4Lx/hnv8tvMHPNKHssXo
3ReEcjwGWAv8fqeftCY4By3MSv5PWsNXz18mLwD+abDpZZ0luXLODVstQ7j1woyY2OBDABlyd5EN
2iBhMD/+clJARCoAtplLrW3x/9MfXOOOnWrHySgQQn1n1w75ISC/1ZaUDQxzPqfXKfKE2lSQWnV4
EKf0tCdRl3Jab5nb8Fltqdd0dOa7N3LKB4mJpWvd7xQ8nDQVdl5QHmn3rf0ZPcUbYiUilDG69JuX
jROWj9TDwHpO4TttTF1R1iDcCPikOloSGiZJlgvGmBj/QhLSKujbMt/m4r2QB1rmLNTD4MeR3oIQ
J/gQtYcMx4EL/2JV99eXH54URoADaJ+OM4y8QwcrtFjayNrGEw+3Z4BM+yT5NnZ2fcZWgsBIxDyH
YOocU9lIqfGZhNhtXpqc5kuWaRqgEYJ9CVxpRfNc+aVLTdCrUMOe4k3veiGk4YU1Ab6FDW5v+QXS
IPer8SOveKwMVPYcITW4sk5NbbV3tKYyuj8H9kmXM/WXUiDxQzYB2GVJy1f12MjZyicd56LUdGZS
Lh4XY9Nz/GB1xIhRX6kwyU65Sgfk+ud7t28YnKfWMUpY5A1WX+M/gv9/9BeDJmHG4dS0SqIbwaa/
6BQEMWVRwc8ZTJjBoDHymKm6FZFDYAqIfpP/FT/rN2ybGToGNbI8DfIIN1Zz/58Dc0r5SzXBO6TA
4FTeKpBEdwdX5uCBlVYiWNojawD/RJfpkF7KgFk3jlxH7JMVgOAz0ZL3VKfeqkwLZTyfSy0zhApk
DgkSzihFL9bijxrcw2BgUhZrdfIRIe8m+SIGYphgTcnqIrbELQlUtgEbMnCaBfUjA6lVUy1VHLKR
ponRu1r3TlcE6feGLiUw3f96ApqrQH9uDrbdygmfL+WdYwYT9nKZNOkFkEPfST3cC50RH3wozBrV
xz/P/Szj1mEOdE+BYhp0iZGi+6OnNO74Z4BQlavjbBj6chMGL57BVwDvNmg4hJt1qgh6Ba5mEoCH
5Ac8VaVCTGyyLD1vuSiK9j0Ag0Yn8DVVUQLiSBBY4ri20cEvHtbPIuDythIsAbrEabmFd9JBjdjr
UGEtoc/ItdgmnTzSo5T4s8hIj44yyaKMay0tdbgCiF7KeNDRIe+WRamn79xfNH8z1Yhd6Q5gybCZ
X9Y9QPmGtXTSDvRKCz0mzPl7XBxfziTAqo/dbwC9S071Wn/xUlDj0HmvuKXWTi+TdnGrhT9TUaSn
F9WaICpnVdhcwlj3r1ARa16JxIRgesOa1c21k5LmCehERJV6YitCO4S7SPyzToAZD7OjtP+jESeM
bW9loeYi4FvTY7xJBQ0M6c7j3zv9HjSmMr0yzLJ8H9DJYBtIG9CiNJI2tQdJolvSqHcEb5vE2Tsd
U/UVQ290yAm4paB9Vifpk4KIDmzpg9RjnwwuOWYZVAfOTVj1GPKlKIxDYiRu4vxRaO11yHAgOR12
uPfTe5B0XCQsqzXYzKyLSRTDlfqXR3Zj7aEzg5+aVNQczk25D6380FBTo5L0NJ++INfqO0TpxSKQ
Iag0hLlnECubi7IZM5KQ0Q9PdBjtISCae3bmPouVe0Ss2mUmcBSdguuReLaZhTv+GNdjMd8cb34m
PzQfaLThZLzq9BAGqg6YdJ1Aj2wHiT0ct0XnKYT/kmZEjPIWqSrdRmRBBLWK3kxV+neCHYNjsPQE
fCfKDi8DNp0I+1uFNntGRZwfCUf6GBe3orM5DPxbF1RWaoJ7RBjon+pzJM8meM8W9FthQg7mlUr6
9f1OA2E3O/ykuK6XsRIW1R8VSd23Pg0k7fpe5spJ8rW2CRkhKdaWrBVDP+ICYrJ66KJjRokxVCh7
sw9hMcsiqPf3Y6/yp6mQztv/b5YK9JzhYAZT8yOjlGavk5w8GSSMuCOphbr6Uf+8V0gEHWkg7GId
AVufMCvqRBWxuQbDPWwBPOtSs95pk7eJsqIenvqiK9fn9AtHNwX1qXJy+ZaPiK2PGxjbF96MRCb9
y9J5B/DP12+orT1N4G026BUyPXHWSY+fr+BwH2BNJycpmktJx6Exi8lCI+rYK7wjpji7MqbYUv+p
dqODxuIaJ29o08O1nmGFcZNkC9I9Qg30oxHBXpU93VIa5e6MhSykDjBrj5h+TL+alSH9hjK6c3lv
0IOsFNBbd6PrVuzRmdc8v5SYYRAz+YpLOwCPejLS12gFerUJK2FoWQgEnnK9fc0PIL+44Rhwz2MO
uyNbODPSuI8JmaSGqxNiSeli/oNVVIiu8F5zCsq/d78lf74fQ+P4Gk5bnufjBOoI/cVy3fPceV/Y
d0gQnns0GNm3oe/smJY16R4kMrt0JgSvHIIjcn/ohJyxOpWJVGXp1c/jXJJU+Vea7Ho0HuwPYUPL
/Y2W4W+Hf1IMolVO8FZjlwc3ANkB8oKemFgxsh7s533lSa24LAbcofqexRdIpWuBW0PsyWszaf95
GaKWy8ygxz3LkLk1qw4EDXCL4mVZFHFaTw11g+KqhEBZydkd6lP7y+783x228WNjHLtK2cdt8wkc
vPIBwvTCM9OzbgEntoqtgfsB5J07na1sS70+tNTE3/sg6RVo0En03GOcgs0185b5upbf+VbQjnkX
o5DnqxzX9UiGiGp1x5eocYh3wGMjkQMZIsgQ7S5ymBozWpTbS8Fr4U8qbpu+xb56kkNzLwqgFvfE
gO/1ellDGv/KmSwr+Rpes04+6M/N7JShvCy+WXJXPu1tAbahP+wHzxn+YpkKnvsXdA31DbCGLOkR
jfy7OCh81+XSjGMjgV9tcdG4aKGKkfyEdID/anML5YKnuKcH08PrmiqF/Ovt8WJQxU5pz2rbpAWM
GIC1T51czdXIhlSh7yEdS6aYCybN/oD78+iradAlnk113wB8LTpVi5zkTycZuzbhWgCNhBj67FrR
IuX1hEI+j+CKDmh/MYrMbqxJxb4UlP7jbM3o/6I+yKa6wiw8oORyRkTjMpjveMAW2JSnDUeWxhSP
Y7A5Yckn9OrOk3qvB7EHoW2IXz/oXDTaETXXKEWeawhTwdhVtRI0zJ+kmHKMTairgW2wHn+S3nWJ
4cwjQgvLyZq6V+dmGEc0GNWjhuAaX9VnjneJdQQducNGtSpenAzojlEv/oIEdVrxPONOIzL23gbg
5N5vbe/w/ZoOx1VRXL7xR1Y3slLtnAFgxl8rn9SrJa0MLHSXF1BMKckqE5Y+w8xTA+JaQ7cKiR6a
/08Gz1KFczsSu2hryuHijnnO1/U0B4Nwn05o1lOxU3oSje+rQoO+pu6Pu7f9qMtqrPDHrHBT1CtI
zSXuJYBL0lYYxb1U+bQbIhfnnZG5lsp53vrdSvWfiYFQyvcVixFprZAN58JNmyVA9AZzxRfk+Uxg
tlObG2NNFAZ4XMzz280prXxphZ8f9aAu1RSnC+2O0TLIhhi04cTakuGcqGXS9eGLUy+DZA3AQJIz
ghx/IlqRv4szpx64/aqWatKkqpe9SZnS5bASjPqJwgF/bEnWve5Em5qkhAGdB0P+Zr67T5Xa4HP+
DuquK9fmPzCN/PLpxtDiWDL+VFHzm+geqntPL73xbrPlSJhJD+p8oFOuakMRibilulK/j72KGRwD
WOsF/Fgup/Gx0fg7EI2kuXWD1r/AUTQ2UJhLkponr/9I0CHf9SJjjN2rznqoYWbZVxdJWnD3RxuJ
FEJNLGjPGP5MLBsnijT4LZthPIEzxilDOPqgbHzJYltu4uGTvwxUgwQ70x2FvFP4nG7dYQ476Ga7
2KbcrPBOZv+xsZYZtuYCETv1FrCfXkPFgCg+8DHcyjWr9lDKH+DUSrnc11w2dM9hkYUDMx/OtJ3Z
r6H0tLS9kDoknPMi5BDd/SWTKGgKsTMC+fj6ZYN4+nC3wQrGPMeQpeMpFzlXixkOF17L26KQpyCv
bqLoNS6RiPF5d8K3hhf4m39Zzv/oUwDvJaTpln+mjVem5ImoHrrmycD5bi9TiSy5BJc9pKyMZb8x
EXwNGphoAkEjH0B+6Pi3XUQSNtkbfdpBhDfvYa5SJ6bPKlAithlK6r++MTDxerDPrfIGMXCx42YU
lnbxad+boehBTlkOsy79YgX6vw1LspVQnguEAQ5HTJHoIJKL36MSD3ZZJ5bS6+6SbBSHSFeD/2fB
2mTG1eqSNtX7gi5cWfjf+uzLv/7IKhdTkUMJT8zGGeqX7hq9WlpN3eXm+WD1/RKiLxk/HgmpV6CJ
lInA5G4WOJYNkWVgPwUJ/DwNKfk336p3d2ENmIoq9VrxzCuu3xfqFhgvzjU1yurjnsCB0AHHO3JM
T0a+5t0NtYAisOQDA2FdbeRlZZpYUpTQKpXdwQqYJ/6EUgHPKgy0a3FJQwKZsxzOovHoEEWapACQ
IevVxxQI0MyhUspAFoZdw+8rM6591f2JiUxlJdzpmHFvwsMnBxgchx3ICa4zumF/L3eAbdOvkag2
NPXPGrWR+HKBlO8IKRs4Iy1mqBqgs2ltLaNifJ96rJRVFxQn9kmQ9wIyt411MxQ2NTpDShak4aQO
nrDBimqf14ZdMmP8UNcXx2/V0OCnjB2FrVv14PjOoh1gqvKT6POIxccnPirP8H3bVWE9m4kpXdpy
Uf8DPcaTT+LFsAenBt5ozHkMOL3lmbxDnvgcmv8/YRCENJvo8xXPd7O5+FQ5uzTZBEmnWEEod0SZ
1HW/PVc9NAudRxgKGCCHU25+XHRsCUnSu2G1CU+/tjcm+zthHbvhijGXM/b0x/V1c87GMI1MpcpO
U5Tf7UT5gzRUmPsJjU9/GTZVw/lqtm7r6X3ngC0Q9sIBecPEJJhkCh1H7A2+VShqYByC2hTe/3Rm
lj4VYbhqfbn1kJSx+MAy76H3Me2KsLuNtdSsiF19Phil+jYI638coDokJgxGCco/vAZ8NgsYwyEU
hZPeLVDAeNSXZYKWHSKJ/pgyZMuL0p5Atlu3EQngK+yyaZB/yArOyYNFnGv7lcHJG07ww34bWXqf
WmJGQAfdJpelHVd+rTn2F/IfTXr3hYrctQXCSCDc/yWmsaDJAbnD9zRPmqOVNIyR5dWxom2KmxcX
NV395fmi5aXmuArmlwh8z5UTYddNM8K4g/neZgQiSEpPurxjZTyZjK56tNqrOE6L/yNXzyc7Xpru
PYXQXi8MZU58jS1Xv4RuwHgCRLQO1qsnvuH3TOBsz4jbYLq1wvIMPhV+t70nUjum9xcXDh7TY5qd
FueY9ekGlapmeH5olfwz66i7EchGARz16xa4ZVuiRRdPKj1hw7IesQzIW5YOxyZbmXfv5G2HGv0U
WITIjWpaLxniRmwiszu8pDtyVaIP6huyUd7IrM3ucjfeBKGUXIKvebE/OzByvAJPjSPAwwHUMZP9
pfpP4RxsqFhis+NP82FWvioO+NWzgMOtqs8j/vS6vfAO/dKvIueFZDQ8/maKxTVkRRh832cRqUvs
eaZoIhdGGpaRwZo0YuE/SFMSWKTWMRFGqHJ+YnuXbPjNnFZySbXuAgiI8pW2HJ1gOfq3sCaA2y5j
Y4an7ciKxNxVGYMgBj2tUHM19B4vJXhdhfC2FZsQdlooAbHdBn+B14z0knzFn5MucQoh/jdaQsZP
6WFBC8xKgWWE7OB+wbEPNAH9wkBs7vtF4q2Y9t1PVHTef5iK/viXFJpDED1arGobx1EWVARKFVGF
/ETMhYq3+Tdb7EFKUMErQ9DopBb62GIxQvJXhMQdoAnYJTLf4mgv+zDyfsaq0aWbJqYM8aWlK1sl
QawOMzqHuiAdbgWuYq2jP9lmWyN3LCR1kWQ+l/H9tsLE8zPyeTPia4n6lo5RleuR/o9TScJUfb8M
sIFuYPIXw3p7hNm2IwhZUfleXttN29UtmAYD4pFCpDjrj6aIO0nfBCW7GscjvUcA6I0k0fNXRzzG
X82mNDlTZSZKiTAuhtIW5dRc2jBYAEJY/DvnHkKvUnerRbS/rdpZzNpviynw65q9H1z4MCYllxKu
Zrtli7+9dBBkAMiNG6/ucajOqhsPt79OCKlXgBX3VEWwdArXxUAesE03YUIRlCSeqMThUKe/1cLO
CCAJvUDLmwreHHVLWrEy12ed/vzi+qXaT0tdQMVgDu4r8b8pPt+UCt1fxP+UkHlD9HXQIqkVPK54
J0/OIVE1ilK8SY15/TDPPVPtf91CXiJ0HBoCdM6OGVXUljxqHb9ziqVcehz7t8qV6COpEE4mtt+I
2YUxE5a7zBiZtQe0l/9uZzymah1hGUhVDmzA8VJMRT3cftQNt3ekNLP+ka3Vl+x10MjIrqz0hYrV
RlG5mqcQSbfyCGj/bkYY+CwdjSyzHOvAccrIZEvm6LMVOXW2uXWa0CuOe2PoZAZLQV8ikt/U49bg
1sBM41G/HI53mphDk7vBGHZurGzb5Xt4sRyhFeVo4K5hf8/j6Sp1oENgbKAW7mhGlRAhqVE3sIm0
MA3F+quvZBqQe/ipT3FEPZNy75jjNlGr20ftBGMuf0+sa0OEIdwjr8QMIedSSM3w27nH7A4vPQC6
MKtrdwDTLV2ExYY98o+a8LfK0H4YWB/4SHtticW9C78XyEDXMpUJE9uW4iVphQrKYeadUmJnTcdD
G/Ik89XDMINO/nQJ/59ihX2m/BZ3reCGNAfPy7/JcCNGNv6AExmm6jvrLrD3fk03rfxFL2MrT35s
XwiPIAYB+A6MJRo58eXioJ1B8LVuB1J79vq0dckqXIgfeh7Hucd5RL1edrWwe2ErCYGlxl2rVJtP
VdwZu5BQZK+sv9svOg5bBm+zu4Nbr6yp3m4nikuenR1UtMoqAJH6qe+zL52TsrxuH/YhsCwNTuhI
KnFfGD0ZXOMrJv47WRzBmDFimYjIsf8rJIivjIHLJ6CaV/w/MjJM2NMFn1ASDwoxqPOFOnuF9l/2
N74VguL6dAfTJPNfCN2sTByVdUcKvcaj0JzQdjDQUgmCrPC3Pg8GksrBTy2wKsreeyBwRwd6ReBV
dup8DhoBNU8BYnqcsw0P3YroZVwSiffnE4VrS7LTgFBtkhOREgGaj2yFJDou9a7Mop0D+OApswPp
S/O1LTq0xrkUAm13vehyHtuYEZaSPB2cRKgCN2nBxGaBuPAJXf7xpV4ZRVmCl4nfOR6eHy2VAeZe
Y/XKfv0FksRmSYgzpKPRI/KCn2DHA6Pw8vjA3Vjk+gQcV6sB0/yNxVaiBwvlGzeraN5PPXVWFda9
hQW/L6c4LQCbewWsFMmpY/AtYCBsm/OCDI1I8Pf+5KFaoKM4E5QhTnTxZHDkW6YdLWEWUKaGixKW
o8m0hmTvVkrb9mZKjC0Yionmv2Kv2epd3+iLsuBw0RBdQuvd1wnv4wk2kfQOsYV2+UBDkS/7liNT
2/1OboF0qicM/HfFaLDOyhPsffafII62nI8tBYcFHYMf7MUEL6rpErmONe9sDX38TXDOV+aiZiIQ
3pGiF7meMuoFRU6eIyYDAxRxTuaNa2MKNPId/7cWcwCtdB0dFliFYAek5SFt7n5+w7jFo6sZbLSu
jsdJtnGEOWl3mM90q+TJgnYdYXe5RFjzzm0UOSMhCCIRhIEOaahfiRAhZwJKN8Nw/A3St6crbRaj
RnjWxfxuyeTlEiMyf8G0mbqknvrUc+fxf9nWAV0fYakL+cOxWY3FKh61q8feDUaTrB1ZMBaxoWIF
kUsdYsYed/30TZEUs2mrvSRozGkbpmjzWNTbcBE6NLctDz9vn/88fwSayvBf2sDMlO0U07hWjN6J
klbS8YbbwylRLX1hm/1IofWIqIE1XARQGf01hzY/gnWz9pcclc8NDWxTUDFUnqH8X21zsnNA4Zbk
yEbNjiocCRAReczLis1IM8O55Y1e6yrb/2lmSxt+33S639uvVZZRx6bMY6Ig29JeWqvqhtBzgMAS
SN0Qu7xMFn9+z4MORnNyWs2D7rae9KE4Qwjr96ZpYRf4jJYB9+qB0pmaWV7v3qgUbaB6a4VvB5+K
O+DZDuo4SHeIkfzGVcumrdMu4mbup0T6b3lN8ieKkkOFee0SxJzXY+zdhGEDyHa/+zXa6ifVWYBk
HMvcmTRyr7oPk6oE+0pm3fumUJ833sjchgdc6ZBWx6Pq75tMqBeLTGBWJG/doX+8vrrjIngSwAKJ
3C7Jxjtpi74Vb2cphDzM58jaKeJt63fj/hXXVjK2J8HyutHY1fkg7PQyP4Lj2XqFPXwzlWCo27E5
pUvcUZwlzO8FsVOeLFbfYqYDzO0CtsFH11QZ2KN3tgw4XMzoqBG+MVDKJYrnNfkZd1WFXYYjQb0n
+9APxmI//2YXn6+bUCI7C9kT/sjNN31NsMlvHup4+MXiZk5pgb+rTIum3ri/uBlJXdnmS/H67ZOg
VomQ6tHzHhUzLikaLTic3SyDWvKjthhEtOpL8A890YLqlXtQJFs8EGPD6ZSnq6GtLgL1fX+SyjSl
BSRjGPv4IGchih0IQFvXJq3eeuXu6oHN6Vr7hEsRHed/ZsEkyXV9VxAHmpkkvq53AGX5hxK+0uLi
MJZ23Xoo3ZJX3NYsq1oEjs/0/FvhHw0sTMWMLgBEVHMVUh1B0ZIEQYugPtkbYJUDS3dZMl860vLt
cKvLhd0ZSAW0URB0nUr0yd57GOx35Hwc2tbMtNNrN3FO2kr4xtWh4zjD+R8iyQuXuNrtxHaFFcUj
6HwMC47dQoMUCwbzFOR63sLJ7yj4an/NY9XeOEkjrvS/Kep7M8hlQ2rh2EqU+6YgnJT+pHb/qCt3
YUxYAJHSPWxfAGErhRQSHOGCYRk8g9WxWC8gWECK6wOHts2yAZ+SrllJNJM+DhhLzkTV/dkButJK
WGjaaWmJ1mGcafi0XIDciw1XDUXrfTD/C6TUud0yNV4vS/j7gzynMJCi+AbQSNa/Vq5tThH8zI4m
timSSvKtnNeazzbQMOIKGPgQxSOlpw/iRwCwkEsqJGZcm4oJxeHeL2hjpTTgODGTtNTZJZu0gRRd
pcxOtM5VrLk1RQeQHa9sOkVGqjOIbQMdsWSzAB0Xt3zGORQZJBeaSszCX4ggl8G9tmzMvbtHhGwa
+6npSerJVgBjkHqnol010fPqzcgbhQ2OnJ4dyi36bir5QOCFH5ar5LtCSSqDqtAuIMBjJCzM6iB4
9RRUOD7xdp1iHPvRRAexknxvFnJgPs+WOWts9abde15RdpmtcAC5OTkNIppQ19ShQTHi7Pn2QXrA
XQipHthyehhtCZWNOW/5lyaxpJpcKiEK+A34fLdjBSwExNSO/+KoXbnMET+z9Tsi17BbL4CoSiNm
k866lx7ni1Mn4gPbBBrbgqG59dSRJ8p0YHAFWP/6S16V9HZnA77eq1r1U0L1e2bWKqXxlBQylfeJ
IxyUe4JHyIgyo4sd8o9dfpEUsmzskAAawpCv4ocAZis1iTGxCwWsJIos7tAqdAh74Nflltpm3kSp
bb4JHNkj7DzXW4UF4wLR8g8q0owf/NILnpscUOE+doatVc3VG7KfN7+YwY1+YX85OogyI2a7ULlO
jQ8pdYGgniv/kW9qSbOBoIIYycM39R525Tvu11XaAhlVDeLxrQKCzfMDdx0dxPyunLCkvJ5W3rls
y7foX8ylyUajEYQzRpQ15LjUPLV/ZP9Rh1wyqir1zyoNb1S3olDasqFBbl6YcvvJD5nL6FjWWPKS
7mU4knAo4pIGu+VUXlYQlVcKj3ak2+MNvwPgnRjetIMZp/Omi63iKTbwE/P54UACCvIDztRl7/Tw
hUw/bh0GhW4A3USGRJi7uQSFP7NNQhGUQbWzNwVN3q2oJoW14vvORD/R9JM0eA7SmhwGbxYRRib9
LRHPF9d75wxDE9Voq/FpuiUH7x8eGZOhKTxAi2h9ULSoQ2B0mH1bLwUbMXbKQ0+sXZ8QsmoFsKrz
WoKUboPhExNDdgoJiNSRNOYvfl60XWE+YxDSgpPt5TL8gDXjZXMg7JaL+t9PmwRqS+3UVNUcYS3G
1EDsGmB4mUF9mhBjIbX18U1jbAWFmEUYhY8Mt/hXxxh3k36rANUc/+ZRJ+YCK4KR2FuT5X3Poh8/
aj61K1XuzNHuB0QvjKKcIvO/WBHBK45srNvxu8JfPH2ORjeWmDhCQ9HNWAml3mhe5V14SMUaxm6O
WRjBe3ka5xvRfbIltbbkWBv3lT3LrBvfCu3jtzhDfGoDQM6cpt7WmDqGd4Ej+mCgo57hqvbLh0NE
qttpVcbnWjWoKvDoQpdSqmwXtpmkuHT6+yUh2NMLUYHldEOhkxfFhPf2p6H1AT6rYi0mX9rOnL11
4419o2Qb0qTd1tGVyjeDY8mv8Ot8id75S4PuBgN15Sbdo+hcBCtCTSb/Aw4vnqvuo5BPohIGkQL4
EnOH+021+Y8eUIJmpKD21dj93P7dbFcKNymqOj9wEDThf4VC477C1Rl9+OIVjfd5S/u/hC2eB6lX
mDbHWjdzWLk3y9nxtPWDRFsTsk34f7TQehD9twDUNsm1Er07Qqu935vJ6m4YZxLkgh2fFYP/T658
C/ShkHhPruncYuB/Jt59bhn0xpPSWESnmCK8darYcbm9L7jTIIs6fOQDiKGj2m/PFbHWVyzcTnuU
roYwGwE1nq6fMIMqo/07G3R3gqO2Gline6JNObiHpOEEgEXEfFvA3Lf2i7hJVMK2sDVMswDwQ1em
gu5RU+SCrAgHHb2zuZLLYZHsEbmPuwCwD4ZsfwyuNP0GsFzcn5vVBB/K+t8wWhOhCIRQV6twilqm
caaiib9PWih7mn5ltrlbDXWSxHhHgqjNIRWt8SWRHQ2P0HOX6SvLHLhd1VjncDUewTZNk9rtM2Hm
SAr4+4m2dygRuvYv3qa5y4b/41+BKQpoNGTGbYYJKBHn/+Ivzje9FujtTXRcyQubncGogk0CelGG
GGm/tPSJdbwc8EZuvtHQ1K4fynyg85JCudZsYA1FF7VwwzMo4yWPasbaDxNxJ6oj6jVH5jXc6iCF
5lV/ZlvK/HY6W9O1uJjI6Oc8MXMg3TQQ2SDVWvfmvTI2+ddYwA6rW4QwRbP4b60ALzGjLD1C9lB9
WKIhB/PWhubxMkypUI82Ig7GoRc0J0YJ90uLa59ijkMQ1wds59cgsJuCQ6lETNXQpG+IoTKVJzRy
A+3j3CCVyW8nwTpwXh1D2NK0r70R5njcah5C3haC9wM273YFwxTpcgzDb3YcYirSYtliEerwLWxV
0BkR1AmXMQrVHWxtEhIT12F8uezuWnYt9xHY9/qTlJgCRk9IPk47PibUvM84EL0jDJX5wO/kIZIR
ZDhhKMHwD4P5lGSLS5AUpg7e1SnkF7lbq2RWR4WT391/ch9YAPeiebOruB4jxhwWto5dncu2On6a
ikym77WgdCM2lwr4chseDNylDOJ6Hf4f/56CW55P8fTeFho3HsLcvVTB5KDEtaDjcNoBYPYJRHrO
gKjoo7NG6CseAKoCkCutV/Fhhv6Rzq3mtNCcmZqM2YzWlgl3zazc9N/AVtpYjZ+2yxrew7OugRIw
ztJ4MbSIex6sbmbO8+pz7VRgPSImQbvMSnW9RtwqvhuZzLIeQXZ5StCXMr2I0Fkf8GnQmKSHZHnS
/y2RWZMDNQ3zMfWT2Res1g0w7pnGNUhgi6CMf4mGNYzgffoZTrN8d9okpSSXIbIhYGkyrGz9T5Yg
91uD1Z/7ZQfCdH+0IU1wCJSeJvT/KGJvSesEn+iR5/gVHhDNBduNCOGglLlHa46SXsjHH8q0NvFK
3UEDexwAjb/+eiueTjYFIdmZOa8YWXZfx91Tru5wcrvq6KqO7Bl45t6pGAX2NzFY3snVInlRnVJe
RYoy6XjjNIhzOJ4gBl5zRhgKItgwc9p6sOoFNOXL6vzyp0tY38tV7IWmVJDROyjOR8NefGCYi2bq
QWhW1nwNhNcO/wSILhH9DQppq7sZzkJeFxsBzARYeKgMLJUJ4mtAwgR0jWRZ2ioDz2seykMSD4Dk
UcGVxhZhZePFIn4LECMVD1DjSsa8eU+3eIY+3QoCSBKch9JZ+OoKCKGgFsFA9/o7/W+hjycGjdtR
B/mnJpueieCPr4V/IcihwDsBqm+/h4k9f1EnyxLiOWjGjOvV7ffFDIZwFsoVGAk22FJLDTLVDFPg
CM1EAIqjsy3JXCicDQz85r13qlPSzr7cuPe1YwCAuq2cKu4bmLVPU9Ur9XfD3RAZ4RmYKKvvyqok
+ZDgJltQhGgFcATK8GWfinsnSeDte4GArTiOAXUR4ACO0kaYcRYjxbUSw3FY//zYdN1R075ZmUA/
UeqxzCAno7Tnfs4TCHp2IUoYKdBFglPT2JY2Bw51ytn48xKkAmdMY4CzKWg1WSCcPRhsr9UtmWWH
OcgSeIKg26vOhFhTgoj9O5ADz/Ll4aZEe5bxVEpGmXOjzIIFM1Ay8t8JG7GYBeEXAqaqG6gDuZJ4
dV3TPGk/cvL3vLgAE8SswX8ABRolA3tHgBGZz6kCghwBF/ESwA+t04qOAV1U+EKnrlX4gViytVl7
mBeaX5XlisGRRkI5rOzRnPhJsTJGQOv4GCtYqC7elTQ9rzzqt4KuipQzpAL2yD8Q8VDJEd4EByUp
cxUDwB0zZd4u8Qf554t/382kEd9PbxmYTn+VEI0M6tXx4UGxpTZhnId6SnRwfKbgCHhMJQ/BdNSA
6hJRa5peNtjRY22RT9kbHMKYtLNBjcj8Pb1HbpWmwqGjaJZZtZtPlwfZo937F7ycJ/Lsblj8Gp0x
cix9wkAFX8Lx8r0LNrgSUI5cVmt+kLaWmVM+H9/WJl4HJtOdEptO3Nl+QW7M5O9Sh7SGLbXJu0lw
s6GRRO4TOPvsekyyX7Gj8uXb2xa9oyytV1eABmK5Rda/zr5LMRXyjerbkUZITlVbLzj5FgyR/03N
O/bkuD0yx31xytngfRPFbexogZRJroQlLktfzFZYlnHtYCAT3vJjDTeevyboLTl4NEPgdI/lk9Kg
tQJ0UoBQkPaA5PJak7fxieW0Gvk8z/Y8Rql/Tic8zzpLjTzv0WNtfl+cLnTinxEv6zDJ4ywuJVr9
L7sjpHpCiVtOYAkUrhzqaE5cJB1RQB+LQCeYkN+RKPCkEDfM1EjS7Zz5nu4wsWDAC9gStW67lX3C
3/S6s7M/UMJ0+5tIRqAIdfzgleC+QYDVPHnhvv5BP9X3TdBltmPImO1BcHsSyvC7HadZxnKuDnLL
cleJsh0p1RJPXJOMHwwCcmdZi2VJSF1poVKAmH/ISOGBd93BiaDjrtKKXyaA2G5H4LVBJZoGYimS
sEX8vhYFlDqiSaFxCaQy/Iu9VvwLgXK2LefyFSN3Bw+vPZmYEYFtL1iRoVxrhwSJnHEAsQ3+arhg
ljTUq3J/z4hfJxqP/vZP6AkLXiVqfJH78N4TLxXcugtP2k5Hk6n7xRbvD2VR92syACyQwsOgtjMF
2EK3I+1BVqmcf+vl3NMVZWbUBuyND5mVP+7wpJAUnoy/oM8tzeOY1ujPGSDAUKAqBthO7DqWQs6t
UWWoxcakLNQ5G7HDnMhjLUGH2B/3Loc2CWT2ADRttbiZdhLLcG3Dphc9Hx0FyBEdA2QxdAbwWLM2
bDvXsZdojyxQ/cr+jh9IUZhY+DaED/FCg/dbtfpAv4qzszUL9y9AtTMXcxW2iR8DjKSYF2lO5oUa
6ftQ0Fvz21ngckXTWVxiUxwWoSlFBtvh0CYkPASieAY9uJU74IhBs1zptPvJ2g3VaQUGzvex7OIY
HSuhVyLw1fqRnTIN2OC+XXIKhIyGQM/YXvAnIlKkiTHlrzmBITkBrOgzLlElyFS6yDysdYSc/qXr
58aMQe5lW6pT69VEzwHJbUnqFSL/jopg/HZ6yjg6TS4fDveUYR6SB4eWTik128bQYiwTw9FZF51X
cSANpmTbQFrC8PqaOGmdt+NwKoUZPjcuTozOBlAFBFc2Qpr0vVXcJMOFvfw+Uq7vSqgDrL+dezg8
J1g1BMaaBbSCqETfbqJ3t/6+teLjVHZYoeKXGNaCL45GXlrKmuooPiaQkf3f0PbKKK8oVsL9beDo
YSbt1Q0UPgxP5m1bBGyf8OF9NyavQHvPNBCrCMjhEpVen/rj0IMQIJxR9YN9DIID8nXXEzZOI5r8
q6otG5+2VnTdxxV+kdRXONsU0/UuGGkeey7ghoGpOLqWjcxlOHP/lABdBXu4N1FU2V5jRdbVQszQ
6sKMi6LmG81qrbbXSwFeAo4fujMP7AGca8HjAqxc0YuQ6PhnruhDmSuSD5p8Ol78O2vhjFFA7So1
S7OpS3ieqZS3UXSW/bGdBQB1xvknDe4vL4mGFTH7hhLeE2XIp1WsZeAyUXImk+KZYu/j7BtTRxta
tRaDhoKP7f9MxS+NIZOSe0Vd9pduf+x0koxHzUc9aIyA5bhOjYQSMkCtBHa/7MX5a+QwNFcL3AH+
3MKGUo+aRJ+BE+i3jzcW0VEoADxaqqMl/S7ixo0TLjOaELX8OlRjPGv343xe9jTcfQuvaBO2FYup
NU6MstQc2cpDjDLZRh8NWYy1saR+h6A03jpLQ9k/KKq13LVeob8jp04GTPJtQhIsMttTerzjaBWT
999eEo69uSAxdE+JNCnCfGPechh+l7ayCzKNthhpWUkqr5QG6nYw7T7OYgQE/7ANB9j4/BmHdhDk
1Fgvrf2eWxob9/hi7Jcej9xxPlksBD9e+gju8svy0FKSJiXYCCfg94AqoFFolrtx8U7dWo0FzTeg
W3CnSWCiQMwsdiiScIcXUS33Y1azh4lVmao6KZ2V1wkgHsuMcoRPdWTQSnyMIPd16qCTxaWPr+9i
RRd+FQzMPqKLJ5QjyuYi87HMCsuLPgPPfkZ8r9265HUMpdY+jpa2UtesJ3/Eke20aPZc6QZq2xdL
vJGqvxLWP8mYpiEiKddkxK7H79Al5PvI+JdPEdQr9+LYF8SLiZOjvKO1HQZNx6G2vGc/pYNAa/su
qHQilzylFD5zEmLM41BTXOj5fzUQ7Mo1n32tZfyU/EUZ6Y/vxaz1x9Ls0t2DNG32Vw9fY/9cuvdk
AnrWzZRhbNurQchXR7lkSq3oTsq5AxVEiuhpf7idgYJh0EY2f/f4iikaRx2zVuBxNOWLAQnD29Bt
i/xh3PyNwalz2G14kAF47Rfj4hjpeF5yvRKTn58fkMaVIOlNYAmQPcE+hcwzaRoaV6UBvRrDoeUo
jvcmPdAGBzt8zXbsN2zuc5rbOQEl78zKoZ4NSORR/CKCP+ZFT52RwTIwRloV6D1x4zPnSVaOhqaU
NMKuWBARup9v+O/HKkc4lJtgucFjKjSB3Oq5Q3lr+UggMz0ZoQsm2S/3+GqWcNWmXLcO/FTs3/76
scO1Wls1CAXw6kQkvOfo9i9p5UiMgot35tJZRLlI+J/UJIcl3APKP4dM2BEEpR/7x1z9Hg3vR5Tf
JMHeuM4lZT6nWg+ihOPtcp/jy638ndqrcbt8l/VBXLVF+Cyy6LWRcPCoDjP0JSz6D87BELCE9hWp
BEmF3D/xdUMaJefQka/aTkRM6jej95VGA2iasrOHoVTjivMAyCQmoZdPT1sprR31bics072gUP60
MGvHCvcK1hGRO5UtJAmF4qBTfqjLZORWW1nWdUfcznM5+OEvjSgundHfo7PXpoB4e9nLtrqfMwIR
C6XYrceAHHIg83c2dzaSJNDIvSZnQM6LWUpbWwTPBqAfFZMRvnQ2WR2d9jbzxm3hBRF+/NcymBn3
UTFBv9p7zyC1MnLlD2LllybHVHEIRCsIs0IHkCjKVEO0Z4XviTHIWYGXOTJ4ZfMI0IhxzvTUKCZC
TyqmKetfYfTtl7DmJ0ACYJeQmSPrFBU2BPgZeOCPlZZ2rFSfBSxKenxGuE0sGgSZoHarW+FVtm/Z
Ix94BrQ3ov1mKjgM0PYuFoqFqfFDvzDu8DJXEIbfqGNlTlMYfsXmKYeTbbj/KVYYcAIHdVFufQeU
tLjz7+16QTokI/dWGvEL0JCZYuIRM66kIGnzS9T/cSIqrXAWLpAogQaG62h+IichkusHeOVQlEqI
QIQYEBPoOjFlNgSTPoyLi/BXEiwa0tvgsbr2n8eGNwYYIGizBOLm7tspyCS+AzHh5oJdMspEMqiK
4WKlWuT6B5240q4vB564RY0QxPQp+ja7Iljrbm73bryZo2Md6L1XjdZRmdsFZV1ieO6bcj2hM4IC
M07ecxxrLAmUPBPi1C3r/ppBWb/qdzNCIEkqq+k9OgXR56MEAxmf2HwJYSxA70AD8kCY8Dn7DTvb
/Atv7XglWPCxInUADfYNjhBm7/3juLCZQ2e3i3iAQ1L1yqFYEqUheJijgox7cuZpvE1GhJsOkxzM
jFbA/qjItSqsUiEFR4LAU9krULMW852pTaUlecWAg0DCvcleRIp49V/kpdr7U6BFT6MKjLEBw3Fv
BcUIHp4IHGLTXvxJlzt/q7EShhvDPolFMSnZ4l4QErLBXoR8tofd1awDYr2k4OKCILskfjqEESni
AJZtBzK7Jf6T+d5MCTAMVnWZen2O7iBptD1O7joBHQB2lO0LibxGltYG7LwD9s5VafFrp6pLNFZ1
MNxh4WhvXgPcmBIk8k/tkRWBqkiPLDFv0YEv/FqOnexp0jTUUZ1WHPtwMq8bwCKSQK9m/PZE2wHI
Z1KZoxQlNavYwkaYOoHQnSeTbnw4ItbaYUBc1CHFK9cK/QJ6sLOdAgr+AOJmvueFJ6YGEoe4EUj7
Iz98eSVFoPryznOiwp7Vi/R60vM5TRHUY28R4GE4FusmPTv6kS+c5Fj23ouQGxrNYCGYLQsScUr/
pmSfpPY0BkKyjpOYabPGSbErr/lfH1Q7UOtwGzlzGuSBYaYWqDqBKEC+7vjjjsuhsHiY8pHxaI3C
RpJAbO/OVO1FDCdHfdml82dUE7NBqoskvlrnUVpAcQHqW91IennEdSEpKKQNPZfjfZRIC+j4r8xw
GVLDvKpoxg13VqRHdrfGKz5y4kNIsFfvf1gwSh3+kMb/cc+dOaIIUStl3HH9VvO94mGmshoxr9Ul
0wbbeslcqGgEj/IFbxypeEeW+atJON6x3fvT4PbQk1OccgvlEA5UdI21lLeiKzybzTD28dbYnu9k
ehdh3duvXG4QBRYuJ8RN10AlbZ3SuetlXmShiycTVDzsKZ4bady07uKj6sY8XjmERl+mNOjVxQPU
ISHtrYsHkcpgXrAi2Z1Vx5bS1QFIOQ0fueZLyNANc1Ceu6/lEeXXiHCLQjiJ+w9xVK8nIRYvJG1h
QE+KAzCJ+0LhdPzKltY46GgarLOjJrcxM4U3SyGTxygLwzHlwC4twmaJ4UpTcEzyFtoC3kGtdLlU
vgxYUd02SKpx9mhlbqt80J4O2GeR7DM3jNGM3SFkCBaC3oextJzGq7gNsFN0bx3CKE/2cnUprNZX
PyeCuoqotSYigpmAiakqLyA6qh10tY4vqZaiN1gj0+Jd6kIZIFuGQ8x5LGT3IJASLcl16PP7Q20k
bGKKWVIJOsJDOYJpo6vf5BwvJwrl5gWm2j0W4R8UCuzRnTx0jPsNLdU9dcOdbioSWorOSvIrrgru
SoG7bYwj23SpeRLlFUk4M/e0vOPEZyZ96CrN6cxmkuOaAAdAgBEzfP3Zc74Rc3bdc7PHHG3fZnQd
ppVK1TGwnvmhRRN45zTS+pzUGblIv/1L2VrEk2KGBviVQEYT4Dcw/Lcs/HRRtBN0tYL0fKya2rdC
d9TVaDsn3BdricWuae7awB0Ln5zDMXVpEDm0jDtBhPZ8DPxA0jMAnrmRNs+gV70WqEZi6Tsfl0bY
42wTZnk75vRV2IsF/izCWuHLyxT8Y1pD0yUkbFV3fbaNHyJ9zg6dvMppyrCMnS21rWCqxDkJc7+T
oA/AnsOxHEuvuAmiugyA8deARTfDVS+nQzHFtd4lv0/+XhDz8MaVnmCs5SfNLVlcFdbzbEBMYsM+
/weMhX3yucFeYuBRHyIeQjolsMevJCJdLlOiZjUFJFRZGOKa9zK0IWcUk2nih3pg0h1MbmCJX5ho
o8Q3aY6ve6HtwkQ/k5eoHsxG/Gw5Abex3c1OD9LJObFUz/jORm2BgOZ3r2OY3EsjUT1Cj8v3DVZL
aV2s08aRHR1G47Vh3ja3qtk8iooF+cglFkmGCiW8HtiZdhBI6uzSJS0Syb0xWCbSIh19JQKFop4v
rlXyNQRZ8bMviKd8Y8TYV7fTOwOsWcokUa37g3P3d2tYhrrS0Q+6RClfXPVGk+YdID3ice+jsflV
SWK21omjXhsfMMg2yDDty5S9z9TfzvN3Ivr2Lh4keHX4gqaIxLIupizNHlCyMMm1+mUQr7aG1QYo
pKj3S1j0HaTbZOPxRFbWeH3erlUxjulrktSjIXAsohLAh4dDzpL7K310alLLX5mcRKXQb2OUBjx4
/OZSCmi7Er5HdTIzZZzSp0+VIVV/tPBy1TiuEk7iNXZbJtJUt8EzXD+a9RDc3ype1aT3fSqALNWJ
f1nLlIJpA/dgXgTBzPj6GokBj5h4isvR9p2V00Im1CWp4jBItWG2UWFZM+FRpqAEbqMpuZXt/AbV
MIcu0G1KQ8r5h5izLpYrFCUfiiLQQz+pGCcROo2Xf73TW1dgFCx8K6huKpBB58AJiWVESeGBiJ5h
Zc98KxMrCbU8aP+p3odb1/1EAzhkA11DCji9mkKretzizPKbeOl01b25xsMmWbYAkuQBasTinhss
xoWc4fKhrmXM58TD87xmJFAWbCsi+bAER41Y9G3Q1Pr6Gh8oGOvDBsNdRtOF99dPeFKezoX+Uc/m
I9ar9XLNg5NftFO9mET7HZe0PCH3+H5DdDiLzaTgFfJoQ/RMAC3SozRyu2dZS12oTeXPdTxRWM77
WZzK7kWNGPiSyFD5N3sE+sR0jlLDD4Ib6aKlF7UmeADqeJn4r8j70W/d04OCKwVDH4wrq4iG+EV/
pU3vmIDlYdzlaPGf5eCV/AJ+Bne74dCAsFcE/YH417+Udd0WgZw1xcKl+iup0+V/MrungLHc6ztl
yCdXWHetth6AsbHzWEALt6qof4yG7WYykY6tWQyG2S34+gegfjwki/gypkwPTpti1sSQZj4OzOmF
mWobBy87No2mFCHrgiQJSvY+iYcJ6DREXHG9YsrBXrqqmqQ4yswsHtn28aBL1KEW2Hu43AaMGL62
M8U2okmrrHZ904Ha8Oa633f5pzRF50QB6n7S8bA8GtZVlrXAxMvk54fPWPivXnH4XDPLww/CmP2q
gW+8pU8AHXito81aoom3Cr2tW52aFueX7bKRTYsopoiU71ZL+YDuJoZtXUIAf/4T7zG+aW/zezvj
eP+QQLIOZtlf+F3BFSsbiRXpHjnTSkLTKPCLnNT6mTq9/ha2s7+uWB4+x7gq8c+HRwI900RCR2LJ
+3nm1CKIsXmXRDLU1SIk5k4CkGlkYXylbpHtNXGktqqm/NqoauOoV7L0vnF3lCOz2Qe5fc060LKd
xAAT8N9ib3UpkjBjCk3X7EUMdnju9B4pzSQvAr7FNK6iOE4aKPYbFTuw4CqyKu1fde71+ybh3aVp
9LXdu9K82JHuwOL9AmRCgtV8/8AYM/fWqa1gxfhykdpqeAfEvc6+X/bGWrSYZoMW2CB46fE8SynJ
BpErxi26r/D49u3t6GrKnEOPcbtHidJjX5dTrM6gsr540FhNqx3QurUF7NiSxQH+Njr/qPqjAgDL
Na3fx/o6UeP/+kQZz5cMQ93U86WFew+MsY8zU1/EJ77P3FcQVHHxhGBBT0d9FPMpi0YyOJWs+WcX
QO1urlvC8+V6MCLDGVNo5GvXUIFrjzA1dV8tZmAasekIdA/Kb2fZ0ML/NitRL5X/jyPCK60JDoHM
72hykH/vVj83ne2Yun3pbzSTEg0ACmfDNmsPZukKCCF2hhavDQJ9q3uxHW9acuVXAn6QKAlYf2OR
jWID50UqKsxqqoPtcOV+OZrMGtKr6eUwfs10F+wefXXhSrlKWjD7oCOwLeKJjG2q9dLVGIEqdjAx
v88FsbPEWYOX5hz5cOVOb18lSUB4BmzUpxZPhE9ivhAqX88fnFIx8WzFZYEg44CfD4eaEhVlntBP
TpuG7Hy+YwHd0PF62HCGMeRVjICb5hqcnwHF4f06iQ0t7PbnBOTHwPlTYwq6/xr/zogdz5RVHBfD
jtL4w1dxF549Y2DpsL0ZK8bFt+nhQ6v3r+ITyttGwk2xTmw2lUrMpil5+BFTqqt1HTWSfNwk2P6a
hhxpTM8PEU/zZxvNId0p5ln8ZS2lFVMTpp9XeMNT0BaKNgMs/Ztos9c4LNopzTsQiQOUKLuinx3w
qCUe5aSETcY92HyzOUX0+ai/BqKiKlKMus+NQe+v/lruWzVZQB3Szh5Yp5wYr83BEN4AtD4wE39w
KGd06ic+ycIbAlrZgBjtkyDnKYWQX2r+oAjtrqdH17q6/gKE/iK/gUcxuQbGaaU9bCKIZ7Qr48no
u8/35uHpL69Jzm7IBeRqsii9JT93+ZtX7x2R5Qdz+pazHcTtpqsz2a9jBLTG8+AQD/lvtIza2syh
3x0TXhXQl2tYPMc6u02rns0csmIVkEIB2ZZscfnszV5rcJSZtcOY9S/wIq5xnzlS8khtZwARF2Sk
csbOWtkFp0xUkJgedXyczUCyqf1coaUY15IkwBqt2jmkBJEw4wkzl3BaB5nUE9PIzfGSSUGRH4Tw
I2qD9JQfRjpOT5z/2Bxy3//HMGAVaXIXB/NI5y7Cca0Wi8CSxrEiKqAvsOOcjL4LFHxBpbVYaOAp
kWTvx1uKPlHzje0XCr5FUvygyxGjjc1e3kHeA5DvPUhmWGpkD8IG38VbiYegoVZ4JOGDlStMzVGz
/PVpTzUUf2fESDPM5ZqnlOJ4JYHu8/mE2I1+i5jYEzDK80HF+TJrwWKAgJ1MaXXYqTQSvRRJDwEO
h5DK3E6QLMAclRaFv9oAY5BfOIT5MYub+7lYcEFXTLcgZcyn30HLvOopLf6klTVBNTuBRqCPywem
LksfMagrt81XEyfrIgYh2xH8wkBbFn2lOkoc8THah7yE07R1F/jU0ZmbMyUp0bbIFDuAbBoGLghd
NSAmw2MtXU4T+jmp8KEcSsH9E04hP+0THzL8zXV8oU8UGm3ezGVt+zlqvQeZ1uCobFlGkzY8y3+y
EDf/XCa4X8YsUM6mRYNX7EL7axQHyOHJkTCkPNA6HiQHfGhWJnEUFgnhY58O8InFLsIeR2JrkLcq
31u9/ba43RrRUdvHYl9no5Lre7yziAMIzCXy1NEhMVWzixJ5ERmZYuPSiwdUl88nrBwVONABguFG
gKlggqIaSjtrrlfJ1qjHl4NtlTdYbiNkHTdKLGhQZ5B8bmGNA6D4P+BLT7CrSWRXtVdDVUyW2Kr6
Dqpuw+9Prc/Q4+pkeO2eQokjop7LZk8/mUeM+c5UYIrpSiwn3oTckWr/pMxf6OCQVimkLhiwUaGA
gLPFC+xspcCqsT4kb8DPWXKWvjkCw3GnXXIteWYVGug3GSqmM85MpkJHDHFTPNRhJnrZ7cFOs3Mb
pH3l9cxGT1O1aSeIDYQRNb0NL5zTWSZwFx3rmK8gauYVvDDaqy5zglUZaHvEAYykTxueB1i8xZbG
ja8+bMiZmmhQrajnxAJ2lAY7RdEtmYHYPZ9bnMAQ94zE8unnm69IVizT4na7b20SFcPdnxy4mHZc
e7VuUOs+hMT2RVxMlbZy6qsO95z5stpVPuy4zJdFhuFxOetSKLGhvCUBc+k4uIB8QcdFP4F8XnHA
+4GorQo3StPIgJg72bIq1DiT3Kyq2uI8oS6XiUXHFT3PMawSNelFZpOxIBFVk+OVah+suGIPKi6I
nVzpHhM6JYDxdpATkOSzd+07ekhE4Aq3gX0x7UT/TpO7NuqqcnvLFmPWHPdnqdgwUCrjowLnFXlc
DvjI37p/NYwOMNA2+CiyK8dH4nfKbvYPGBIGOk5MorkH5iOCFSzQAA+MY8HPAq7klwGiZ7oMqc4H
BzR1NbF5nUMf/BQVdS1MLVG/BlrrsBUjICyEKRlmXf5LNAmtuquUMqYvjXqSQgms3W/V1PiQpjAS
KMzq5jW+NomVdbO5eccCkwbiLef/2DwprQteZ/GBZ2xuanauq28DnFRGn5ELv/lzGI2QRYXoCpiX
8zcQk8gJRcQkl2eCsx/Atem4jzfEgBuhuKdoxwp4H8Cn56hdY2j2gbRYFlxSoKrb3Luan8zkjkoq
zq6q12VWksvESrtU7CbjM50/Yj8AHnLSR+5H3zhIm80dNoTGCGeOgBlcJn0kif/eVy3NOLMhT3oM
7tFX6OLu3j7J76rMbZxFoQJ0qe7jo0mdKrmwDhI4mJAoDWnFZx2kX2fGLVoxiqHVuqAN6XGTl9yx
g+Inj7D4U0EI1cwRuRcXQW6Hr/30j9jjLmzgHCrZqZp/CDTvhF9egT750e7494zA3ZvgEU8hNWaD
wYxyrxryov1KPo1peQCOTXbSc6QvPScj1b17DKK++lmTEm8BRL66gQKELGe/7tUMeQ5OWaK8PdJg
G4KU4wVLvHb+qOtrjec6DuNdwZprLINiAZYAjoDaAZMIxcXO1JmOzRMNdWUiJAs1H7qrsTVTuYOh
A1G7juLifCpzyFLVupwwDEfkUO82T+XSQqObaHKQIF4dKtWqhiBIyjtG62om5el8LpmXSMUDtH/u
o1+eh9MrtN6FFLRuYwGA8eanCuTeBAObUwWKNlvCwIlbl9XCe+YnobDAubbRSRM5bAEqD2JnSS54
pMA5H98NguHTHGQ6MnZ7YtAMiuF7kNGgq4/M3QmsBmbAtCHohiUKRoKie6J/7ntqnMdlUHDFrjL2
HNuaQ6ymPiw3YnkwoPCjnvRSYdZxKLxYdsv3uOuRxJCUR9lxw/POm0ez6U4K+5saQA1MKoOb64R1
h6d0n0ey1ZE++3tP/JrcxPWfmeWGd69JVlDoTeQQoK+jEObpNspmmc2HrB6lsS39UmYM+2ePHW1A
+DKa5L/MSs8QKSoIcF6fa+GvVdI8me7DBHqJTSP4idsAYoV2fJ+umtrdiM/hdtOhxhNyZOT+xWfK
2TQzmUxaJUiuma5A7lYbhBzE4N0moEUpUC1Fe+YyrCHd3LWyQKZbGUuQAXi3Fkuz4e/DvwPjiS8H
Bn9mpZeyWsFm/Z5XtRu3U2Ox6FCFcNFGt5ay6pTo3nzNmnW4kcsbH0uoHkzOKIoK3OeCOWNey46Z
SHG4Dlcu0evErX+qmgrZ2bnqzvcN258sm7+xWGXAKGtWK9dgum9Uj5V6d5UsuzcatKHsuiH29VCR
lbeEBCkgW99cWyc4YDHVmlggkRUKEnBzrAuckGJy8hqe386QuNLTlmcOP6gcNerxWVKXTh83sVh0
/sof4us1zyzOCH7Ky01B+O/DkxFS7I1LpsC5hRLb69bNEGXL6IL0HNsks3YqIR64FYf0HXzbph+E
JOmgNCBYLlPDy6qYHGzS/BfRQ8ejQUXfzpFQkoCIdUyFIDvpHEQOYsiFFvcb/pc1u3bUX6gvH/Md
3ugRyp2OpYCQZK6r8bbXHnDCy0+PM8pH3ZdyyXVwcO/oiC5jxydPzJYs6gwCYpJjF2sQG63N7WX3
TNNx2Nh7Ze+5CtJA6ZNF143qugvIAmfeAmA3LNm3OuAHqDHMEqJLS0yaM4jf3tADg+9IthCvMWw3
/9cvoDu1z54sfetw3aoqFvdz5/rREMicvLTvb3WzTLZOgrA4XRnPds/19UG2u+9RrJwhTl3ReRyd
4YsOl4MbUY25+vhCT3X4e/kLID5nNKcIb9K2KFeqZZyeeWjoJ/xGYXYwI72/k085YZnBrm6RIRVg
8Ptuffvyiic/y/OE33mYgD2bVwexuiHFsH0lf6w7K1yssb9h/a+7LK0BhXia4EsGCRs4Oov+buY7
iRitZNqfuhwga+r5E4nexCY5DV8rUuD0QxfICTVrt2ApAE3tuiHG40CxlWHKaY2HowjJ2B6QT02V
8Ht0vFpwOzQXTCj0WiIFxAdxtCSs7qM6F5fS4tXiZ8szf/XPEHEB7VZO5GTat8pccYEna2UgFqKg
SuI8IYNV5vJF+tgzOA7Isq4zSYGONTMqSAAdbczE3dh6e6BtFErWr+mEpIZgV3zr+Oc0ETmXpABo
KkvjP28l4ITw3r8WPkr/1ImYJu+/Wx7BZu9S0T+GR2YnBtDWCfRPhkL80v/0+6W++jExaE6WkZE7
BEfhJ2lrFkLaC1uSWDX+ohvyY0qN3dwiuW+q7GtE84m2nu4Hbo1dR8Ce5d5bduxG0gCfKuYy4cXQ
y5w1I6G7OlCYvQeDDzLMcgixrU/wDad9mf2HOy4Ds0UrjG2KOwRdw77Vg91wQrddcI28J4HUBxSX
l7nVI2BUW1w0P68GyEDUDTh1C+Gz/sise6iIiGiD5+95j2qHp/n9TTkkq0Qo+8Dp+Sme/8gXIh7u
BSGz2GJrh+XcGGQk8STcAh0nmJEqRf/5z8j/aOk7uVIitXfDjEGuVfn2N31fUTww49CjV3T2x97u
lMb1i86DxoVsk9iecCh7wWdXwbh27Hr7fgjpP29uXiKEbbvGH2a0Y/fyaU86b7yBcsleLjbnyv8J
f9XPieOwZOK6CgY2082MoSsbPii/cdlpmGilq/7LZ/uSwUfSy59/DvTxutWbE5LqB3ZA75Mc5l/J
x4rAKuXGbTC1HeW6PBSQiebByPWNSpWBzRNrcd/DvxOBaJp/PnVyNdYrRCHPufb6FjvQDU6kV1cU
7wPZ0O7SotTZi65g4Hx8q4ozXPICf+RCZ3NHuJQArOK8KTXNV/PD4FBYiddb5lKWhvMcdfLSvzh/
bCwGlU5JeiQsjxeDiR/6gg/whDlkoxIPCEX57RJrE9QQw+l+hxfuUvNBtB4GJgdUFoxDAJgbq6tO
4djBMjmvgx4/uFBmDhMUAKRNzTS+W642sKytpG4hZKVz6l82uqJjKu6EgJEAWqbd5X274v83E03n
EUBc5g8kuPXFMI/kkwIW2qDqHz7DE4JFSy+uLFb8U8QuempcAgfP69nHZzEdzHEPxsFqjaTbk6AL
QCeWDSyZNLdb8EBUFJrF0PO6mR3BoItycXCYw/SiAuQcJVcjZpETit/IE49jkgd+oPvbbCi6b/7R
M8iCa/TX6qFH9Sd4yp8R4IwpgFtzzQyGGG9c3Slavvt4Z9MClDC5g49gon3bIhfNce6HJI6QSvIc
vknCyQ5T5Qj77lDDStbVYHAhx4Tf4pzCQyxYsha4ZFad/3nDo+XzjBjJrNEJOvfp0MUgy/891NJx
BxbaP1IBph1kvjTO9s0vZ8uN2DxaOTOlP2h+QdABQvpEY1V+J/2pvoLtaYCqHUCGF0u1hU7ZjcHi
Ghwh/3kfXLkafrqpY5APZRwGFRpVOCDwkobYr9EEAxQ/7RjvosA3pSfJuVxuBCHZSUhC9wOcC1C/
Elvk7bwewWr6ve1xxLOJ3KG5BTSP97ppy4mQg76QwwjFWgqNAfyKdRMMT2ySWnHNPJtpCx4NrbUL
duEktr0jdVYGPLz+UsV+8R1Z96VLHf+CnhS2xuCFRmih6YO6z+31esnE8lOpe/C8dyAv9Qr3vqYO
4ApftcJb+Gq3p5kLFH09X2UWtxQb5VE2/+MttCAOWTn1Q2lDc3zW/is+YFWOBqFoVLnrrgMRKmwi
YTfSFQC7dgz2QRANYkHIism7L5nY4bpq/3cUnk860z9Hi0VLy7aNALj4O31lNqZj7ZPgYXllDtCB
b94qAKzP7P4p/uItEIKel12NmvnZhhIjqEDDHlx6sQdpv3bBJViTyVyfcvBT7bYkwOrWkeuDEQPI
dLC3O/CnBvG8HEaoyBqDljQlZNdhhVvup0IoxnklPuXJF2bO7bKtEj7QukIRCaelQdWGsyqVMN4D
wD+wNIZIBLNlHo+Fzo60ZvXBl4/0gz/uFfCWEEaiOdfbxHznI6SBqlGNGCyZR21eK8ww950aPniE
KM1W1zo84wSMJ/ifVgZBmRD0bNE8TATGyGYB7Ywd+Y2O4dHWEFO7fhsTm5LGmMmQGrKt74lC3e8/
RudDq1gq2dW8/6aFU0UwgcPwGiZnkyhgpuPDZCYNXuyMlPpJu2kUYGSOkOcf37O45OahFaSqqDx2
TZUD7sZxeY4TUBCjIKGjPR+DBkKvJfzsy7r/2AzcGNe3wNewWPu1cd6UTd85Q8gQd5QQw7IcYjl9
pn/ZSKA4J+nw4PBQfUYVPxfIbK/2QiKNtmM22m4oUgOd8EpAvXbt9KQwUBlo0bp9Ydxx5OKH5fmm
Z26uVdDJm03k/w9OQUwPupQA74WHk0zozXHFiTYD+tUcQssv7nyHr3aIj0VCO7tRnwguXCWwxhbX
sFWmBGjZK9ch5NHHdLoLGxyPKBniKFx24SU1W3kX059o2sJfcAi4peKWiMr4ENVke7i6KyLhE0cX
x3O/YLZ70TlxohcUzo0LliAzpkXjfGul7Jz/utx0WMn8RjlvzM8r2lDLaWty7WS2UfHE9QKVOpDw
65n3Ym2SilwvlAIG1HwBNioOcW6EFQ6KDAfNEuGqIMQ3MYiN9V6Fh9h7KqU2DcBHTEKkF96e+1Y8
j97JyVDDN0I9zXlimRl4VxuSPeBHNEbt9bp39GOLgGPRd3mBj5+6FGX4+XRXSTPKixCz6ke8nnnd
1TH/GCEZUTRhgYdmr+wFEpS/I+weUpWlb+E2tib87T+Icw/SJy6onPBWpWdI1IGSxf38VRFtTqnA
6T9H/Zj5bmrzuDOl0B6WuDAXoy/pVhUL5b6Wtqkly7CIRt2LZwYhwDb1k4Wp286KMN62KKfTqchl
4p0YFV1uvrLA1i6NIZ3/OJU5gr0TO4thrONH5SZpBOGyaY9UcGV1V0ZCvAWLmFV1mCAWcG6F31mj
iwwmn9bxcGkQMcjDXC1C1j5axzvDBnPcg+YfjQoFbt2NWjERR67UWDME1xJHRG/Au6TFZAnlNbyO
C0gdYN4ghfgoM0hKn91W2BOYCVnepvPanNTB6HjRK9PvDUK6FEN4artl9kYaAdx3b0x4Ty2fE4Xr
NE8ymKT27wPtz2aoyPGt8OHyTCta6cu6Lf7lvHg0zMWnZeMiEzdLoxchYMXg6YGYq23bfi9v7vU2
sIIzeFwpU7OFbPsC6KT4uxEbwell4cWzNpETiCYyfsC/SxqJjQ1hYu317b6LMZBA40LuSAC0g3iY
zWvmHuJCrqZCznovEv+xGmlL14YscFT4LCuHg4MftzkWhNeeeMqn1dnfcIL2o4h2W3cpQTPDHBLj
c7uLFHGZ8ga2FqcXYZymScIBnVtshydzp9VABUDzJyPBeouxzPHHTAlgS4borkblLn/LKOqejTty
mWnam+OxIKGEFSdgXB/kaM5GeddU0/hOmKSK6OgRnB1KxO+OU9/qtnIp51rRICOWhT3Om6NW79Ev
1mzEfWRRSEE/hJDq6AyhGZvzjgcDEFGa9uVQKa/156n7METeNC+NJ893AISftTX5CP/WuxuSQNHg
tdBqYhxYYkjFSTTE+6J3PoRxRfAJRovOkoF1jjh82+gFsEf3WO9j34rdvqdXpI/b3Jnwq52haSON
ewR6xdOryJcN9O7IC7Y+A0EPrq72p00PG7OVDkWr7tYnu8b7Q6GsmyYP4wnmOKa9OYlMISt1UiJn
9TOtTIpY9eYnD/BZKuf2KZj9oMIjchES6JrRnWs5jWKWZf4S5CZwLs+K5DuTP1aS83J0WIzQc1N7
0Gn1VSs10TG604w+7rQ7NoLeKBASgv/JrKPgwVESo9K+pJDspLs/w12gNbQXawlZDvoBlus8BC/F
xKO67EvY5jllA7UQd7IxA+0CA1ZH8V6tbLhYv994330Ihr7oOkFiil7/h8ec8Rktk8t35KqCHHud
kM2LkrUL4ZNlE45rGPF39iQj2mHEBv1/YyufDhji0//mZOBxxNseK4bbzg4Nx+qDxilPLnVQrVi9
hcmNwwlJaLygw9/ek7CvnRX5hnBDsL1uvJTPJMual2J9UaDoFdU4OmrrJuaNELq2iCvX0CVkfCvD
kTt4HE40QR6irPZlNUMO3rFXIQtcwiJYJZCslfyclLOuXS6wAxJJVbwBtDUKnS3jPOdgVUMXg0BO
OYPUErKbvrXAUz+g+W+auM6iq23Yk6rLh1CcIjGforEUpoHTSutgPQ32RRM9sZXqlNzzckoYQxU1
iQmJQ8HNHHlXwnF9RcgmkUv1Ergg4QAXXmmxnJAYsO+rSzelOYdlKv+53Q8qIHgW18OTDU6i4JS9
CEYGXLMtYvSzuRCR+AOoJCjUpSuo3qUXmRgU2xGNEbnGs2JwWBnK6S7Nm94gEPitPA5F+fcHDvHq
y67yDcmwbSBJn0vucS7QWT085vERJ0hRvD2gClwALDSrjzYw4sQ/fOf18dkMnKOBsukSsQcE7mca
HTf7qHQO26QisAqleAIJl8m4e5RelUBf6ZogoPpVS1QtpPj7YaHKKRBpo3xk66T8u/sqjw5T9Ier
IYoCI4ChM5uv6GiDXV2qt6Jp16t+0ZGQtbiwCDtyrbeQQhY0iWZGOtTlut3OehP7QeB2Aha0OpZy
exBrGf78PhUw22dQqKZnyAcBcsDoR0XLcM14ZZBsIxa7UbPKSW1IkiIaxbr/HO6yY3wFPey+ughu
ISBIeZ6NxoEBh4lwQRj7W3qATBfF0/eRURu227Cb8FZRI6EY4YJUXfvq28CraphLKt3De7t4FDIa
Hv7oh0bgRAxPUMPjdcDlYi/snq63XP6hKrVN7+hsNr+DDMioGvVIB++fDw6I6hYUq1ziCeFVcHxB
bYwSnkGBT+JkESA6j/KaB3jvO75+f0amXgvnWxADtwsYM/Dhep5MM7I4hLbg0uZ8RiFtXFbespt5
GYNTaFRtsELRG0yQFPMrafok9RS0v7DuvXSAgZYhVytxKDFjaZFrzhx1C7dIHfrAkkOVAt9mFNyD
XzC97eZ8Yr+yHYM6t3winLgOO3lzksAFC1PQqPe1eMcLbK9kIRN72XWQOq/3q0PvONuRIc3snzP6
TrHYD+9CF8V7m8vZf/s4NUNA3aTtbDWGsJjIP3TF9Gur3q5oPEJe0nVIszMNy56+N+yckMtkXuNm
pj1If8MqvLFGbgo/6rafY8Dk7APxlAszzX7BrGLGtPXu7jZNMEfgbqkQJvnsUKtobIH0EwJ3k0xl
Bl7pzLJMA+4Y5J6ln4FFWjTDx04AY8Wt4a3XKhF2nMYEwBcYLzsuqSAGXdTv5chDUb7XQwAkbRgX
H3L+2skd0eydoCO5XGFmP0yhi9EypQoMHaawaQmRb7/I+4iUZsBDa+F4/JhsthyzuwIeO0wOxcxd
2C8t8X5HpngoPDkzHQLHEXWC4o61EMfU4V1C6WR6FtZmKHB5puBLZqZ2+NK67R3itXVUeuovtMZ4
TPcQPgGsuWAr7ycyNuBIfNrp3KrXRNCs8XyHK5Ai51ljONTfWsWB5mEd+J7+lfrpm5jEfsYDpGWU
M7ohNJsY6Q0wWGRpgSt2WgvklX+fDqmNecAI6FC7LpYfZz0gyG83er527/SqJp7ePOUvPXzLKbIl
bcGRgfUNx3We0mxDMXSoCcdAV6QJRKKbst7mHb6Ak8uHyiXkg0GOFfWz0ox+ElGAfiYbmAkanml6
8+qOI3BydRY29wMfofNLAFWWE5GGwWTywsGqC55AdjtN9n2KIw1GxS1vCuvOcF4eYc/fPUmmxFgt
25rKGSR58pwgtPPe7sa/NMx/ar+Kxs3jz+kTyo1UeMhwOHvkEPSdQyEsKi0KksbZFT2ExszpXU5g
JBNCjvV7QrZdr2bNH8j+dEZIHy9rZgEPpn1crFcM6vH8csLeTkxazIhhQIcxnRdXfKdXlyhbhNpt
zwrzJuiy2TkVRR7APFKy2NGWj6FlEK1zotMmjNIq/Nmm/TqaE5e+oj+f779V+tHIGxSUVpdk2LhJ
AuO/2WcuTL5tvNo/uSwu0i9aZq64GHM3mrdRN7W1b/MD7YIukROO7YyT3BK7Av4YecRiAon2pvlU
espaQZsi0aXuS+7fIZYPO94SbSdscD6PDVC5EFHW/TyfGETBiskfSqd1OoabYFcOYAf6DFFfxW/i
3pkDfcfCgNf5kZ1oAaDk3mtPUHas/LLALVsn4Z+4vNEBgApcdkG0+xC/86JHHoK5VEbxx/iZjV5O
8l6HlygLbaERDdcspyiyYIwUw4+WaiFI0h00QgZahW+QdzjuDxa6uKLhrOhd5ip3Wp4+U2eme5FA
e9Q50ynQQmlvAiw74BjgtctxWAv1KXFasi3MCXrc8zagfOyfGO8adLivjiA6SK5C1uno6DbPJ4TI
8LDDbTRAUWP9bdZiAvPVCiQN7bAra/1WCiLOnYjdXa6ioIyBexn+dfESqL2KsYE7G2v7rhlntIxu
y35M41EWvt9jre5pQhY0/cqtwDKuQGhYT4hUNKZV97Rb0+AMhumXm+vIcOC20JiJVEA2hX66zOVs
ajgaUK/rCcrbBcvIWpZyYWOD2h4ro+edwZZUZhM7Q4HFvFtwcxSJItFEp/OMkPMS5EbpkY8TVU9H
YRcIFygw8hWxNCUtI6Qy1y70EScrodigsfeWBTFbdTqvhNKuqbRmHCZvvDsDR7wmNmbCKqAUTHVt
/8I/gO47hDMIRbQCczYHUP8RX58SVwKGydIPIra9Iy1MS48/XYRI5FuFrdphmaz/bcmxUGB47oTK
/8y1JbsklymmSmb3g4h+cKSpNJBNTpD8An1AcM8Ef3cDUTJopC272KhQg6JJG6SPYGS9+Yl91rNG
q3w7YQSxjZQ/KxmhB+jaIze6LUsUrQh1Liq6PXOMRU7nAndOLpK43MgR5stXfRxpQ32QUu8Nie8A
G9Oln2Nyk/U15mfFEXIsi+lr8q/LUdewDpyZEBj/X06kB+VCXa7LKHQi/h5F9Rgu+8ngvpKYnNiX
DstBjdHF5NAc5KZOZcmlTiNmaMLCIjqG0iLl2oEn32Wl976HohQNAf4o9NBRm+U9PcXyEI3Dmlut
BbS2/5ziK2ATO9cjt5iheb0jTz9KjIoTRWnNvm2ONmhENgnodOYZ9bA3wH6Wldn98GwhRoMXRLFl
c8QCYJAvj5O8Y3pQiI5RbIzd15C5tjFKA1PqV8YJvjtdUNsLZmCS2bRACotsaKnGhn8kJpa34Eal
EUSTjftCwNX8H+WyOESGj+uxqKQO9XNlLULbSqKeepYEGvY9F71DavgznBtA50wILSt0GGe4URkG
6TjECQ/GwcsmegPXXCaJ9QZgmeuhL13zIai/qQY6JbLXFCQrpIA5XTK/44+9MF1prswwivZ0Ez+9
a7+KcQw2CXyKl99L/8vFu2Am2/RxOYvohc1iAtb8XcqHGPOmx6emtPgNysprh4KRGKlu0MfHrL2L
NSAQExdt3jT+tOWginfsjsjGP17Zx+dagMdmfNWZi9CKC50J7KMzAzj9T0QLgesmWMvKvtspAWqb
i+5UY0x7MU8Zc67sgEtDZFxqZ8fAMfmStVGdtxp3cgJUgV2byMrq+OwfgWjNYJXySPKmSn4cqboR
gi+TIrrvvhfKJtJZfnZCJ6CF8D8WM7xGl+whHAJRvqO2kADmeSv91E9YWmYK+RmvVJ3uqktzdAFR
xYL23o/kEV/gNjJnE+J07QWwseJmOnq3si5DEjiMPMrgoLGx/YK/6XHzkYf8qZNQ26t1ZGkP+rJS
7sBJhBex14n48a0nLn7W050mNEanto3paJzXdj9ggrhFsy4KdmGXjhkZMYcD/LdDDpL6xzoRmfzk
IEsRj4n7L/z4X8UxTdIXLqICnDneU5jpBDCknA4V88vtKXu1zZzUc5eniWYY5JV1WuOLHXXBpSHx
7RhoLKG9nknPAoMTuPK8+MjGduroGbGnemgbF0FjOyI08J1wZi4n09EAKDvo0S82FnSc7kJ3ZSAi
OJPNUd3XJ04WAw30IN/n4t++XHrhvUfL2qJxTdz2tRaLOV2uiitgYv6KgZjwCPKYei4gFjoV12vU
TfNLvDegeVILxaPpH9C7QSDj4aAiz2pLWmDN045xtA9pEaREnKodDKdqS6ZYZ6jwTrPsaoringyc
ZVSY7aLe8SeN7ZSsHOcaMs7mn3W0AwmFOVeF7AYHX+iLQYq2xCePliCj93xrGh6p4R0k93yJI1EI
GxcPtZvdF2voSpGS30GVujvW8yNhmOKziGmViyscaoGf1gydSNDeapGlwCTGqjxJibE0foB12H5J
ymQe6Fqwr02wm/+c7a9grc+xrUPw7Ncgkce4VQ6LJQp+UKD4x1Ls+/xy0tq0awFyuLdT+2TVkfXx
UEnUEdUbuPq1Pv0Hyk2iIsxL814LLto/MnOsLz+mRZpU+U+mN06e4gB1GwLDWp9uWK8b/do/j0Sn
LfUH4m1V24tpI2hVvJOf5wSR8phlGgkDUTo6nx5F0oK/4rXEEODJH+kfI9kio4c063xYs4aIsMAV
gKu1Xe1suRa4chpVRITxp39I0Vz+pyQITd2nGMrDA2BQt6yRGWYVVIxc1bV/w59uwiIuG9BtG/lk
byTDxAJvYUJcNRq5UkbVVCOoWcsO3+ftHVIyCBeyBn15VcYkM0LavMGcefMIMy81ojcHZ1H4Ix0v
ljSpMx2LljzxZ176uuocSmnh7z+nRA0DhtezukOkoL0GhAPCOHy1WGDo0tpfT/EaauV29WOj7u91
NJbxsBpIqK0zzizkrVr2zftjnenVRPeP61nF12V21rynJohoX+dCBYcWUIMef0NKnXMb7a3/jxrw
jH0SkKWo9s6EEGZ3vxLhPbIVZa5hq3aNEdMELfrB+63dhpsbGj1eYMMlbTb3NzO2AEVq9V+QOJXE
7SliZXFrAwb3DzNK8znESVCbog2xNUUzmCNlo4Lt0GFRE09RRxWkig6d6FtUNJ8e8m9t6OhvU9uU
02xrB4axixviCj5wVDDv1aY8TNltE3uSkh2KlU2dVyNEk8Ta/PELEtFzxazDWJPS9OarTXAcpyY5
V/YKtYcHqIY/MNWKZFicpx6JABVYqgWSEuIisrNHvBOQMcRV5jvhG8mtjWJsVft7wWUUhK1Tf0L7
wC+N5yUySziiusEmzastV1pHJcJ07BmzGu3IYjgK2HyH9zHxOPPihrupHgcn7AJgwCOPdj6M55tx
qTmM48BE7zbHEGDXBfq73mjYzQXl+4XzXTu7z6X0NGa7JZp/mtClilnZ9U8EPpHtool53CEwQe65
qajO1pLvmO//uwvrGeaxAk5SF643BXz72jKtc0ZRGebt5RK92ZyGS5ld2FDMMWt1t0Wn8geJccna
5r+2cN+yJSXHgtJcfcEXpn1eVGU1ZwQ8AItnOCYOrCD2C8zhkMOGv2Lc/uHyrHTXirv6/onglbCd
ogVRCvrKGeGiDMMUtUxZW0bFtgPlGIZcnpOe0fdQcYSUjoWq07GHN8kmjikOffObqbnGcPTwRhf3
fLuApCeuVOw1rZBmNALG2oqsIbIhWdkV1uEv2SCcTP5not8LInQJo01GjJ7Xhy0FrhUnZhRsYNGo
YTj7EFnnIbtBP2xG34kWZIRNmlWDpkX5g7zHjbsPORliEOHUTiTEQRU/1zFWqMk7AC7x7nvIyg+b
IWLbCdXhbhipmqpWOzohrDuFmlpa6LBEdFaS07CjSCBtdnRUTPOep2jfp9VVNPlV4vgpkGsmY6Br
PVelmWPKCOAV8HdFOYaBJlQR6XhtfTjOs1HDppX3zQDzg+Gknjg0GX7zdQS6qp5UPMS6ieJcgnXU
/sJqWs4cwBoVM7VVGcr+TR8X6ifXRbdZzcW/vHJiLZSgNCAdPE+rZa7XcnTpmuMGcRWLTdgcu1Jy
6M42N9wnY2eQ5y5uDoWJCEGDFASXvybFE79nhbh/fRXWGigGaaZ5M4FYflmGJCkiCCNh1BAI+NW8
Rl6rF65DyROiFZNEs9sjJUJWlMcQPi21z7NpMFKSPA6qEBhDGNz0ixo35do36ASzZ3bhEYhTw7Ek
6BGq5fhx/RIboRE7/2zUSzYivVTUVjZBcUcNC3jUF9oLDkm5VdUCDUUf4T3X56li9VIyKPqYTq5C
xgSs06zga8EHbQgBj/TRd7gMXfy7BheGfVWN/IrPdpKf05WXVZsrEWthsSofjPYN8RROjzr4A+kk
BpUVAuSPKWH3PVQdYL6LiQOozscrd+RXE1wObmsOH8d+EeRukWWJjma9hZPtjCLpy5T8DtUrvInG
HQ295tCGMrB6SZJkyfj2ae7ggCPegxsKSe2nTNtKKKGV7BV/HaGcKd+U3Q3qS0lYPDk5h09WIpEx
sq9QB2HTZ+5tLs/7IrSS0xU1fSNTUbev9PsNO/l66LEBVwpNGLS+aWyNAw89quMrQ+lcdexWblJ4
1kcswwJf7S3r/C7U0cmnHgNtII4nHCYZRtRI8e98W/rsobDPwkmvNpNfp3Uig0AwO9MTwDoiDnsF
JLEleaES5zMUUEJ140k/jXUZyXzHl1qgP45ICVkvEBm34s9cUEZLuQ/fMC3uY/Q1FM0R1ZAOvp5W
VZLxBkTaeFAt9vcH8ljkYbkSEYTQ2GDLIBBDTKhb/xmLg2L4PjvotIcoB39Y/hTVJHRNZfsaDhpQ
ONh9L0zGjkCB4TStYLbrAlmFFwuy7a4RQZ1ICg6FjkjlRt0/6+T1+niZEnt8cj9eIQNsDPSZmMeR
N5eOHryyWIG9dqF1gn+fOT5CCfybKB6RlU8HzH4v1C4+HBxKnd3MZLKb2p8HfYGbkqzkKLoVQ2R0
SI41d2Yg3/OxYEcn6AdCaUZzGmDK9IV/f5D70iG5RA2i37nmBZ7cYlyyHRm/Nt9lEI1OU/RMIPES
p4Yd5ch6JWKlSAQPb1v6d29tfTprnf067i9+5dSgZ3R0UUkIDRxzOSZXmFw2cnOPjX5euvsMgiFT
2r3cKjuYaTa8WCoYZFvcd6JjX7bcU4oUAG4yjUHmDlTBzcG1I479Zz+gahirmcjp66cK29whxBnp
idrCfHvC59CIwjGhhgcqowZaY7WIdNdXXSAgY8t6eTnv3amgD374SPyUiVQ03rUMVVN/YjsOJxhW
KsT3pj3p4tPyuNFmL0aHSicXJX6egeKe7QS73nlk5n1VboumHVlU+9wEsr6vpnAICQ61Tfk6unWn
wxHhrIGF4+D+mVlu/OulL8G8BmQsywwNz5YC3KJsv2H7Lywe8OxoyvXXYS1q6ef89F09Hvhns45u
xm4RP1y129bTTTQ74HcYI73CY9V8YbqhQapThmBAY/XcYiIOLCbV/iqIEioQEtq2cLiFz3mbnD65
KDbG8PXiSAERdObtRxlRXn3OVRvPcUgj8/WrCHxrm5qDCaR9OjbntHpS2ek/y1gNtY1yYlzHjNpZ
OH5CIaOIuqLMWYnuBsTTkirMraTIno8Yfljg2eDAS5008ErMiprrB3+tp5spm4AB7kzy8S/8nQQR
h5oFqw6+zfuGuo9zkvsFCy8Ftj5b66KXDdJxiDpBECiuNrfjg8A0g1Wo116+M9w5biojFBueqLUE
1weQ0llmUXP1xLKAVUBJWafzXcGPxQDYq8ghoFDbWylOO9P0l1IRDwXRz8nUdvhCoa3cVk441A/6
+M8Q5NnA7BHVBOt1ZPb8FbRCsWQcTkKCNG6k11QeamSXijT/TNay3DYQvsfuhuAs9HxfmU/iQRdv
HLH4KSrWv/9Cmj8I2Do3gEwABT3EEO2oWtm7IuQNdKjKQfGVOrnpAAikTD88Js0+9/2jlF4xG+sL
kbFVFERiDMM3BtfoP4Ry65aauXTMu51EjOIv30qMEITX95ePZoudpxBPbvbVaGw3XgeMqI5+kPeS
eJPwUMP575uSkJ6kWq2QlSRLi4jNyER9ys13SSR9u8+6zB4mIfI/s1AGOwVF7WyAuUMekNSa1wPf
fKBwUUBzwjvulve6lxfeDl4wtI9rJsG9pbvCd2mytu7YGfFt+Bk5fi0fVtBwg7oRcdnvQyxntC3I
+RX+KS7iDHaOQg/KcDPUYymkGbR4A5+nTho9+7IGoe/d0PkWd/bmOfhCLaJgaB4ZenfTZ73+vQa4
bLeabLN594jmOhILLOrchUMhyLe1YF8r9rwWKTs1F8U6jtg9bq1WJdtSdWs7nZuixnneVIfKwdVp
aOpfydpnVFMhoPzoCt6TZ6M0DtisDFBqWkJu5HdB84l11S4WfyOJBATbvb2J22ASg377sqjtSrID
JVn7L0kJMGgQAESCCYs/jy3dn15Nu7dD0FqRXo5T5gOgpkxZ3dYh5s0zHe6vf3r+gZPnKD5/tc2t
zlqyrP1i+ZETyBvPC7WrnPgDz1Sp4U0axNEFvDD7OcjtBIReoThilFEti770lcPZuqtq3jaGX1pz
j3ZZTtt0/r+KQxUM/+5PA0g6wOINab2zlx9lDhea1YDdHKgnC+IHinflN+ikjF3pNyehRJZbz5B2
nxDTFGHglbQHMnCQMwEKPyL/5QspEZkvYxYtQE0frOHCbEXlpjTsa2/2rEiMnVQ1jshS7VCGsSYo
qcbWeUfSzsH9J5U8J9hyBj1yfqOcYp7xUA+XDiasiZo5mYTdWTksfP6/OnBj13cvE4gU7pWSzmpd
bLa9NWWDv1uZ052cQ0Q+lE3pHHyrUY03lGLiA4PXJ8eIChxq8uBe+luc+DXvXz3czPpFxjql581P
N4gjxikptmu3hT9QACoY2+Wjw5lY9TPOunR8Iumj5RYyFDOcshpbQmQMOfcwhDPqNUkFh/X7ZGnb
pGWA2ILA/1I6wiGushkutiOqjzFnNRlggdy9J3b0P8PMAMtfnkN5ErAGWxSNfQ39JM4ru+hBF4U/
eD2jCQfOuwVjX1cE8wee7hS+gGh27NX6g9LWi73qpgvNaKwO5SXqASPjZLWjHyXmNFMoMEC3yzd4
K0beUdmSbQt9xC4JXDMnKURkq6JjpN+eHkV7Rnov48wzvFOdLgR+3G3j/NUS3kgiCU6d2DqxEhTZ
2mhyWnYZD0G+exUWn487eUnsBcC3unl49mTj9lgsDOltsoLjkHxi6BUzvZUoPKqsTLjMBsIhgws3
kav9gGztFsQMd5MCbAyKOf9vymfX061m2JRVcr6YsCwBQS63XjOQE969bxrFOKi784lNaS+sRp3C
OG8Rf1AvhrShtpK54RuejiXikCrQbucooblq9pev0FwX6c9wwITfDk6u1ERZMh3S9a0ZUE1ojI+u
oY+6IIKqHmi7PWFKGYpl34ipwjGvY8mCrXc9xOdPXb3X0vhZJI2pl2iiRXOJQjd1X49al5IMjVrS
hPLOBsBIpyFHCq1EtR+xjetVjdrGYRbSVE4vnSpss5a3pm04AiKeiAT/cSIJWQnVaKg7O/ACXrSh
QQdX2XBUkWeFaQ+ZNsbjBdbEEu5DvBCq9n0NTissixxaLzaiuRdcDLNeSFarw3KaiB3VT0M3DhSm
0ulaorr1DksSLWIy3W6tqvFVPBETAJe2QyjQ6Ra1GmQKEEk4y5EFE1y/diqOT07jR0KLmb2s3KDX
6cQk7mldogav6lcL54er5fOvoBmvIR7wOLikDQQJA5y+8KI70DAVEA2yPurv7a2z5pgXh9lejj+R
caRqldxrGg3+FaGy0h+BlVDy6Suk+bBj1pOp9sdmPzNU6Yl+OjW1eRu7OLpudrMqZDYukf3GHjQo
PJiALJR3Stot8cta+SUpXJizQmQxzbUjMQIBBClnO3BPzGS96ERjubTvLMimJxWx2Z0NzdEEGM0A
eUuTte18k8xIIhOvImNRx4WUcDaMwl94j+LE9jiIOqrw7AKR0DIAAZMNI4JZBnGz0wRqTzV9tzTS
9r1gcgFafxHQa7nAA/Y7TVV9ODdpvmGOfSY9O2K/zq4fhVPQlWubByOI6C0k5qduD65/faZUbi0M
eEM1C55fMowwnzFQqSaqPe8lIj/hdaV8LF8TY6imdIEAlHH5ex+FVUn9BxpPyOcW1XTkKxIZcNAb
bfVpFNYEU96Xx6SEWLrw+97dY23BplBiVr9Gj3HtRCkMb1FaiymH9ts030NPtv6BhuzGfIB0T8pz
h4AvM4zTkB6XohGhQxuVe9o+tRJknL0JR5CM/5UK7x61wVJKmo8DDGRz+pPK83dj2Em/ZKNVhgfF
IgGOMa2q021xfoSA+qpKfJPUCL3JHwuzbltRty7n0Jii+S+JzT6qoYlRfkvvL2Jt0C/C0QryGKrm
quW4Ew7mjgF2VtGciXWNNg858gB/5s+NyirjoP0iV4h5lfgjpzNzHtSvgGj5+rITvckM+kL2EtK8
y4LKw9KQtIFB4C40J6beRqADHL724EL6R1/2/lyjjupfbQ0acpWAvmDjbezz3D242eCJugo+cqt0
R7YXMYM+dwLY28vvoSXKOAgodh2ksuKIIfss4pzNtgq1gF7BLhuB7soGYelRn9RTXZN14sE5oB0W
MkTOuFNyrPhn/2BIXhBRgtPqowyBdUtp4wWvv4xRHfTaXaetEq8MCZTCPmCLQPV0jhjDWaXplEw4
JuP580pcgzIUykPW1sPoln6YNYVdhEYpk2Rje8Rik5YCMTZo1y0ypsucIia5voS0d5ndyqttruga
EwK0HX19OrfxIpJhUHBDV/lS6XLs9pqRvLJGZSd5NaIK25kCarVNne+iZnkab4B+c7uwVl7FGmvf
DOO2dH1U+jji9sKo4x1Hk0lMlK73tgiMExFFkUn71K+KhCtYwlKhfoaCgAx/hruTopb7dpd0RO8N
rfbgXE+6/PgGp9gDWg1jH/TmQwnidpLWMgZwd4W+sWUW9uWnlSNXIDXQiUMJlMCzZ/lAyOHycuWC
M7WkIc7vV81IRqHfRcCa0Reya5a98bb/muH1fg9j4RdqXmo+l9YglmMMr+wYzhHgG2xj0EE6J+57
XayUx+7y6dsSFxqdlTcMGnAvNv4mBVDPrzD79t6iCcKIXOUcMH4DEr1SVF1p27XEXr73cuIXsse3
gX3j8TNHdU6L556FR5nOBh2MGLMrNIOIvm7sRidkVFISmkZU7th0C71lN8TkYeXUTuQWRzjHq9Of
17OC1lkpEQp0PJJ7cXX0f6+oDo8WXnXBB9pXK1TvaepSyuLhGLZQuT8PlqBr5T89IMTlWu9S/gh5
nyX7pTPMvUkPTuhSjXiQtDosk8CWUvFEVU2pvvId01PPWwZU0DUQehniU6vEUKjb8fw+RrgJc2HG
QuqoOYH1KQudhDsn92a5hKi/4qwFLpf/yPPQlk8FPetnHwMcBglshPg7hMqEI82X/LKPwyNnNxlp
W3VtSenBjj6N6PIwQ0/1IkEMl1BjknPoIK924IRFKNSIt3k745GsE6ZfhHCG8+RtCvWVarzaelD2
HbR6bBW9SKmBal3KjhW7KkHJZzHMc2QDECdcokJQvMTnmptpNfqI+L7YaOIVHUByHA9HRZzqIGDD
PleJNx12Ddx90nVUtayrjTiEwkN9jVtm/Oz29FqpEolwcSG0zVrHJ9hSjA3v6p9n/1Wee70oCXyT
sasG+CJq+VY5JIEpzMDQnMCksLRcoEb9iW7jCViGJ5kewobxMBzh3PNr4pdO8mf+avaCzg4r5viU
ZS+0MF8x+mDtiKJYn8SF8q6JqewZ3ngUiOlRDCWMeAAcsFl5dcDePH3cOdZfarg4KRTX/N0HNbOx
aL3XZobHCktpRvdq2aB05NCebn2gw7cQmnq/Kj4c0IPYhYtxvc4VgY3fLW+K/eOxLD8q24vEfo1c
3njVPjyVcMbqwrLUjj4WOvypg2mHToBSHkZROZlvglC165V0N/dH2YUBKRU7s5963AxgpU6v+TuI
vHXl7ByO6EZDGTmHk7rst4BIo+EfiR/hsRxY6kqCVNcJHtDwx2Cni3ZqWpqpQz7hlksK9zADpmEa
ojA+WnpnRXpxZurXDkfPyOywfYnoRnxVLgUBoWXXVbM5II9Mck9NXPYAi3U/WsFt1/ZrhC7S6Aeu
DG2MDKPo9rEMRAp5s6X7lgyf29Hvgr61i9XhqHdvVHQSIqTU2huCX48e0a+ns2GsNg+cp1++o22q
0DhIDOSFNwFZMLo57W6xu9v6Sg2Z/xnYtJL8VkVO4ztr8eryCBZQ8CLCAnIKPxQNUqpAtMK8Uktz
er0P/kHIYobkMZCkD9rJzuml6EbrA5p8kWamZsxWNGFoCTISbX6eSKPa5RaVUHaPb0lgbbonEDwR
zZB+dCPOl1Vw9Orc47RhFKj5cqBfrEjQlXOyd/VZ1ajm46WNvOSoq1EWnMHn2DpLeFzidsJRkA83
vCeYQTJUViE3NbYNJ9V6PaKUZ4SzQH3lq7hrhvj4PKRF2EPwD3IRHwrm31wvjuf7V6Qhv/p+en6u
ngE5O3cWuvRT7ptF27eb0rQ2XnVoWO/Ut1uf93uxn/sJhZNA367ZlB4pdbPCgSDia0O6IvVXvHkj
Gj0oOMuFH40FkDetSVTmZAFki1CbDJ1AwN7C2+/G9swNLgqTWcrZ1qmSe4uNc9S7hMYxWBqOdjsJ
HJmMnPWBZaLiYNx0vDu5ezkpC1t2rPmOXlL0kKqDG1hBnHdfKLhk6L9h3WA/WAE5X60BBLuzKFun
NAovpzhPCN5+F1rqEn8CqHbdwvEusEG4fLObBOkSkg1874lAUVygyNjWu8XiakFi72fFh1s6vQn2
P+0XBQkwG+wGt0VDjrn6A2yYjuwaLWNd0CPhcK7RAOjApDbi4CAY72Np6V5pO+mrX5IeEyvRmQLu
/4aX7H75kAzR0Gdup2dUl1uTabEekGafR6nt+LWoteLuPHUH0jrTAFk8tMQ3PNJO9l9nYHqvBFEh
t6sZ6xMsk+N6LVY0mJPhytj+xppFYNoC0JbJc3kXhrZyBWBADmiYhTxSIN+WnKxJz7ehtgGYia9j
Yffq26d6PIIQyDd7U89aZeSZ7giMTcMwcDW5rfc6PN5pqmbzpcGej98vuyX/o0nUKiBQfdkuCX9l
5th5LcXlI0rgeOJjNwmb/iaKDn+w7Bmqwc2ciI2KwJD7wpCfqyLCz33VGhJFxqy+qkIoI0yfHQg8
R113r8xXL7cUb3l2kNZOdQukJA2gVF6z+u73pHuupxpQRf9xvGS0yTVzIoMQ4BJ9rj3oI0WE1mMF
EGxWRRofma7BLWWRcP0X0ASwoOJWZotMjGYDZFTVo9vPcV2uaGbO4rwtm8IUQBJNt0zRu5gN8Z5N
L3bpxe4Di8pFMr0pO8H/o1RZ6+TRsYNwU07tEYlb1Xcar7rNYPazuQscytbFs6Kn7QVfGi2eHtEc
DPHBdYWI0gMxb4JjTkb7Ib3t7gxvBg1t+niLkjksnWNsS5t9Tl9jtk6IhhHEUKFHQetEnaMyAivX
oe8Lc++9eDtZW5g5QRzdSDmoTSSjFICVvcvter+rDIrlCM4kER7Des1VnYZGXACtUosjeI/Be6wC
WDiVjhDi8042sD3E1rgRxxrLhlb9tPmTNcKTrNAiRpJdS3Vyn7/fs+i+Zx4gVeHJ1jU+bH3QNmVE
jDqgG3oFR9B5V4AFYe6zpy6q1pred8OTF2ypLmdPe2oeNZwBRny/PBE5lMtUObbvQnhykUox8X2j
iP3b4H5LpbelZKhdCWIjeilHbGj6KVG6oCRALVvNQHLPuA9EfZZfmSuC5dmTIDIQTsexcrDdpvbs
2x995G5USxGltQ3sI8w65Qn6PeoQVivAjblnYj8pErL1u0Mb
`pragma protect end_protected


endmodule
