`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
nYvLUhHhHZon/o3z0C/MVyNrDfXtbzXtl9mqu4zDU7fhnmL4e9tK/tHqvSFnPwyDkNgUcBMPbjKM
2ilkuJi56XTEGlFyi2WPKb87bQRjXHD6H2Je3QpGAGKl7iysx1A3JRvOGluv0YFQwp4vLBIO/pqZ
5pb8L7J5JNAgNXtPpV/Gozh6l5mF+dvg7IJuZn/WcLTQOCRaEomF/UwrRRyhqBdkgACtDjMeRlfP
6Zd1NjAB2abwtEq+FU866//CkNy6oBbizDPF3gqwdes8NN+52jIR0Evz08nzJTC2mVKv32u4s8P5
Iy97Rk95AdeR6StSeau70ARlEERvNG9EDMBSIg==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
EUp+OTZ3QzUVVUF/vGAxHhJ772LJHZMyga+iTVpGDCkY11qKMt6ogKh/zE2zqTNc8aTSaZGnVsc9
AHLKGS/Tuo63F0vl7ewP43vPtms2kN3JInGrwIZqXGZowP/93PFkzkO4FVrmQQKWfhErqlTIPt1M
sNl4QutfnAvaNTQQ+Ms=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
mVMyRAgHVldEOtDusIK1Tt6+0yoa634d0Hgv3JicmtHatFY1jmtLz85hGUyTr4UDn86b5lMRw1As
Q9bj7cNoVRTKjAap9Xk+B74SYiuRR7V7+uBLCw1om/txd8wkDCu8VvZYsTyM/x7m2pEDvzmUFqIg
RcAyvP38uovqNI/o5P0=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3056)
`pragma protect data_block
567M7fXAqXCI6VVHv601eoeiJpZA9e5cs9N8rqca6WZt8qjkC2Vx7jY8lui91iljMXyrQFd4FjS/
Q/obpp1teArmM2ljUNm3/ow3otDp3fLanWBs9D7Oo+3PdT9ssBA69oGeO4Yxpi+6KLmgFpEN76sY
/Ox/feqAMr/LxuVA5E5bNAMdMsovrHmPZI1Ddz1maBpZqr0eRO8D0Mv2hrTr68ZNHb7WDKqldHMd
FpU1kMsxjN+exgoms5PrE3p/BPASljXnyv9/kmk7LA5p2FVMvp7SUWt2GwczJbvzXT9Aq87t9OLB
MKRvT+9YNufZJTqSsBqEB+bzptzbqw10y/gYj0I/AO/A8eWzbMM2L7/w2zBZFS+CzWF5nT32xbWd
8ByC+hF2uyK+fKtTElVfUEp760bQUynxZ2ovutMbLDabDRsraC922W8czkYaK4VnuJltgQsOrn9s
7fzLp13nrvQeyVPtocFPIy3YrlUj84CjKO89r+2k7mZEue6VZJsLV/B+WT4K5Ty9AZ/Gg3AIn9Yi
X458jsHc7CTx/FiEwzniZM5aHAqIpVsLf/UlHyHkhuXUiou21069+hw1nNeEMrq9/AQv+Sm2yEGV
8hYsFH2GrEFtV6t0A3spXnogP2IQVz2VXymwpI6j0fdqx0LX1Og/WhrjdKB03PC0/yl4v2Fitz6A
Fxp2nyGs+Tr+WXXYlKc9b4w3CG2WHaezBbbZav3F/IfTYKvnLwqJO5pOg/4tkj65PIOKfXrWY0oB
sk4NrqBfhpm5RMEvsU/iLtZ1fAerYNCEypIdDw1RAJlA/Xz+11XP/kcR6c9a3Aky8dOY1fnP+hEH
tbThU2yVBDJEBiqY/jS4pVyVeOuZcadavr18ohWdN8oiEMr42oS9Jv64+nj3/EjJsOBFgzwvzsxX
R2Ihc14Jsruc0Cylj792WA1tiwjUbuYegFnVg+nh9S2YoUxdPn+Yu0DM9xnnRJhLSbRGUO5caoDM
vF1e115LGcBxob6NNEVqiYuKMrLLMw3HKbxol7nQeXyKhfsfOUh/5jaHcV1Sot55dn5ramOxJ0Kj
80v4xT6Znjaqi/yvDyHvEBHPj/SAALh0I7jHOhPndnJrclfBJzLxZfq//wcjTl//ln7Nl07hTYqI
LiDu0qDHkMLWSU9K5EIHHSxOp/RYK+SH3p2kJAnAwrMnGU0QhDZDpabE1Hqu2LM+08Uyp+0ceECe
KuAsUFpHfRKYeTNMcs0fJ9n/Uf80hC2wejJVqgaefYG8583OEqT4rH1Rgl7UGrXBg7rRSfdIvwKg
vgd2lG63YF1ejVVcJ57us3wTDm4eD7jVz6Vx/Vil3ScbbYPu1Vb7Sc+HAK6Z7ZrvGQHmbuxH313c
3uFNUB7+RIzqKzIjKeAEUNpVsWIj1Xh4Eiy76Mh+OLtf1H38roWnwinYOx3gQIy8xCToNx5p+NIY
ZZnMVko9jrcknRs/hy1wwEKV7E5G+JNKwo6uGLSwKgnxpuwrWhL0esCBxWriLiIwlcSaTiqcQMMW
THJo3rgW67SiawI/WwJM27OBBkbklwT0feYq0xzXrD/VKOElR1GlNTJVIAet0oeU3LLAEekq0l+5
Q7Hkp0UT+l5armqJoNz3P5cR3GfW+Va5jlVbklC09w2Oi/iOoQNo/1WPhSyMMOWYvEdu0MMVTyCE
zyXnw2a5e5DImEMdPa4RQCQhFeXkm/Pxwtsv8HPtzumF2ir400N85gcF32tQQJfFf20swZCGa+JM
StDyB3cvYCl8jJ2vP5uys3jx5a0vTWxmgQghx5RANzeSXc+9dR+jv0TatWKD/0Xc9T5d/OQnIMTn
9ARCZYcm4iPdwAo2mtr3r1ZHl/ZKu5u6DKGrFmsa6zJ7gf/YiG5J7yBRZmHYlyVVyKqBleN6nldE
ba5079u+Cde+Wy/m9SQ8y2e9mRHdbHhJaU7k/xX6pPArvAO0DjduvI4RsNatJyHFlmePhe/sI04h
gpdjbvdJBLakq09KGGVVsdJ89OYNHJsdoxaApZM6UTGxCJ/huoQZqpalpOqp4WXnHrCI7Ac82inB
8tArlQXR41O+xTbf/C2yp+BbzUQGMTOjEFABobjLQESCbUQqTtkUf7MqQ518Vlsvxb0VGTnKMzk0
zfUsCuePl6BhY5g3GewSMJmVbUVVHX6an9GHofIIpN1WYVSlbB2J8P1NTFxyDwYj2dMfF3/pNeSI
pCZkS5vNp9qvQsYqXQY7T2N6RJzFSYf3MMeWbxo9w2zoNPo5KNoLGiMT4zbGO6Y+IPAJK73zshHh
ErXXNOsg/uZktXaDzRsZtKXkIGX8WNPVycRO62l07OYY40/MGoVI4fKsOvarQyewibpMJRK5NHqN
z+4nENz+7DVWPjIL98povO/ZFs/His8oyN1KXzz4XlV/pEr/Y7yl7KYK93Ne8IO1YR0uai8/4aRq
HnSYHPJbGjChZBuVmM5JdV7w7cH3euLAgSCvsU3qWTyrwTp32Qni3NS9LKuVdajpAQh5VEPv9Guw
pGjl3ZRq/eTyEa+kEC0xMBtJono9c9mSHGfpsoNln7LgjuzAeWpLYdJ9xf92XN1rGIHFQCCGKl+b
5pGG50OC5uUsqbSe9sXfNl1+jScoq4OKDyY3blgm7U8h6woNUJKbQbRDLvkQb5r0MwZTyWlctmlG
D+0qbFRDxR+5gUtn2uUxoL/Ou97aGBwRjNZ7al4OBIMMc4Kda45JQc/rm+HW+muYUXYa6HTxhLhh
FiKZaB3MXQijsidGgIc/3u8tlkdN2mJlN4jHOlJxFYeCmoIo/SiEZYdChaXHFbrbdKqG4uihMcX0
mCI/DNWnbq8lTYPv7Dmz9Af/HU0cHhGLnsZqctVkY4vYuBv3WyrqOKgm6H+1hlzjRsVrudX8sQbd
aQc6PruCOvDnneqepAVza9UaYc2Ewz8Ojzd/tDEBXPM99DMQYwFDq/O0ISyQXG27rk1CZSkVbz2d
rUjVRhFLeB82ty1yUv7h6b9cKWffHID8bG8kwUyxis6FE3GptSeFecvIDH5BCWThEqfPV1BPf5k6
6ZOt7nnj0OuexhoOxnKlRg8xHzYyBmXO+/UspqThXAIcrYM7x+lKmFz5Rjz8obazRLHBmzfg5eaW
TZge+6QF0efnkaxY+CWi+Pdb+vcKAHkguF73GyjQxMuq9JEGsqz01mVVdMyOv0LHpuTQ5I349Ai/
1TCbB9Z+E0q0+Zziy9TFRO20fSy76zg38+o88nE6AvTLy5VY4P3NvRlpxYTo61RcIaMEvaxt7G3N
cwk7Qm7bg1PQwvCU4DxoMYMzu9ozLso85F16qfb8CqmakYaS2cCOgCmytZmkYner4OaWIjAUomFF
auRhKb6eh20B5P230fTzPBMU302yfYUSlegzVoYkM1QDCEuld0vcbIBRmFXYDseX+zcRTtKORN8X
rZkQAIQyJ+q7Qda6XwuSBYiCrGjY5sECqVMSXs7YmXhTWK1yny/ScOxnVWcA2HsvFfT3RSyR1YqI
r4mmyjdXJbFE2q0YAH+NYbEgP/lDSuZuD1rG9WzNtV7prTOEtGmpLmaIM6uN6+0Tn9h3hNbAfg7r
5C5pVyOHMbYZ+cpiAmau1Eqz6oCnPRf359JS5xytci9aPeRQGRNEL0sPI1mNxENrAQ7UYwmzY68A
F9LD2UiLFjHKgetdfY/t+7dMQMb+BEAKlDF0vQ+m7GxstXICAFnXce7nrEELWdbKJUa0Unid7SuI
K3wnoqFp+q3pA/ZrGjnOM53l5UmECouVJ4Ui16hzi9BOf2T2Q9RO35n8jHa/AIr2tfWcpJ6aOS6C
XrSWjmabQ+PXYLNIWB4exTTSBIFJHlLI2p74YMXnzNe6GUk/8Enp8fcAcC7bdVolegq1710uaAxn
6mGUNjIeTByO6JNPEKIPNKd3zofWtW0pABepSsGD8gBaMleZjdHP1uSUV1HLY4r+sOuIUH2WpE/d
FhbltsnOLwsRLoTeiw3yz/CxDKjM4hqf6/AbPV3uz+JZ/R9883FZwyyMzdc3+J9QKrNZp+yHn3An
/V/tJaYvwKBSgQMRJeBq2CrJvCHAWqxv13/ddRqczA6GRYg=
`pragma protect end_protected
