`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
TOKqyHER2xsCA6Tn5KAT4vXwlCevyP4WOTyY0dr2h5CsMMZYtKsnLH5odvqUetRpZi6m6mOae1+z
aQnZBjMwGpW0b5DDGr+2Vie4iz6kFjST1UF9F73jhRFPM2cwGpENJrBpId/rGgnbN+lvs0RVLaql
Sg8r/Tz+mfjc7Cr4Kp9l+1OOU7V6sC48PvxZ2YgU8HuGOGMYZQXKU8hQJNyidzYBL5XTq/iwDDN1
uH6WLcen/9sZ7YO9S3Cl3PGEaAcG+4j6reN8pMnkg6APsR1x46zCd3YmkDRO3ZVSY5lPgVJWu3bT
SgVHn6o9tfPbX+QX9VFrKqc10V6d6Ih8yXDNyw==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
Tao2K4374vPiUEEO9W9TTxyLbyk5Zxyj7yOQ+jQ0ivrJZDSCZbHd6ZWj9tMbUdTxx1cG/q4OwEoy
BkaYM3cpCNeQJxrtIqdyQGlsULOnhmLcBvVvc8Dz/Mf9OHgjgOhBboXvRP+5drChjkqiAE6IuHqF
glVXwEhI8W9pqb95Y/g=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
h9PyGesaOdKzbkZnvqidez9vrDGfQzm7VhohPAPSCMmiGwC7EmURC3MyE3UBRmbhdFnMWyqSoPZn
m0WtNXw4zU5eYHCQfBVAXEs4iYF7wGWHvL0HYg4rCIPpm7AZKf7M3Cnd25O3jRcCwMJbVSqld6yC
7KaBlmXJm8ASPfGqEI0=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3056)
`pragma protect data_block
EKcI55eMo91uDrQMiOpgUGT+rCsBiSaDqAGhvispNFcuGSd/dbDvtHExlaqCYdrg75gJVXv61aun
OX0ADxkQD2DyAYFVmC32q4VpO33H6tkOVv2qgEvaxvHDgwClltK0VsuafY+eHUgSaPXgl9FlqCnf
sYn+USnbngXP2vBuCz+RgT2wqpediXETTQXGS+F3yeO/UBKFC1LM8pYS1BQivgpZs/A6uSldLEKC
27TCU2E4FO1hI/WDKsIXRIRlmPyPkl/8vk+CcmMM41/c9WHZp94LdlfgesUTd6za5HVdaAgms5qY
tBr8HwJKGGtje76BzrJgBBDLKHo3OcLdthUJs7RZmCVVr0GuGGl7RxPrMowb77OSO3yyoxfCiNsq
1Obe2xN6O0tfAsmftj4aMqKJzcNPZBz+Kj+k6zB2XmfetVIRnPxd1JWZm/ovk4JLjcF+p115+l19
Sq7WM2fmgMQJvfVr2XjIxY+ru5eUI3UUIWnMYpj7EJRCz9E5cDCfhBc+yt/Q90519g+2SeZtWb9I
yFExpk97siNEhr3VurBBVisoetmQlyErhpo4qXBc9+24ZNnJ+3ADB5W0ki1ZQOj2wxbtn6dshicW
RpV505vd8M3UZ2VIvWr9E3dMur5JVVMJds1XRCmJrgYNvxIpWybyTqAbpdt6QG+8V44g1/APh6c2
2+6/as3kH+pnFXjvqHo2IegK7LjJKK9OAEpyUe1uHi/EsrYPFvrhC9VK6qoijIQRcwUFbB1YJQ9d
f2qoO53NrzjRBWcKldnRR75bcLtBXoLxyu/sVQWxAAm5hM2UOHuEjoTl1DS+4HEG9yTBL0OVbtKY
D/xioHRk8CtRZKu2m77gNW2HionEk8Wzyf0qudeawWxjprlb6X2D512L72JBmORWYdVhDeFfQu4O
2EWxdIR99GiDZX7XiQ6spGwSTZKllA6KHmdAEkRu+xW1BG/L0R/J35eiq8YT3A33/XrS8eNxmOO7
Ay+3fMmR2bW0VKthv7GXE3EF3+t77zNSi5yGRb8JTK0+eD05aDM7cptdw2KgmNVpxQ0cDMrE0NW+
0yFXpJ33M2olSj1JWL4dcPIXzPCbNDdZwEFB0xIQoECgtS3HXlbSjptLWVw2/ahQ521AUIQwmqRV
cCNjxrCv15P2yse0PRkzdaWNk/LCgv0biOzKixsSZ+1LVMOgZrSOt+XWLisAQdxYAEEqCa08OLXs
OD8aiSsWQNOtfIXO4Gzwyk5ljOV1VumgzzCwvtaNZVahyuDbQCFGEAl5MN8GfHrAfOkH/HN5s8nk
q2TtGnx4RNSKDQqaBWmBJUniTLtAGVopsnBWAYDuvM/WaXBIJ/qXiMfeyhyD2L1T62X+ySq0nl0h
zC4V8Q1pEcHEnzM/eF3Q3XeIUP97VqSCM7tDu5UZSDJXMkd0OHP6WSO2lCT6TtoVzdwjKasyrHhu
81Dj93m5nhrrdQSiE5xUFUsHsalfslgp+zxHAwL7f231rys8w8MteZR8aKmiAm7Gy2kmUWiyGdet
VvI38ICBxRL274uz69n5Dur+b9k4XgJtBDhAl0Gn2wtl1Gl9mmnnyOocrFXvhye79TIUT5ynZn9x
D+xAzU6vY/+sj0x9un02YkgnwMO+Rbipipp9Co4+8MYA2Y8ifOeH2+hlpcdnY7SdoZWXFff+3zR4
dcb1dSlxq8ZJMQObTMTDK+FgYJCcJ1WahmgEp7gDK89QusKmyv8XvoLSfj+Q5bNsZKpBf45RSshu
nxmgwWnCKsAzvTBvKPEjyXB8xvlWjqCZDbHkARRRPbkMwiJJL+OZXxQalikfGZ1FtlBZLCNduBmL
rpv8oY7rvxev1t2q5nbdLgT0DAb3wnwLlnJeK2oUVF25KiN/+7r88xRaDaadzOwn0UUXMLpowRrq
v12vCYog+4OEv0tCjITsTE9om4nZJeeLhcSUp/RzPvQaNlysQ5BENC3qmU4sTpeP154BOslV+ye6
RpQjiterpi0N41M18SV9/VDkxD10ZhD56ajMryc8z1LWM4kCmYpzNEbozwT0TAPhHqObwSnRROPV
nOu4cZ+NuOMqnhfRrUAQ/WU8BR9yS/TEOhqzqcSS3W3l9Jl2vV8PDWJTlE4vrIIUKAtHbA9V4My2
6eZ80bQYlHuosR9dd0Nr52iKrS6wRPMUAXhKi/Avp7DOxotgEwC9Gs4YZd4gbczERG4h+RZiOqUm
j2AI/9HLSB8bEkRogdZqWqa165NED7xoVm8ncoPccSLMd7GRBGxNFgYXQSvnbzyYXz+3Swqbpl1R
M+8uVnbSVjt0cT5y97eT++xWc8udH9sNGwn9yIwI+/rZi8rdMHp4zadkM7JTLrPwURPAWFrwIiiD
j5ZeVbSUqXePfaByOQwY1X8f4yogQn8jGbGVPxbNaw0zgsWRC3kF2dkFGliLlaIFQLlrWiCNHGog
VmcqDDqaHw2OwbC52CjHNN6c01IkGI5Wbjl0vyGHO751Jd4S6NyEQvLa7nBU8d9jKM+REUpPxvQC
rY35/EnjYyIRscGvxhgcpkdAH75u1nf++vhMo7pffflITPy4TBaVeEonejmFg/rmaEQxofunxuk3
23rOh0LqXkWy0BG/Tz1ws+xZfRdruIOiOvJYwnvGrxo1ADOgiGpIBj9hpomywJGj0h+oJbappam8
KcLQW2ngtqEOXGJTswjhQf8td1fRUaMNtmFB4J3HjL79UdPbR1MFEmeU2opHElUbOfUU6IjueKVg
Jq1cAzqpIkC9B/RB/vqzRn+89ERNCECEjjvCt2oPYX2ULGBheqlM238dyeu+x8qt+BWK9CZ7fB6n
+a7kuLUm0LDmRwDorpzntLee/dt0g+ObEwukycqDYKxy38UHXauEMqyOUlFFN9A05dZK+wObdkK6
MhmaxtJH5YrHytIOuWGqUnXZobPXNB4Lw7o2z0F3qSgSXfg0zrCMDZYp3yccW3mJLmcV9ILFjpAI
klraMPwqPpOf3JmUQVoq+cjdHaOblNoVFMJRrSn3rOAXFat1NNDoX0On+2zHh0ek/NwQ8M4iLC1/
KTA+t91zxI1uLfBEN8e+/EXEG3kcJWXuSlV8XP/pMb9MjU/jCYryyo75h43T3C/bh0zwdBh/dNdd
mg3316wbqANRL5OEkil9a3K/78SX4FvJdGQFU3/ZV9U+NjE7uoOuKcvxqe4tkNdisIt4jhL03IQ5
+7Cq0jGQTbEt24wzTU4ctzlyh1dNWBqnwUMJHIL/IvhmwWB4KAfBUDI6JCMyZjS780S8iDLIYzIV
ESD/Z2XTHyylzr12Vut2FkgUKnfjdamcWouQU8TNz9uuGdKdker7NZvXCo3U+oxpHqe+64N4rZt6
Mb6tPVXBASr2uCioBeT1rHGwQg+cwCfs1LxOkTUtEVXgdyhW2h4xEojSHCrJSVCfDUu55yhmMAbG
bupCZtpH8NvUVVa/JvPa9GoIVTOaPErQz6tOLiGRf1edKm0lcwYTBcT+aNjOzWfNk4s14xP/0Vn5
I+qNMLXwE3x8pj9GngPuWvhHpn0dOKuSKUiAAQrbY7KUzmAzbQ4lZUlWZNCuF6vDHBOVgIUyUalb
vWztqWUtx/cAyLE9VK6mGZ4zzhB2HAzv/Tugw1J6Yk+ZGzNTvTofMWPhle7Z0g4LmNt0naURhxiK
Y2OjWXiq2SMTgO8AbZsAr/DnaFlC7Rnfj0ma5fqReDeLLhKr26eCL5m8vkx+NLE63CKEtItCY8Ej
mjbTY8x4c0MTqsdNdR06E6hh1bLKnV8H6ta2duOtD0M0SSBWmWEOxfVKiLTW0mVU8KOSUo/43Gq9
zKUi+XKxEkpgVG07JGkIMIX46uAb1YThfOZuWx/RKQdC2HLKRTLfEcpfqgXIJHRnV/ld57S0fhlU
AIfGn0il85FVt83dk/8qgbrvC3lSQRCtEICobPWcxbBzxQ47IjMS03LdWdH5sfEOacO8h8eJAuvh
En/2sDClCgrsl0+DkLKXc+xhlBvaOXsaYJRoGsiJfNJb5rrJx62th6wMHtJsF16V42RqRfR8zSLZ
6sRE6dnOB5Wbyoj9Dh2Rh+YQSla9ArImtKJVbW8spTte8D8=
`pragma protect end_protected
