// =============================================================================
// Copyright 2016 Amazon.com, Inc. or its affiliates.
// All Rights Reserved Worldwide.
// Amazon Confidential information
// Restricted NDA Material
// =============================================================================

//--------------------------------------------------------------------------------
// Stats interface registers
//Register MAP
// 0x00 - GPIO 0 - read/write scratchpad
// 0x04 - GPIO 1 - read/write scratchpad
// 0x08 - DDR is ready status (bit 0)
// 0x0c - DDR reset (bit 0).  Set to drive reset to the DDR core.
// 0x10 - AXI Address - AXI Address for accessing DDR core (refer to Xilinx DDR specification - pg150)
// 0x14 - AXI Data - AXI Data access for accessing DDR core.  Read or write this register
//                   to read or write the Xilinx DDR controller registers.
// 0x20 - Write Words Low - Stats, number of words written (512-bit words).  Write to clear.  note is 64-bit counter
// 0x24 - Write Words High - Note can write either register to clear entire 64-bits
// 0x28 - Read Words Low - Stats, number of read words writen (512-bit words).  Write to clear
// 0x2c - Read Words High
//
// Interrupt Status0 - bit0: AXI-Lite interrupt from DDR core (refer to Xilinx DDR specification - pg150)


//--------------------------------------------------------------------------------

module sh_ddr #( parameter DDR_A_PRESENT = 1,
                 parameter DDR_B_PRESENT = 1,
                 parameter DDR_D_PRESENT = 1)
   (

   //---------------------------
   // Main clock/reset
   //---------------------------
   input clk,
   input rst_n,

   //--------------------------
   // DDR Physical Interface
   //--------------------------

// ------------------- DDR4 x72 RDIMM 2100 Interface A ----------------------------------
    input                CLK_300M_DIMM0_DP,
    input                CLK_300M_DIMM0_DN,
    output logic         M_A_ACT_N,
    output logic[16:0]   M_A_MA,
    output logic[1:0]    M_A_BA,
    output logic[1:0]    M_A_BG,
    output logic[0:0]    M_A_CKE,
    output logic[0:0]    M_A_ODT,
    output logic[0:0]    M_A_CS_N,
    output logic[0:0]    M_A_CLK_DN,
    output logic[0:0]    M_A_CLK_DP,
    output logic         RST_DIMM_A_N,
    output logic         M_A_PAR,
    inout  [63:0]        M_A_DQ,
    inout  [7:0]         M_A_ECC,
    inout  [17:0]        M_A_DQS_DP,
    inout  [17:0]        M_A_DQS_DN,

// ------------------- DDR4 x72 RDIMM 2100 Interface B ----------------------------------
    input                CLK_300M_DIMM1_DP,
    input                CLK_300M_DIMM1_DN,
    output logic         M_B_ACT_N,
    output logic[16:0]   M_B_MA,
    output logic[1:0]    M_B_BA,
    output logic[1:0]    M_B_BG,
    output logic[0:0]    M_B_CKE,
    output logic[0:0]    M_B_ODT,
    output logic[0:0]    M_B_CS_N,
    output logic[0:0]    M_B_CLK_DN,
    output logic[0:0]    M_B_CLK_DP,
    output logic         RST_DIMM_B_N,
    output logic         M_B_PAR,
    inout  [63:0]        M_B_DQ,
    inout  [7:0]         M_B_ECC,
    inout  [17:0]        M_B_DQS_DP,
    inout  [17:0]        M_B_DQS_DN,

// ------------------- DDR4 x72 RDIMM 2100 Interface D ----------------------------------
    input                CLK_300M_DIMM3_DP,
    input                CLK_300M_DIMM3_DN,
    output logic         M_D_ACT_N,
    output logic[16:0]   M_D_MA,
    output logic[1:0]    M_D_BA,
    output logic[1:0]    M_D_BG,
    output logic[0:0]    M_D_CKE,
    output logic[0:0]    M_D_ODT,
    output logic[0:0]    M_D_CS_N,
    output logic[0:0]    M_D_CLK_DN,
    output logic[0:0]    M_D_CLK_DP,
    output logic         RST_DIMM_D_N,
    output logic         M_D_PAR,
    inout  [63:0]        M_D_DQ,
    inout  [7:0]         M_D_ECC,
    inout  [17:0]        M_D_DQS_DP,
    inout  [17:0]        M_D_DQS_DN,


   //------------------------------------------------------
   // DDR-4 Interface from CL (AXI-4)
   //------------------------------------------------------
   input[5:0] cl_sh_ddr_awid[2:0],
   input[63:0] cl_sh_ddr_awaddr[2:0],
   input[7:0] cl_sh_ddr_awlen[2:0],
   //input[10:0] cl_sh_ddr_awuser[2:0],
   input cl_sh_ddr_awvalid[2:0],
   output logic[2:0] sh_cl_ddr_awready,

   input[5:0] cl_sh_ddr_wid[2:0],
   input[511:0] cl_sh_ddr_wdata[2:0],
   input[63:0] cl_sh_ddr_wstrb[2:0],
   input[2:0] cl_sh_ddr_wlast,
   input[2:0] cl_sh_ddr_wvalid,
   output logic[2:0] sh_cl_ddr_wready,

   output logic[5:0] sh_cl_ddr_bid[2:0],
   output logic[1:0] sh_cl_ddr_bresp[2:0],
   output logic[2:0] sh_cl_ddr_bvalid,
   input[2:0] cl_sh_ddr_bready,

   input[5:0] cl_sh_ddr_arid[2:0],
   input[63:0] cl_sh_ddr_araddr[2:0],
   input[7:0] cl_sh_ddr_arlen[2:0],
   //input[10:0] cl_sh_ddr_aruser[2:0],
   input[2:0] cl_sh_ddr_arvalid,
   output logic[2:0] sh_cl_ddr_arready,

   output logic[5:0] sh_cl_ddr_rid[2:0],
   output logic[511:0] sh_cl_ddr_rdata[2:0],
   output logic[1:0] sh_cl_ddr_rresp[2:0],
   output logic[2:0] sh_cl_ddr_rlast,
   output logic[2:0] sh_cl_ddr_rvalid,
   input[2:0] cl_sh_ddr_rready,

   output logic[2:0] sh_cl_ddr_is_ready,

   input[7:0] sh_ddr_stat_addr[2:0],
   input[2:0] sh_ddr_stat_wr,
   input[2:0] sh_ddr_stat_rd,
   input[31:0] sh_ddr_stat_wdata[2:0],

   output logic[2:0] ddr_sh_stat_ack,
   output logic[31:0] ddr_sh_stat_rdata[2:0],
   output logic[7:0] ddr_sh_stat_int[2:0]
   );


`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
XgJJf7f/7Bmaam62fYnVZR8KhK1xQmp+NT8t4cRASr1tdzyNz2kd8RksEclTeSvLfZOp9z9rrCqc
i6lSc7YQ3IGyrDbkC40wPkLronBO+0yFW9jDtrKvadujm1SSHvpD1Mju/5mlLu5zs8w07Wea161i
zPlROoJKxGJfO1D3WSE+JZK0DMp8hneJXazUb7HI5FAg8f5NxFZ9uo16+6lOFgnud1W3NXJZLViA
Cz6qI3MQag76nelwmIB8XpqZfGtkEvVZgr9vFhWUDS1CfFgxBQQr/vc0q57Iz+QcOtcTk7O1cqjE
4/xOSqWFuKC1ajTal5f/3K3VNvzTjk+A3cqTwg==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
qQIT4dtpBZOt6TBOy55M5eVZZ9u8yv87mE+ZkdO6VWXB3EJZcxu5NLymAoeTMA9n5K/wOSu/r9kb
roocM2aVNsMoLT/9J/saj4U7CFOIrkpChXnACmW+/HzaKkbhnebThtWejJKES2u7/OQDcNcRsFCM
jQ4FaBwVb8JF9VbKEHg=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
BoWrt6RjW1aRw1owomYdhgdK2ybRUh3sxoXfanvtV7FNufbcx3cetHssHhxDaX1wQIeVaIn6VGdr
ecy9aFAVwiO37QA0NWw3PnSnsZVVsaUJ5wNz+xqucCF5wwxSI2iWusgXm/iJa1XOoOX+dP/Wdwdf
5GxTuCmhZ/X2JvVABjk=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 35136)
`pragma protect data_block
/lksjp9ShwBiu0ome64CBEK8rWI/qunh2rON0xRNBulYZYJaLdc8CsFOScDgaJGd8keFVo+znLbH
yJ9SFoQLw+5NFOlrhwZpbFcLHH9fytEFk5/3WS0+3G6ykZ5gZtREkXOnlthFUq3o5opOnxRHXaKn
dLknmH7AcezuL40wzk+/CONOz9JBes3r82oGOHMEDmK/r3s8b12ojOANeWYocjFdOD8TH0E9dndq
AxFvimUgHU7DgacoCVwIcvzpAMJiotpmj7nHZXI1vFCVEUBTtWJIompLncURQ+3IeP7nK/bv0us5
PolA4Lk0rweMwF/P7qYNlt7bBFCRvIxbCB6nX3MQJCdHyw/8Or8RhVvFWlTUkYBqO1CXlw2655Xh
IL3mUAQ+16id0Us0RajoX2Sv+sZrdhnYcQvmFkuN1Gb8nrFNR+6WbUq/u+DeQjizhbsgLiV/iHY7
23wAPYbBw9w1HYySS8ut2xpabTbTaALt31atvQeEMmsKaufgwCfvniuu7055ESxqYJKINqLSePgN
HzCiJZjuBUgVdlDaTwCPrI24gZIuEPwtYUA5+SXGcMSXU0Ycul7WrqWHJq9uUuoLfYVMeA3Xa6z4
fumMxKpFBccrdR9DLHN40D4Apk6aQOLS2BXxHahj0UbbIfJfhpCmxTbe1rgj5ozNkf/F2ivOmvlA
vrnBu0/iA7Upn3l17pslA9RDrPn5mF9m9epQ0B8xRoFezDvTk80O8hMf7F/Xd92ibM7a/wTPBje7
hqPy79l3xdLQmKfB6ytkgVPp+mWE+gJq/aKnmi+USW8yeblf1EER3B988Jox5sm6HD/wOrZjl0pL
QwnfRtHSsbED+6Rh5F2oxB4bN/vKZfeBBLmdWr+Dzm1cqWl4Isgqw8cls/UFKrttiYZne3naXoSP
X1Yddvqp6hFi5oSqUSvpD+ruA5dac7U3xoJAt/TxYxwyo1ws9O7xUIILjc3CUJy5s7S6vSZvsGHr
sjIA0iPk4K0QXdCiuzRtk9BSDZrpeqaXUo8IdgdYAXXQI5rrzW1LWI2r1OKTStdZPmAweBU1uPYd
bJ9WR/DrUxIYx6XcVf5TV+yvC0WPhrYsddY2pd5j2VH35UOyFWozFiN+cqVndtkk4J9viHYO0bl3
pNMIsYJDvTMrGDOY2DFY05OPJlHtTPyjfBfme2PC/hchjJjKXGKT9EWwmdrmqM0LhtApImfaLwd9
lJpbJ54pezR1kmp/J0+woiQNH8xN8fD2x798ZDphLF+EHLRyJ7W8niHkkphcGmZnBDAWDktz3dRg
2vTC/Tz/r5NkJ02gtL+xVxlw0kO/l0It5YtSrmbnAWz+gEDOY+1v+aHZY/2XiJURgEU4LRVhaYVZ
Uk3TRJgeEJhJAOj4olGtFqCsSNTTk37LcM74cQUKxnheviSqWnIqovBb4cXGnxSabl9qEmd1apiU
BxAWRhhveRDTRoyHFV1nZc4O6X3PVYBxhkIO/wLO7MliZVpy89pMQCbdcRgy+/+SJGGKFXWmGks8
gxt6NakKhB/Vo+/e6UqqyOuqYVFtZOYRzY7gU+J7D6yiRhT89WsVOSgpCcbX/pyaBJalKOLsdQQE
dr+uBKA4FwC1krmpqgjA1EydbK0PxdzW5mg/DetqqfTXC0LG/FOU50kaUTmqJiyQmVCOpyoeLg9t
VhIipeoIjMfTuS5NXnu3ApCDtYa+viDiXbo/BKSNUCtn5bIXlhU/vz8jhdodg3VzOsGsUuRkRg+c
lTYBFBSBVtWmCOGxR1PwVpRMtcEoKd25RBrScbJsp9Xl/7vB4U8D8ES7umGRYeYi5myY4j6P3Pr2
FbqilNcjF2HhLRkDzKARhgd9ggpAb92hBzEeF7eX3nJS5ZrVOI29O1ZbDEsU7f57teA9sOEqVmC5
OsqnPyJp/JOHlqBFKmhXAAD6irneQGhLy/Nfl9L9HgRUac6lBJ95whFqE4Ys3vg2i+pidUPJxDNH
ifhZFyCch8NFYI6vK1E+oSEHHSPpWcP2RXpqbg3UnipXubd4Fe+PDRM6/kVfQ6Bai9kjBxm1y30z
DGcMCJT14Xrqs6FivK4A988LjhHhtUsHEQzpdTUhYaQgAWGKElHSe6/cmqUeQxnGT/Zh3e0Ci1ik
IaVoM7w8XVtHKzpU7cQEbwvC/H/sNbAaofzCD9gcWcSiv3Yod8N6q2aLmp9Z2EbENc96UgtUcrQy
ks+ZxMBz0WY3RWuvOeGysEnK5hB7fmVlnxBXpxZJk/p8DDVIrWD/PB27j409MwgFSNnIjO9tGLqu
NXDpD3cWY7dOw9wtbQFuzIZzeSYJqBLRIxtGARNqwa6pqoiAHA1sMrxh8vl52QQXxSv/At+L3OFO
Zu80d/D/o+NTVlTxaCSzZU91J/2fF1/PollSvF8OYJr/WHiEJgdFji1y7+nQ1lVzsyoQz0wT9QaJ
gf7c+q2HfSfOcetUrh8i/0rKy1dbBIqdOqUNedMyMfyGs9Hb6fAt+Zh0NioQ8ioIKBjwmzalpDMi
EAdN2L2oupdfwWXMBl1EV7CIvx8lefbFrufzLHCNcdqIIwtkMqaexIquCSAIxsOTTObGhzg/+3wi
y1Pf+bV0Lo6hFlzR+Wc6pXj4UkwwwsMCWl3FC08vYtSmzXNwUbYWA8hPg/KjsnMH0WhcTXn4mRay
ZEZrCJJrYQo6ZXD6pXSJtwxCFQBKfvSP8u3TUI1VOIWa9sOqEy98oqLAB6pUTsb8qdh4k6xCoPfc
1TFxCfruTfLFDaKHWMQI+sfwDgD559KefmkPq8nXKYXBP/LSbpTuq0JwqKo4sz4AFO9vvXdz6xVl
s2NqXZnZE1UeA5Nu8GWIpgADbA6U35J8MnRn2JCQCxSxqwQtd8pNLrufOo2ByDIMvNT3OMu461F8
jP8XmtAcGMSenT36Sim0gVUQZf2Zy6L+NZU8w8L2av8UvrDXrdts9oC06ZXpv2P/pj6dyFbK2VIW
bgAupSrcJs8/pVPFIUUjSRZde1JGgQJW8R2QiEaVB7ix7tFXW4QobAtKSiCwAWvkoywWvvFewtWI
97udy7ZmfTngJFJsUkF8Qz1WtHJBzOAhSPHq3beYVUUo8iXQCxV6xZG53NuqJSmOlVVxAAFaJpP+
QvLjya03o+nRffvILeSHdNIc8PIc4hgjbY2uxxRfT/pSUAwJy0qxUULSJtDULLK5MaSAxsQot9H7
dFr/FujLJULbpz7cvlTjowt4sXKZoYM+bKZbak7G5Ie/oXvx75zT8K+Tm666CeTmYKWFN/H72uGN
3hLBZFe+X+l+nWKV0fQGRnaQv8wJzk95dR9Jk9BqQdSwWeWnhJj4nz/bGvkXsvRXWwrkQtXnGf6y
UvrXAxk3WXSS8MCRfFr7a8ACUgG9ioo89YWALYoqCceo8tM2nlpoyRoIveWTzpis3gVr0ZCCR0IE
WhX2Jk5tFlQ128JGuVSASR7fhK240B1vIufof72bPhw5LKF30AiBEDSHWFN1YXuxlHcfs4Sop95U
Go4cxUKroCFkfXUtxRO/PA9o0xM19EYLxtqFMnr1Z3S7H7Ujgl8ZSftCvGrJmKD0BKTwuYt/+Ycv
Hh6ttz0fZts10ldP0PeYd3gVB9QCVaBHaHsJJUTLnS+Hm9mp8cb78h1L9PlUDQyeVfkikLUQe7xA
gF7AvPYCQMmNLBcyQOHj9UC6p+MgL6IG+vXfDPsmV0WFTtiAtspNE37zOBpH81zpv37bm0mqSip/
YivTMmCtuUUfy0I2GVFaZgAM1DlYwH/VQMzkZlRnl7uUJ5OpEK/KAzyzGcowhMhYO7nk7M+y3V2a
iJtNm3ZeOJTnwD8aG/ix5VJHgpfcH3j0scAsGl/hpVr094CuggnuXyuYQx5rg0pdg+6VaBwURetH
i+zXRVsfJ375IAKk4CqzqGZs8V89sfnD/8QqvbrBl0wo9PH3WSFe6YP1NhNuL3RhIGD22NloThs5
Ax6UsLVLx0yRc4jLafUs0nrVk6sxiYaEsEUgGrsYMZwKv79/SCTo06xujZgow+9OrK0lWpFzgr1x
5u/YoLf1VEycMNyYzlNol1KDHgAAdN0jcYb4iU5byRLBIhIAO4/k3Nreh5sqVRFXuY8umRMs3B/q
dyJR2zSMD6Z79OrcaJ5DzHfTLLvU/a2GasFXzKKc8Q53PPcKBM904F2KsXwi5PIzDKma1E22Db4o
00PXxi5wemZJuE62y2aTqLMLCUYIIoGk0nBf9SeM6VNN8ep477kKd/Jj405If30L/nQZcStR18mY
OnZNxZkkR4pC4geSSbp0wqgMvRVIRH9FO0CcpI1rYo2NoYv65KXypvFifemPoVIx+sakzZKMXFHU
86xmzSYChos2blSbmiuPB9bp1bo+mauxVot76KKqDKSyOUrK7a0a4UI3VZMKapaZVP6TefsmfXu6
tY8qiTfRiTO9DS819uKdOlgO7NraS78JEU0fqXkKPDx6Bc1DYwtiFb2Wp8aVI/w16oHF/w7y35+t
ClBmbIWEtGOL9/+ooVbyTFhbGKHx1QpvAey63o3kz0GFsLa1nrHgTy28EskhjLVbFhUAtKnn0tnF
Xc4hYapasMtCPZSM2ri39+diBGgAq1x/3cxjptlfeFji1W0+eNBJAyfwTFlT2MMR9hYfwS6pg/hO
+sQist7UKBTjbh6+7Mgi3gyy8xH6GXhyFlcNjR9IwqaPqjBpYSWmMFw+XGg+wKF+Bl2OJXWowvE/
G8hvsGiJOCLXOiGF7SMviFO55w+IoDSykDKIE9OUOIKPbtbC5Thgw9bEf6TBvUzGjfB7HV/8GTf3
JhsimCJpx5tRPmYNwKZyqJnbuUupYZb4jNFFYHcPMzd2YcKcXBZTT+oMA2nI/+dj5aLL18RXKq9m
z4juPa3MXRwydiAJVipuuNT+/SiYKB/lNLod74bqeb3hEoi/vRxnyEICx/mf+eUjfcbenxBLaxFp
/fxRANUf+cXifDOleGsI/h22f1uWPgHBEI3y/fsM0/Y/4HEC3eSaU78tj293RWeuU525nUm/zhGr
770uqov+tehxHHqmaXM/S4o8mLzNm8yOE6c3J5WjQQRlm9gPNU2B7R8gFm+gAi1fDAWB28aES/4d
MyC/ZAEDeeyxA1CJM998qrGE32tZh3PEsMNsYvQH/YkmrJxXKAsw5j5hynvomx0wKZ9KHuxAGs/P
Gc9Ftft38Zm/TScB+iOnNkXzxYbRhivpGtEnkyO33GW/zkzGBsuv6kHttSgVKo87MXJw6Wc7JskV
zVvxfgYUYlu7mJbLujlmRJTJg3gH3y9W978Vi0XgGM7yYIW5/7ketJU8wc9XTYWZI9RDjuq4Lrh3
5u45cmw/hZZ0aw0Gl2F37hKrOf8agKzG07EniXv9t1gMjU6xpYkLd0vIZ7r8DZPNaK1NAFVZMilg
8AC2MctOKPYwJGy5JvPHHVc7XxEdvrxFhmNMIDon+fBXuH5TpY0mai3bVUraPUcHvXsv8BqE9Gkp
yF5MjQkXU5r7rzh/FHtmLA9XlP+JsaioSlqlRt9Hsf33LyVRrlTj5abG2+FKU7T+uMX65zxFEEut
WNAiI8sQr0YDWSg4zZ197CbWeVqvfehgcbcB4vz5/UwilkhSDjRmJgz7rigYBQdihR+miO4h8WVg
LxaBEgNnTnpjm0/2YjwbIbdVAZSZgUP2y6E/OcE9FgmdNABot+rj2drqgsAn9UBGR+KYOEWk6/B6
vaFG2ucdYh8/89NHZSxJrJaNbWbpnBf5Sp30mpQC4dbKBX5ZY4Dzgfvj3KzyorM8Y9+hJToeCsJG
x5eaLhUr/tAv8oaXwzIyo/7of99ohQwJtnkTndlxshl05qA4w3eod7ATBmepAbb/cu/161ZL8YHd
EgPYuhro7RJ0dvNPT9f0j6n/O11zQLnx8/WjiYMiB2LH3kCbJRhwDRhkX3vUMfhpkYHl7CiImBou
yibgnC+6ZTyepFUAhH9pdMaoYkhnJphLUw/N0AHdUkQCUhXBfX9pmh6sKLv9r5Qi/xUMbOKF83mc
u4pVKVi1cpvGbvcs6xk9IWh37148CN4Edp7F6Xyx6e17LXHRvakItYP60cilEvPU19uODlRCQf8B
pdqJVtI+TyLARK/b3s2EcP039OJO8GWEAoXO7OUgcFgPNc6z+9PAEYHtqsSsZxYcLcXrlSJlht0g
R4CyOGeZCeATP+edtqF6l53+zmWSAaVjCrwNcWVzy4Bb8gzegV+GvZ6IAF4ZJsvaHvH8UehnCBm8
eM82WIyWea/66plKydj53GeSQ+bhRO/njt09eD12NpjwBcaFwYABc5RM9ZZ0tImq3k2bQpqGphtP
zTkRIXn/zgnS6o5j1yXikrD8HtcfuU+VKg7yUK/zltgYxj8PjIJHJqRmt3AUkK8RczrbESSrjOcd
qFKutCwlTvgAAdRoRmksdFgdfHGbMT2JFQBi+2INdwUrKNkrfMEMIBjIXVZrgRHuKn31ZKTdMSEb
T+Xjwppc66ZBjBN3MPpMO0bTEyzHuJgV2v2//CFKZEBxHoLXaxynwyHEHez1ldJIqPGo3DS2cnYZ
t3k8/pkqv473crVScZXm3gjpaq9WRerXPo6ibdcDQBFw4JDVkm59t3eiKjJBX1aY/ADw8vnAHnNC
Tpk2Od6Jm3KitrIC54t3pY53g4iDWC6kTH1wYfhQDPvwu0qBokp3CbUV2l/ySjgf8huBaVKjWFgy
MQFJIzrsg8CBvW1UiGATuOS5/fpOzDZ+4BDm8alHkYQBjlNQBK20zacj7lxpIiY0oiC/B5a2vdia
BeLY2tNBPo88E6k16lcxuZWY3PC5E3suFJikzlLYmacMuMN7fXvA3AXFWCYjZiu/rD295glQJwEB
4XmI1wPb6emP3aLZA2q7yIvRJGadpZgOiZPLEVubuYHne409NCBrc8dO0UYCy6jc32iv9XjAiSqy
6BOZJi0O5KAJB6AfIVSjiI3wIHIDOiqZWZJtqmZsvZlPy3Jt2BihZNonS2D1GXrUev0FImmomJT8
iGY5Nw0FBx5NWfXHT5unj2AW+0Ls+3OZJfhS9B1BZdMTlGZRyV+6uyUlWROn9uhd4wjEvGsqLQbZ
ZiLzU0RvLXBeX2tx7LNqhlVzYeoV5gYWH4CnMqNhtxsn4lBmWED2Cn5t/iWozIqe1iJ0mgq1563M
zqGufxhjr8JYsN/pcLtWIH7+x09sFpnlsG5nr6y9nerI9YiyRVc9eNPMib2M/bE/h4zJbvkWsx0B
LkHQ2Cr0AFlVZD4tCucqA+Kz65QbGd7K6XPU7VH/3Rb9b/qu7SuE8E/U9JxFvhRd4oD5eC0ZFqiM
3T7tt5ejPqkOKTWAp43wdeQo4kiUIAfshsSDaUpLQmju4O3VWmbptVXYvYT2j8orrpN7I6MEZEcS
n3UXtu1PbLKp9ARAOdu2w4KI2IcFiLOQbljdvu6nY9CMaWdGnMvwKBsK5xcdD63Lh2+M4rL4RODG
eyEuJFzhEGsoWO4vXSyuUu4vscMoIrU0PMEWbdQd6zMJGS4ZE4cP8qD+zRK/AsGmBcOlteNQWl7e
wDYsjdlVyB64vuMBhfCEaLBNvS7ubGs1OSVWA0Eb/Wq8qUHa8LDPGQX1LU3udPFKHvSv8ALDfSuM
LkAGXFe/51NkNui+DhoAR3dy3/iBFOHomzU+LxYtMpkrTVP01wpT7hunze2yFYCeKkrgoQjKkfRY
pVlWuTw4uUWacPB4mm9Y3a5f0pNCsKssQlL6heI2Lf3NuzelUVifGl5Mf1n7CD9QrWWz/OAs59ln
b9wZNiROV59FNL/NYvm9wn+wBT2UErWSHeOt0nYzaDN6+CV+YkRozYWsnoz3bkbP8o0PhOOyyDL1
OxSQsWSRRuKx2d4JcTiBgOr3QCzMUE/OgAjEIfiue8Xp09rY95hDEJSC7uH53E/l0FDaurWJ+FIU
FbNti6fLukCykM14y381egwQ/0cjxB5hfPbD1OHYxjPz07z2TDwdg6MzBjsqZTGKeiHgKgNzxF2W
HSfBVABk5Y4NqYWcMGk+kZu20HlHYFHrWrNR/O5Q7aFXw7eyiIZ5Od/wwBhwSjDWUMKXxF3Q726S
UAmquzHY+Ummn1uQRB1e4rcHPu7p96aR4+lVB2oQGISUwz9Ef3hZtPGPCeCvBzFfTCR509ACCC8c
E0ayE+6X4xvTIzDFvVA+Dc043DzdsFTX4L+ir8mWXt9q9ZE41Oku7t8RWyi4eacRbpZb2zL4CrF3
YjuXx39G753vWiLLwwHNZalEVujQNSw3mtUAWWvL2IiWYAw4YT43h53Npol7h/QCLJKb7h25YVtO
mtps3Mbm6bwZKLxtqAzlTDILMr8hKwWVqG0lLhpPWEIE6N1QfewEbl+dOiHkhYbxAjUuqYisK80e
2NNAJ2KkiKHoQZve6UWLdD/7GuVIUutoaGhGd43UwQ+3Rcp6jfrlHtuvkZtt8NDQhiIofC+gEmlg
73IYcQZqfVIBAKGek9xZ9YMcn++Gl4HSI8/4OPktNDrKhadYPD6RewXLzK2HGzDeBXPtaiJDv26T
yjlTjJnTcvTIBSuWAox9b6pEAam3tFa+FBz7sz3XVW36Qi+o66ENYdJdk6rngZ2xlkXD5uhXvUZo
GDkUCJeE8Eq9WUtZ3TCYzrjfsx+c2KmNuhb55yNWY7EPhz+m3G50upBZOXTgWN2NHmXdBl+JaE8J
pvBCj9jrEz0mvqD2I30/28TCApP4kQ6/cJGoQxJfbBrqE3bJj87tV+/LtnrP/8PV/+ZBcIGz2b2E
z6v4GvYeH+t0kbIMxmOFeoROGIz71CvtkPLNs1WDgwwPqa8cvsOFvFoWjb+uO6VgxKiD4VyXVotL
8uPkQaqlVnpGQsrXSJxp46u3nQc4C0C1Uh7ONScBJF7uGe+XKaF5sVwYKZEAkvK3Kr87Cj0jcG73
Da3Yi/ZTebD+vUrSBDMxRonQtmPqGSdosl79JBYqBHlIVoLJxjt9XF7i4tysXD+RMHaLK2QtC7+s
zDIp0S9AS8UG4EPOtuc/vnEfQe8fPRbU7ZTalxIVuqq0l6nVcLraowkDonKoEsh9v+ax7kHuzQBJ
6/6pGUvdZBt01GwVjBfd42inK3EHx/sf8lvMobHWArsGNTw4oOquBLS/Ulf//o1/BojYM9okbTsj
tAD1vUXGIPjpbrLOjxOQJlM2F9Aj8Yj2BNTr3d06ssf10UgUVxBcnBMtjp+SQ3vIwXAX9MUnLuMq
uDSE2NZIW8JIJneIMZtnJB9wnPjqicS8VILy5qlt4gseLE9dnUNSYCqnunTaGgSC4a/vmBWw+sNY
4XDTWxoT4oZg5fNQ9dEHwO0HCl9Sbb2/A8D8CdkOXI3n9/c20Ft3kPrg8H3Da6fxHSsfDv/BjN6N
CCWZmMQ7mfTlf7D7oFyKE0NTFELLgSFIfg+q3AK17s9/bTMDRcfomwoN8GLE/7U7xmsjlC/ulzE0
FerBxA5nws7bnbBKmXsnzhmumsBOWRV8bTEJr7qhegEYwW/ThbLg795HkfkRxOLcVSgBm6jp04u4
wg98E6V4JfsuEBUGiczl4WMfyrhRNUoe5lb6EJ9j8SiNHBhE/wJEHeQ05Yxtyg4Q+BGnFrHiDgyk
Cpz9mXSfN0aC/AcatJxfIgeh4WvqznGoCcxkz13o/kX/qz6YaAZ/eKLIcoFmKCJzS0JRyjw2XRYr
xgQYtirCiVgW3Oq7xFfAtFRmp63bGONjWw3ahAavNon9H/kbxhdkqQPMAwCCGOY32i/NT393YiqG
sZhqbEpwOoijtvvBvtgrg8fVohDyyNfpNnzNLSm6YGsyuUAtluk+OUxvoj8xU3dYGv0cPxNlGWrZ
sCd2oB1+HlbPdg3Rw7ikb4IQAw5GHosmrjNQFRv7GKhY2nRY264Zx8L/8W8wWooA2OgziEA011LT
o+AtfUuCu6WZ0qVj/Zb1EAZv6fnK6ihpS/8OJMNDwH/nbbFDD9+qDMDB5BQW3lWFihL+RgRxWbJV
tigS/7JR7SbAn/YCs9redbouwtucFpzkPny8EiFPvps03D5l7XgipGdUz76ptaFzthQ9HguQg9Fb
Z5Q56+Vh21jbp6pOtze0nayQsjXLq6ICWUnBp6kuDT2YRNzW62J8JQEoElhqciQvdKJR/6j1Btm8
iRDB1OCD46AkxbcbQ5y5TKoK3tZtol6DoS6qy4yokyKnR95/OtnRMs5TwpQcU+NypUkt1tT5zEEL
b2RMYRxt3osEnLdxipTpKx5VFe0dHrQXWn4g3CFPoNCfTXmSR1vakGqUbyCn5XQvCgAWwjNF0s5s
CZDiERWOvR+ogNbLnfD2iUL2W604yv8UXXru6uAKUJ9R+Ceo14kKCaDNCKZRfHdbzntfJAGL7oNk
pX8+MLmqivzf0WU4rBSyNE37AlOCbjt+R+K88jiJ0We7oO0xi6e4qpfDwyrVup/Ev7dLJ2ZIdTIg
Qun5or8DHY6DL7vZOWS4HMUPonWSDrgpnwtDQ8WpHsk7uxKhMTFD5s4TPHJpF70YYQF0w7tmuhmF
+hsXnHlydI7b+/owRUseGKvCfXXehlgVuwC+mSNXo9ZAcUqnNbkg1EbyH9y6+p2HDXsAvuXT6hwv
VEWVBlcLAomZVJPQ1DzqwKhqnHycKXXQvZU1im/+ZB/racoLNC19wQEPKG8Sf1G/YPfFUa0IkyId
wCE2Y6nQGLCfh3fveI7sH3/4Mmc8li0Xibw3NcDjcVIVXiDyZHbV1AvzrnD2tWz4+H1vwAKzNztW
CLMR5Qtvdpt2Xk8kXZST+QWoz015rQZfI8/IqS+kCsvEHr+PM/HjRSYk1pOK/9Yizo/KVnBhbGoI
gPNC8IXWgrcTCM+Fd+HQBGOgd1CAQALyVZ7RhA7eGZJ/s1wdT0DcxZoy1jYybxmbB0tUeTaR52oC
TwlhHOraLU069a8y7pREP1QPQfw0ghx86D9QskOvHa0A6ZixK4DudcoeBLAkqU5tTKF5AaPKNPyb
1lh4P4AKhffWKnIW712Re02tTwWnD5dm+7TULKY11FiypFquIKwrZ79juJMTMHjTYxdn7i2Xuk2u
N7aBQu3wu5ab1W5u0s9sRdOyOde/FNs7Gwf4yuq0/FM7Eh25eHnEDSMY0iuvIETvWechh/wn/6oy
QQ667luwJETrqHNhrL7kujrht7WQU7yQ7CKDUF5zvx3LAeXZA650uLwyz2oYnn4A6sT9VkxVZ5mJ
aQqF+usXbHczvNe8dX28M9mTzvwCSgAMNVfal4fYKz0lEOE0YvBTZzjQCzace9RT56zOLyZAFJRv
6ffR/B2Xjqq/ER5HR2dDiHdhDjqm8ei3auQXvZ0orkhb05uZkPhnlHJI0RfGe18V0m03NwWcu4sr
hv1UsPLUp1CWlHz60WxyI92rHfDC/lNdlkcFbAwUGl9FZ99shMCOZiuJ/2FvjUvauUtcDJzfN5Cn
xmycKG8RDd7qf3oLIvazwbUVWEiGKVlBA2MA4VmEs1k5rwvv/bOPEOwRWz2yoG2tAw9RNvp3faW3
JmBWy/wEjmSXwG70sGWzSWdOtfDVCP5wK3SrScas43jMwMW8kJsADiDXkkLWjXgY4q46rlotWja4
oZOYWxQEvtd2C2bR0f/K+e/thsOatafYYziFs1tkaVjQlDQFappIhFcFcpA9gu2q7Yr4DX3h3ZaF
gf92/UEKNvonPdeS4tB0oO23FPZPrUIk9dDqw+/CDfY6xC6PvqeBa1ztr/JESsCjThSPS9TiUm9P
oxvXd52cpFWSts0XQHS8260g7wsSb6G/spOyvHXruqQ0/yUFlGZHGA8HGqTNEYiKKEqaGqVpL75n
E/knpkMpnBhNZ/wDu0VmMCv7fogWcX64CDk/gPy8xcYhFaK73hn+rw4A3LMgm2/FSYBFiaLXSpwJ
kyGbHGWFKS7yNrs+A9cTJxD9yLLcHUykE6qfshRgCD5ybpeZfz7puDp2cnRwVhvhaYGXcMowQTT6
sZAy3ogsnjzoV6IB+3ZU9kazoSO3C1iLop9itFYCBo4HSYcswEqRtzRwfTW8RxrXB/tpBfkc9WQW
sz665Xw2xHd6cJYdyvqSqQs4BuRA2WK4xVgmFzZGJjSweydt6geRZlUyIyE/5AxqRgoCpudAAyPa
wFLo0g1IGZHuRSy9oociYoLmP8eWz9y5L6eHef14T6N1awoUfV7osbmmDGgEjo0M7shfkvOOfdNP
0bLlJ0vVvpabTV90rVsRD9KlGPl3GiJVxe85y+owdSfgaZETusTpMlN8KdmS5OxRGLYHI1Q2IVnD
U1SznKV/rmr+HEaWH0m9pcoAzJaOwYfHDMs4S7sslNzdZhLre4GzB3G3grAGbanbOTuvWsoDkSyF
hm1Umvm/Iqe1OdYhM495DxCCI2n9E3LAQ2PtYIKCq7eNvUk6Bo1vI5aewzfs/qjgg27j/deoNwD9
mhnUgoo/nZJ67AXnDHyWJFrDhmUbArBtlLY8h6Ql3YVkKECKAp9qXElaOzgKokoxdcszZ+S4kf+c
bV7F+4OXED5jzJn/BnCjQiczhQvlWLOouq+1Y32Ve5r54l+nWbcvkEvD/IJqyVSXgm3HT6SNJpmD
kM3egnJTHAgyGUzce4Bfxzi8HN3tcG9R8wAR5r/VTpWX1siIVrBwWlthVc385uwkfysAw6tv33E1
vwSYAx+X7VlxnG+fwKgaqPDejMgCZfQ/PMvblnCUn3tTv24dQfC3CIUoq10yBhDkTdSJMt2QElI8
9UZTRP4axDyV1xaOeK2wG6aBcY9XStuEnjXm1pvwx3rLYQwlyQoZzX7ARIwKU6d7/NUpAqBY3mVA
Bzfa3ezHyHV+OO6tQ8OGdsCnJcHpDPB5kaO34qbg/Tp8kWz3txJU/vJfjPAyBYQymXivXtx26nCB
p6e1LSfwDadaoTEGqnoD+7tyK7978Qz51tAdB+VdEx3uf+NgPyLt67WyNFgVymoo/DbzQsNH87cI
/p5ViuhPWczIhSzofvCzJv/atUoQRCnObXZgopJz0oeqKL91vimmezqF5UX1q/l94NIVmC+J0l7m
ApC6une2Qi4+YHWLc0IdKVjtIPGqJ4IZmbxaLDqgEIW6bec4WFBzECLygYl4cQdF5U983sHwbkqG
VfDy2b0Uh1DLeLfuaN/YeiY3MXbDPaLPn/7n2nQ6YRB+Ab++xJgJphZwnmWaLZrfgYWaI4cEbtk5
K0+CMhDYBUZj+1gf3rXMc7KFU40CfdbiOXWxAqLLf2N16HquqzK6HpJ9XFoYkqdQxP2F9cpOhSoh
z1wy9m9aC8b4FdfCuM/PSB3h08QS+hfabDunbkQWhlXQuJo3DgUJHkqsA1lV3qB9e6Dim5vySCdn
11jtH8fqUHfRApwxtonbqL/iSx/rBvRCxXC7geOkbY6fadIXROpjx78hDm+JZ2zKhq5ItnQ2bXe4
CIb3Xf65NZnXVdm21cPdSD4Tag5d8qgR6Dz9UkyIyIxXJPzsYrgJi39w7+TVCvnpZlWnI3AQxYa7
bPfbnRYuFY8j5wTFdq/Ekq50X7Ijs6M9dJEL3QDZsbIp9OGLQzusH5rCv5DYlmv33+eY6OTrz6mh
7zMluBUdzQucykcfHCOT5VIxve6kUHuCS+sU/KVKiXpSOudfQK1+4O2GLmZT9r/w3raSuJZjjDiH
MS0m3wriwHc8c2DwebmKqoXInGxMyoY+ke6yYwOitIdzS7IK5vF1R63yNaB1mkR0Hr8l7tLmuDdS
RljBPl9Di4T7L7N3Jhs31IW4M34rg/fQwoev+/6MSSc1KiYsek5DHzxU5Jwoa5DXvBauR187OnTA
Pc/cVHYb/vctc9AD5cZB6u8BrQKdG0OlrkF2lYMOVGmHXYCIqLT6jbI/P1GZushvlUs9uiXhumEp
TEoYW69+GtkPlqdOQUWKMqrwVxCofMMGIuqt06Jb0Ph5HOIxd0XyeUazrgqKiRzVBof9YXEwfOQA
xJ7FkOm26suOPBtC0UkTOyWbXcuHMU6PzG+RmXamXNtVOSJg0hh48TqGmjw5Y2UWXn4iPK9JqR1H
9LtjttrUK4g5U6W1D2ZdAEyGvD3wTrexbySooFq7ss9DoQ1JIAksTinK9bqRIzPdv8GpqyecXgBb
qziGcIh1TNfcRzbv+rLWerB7NwIA/Lc/BM53h1vRi8WWGD/PQeLqJCsmObO4vEcXTphvT+YeK8rJ
KVBAcKYRAA2whYUFUrifVBslZyk9Lii5qCfg9R2tijSPkTONHgNWcoQpy16OD9DEeyyDS3YhO19i
VOIuvJko48uLdjPCcvwpbazI8QUaQIqa1rp94OhIkXcMGXjQuDspcTtGG9jVD3u4LNiNDWWBbnFD
8h3m2YcZb7LzYTIF2bs4do2n/Fbpr1eOwkxgHgLhz6+oronCic714IMIStqDLyM18LfbveCBA5RD
+/v6g+AyqzRofwWtBd74OBBO9xvZUID3ErfvxC9P936WruS0VYHCJOhknioNQUGIe0fvCfBbAr6v
b6NTL+UyLC0LjBKorCf+vcXmAdQgE5lvmLNp4X25evdyH5MhocPzmus9/butzFadW9h7LYIvMBhc
yDh7XSs8pgtfPZQ0pVS9twXT3YLC+5zHYqEBWFTcH5r1Q3+BVtMHKbO8cHWLSimHoAISg0uis2m0
x6Pv1hteY4koxlxqmaCmY4DAvAeMUj4OgU3uT2Giqo9NsnQ5BWoC+wqC7VLeBly0UJ80o4NxJUhL
oigVLBkx6rfko4kAciRUTe7a2XsAlVcMbsUwhO4kgWGE6F5F5cxKnnBL3ZFp8DHPqEaF6p327DKD
RoNwcit3fyhaXlct4Qh8nf1rKHreGrv7OX/zNnBe7189KXTN/Vet/+q8CJzzPiePgv8fN60+0sgY
iQkmaNqnmQ6u2fnHK2zdofgS0O/sHXHRoRl7MA3Php5atz30ehcSyiK6CHOtAby2+P3o/bC1IpTp
2jWLpdA51iJLjhJIzq6XT1qPdv5/GnDJSbAt2WpYpdPlUkJNlQoJ7GUR+JBGGtKOMtJ6Ccu4Ahoc
6OOYpTQrZeOBfDyJkINZJlqlnYkzXy3tXAQHq+aw2/v3TD1dcq6iXOEnVwPORJpgQy+7VPbM+W2Q
JxKpDZnIljaSK6lsgjzQV66fSXpKezpFxWThKg+r2PG998qy6/FbfNiJQhbspBYoeDrmonGNmI5C
li8PZ4iwbTadYn9j9VNR6CMC1icHT8rdcb6MFunKFQrEXsH/MgXqT8l3iEQzu5ZJoDnx2jupPyi2
3NqQC2QlSJO1AXTsF7Ko23b9661Gaq1GPJ+UTGD6FsKkC+ddhKS10hDu7T/Qk4Pfh5yhNJpXiMBF
z8ROnOXBZJ1YBOS7PlH1/5v8lYl5tSfpRKis575p5QyJb80ttRHhawFu9usAw9qO3dP7DWwYUaey
0heiahYYpQQdeslhOFBQvMn+IoM/LfMgU8CTqw9qZBhO4lX3XmdrQFfKEDZlQY1v+XMtvtbUsKJz
g01HDQ7Esb7Wwmd+VOcHNqBQHWoMHYHXVrvh3FCT6qmrckWVZnkZr/RwEEkFxsZe6+xRcO+3X5qs
mdyxLY2wX7bZXflo6VSZwsiONvcvoaoWXlVeOwPAVuCb2WhlkRpViYyYSLCUbFgsI1/JOKAFUkLM
O7qxCl3+kzAInJT0Yzi4rc503cRRznPUngHj12z9Tu4TkVjK4Zy6eBtCo/nO/nuLrLNt5fYMbzDj
nOzPlxEl7l5y3CFOjAh1+V8amMMnK5VJIVgwSpYdCGSVR90AhfZNEIlejUavQ0HJ9gIfhUPRAwHF
NH5Q7KGFTwGwQChaSP7XuIdq9ueaUWJkcYO++HRqYf2QndyE6b6y7xFu4Ake99IquZEsb3gQedvS
ab2DvExi0jC+nzxq/aTpupA+hHH7v301cjCNIKm5kPAj1KLw6FqnWhJM4LxezT65nVHl9gvYSKz0
JTmn3359Dx9HXShDJoI72pit3voZqNepCTiW+5rt4VjqSaAWEW+hnXHyInwmpZVP/QVvHhIPJpS0
Lo6414q2jQJbSfeYAwwmSm7cmVqv0x8IjN6A4HeYyYqruaO9NAPSkfaxOFU8uOn9ZpSgiPg/8u9i
OS+UPFzVx9hWUcTmKjEiPcnAj1V8tpsreP6jpk6Fom00W1tboHPiNCD2WUP+dKta3hNA5+Qsi2B4
A0QW7Pr3A0e+onoI/xj2ZV/3d5lJkYxPobzvkP7lxBxMZoofeenypzpsFmEDdnraKluqjJWgOJX3
A/XoGhol1RR/NMLs7AKRGAnBLCqpRqFOBkNdtVgbGHWX/+8c/yIDCshjFDjiNHThu/vqwhllt8ly
HTu4lLKrRPlUQgB8ySKn5M2fFVuv3x9w/j3k2/BJtYLEGnb++T7m6/XccyE3+Tc6iuRXcJcx977y
u88QjFtzdbRlfvXEp1Im5+eX+StrqmS5Oij0if9waOjRZSnrMrC3O+IlxweOH1FxIm6joJOjTwQb
CiMqDJUPgVAPXUMbIO4xPaPHF+cQfw4XxjV/kZvHXaRDMBrDbuJml6ZT3YHNam0H1xByNMpmeaF+
ahuTBSFC/YQH/xOhy5uqRQN60UhuuVH3uCMnYzId2sF/GUE+dslQtVc8ylK96wYEd5d2UZZXaUZb
QUyK9i2VPOrbZ1tTO2jojViGwuGvM5MRUYAnWSlx1CZEJ2AXqdyQmRhXyoV2eTbmeqTkcAXYAbFh
WtCAyYvkjlLi8F7Um2GAqtQHLmVIy37gIIk0Tjc6GeyrRQOsC/kBdnXChT9zZ+wlHmTp8g9l/0e0
5p8lkKtwQeHPCKohI+2rjsAITSWJpQzT1kvPNVyEFhD4Q6UhGQuEGCaOrbnGUivv6A/qS6Hmuy8/
/E/lDH5nXpy/jjsUX1bIeU55ezRf9VT81w1cQC4BSFWNl/t9mzG1eQDx8x4h+5wJ24AEyQfh3Uvd
Q/yz8w11jxRno4NwjEd0PC5Ter1yHsyOk019e4cU7XdW26hQKtQ+XM+ZGXvPRhm2DpM8qTBPtv7z
uQHhxJ2cgTh/2O3A/EAkWlJdHXn/4fpoIzyRwfHcYEjn4XLEPQx88NhV4SwdHgeMISdKMa813JEe
4c6/AP+COc/XOxSNuhYo3RTlsn35GHMznA5Ud5h84PwFFENLqMg2kWjpy2LTy3+/blt72NoVlcrs
Mqq5kcwpsKDt86n7iJvlKEEciFWCbyzXmetxIgVvR0P/7zhSCVcCoJtMpu0nbghhhv9cLaQc526W
F7wJ2wFTE509fmolS7RPM2miTTVv2H0euPLhVJlvCQPsY/zh33HyqVpaMPWnNXi76IHURhMT8PUu
Na8LoRGY20YgyXp/K8wLsuAcSUEI5WxqM1A979uF5Ir5RFBW7rYrMzzzuuKRYDtiCxFZe7h/bBF0
ZaDmFGQtuLWGkiJpgahiObIwEy14hq/uv9TNEyPynQsAeOVecO4AnhPRq0v36182KQTQRffMGypC
RZInGt6FEDE/rZtdB8vAkTfrrIR2fN44JfuCCfmc2e2chdnfQlf42XqHR24m2RjGPobxeoRRtaBs
F2hEMRTn76nmsZtlhaTXmLOK4V6fSK98SzLeI7QWdowp77I6wNACDJSqplHgGCBnj6RFCz21NHFW
x2+3pGpndU762/x/uQsUp+luXBZSZ7UpyQUDo6Ja+s0L2+Z1zXU8QfMIvCqIY5fAPyuzLzp7Mafx
7BajjGiAOkEX2p63YlsXp5ISOvwE2Sb+tbtl8qfBvj+2O9nR1Uiwhn47c+FVTpuRrr80zYDUOY1X
s96nVPJI36ln6EHwyWFYjTyOHIQIwArFcxpvAMPCFhaeL0dCLegCRRdvn12xWoIAUar/tw5YbMbf
0ylEFRQhRT1r84rRwtO34tDo2FezprS3b1ezCFRe3C9rZuUae/aqTmZp0hNUJQRJa3k0YPDyVh3l
y7FDx6ElD+pt5M8TQkbXDWOVijriHy1dub1DO4C/KwcZAowl38lXslASk+Vi6VjvovhxTp8ksR95
7+abv31owxKKn5xIXb0SUZ3Ixmne4d080svylHQbGYc+txjKdAc9RrHWCcR8zYlG6sAO9uy+clme
xMHnK45Q1xzaAPT+Hd5uvlNyC7DPD0xCTcF40ZAzuoxhAjJgKRlDzvdHvj5EoR4LBCfyJlNSPxR/
ur9x1jztxgVeSJVFQyh3wwpZd5STFHaolLF+ZguUjSRK7r6kXpCTeI2ExrIW2TduPZ1nqWGA8YrF
SZbJ6g0c3EVPxgnRDTcZ+Um09FPoZmvMoGJ8au0mTZ+FnOCedA4tC4TtGazzzkk1SbkjHR9krY3F
ob1n4vEOwJTodVLk6Jt8cR15P5RBbxrDDNuLv/3mzXjeR8NZ9v6y/zTl6SNxFWi0Fseo5XrizWF4
YGBsJAObfy9oShNC2gRdhfD+/z9c8MhHs8XXM0ZUnypUAt9fZC1/n146gR3KBSogaQ73Sa9VIXMV
H4u0di9uhDuZ66KYmzcRN/YzDzsve1cLbh540X1OHXlstZvH1zzAU6Bmzsl79hgA6YvqBcrDq+GU
WsV+Fv+cj2Q5ZskLabPwtt+gWtW0E3xiCbH5NLP/KLAasELt7Jx8q8074EnC8Izx1rVpWeREIAMq
hJ7as7cJYyuVnshPjT/n4AnP4uabKstVdB4GZlITCLtrxtPhsOC0w/Yi7/r/kTvj1/HzWG8gKdHb
rA/8s5PohfAwGcUkcGRGaJnPNFT2HQan8271euQSre5jLr6+/crYFg03VLoC6EGz/nKKdgs8uXYR
NZLUnRKbhxHl2fNIMO8woveLMkfiXZcR0ZzWwxqYXfBDngjHitxKzkJ3psM0ismCLXdEqkbE9BU5
v5lOltJu57/BbeAMIid+SeQw1a3HT5BMsHPdBi9t/kS1STPaJOqQba4l7yXZDNoVOmwqK/YAIcfO
adlXiabSZzob4P3bK+cACkSot2FR31pJcwH86cQV/4aokwUXKTqP1LQ1dN2K4RrSG8T6HWMhSdWw
RRCKugFVcfBETjrFTaKgcDo0neTRHuLSUKmGCWBPIaE6Z/x/VXDCOWp+qYTyED/ZBF+cqjQ+/i9T
d1z7tFBLz4uMGtdHLzPOXxpBABPI3CZh/4bC14hiUgMzze9Dsb3FzCoo9QLNOt5HYXmbvJkMxGVU
WUJ+OEJkQLrp8FDA0ZKqUaOrLCeCvBx77Kc0Y/aF3bFjxdglR/R2PYRMHyv31/MwrpZOFUxGEeLK
VVrLT8ArhX4gg/FVrtYg8fMyp9W9gNQeFkQUm66uw2+x3iwgNMlbXZ85FBNLdyijD7qDUM/+KTFV
WHLzGYihWo20g0HH1nvHBgSXTUnKFwnLJdmJivjCIEaN+NgzSlcDtUH18mjmiDmi2WsCaD76Yf1+
75Y7xHClBj7O0dYty+7yxwtMi/kRiUtf7/tQjPfL83TKY7G0lqDZxBD3HSNmNEQc1o+7d4hh7UDT
7vrDM076lK4x7aHWINhL7QBarnGqlSGDRY53iyhrUi1lI6L8EqLcZYakvLCooCl0vr9WY2vPNPfX
dCILq8PfmSTJhAu6BpAM1z4X26uJZOkVyTyTLTjrAkg3yeM+j7J0wYdnlsfpIFboTF+Q6HQgfYYm
37h4cevylqKGHREGQ4sfkqmP/atMxGc2Jg1zjGlttpyr/askwvmTneBoiv9XtnmaajcbuMRl2pL9
CH9iEnQV/BhU4Ne3KatfOY/97xpKPTkhndqCLNa8oeVT1JYP3xOjK31b4BEDzcW/DdZvK/LU32Iu
/z3Etk8+Czfe5DjEA8d9xCMsBX79Gkl4v3VjZDcWTel2S2T3jKpYAWkhXRc8BEvvpIgd7npT/Txd
jHGor3rjeT0pWeQmjIdtu4fRtxg74bsyuOkw13wcLnefqSU3vh/5yMRLzJpKJcYXGHcWOmxl45DS
Y8PaLmRRw2Ij5j1lJZLYZuVdxNsw1KX7tpByvrJaIiT8YhDzOFp0C36TpkDIZGichray9U3PiAKu
DqyqvMzIWsaUvH4iXScEM7xobjXbmk8Xamiw9ZLZz9PiJxI1oriQD50WM5Dl7J5sFym/defirgmo
uNNAr5hstlCxluDA3p8jJZt3Z228vTfrxN+HickH+kCQpL0XGBM+0+JsjiHI40LywpA8E9NR10+c
Y1CMAiblHzmY2sKJ7A5/BSdLlil5nudsenKwM7rgbGtj6VK5Yc7pqfsQ/3c55W4UncQS5Uv/DK5Y
HXxmWqJMNLx3RVYHuyD/1SMpFgqyRU1oHgmV26+xAxLR5gA/fRGPVioeNx4NLcULGV9z6QBkhh6P
TjB8/JmC1KvEWP4yJO//OKsF3n6aa0cCB9Tl5aV05g51bzIEKpnZr+haVbeCBSI3IUYkiSSju29j
FpHZB6smbEO4pRNZwab39sSqDmLOYuXqe+dcWVgY9WQXEtgr6O4lccAygY/DBiu4UCK5I1KPNzw3
ua34Uj1tftpYcUD4Kj5ebNfeR7UbqpbXhpIShU9MpSY4EpH4CVh3JYMisF0Z6jKvRBxQ29P13V6A
sBwNSHFssQqV+qzfMnn2ry/PUtmzT2FzX3p2TBEWbSfnyijjBvbnPdq3lV4aHUZalmhTWKDKUnmA
CRnXLctgF4yD5mptn2Oeg2+VGIKzS2FfNYVPid8t1mCeIA36sJZ3fVyM8umc2CIDxbYmvmMjeMgT
KnEPEkt5LJhk7aZnrKEuW7bBxfavatjsQuy/X+rVPxj+XQZ3K0FHoarXfFHY3lX9oaXPQEWmlrHa
ekJvANlwBERH+efdx1rZqX3Z33s3B2yCLW2k0WyaSO4rmO/ySu+cced+QhuyKx8Xr6zmOX9vzcVl
nb0b8ivfXAfUsEhKGVS/q9/d3EST9K5SbDNuUCxKPK1m+/Ma1zntjB4Txpxt2Ao+vB29KShNhu8K
RuPGjDXSvK5aqzzITN5OlewBuNa35io4+gkXWgR1weJTHxXRDsPcQZc7mue3SlyYvWsvKqhBnMfA
SsCJXRt9IYMK6V1UzoIwD0slZNa/43bvQAjuyHU4XI/paELbyYRse6/BcfXN4DvmeRw4eboWAObM
4/QizXnwVckieWwlltePLT71t471i1QC7fAQ2E1b363/moc/wl1VtNPTydaWGeiJfOFwkirZgg3s
LRFIpWC/3FimjzcuD0Z+uN/LJ+uIXS8hCBBOb29+5sprgoxM75zEAL8QWxVPQNYsymKQvDiH8Nuy
2+N+m+ydweyEb1Sw5rH/cjvpd1s4CjqLKhbR6v0YHvQYOKuZsE8wlNEFs8bfNX2VG3GBItt/ZRhu
ODrBybwEFtrA6hJ4nSpztkxyqlSLjmPImIzx2ocodpSS9vUGcEFkqVNOciXrLgoMpFDZlbieAfcy
RT6EnEOTCRe1AHZBq/hpjLlxfdKGTZ6J5keSejgbYHIrdGKnmF1BZAEVDL//auYXECvSzqMqC6YC
/ksqzR9mPhlBJGQ/WtBtQT7bFx8RJTKNTit/Zj3Jrk/H40MUSQYQ/j73OBz+KTSBhgVHKcWyQYBt
ATDGWaZ5Rx3isjoCSB3S7nIvrIEI++LkG0XMgzomSEeKV0L1rsdmqLP7Ta3oWATDPWG8AChTACsY
fAG4HJ7VuutztTMmnJ5HsVvkMHFs5HPs5EBtf4GFLE6cMv4hW1V7DZbStPnSfyAS5VGeaMJd1kHA
ZdljWjIGTfIr/kFxXxAhxrBYJcCP8Aze5sodXpRFuKKVVpvFhXxj62CKTRCs/kGv7S1RYdr8WibT
7ySggGACuAigXJqaTthwETv896/mfChQMTePR/qGRORlKkMAi+D2F93eOsHyTpPdk7fIz8fce8xf
oB5CihKARDCkWaj/yZGgkeceNKVi8U7W+ehH2Ix7zUbPn5vxQWifmQJCb8RpSAcSaonIurdxNTXk
6r/GHMBUc+lCYM/FgAmMapGmz7SPq3T6rEZ3nRFiY5XHuCSXunXFbx5Iw2a40x1exgByMUZxQQKi
fbLLQDyNYR27JnPtuZe2I4gCaiskMe4KKCiHJWYWofizggfHMUExqnxubgvzN/f9zZ0PynyOoAJS
ecwAxM3lJ9VP9jsKRI7e5lcaJVZv0XVN7APSv6ieDjRJpis8DJ46TdM/+lW88SRpLX6LQRYitBPO
oWWyYMOQa7DUmZwgRkMn7JTcWZtEVS2Za5hplcDdc8Off3REl8TaXcY3N4WtHh5SPnpugnGV2xnL
PQ6V5Im3pyqJshREH2321mrdo5kjV9/2giaws+g1bX9VYD7B/Bt8u0YkeOtT5TOydgRiP2espMsD
XeAwIXSHww2XZC9jcN/qBunZg4tSz2vybMpiQ8ufjpUBLyDi/Nx6+zaPwOy3t34D8tcA++Tgt+cD
zl/xZF2iEmL9GGpajjexZgINEn/kdTYZQH0uk0kvcxjFmWj2bDwt8G1sUUrfkOdniluu0BVehlp1
QxKw6ZytxtkmVULjwSKBqnJgYFDGzI53Vn3HTSSN26DsCc2jJw4ehvjqmElapkQ3ivPuN4g4gkRS
Vqxng6V4Ot7jG0ZUy0LEBu4o/V+WOcBzbTRzzhDhSfv4l7CnBVdBe7qpHXCmZmgdD//iYx2xW6bC
fcD0gebFwNi6Ulbp/7Z4hSNKRqcZgWfhLqVXgyyN3rDyk+fyDFX534YbJJBdfQD4QtLDb0iEs6im
p2Ib9w++uYZcvveNKepDIaBnigNHmnkfY1WUlcfpcyvY1S+Cy4OY9rt820UbKjCl2VBOadEHNds2
5q7YtYRjL0soEHnyEcBm0IwpIdkdMDyal21IwSQhfu35dGtj9sOf+DuMDKC+1Eq1Fbtfx6rJ5qKO
IRwVPOlpYQGbCz6rerIxc6zulGOGJi3dkvnBPV1wE0aL3H/Bf377u2SLGyKtSEqWbWdU1LckvEQ1
wGEaLXBr2hLGz8om6AAHgOAYiSK6JTGNKjPXiTrM7QgbeRZe3fnu/X/CixwOt8re6W9smh4qkzdv
ZdtPsnjwth9+EW65EF3fVD36ZZGKXpsEt6SEL9DUlafA+otih5DM9MGH3CBGGA3Vz3lgcsX+r4k+
drWsT248SdXTTS5trIBOkMsSFZyNR6U18EAQdd/xRc4Tp/uShfrX+MWF4MHDKrrgdzDyYMqZndFr
KNTxeZdlp8K3bZujVuAKZQCbkM6hyHABMM0GQAZ/qt/QhBI3TS1O5Nv1mqXfJgoi5aplizHE8I7O
b2NTemKseVR0iERriq52chOWp9ZAMU5Bo8C5ro2D2OA2Nt/X8YHM7TPU472iE2ACOu9B9cu76ysr
NhyUNrFVI0E6s9niRHCkbPpzGKeMhpqg1j0y5P7SB71AZZugK0CcwLPNgm7VnWr0tpHb2TdsixWq
NRhnwFsi8LaS5seRb/9f0mEc/HU2br9b+C9Cj9zPe3nc1HCsGkpnA+Ls4XzXeonFkIcQbf6vMKiy
RIc5OdO1lEhoN12yMiA/RR3rrKhcMSmdNSojBO1Xsvb9VUwGs2eS0zE06Vnly1fglsPFBNQq67wT
cpsrcdo6QU0fE54iyrI+6fSpsDbVkUFHAWxcJw9Oalj25TC4p2g5nXumYrOA1mtBcDzJLMddFHqE
U6L67kMWFwKQhLholRQFhk6sLURFCD1r3zwvjon2zhJ1A9vQXZKcErDVpnWzOo3y0Vd/b+vELR3n
hi6tEgMDCTZ9BtIbvNANcTGPRUVRcC4lTEMxVEDFeQDynETxC/hJusiPAgFHXtMmmSjGaBVUpRiz
LaOv+JjA6gBLV4giCrRQUbr7QwtvFUSCLj7PQvmEukipfiH/CkYRFhoLDn1iQrnQe0G7dBmbslZ2
yBmqQ+YBeaA7WIJ2Ua62LrxQsjlocoaTY/dJ6DIcR7HcbztwTP1virufWLH3TtPthNlAmNK8SPel
Dk+AOVAOiKAzhrqOonVPyZ9feWskk/KwF6/tUtQk/tQO8hV3xx/F0ZPj9TcbTaWvQI1aSd7wL5M5
8riEcbzaQQV7BFcn6eFfYKL6WU1/THlyiOIDMYDUzZIWbEahXFyR6htKnFQc6KHIF9e4aaYgo+g3
Lng/7UzseezutxnoAWHpKuW/dvgc23AUdfvHIyQGjnS/H2rxdS3bBJ+6JGNXkmtANrP+pH+EMtQg
f5a7zQsvy++HYQkHpcBzE/ff1AkNxNN/eJzy+LohVx1b0h7GqYpxcGXZOMoEktsxwG8ndCjGNrla
LxfbEgCW6hE1NM6+NSokYvt8OFPiHARKf0iMCVYmnKpcqInaA35LfBU8b52coB37nV+NuYtlOt6Q
xftLEyZHtVeF9hrA/42QphnWdTvKLU0LZx1VpO8xG8j0ntWousOKG/6bfbSZAJ8eN8N8kfM1uo2M
eYhfYXTYWLKljXtLm6c13UrCxhRWNqZx1ivaJXXR/oCWUbiGRgdH3S1fFHB1GT9/akTz6YWbOnTR
BJzIH70RQ87RsHJD6C7afpBusFUQeOmG/Ob6b/isE66+LijFE7iDsBgvWmYfdd9b9Jdl4VkdLlHS
OtclTRDBY9Bo3imKQ1aCk3ubhv6zRvPemFmA8oF0nB3okR2d7+jyNtqAcYnN8I3uPEGj4LaFULDa
+/ASGNpThBWH1YGcn4wks3/Vt/0XSpNSgNCIFTHMEP8prPdoRB6y7DBY1ZIWOUQQrNlXpXdrAi6c
/cxBrIc8XKq3eR8Z8i2lMtH9I68B8TxHXstulLXmgZjvbFxD1Cb1OjyEiIvMCKEx8Z1VdFWhcjF9
8bX/a8hvhPk2fO8ewrcT95kEbtS5VYrK3dDr4y3dIHh1+Kgy5iuZYppZ3uRTKNFk4go3KCVBjAC0
twJ2KEoHStgYEQjZeGoH7cMsSSH20C0zFwV6DFmuA5kmh9b14Z7PRRsXkzC/O6Uo0YplbMtYLd/s
EemJKo1sJVI+qoZ3uWk4pmaQPQkX5jLP3lWFAHvibIqjNHt/H4nDyBJGwL1DPk0QIrIwUbuNhsrW
DP2M6oqRQm7rj4EJvnrs/nmJZlzA94gX0TZhZToFJHUlz34rtbq0+2TgJsj2D8Ueqx7GJJKlGEX8
8fvnu4uU+xt98kTSZVuSQNS3ydStlIfre4d3Jf6Ce5vFJTAa9lhTvdqnXU9GEIMFDnhJt34GWeRT
XBCzouSMS7DoURT8XrSsiFbqDCp3xU2eIz2Vfim2Ro1k4eKuooc5WrJwi8GNPc/zlNBOpYAmTsra
YAZkyC2IacRklRd0vHxQzcoR2RzSZI7FIKAmquISwJDyFuwVaclW2UAKIn3fcLzhYWE179ZwAcNT
Kb0RWBNqVQuuDbiFlGo58qkauRm5h7lApQKv1hgMEAxznexAz0Mmp/03OwAt5ZZUyp5J/5p+O3N4
bDSKtn2XkbxOXDIy/BQDI5+uWdumJ0fc51n4bVt0Rz851NeMGTePIQx/9l/La1jim3CcmpvkGQRE
wMTzoGTcz773w4p776GD8OEm38nHeFg5OdxwhvtSnUxrEyKJ3ODUJhdRk6tmLM2CCVcI7efQ0jFI
wE5ZxTkuiGsZYZXaUcph7MHNl0ECbLDZnqNIqIAOXhx8aTa2PJKWsrCJEW0gWCUzKUsxR9LTWmoM
gZXNQW7gRykE4RV0XQMOUCD8AT4DTKbCdKqwMU8X/4NwE+D+/uwLMpaoyWjnMyRD1ocrb3qzdAF0
1jy503XnCgr1He5Knna96/iMEDxkJmnOsRTq567QCtC8PyleH5YyYPU7P2e0eEX+pmY7gxEMmz/B
4+A6W2wmHT77+hzxCo+xgbSEIaGDKjMEFDhnI9MVLvMlobgp+aK/Jk7uHILBprjmNpzH8J/Kv/lj
YLLa8k8n1BBZgCdlSmBU0QN9RLlg1VrBHFpqeOd5bVf6Ha8IpteYjpRdn3kOU0KM+vphAkC2jjhN
c+S4XQSBsaRM+fg6gqglE5kD5fMmRthBDL8fVX0sQd/sRRD00qhmrnQVBLIlBqd31upQsdPvIGbY
45+vrCB5Pgk/JMwshS8N9Lqaq4M4In36dR87oiiIC8jMd8hW0n/LlvJ89S4g1GuUN3ZQq9+F/MA8
768hPZB8KBrHArnn3vDJ/65yJJgMysv/c8Q+vT/bKxUo1uv1JZZGzQ7NgYF83jX3E1RdBgYHwjk8
BpLwQ3sIYWnn8neEr8B0lejokvcVCEpH8Wu7D1ynbSoLFJpb4nWXTavq9rKql/ctLWGtEkRkpwC1
oX6QzinYqVocfr0Cuvx1at0rnx6h69qkq/EFYN/IOB3CZU7CEuO0RxvlzLIwiG4KROtGjTp+yFzA
2JOhfZ8jAQgfrvEt2b+I6BAivx+VO7RGFNLriF8qVKefnKfsXMAnq87+3BIGqle0lNp+8ahG+cA+
ZDZQcYtLsTEpYBwbIwDit2jXpgInEhry9NnF3fpUNyFuLwfAgnarjOhZSXGvpGI62osFrzjI1o2t
vjO0Nm5N3bpXoepptJH9sHlNMs7hctxgEg2qhWMt00kmOhvllQR6dKfqloN29CPzAFYKPk23m1IE
NNT+U15nZQ1V7ol9IfokLIsiD29qtb0X6GsQ2bxjEYIbShnASQCXFF9QEval4G1Su4LMifzBB+I6
Fwdk9JpHk7NsETc9B/y19zjGxLp4V+y533LQTdY5Fds9QIjFjVmP4zZ34DF1eunHoc5O7P406XoQ
OqqqBagu8XLDh4c8B28BFThong9kHrHCP5nVdt+M013pUgU52tvB1oEC8YHwIOgnov+uaKrzksZ3
i3YJ8KlC6F4VAHCw44QN7acSo66obSlz2VBbyzOWeLmNXOg+gORkEksFIbzOC5Ffm72OxMnW5Tvi
hII60qvByThFhaG5NBeay9XHqCI+flxvGOqxOiDWel4hTw+8FxoLSj0KXmupW9U3ls6yClc7Lrkf
1IpA+A0bsJJk/aCDBCklhs7vfug/WezblH0Sv8tWBAlx+uOtPeCkF7CWXnWWql9epwC2uGkDcuK8
5o5YvG/ENJgLi5irMriH3ILgJIfSqNU6FkBwMHSzPmedYdOoryKlwwEFf1X5u7+XXuz11LrBwXVK
srzE6E8OCeIT4SaulY4qAuO6fa0x1GG7ViiobNUx78389bCpHsbA0Mn+xQwJwk/y8oqehEmkWzna
FcaWlMVO9iWoX+uERIluEcayCwC5BYKaiFbjEuXUZYn51CryofHf73J2rD+vkGxYQJI3con0NCz9
4lDLrAjcfghYkRwSY1s/Za0AkVdKH0fH0B7vq4V4UdPfsphLtY9MwZ6qyfJWFP1zgTxsIIoLoahS
cxHvqRkQVVPxA0hW61iPOKr0+/aiJLcrrD6wP747BH6fHoMqcYAfFWjTS/CIYqSCVHedYdimQno5
iWjpUExCSAtOtmghymTJW1txWt5Klc64yo4jzXq3WgdetrA0eBpKfc+lGUJlvETv1Xt4RpZHBWjJ
q/RBGFElNm2awWN6Azil+k+xj2i/Q2cjV1xC/GCSRU/Hd2HtcfWSyUxXaAXbJYcqNw/pnNe4LZS6
vM88IR01hQq+wl2VL4yHDbxvKEjj7ccPV6bz+RVxnkRE6Y3BorWbAr+Dz9tDAzWdKX0ya9Xnhq3C
Wn6lZRpwFgB86wTb1Xmck6VvdMqvLSndvczLnB2iOiro8ThVX/HxZXic7ba+dDhDQX3igh6PT2Et
JsJdiOvdvlMWlT2MNGJfV+W5kjFUlbYOqmuMnk7hFRTWV/20mFHthzLR4ZDVv6L4o26NR9qWTjOt
cd/T/u9T5gwfUmsbe7lauJVY9PGQua/E/AD6FUfHjmOdExLMg+CSMoV5gcXy2X4EMo13VG7BAsUI
Tc1q5XQnxawYa4lCFa/wkz2rpyg7LjPyCrif/Kr7cC53g1kwDs4rcsy5n0sZIeL91mQ6t5LL4GqZ
EK0nwgufUqxInjLwunrNXAJntCQP1siUQZglGIUKXTXtaYV3mi1WiQXgUdDvgwxNKghYYR9WwJ8N
+VSE+9gKTkf1uTCnIc7i4nXxSSa6fVEHvoNOMDxYRFei6L2sxvmW59YH7oyWTtY1Tlq/K2lrK08i
TQZgiczz4IG9BIE/romM60NJheDblxookeGYmagfb4X0tcRC75C1Fr1HBCSiC4k/4dgnbZ5wlEzb
ufPR9y4AHz7tWELZH6PMPXSyOCwzt4DOAfnD9x1MGNOJQJysz0aJDzdbPS71oZCA0E2BkqGVIAiM
pq3m+T3fMh9S8bar/ZrSj9vZSnl+PTzmTNZI3Jk664d/bQbXuJqP42wvOwiPT+uhHIRXx/BoTfHt
0jC+Q6YlctKbWsavUHEH4Y0iG+BGoAbV4+EVjxS8oqa6woBuyGz36ApbfyrUm3eioqigDhfMyKKz
wqp1+hQCHReGhR5ysWiU9/UrD3Qlwcu0TuGz5yZ/tReKf+udPkkNC13uwffwGNRWktLmPKERX1p3
ufa1m/OjcKIgJJFPR2fO/g3YiHOrQavq6bUsZZqTM0ViTg0R0Jq/r6IDDB2xhFbYS/envBza2Ngc
0tiyxXr9g1iJutaqUJNWsSemYSF63SDk1DZVwOvMzG8LmDqgSv3iNXIJRnbq3Y1qbwQs7EE2LzIh
twq4IzQfMZyxbuWHeSwD5DWvwKefCOQo0iveXs70mijDNSDr0kxuhfJvnRSGE9R/1MJH+v/tc8wM
atL56u+FIbXMOE2WHi752wMxSeH7gNB0Lgm0BMphHCGtgHwQfw0DShgjWqCGxcHJrKuiBC6av+DG
6NOVS2xkF4jl8H3jU4lj4lsOey6N5WJRRrwExL2sczMTHh/DELDDl27gWBwUGmKCFw35p8gjnUV6
8ZHkxBUnZW9+8wn0xR9k1GfZuOlz9OSRntzDlVWWlLQ4kIU0HM4vzXfa6j36+gjeVyJ27N+Tuzln
nzfmGulj88dtlNlctXVW7MXfqVFPKcBOZi0v7gFonDLfDJz7rOoR0na53CWr23+wNgoPSFbl/DGR
uk/X17CDLNt0LFOe4TjLvUbSlxLk0JryHdSHUt4DKlecUmmEgPQWSV3uYRfZHBkT2A4Dx15rd3+R
y+TvUkPIkjp0+CAQqzCJsm5xw0AruL9uUCgR7BwtIZeEehodTJaGdbq5XZ+maN4uzxHSZT0q9lyD
85V3gLRfg41tbeY3+ez+r2dqjQ+wjd9XBi/p1p1BcuPgKBuQB80OhwmRfrrxTqCtGe59KZno7Tmk
ORuxdIK7Rx3zwSMCULPKcdP+cWFRQCGZyFgEKSCCBB1JGZdleS2buluZeG6xij7ohUxX2W2SODbB
JtsJg5ugf6GCn4A0pdL2bskPA2WpVoDUnPECB4OyWeNgVRTceTTTEjFniwVjkCnixCgD65SKCtrW
ecYYB7p+t5XA7Bn+i8vHjeH3Zq3ilu+hThoSA4frRUuZfIs45ZrCqaCnH/4wsc1gO6O+SYiTDVDX
BiZe0ffBMqbzTibtIftPFnsNKuFKBH4MJRNhPsBEGdducKoNeCdiJmvYSWKytP6Btxp/lTCUCRb0
TE3hO/g/PVxIC6M0EAtAviGvxYykrwlIlNnSjm0AqeKRDtdL3NsfiNDss9yhJq8ciJRxIGdRn9Ad
4G922/ZHkeK7GxkC3Dg0GEki6ntICW1WoKwfkBeHP8VjRVb1d0zFFisw5vL7jqZOlRIMwrerAYNT
DaSydQAmlsowQXWi89/fzpQMMXuspvz98eWQ2qR47CxTjBBa0Bhp/Gg7qC2deXaEzP4odY2qDlcM
z25b2MmnR15C3Iaw4BTYUQhqpChZtL1McMryaK0pTVCB4sjgYjMOSmR0BSr40mwiRU5X9hvcFfnp
hl9J/5TC1T0OAfz+d6iI2bMZ8ZWPzNShey/4gZ3DDxLDhoQfWztfsKxed7ZLDTo0hGxpHtSEnn7l
bBLoTuA8VWUGkWknS0nqtSVxh3Vj9XepY61/FY+Y6HiYO0AELXFbdaXiV7jpOJTwqGugejFjcRiH
M6zN7F9nuLxJpJ8PYoNgjYRAbCbUzKYS4ULc2CIlyoKQBUU1LJYuN3AQlDQj4G/jsUhiikIYVfJy
MXfWwgotkAIUUNoHnQet965b7y5L+dP9tTcW7CX7BWHmc/HMh1+pkv64lpp0ddOBgv3Oz6GE/wx6
ZZsfN1acYysxeRNUaaGnHSNTWr6nYT4LHfMO5Of40Utycx5zMUfhRLX6FNlUI9auGHk5VCwi/EUT
IS27RnB7KUxeOtHwS0xRt0exa++Il9kIVWFoFdGUaWoTyYA41u+WVbaMXcVEE2TwgeL3HIbDDCEE
IN8V4hl6ZmBIC6E2ZrhJroL0y/vr0FsrJFQNwMOiGehV2K+1Xjga8iL1E1LUoJeCqlwKhbM3wOco
ihED+eA8i/r8xp69go1vxbsWQaqTbZft+oanLjPeYRA5BxzkuC88aJp0Qms/PKFlq865Va4csOZq
AgeACJf5qdiXp7WqETd0FXswlYUVMeUMnu1QJajEvne1/cT1PoBkkjxKcs3e2tilV2UdU93Xhxxt
0l98bJIAsFS9Vv03Q6gkKahcFQnyC70SCXgr27luABgiJfUhGrWZOGSPWbWIdPEglWXtZR59vN/Y
CHWhHR2mZ5EzPHLcDs6b4Gh2s30rtXmY1O7X5Fo7LbUlRaAp98x5KgU3GLhNIuu8az5pg9CM9Aa4
ndcxpxoNkpvlVry30lEOKOTmbvb5YKoqQVlK2o6JGAMSPlDRiaoPWHxTd3SgjPz5nN3BmmY6DXf1
4n/3hCmkCYLokuS+wLo/slrNo0mqoCQmX36kqWU4l7l8V88yZB3yOENYUgE8K4nHUpuFpNJ9wt1U
J/WycIdzTgUNHjgbisfUjxyoIrjGaeFFZDQNGsfEnHWEG0gUgvR7LwNT3y56gXAD3m6oMxKq6PSg
RBJfrWyGKDtJFj42AULswcNKlPOo9k+dcRIslJ6p9n+CRb6/Rahhli1ME2nvQpdN7vsrOB7y2Ez7
48VJ9PTjiFhSEnYnLEJLZhzeI744FT0h+jaPwi3qQQp634o6RL4wEwdzcfQCuHtRXTxNZoNrJDGG
YTWvbldjWVCyGoMJBDHvvCTEBluqF6qahWuZdA0H1BN3UZWLDdXTTJ7QEZmRJH0qlsVm34nz0KF0
dRclXKK3cu9TUDk4M19kn2x9G3ibkAruHPKXlUCmZKJIKkPG5ag9tCaAhwuDq16fYzx4hgvAOq48
ig9QfwyjBO0AqX7HRKtXyH2gUonyPrtLfXc+nz8ccB9jvqqwkXwPONd5joDyqQk0tYT9w31dEfRD
rBRuxU0iXSRKAg5yFEzajrf9UZLdYvY/rq6MgEo9OnLZLXQ+xS5ctJFFerauz1N8UUgMevyy6JJ2
rtUc6//nTDLpKDPxLJQscAFQB4WKUG2DSFWW/XHefsW8qnsgnG+6OJTQHJdy9WRsQAJ+H5m6rGCa
HSpgPLe8Ok3Kh9CxKqp0Ocj+wEnkE03ytEbjhEiyUYo4TxGOGvd/6KDPioTjYtPVx13XA2D+3TbT
Jq6qA/lWWhPImsRMpRnlLdbXrWrwHagfwje8bpjHNLe4FbbVUPHPG2zmJ/O85kcr+fy8ZsLM8zPK
+8p94eEXDqhDi/paVXp62Ry2pxzT8JK8a2g4EDnX9gPJom3ywQcqV1hPdEVTl+TNmbslJmMkCh7a
JE+WCTbAzjj2D+yFUFijSTGRQYhND9+bRpBH+7Me+nc2eHlUp+SGvq8oQ95WGVzjun+om4yyreG4
EFrsfjFoExD8lkfzEvFkWlNkYGCFCNfxOKXJikPcBpNzejDHv2mKmOg5+VgYK3ZFZOaMjxhl+hJ9
whxQMlmOsYXEM9gN9d94pntyYw/YRQWmCUvcqN7SpPQjjmwxTIX6eqjVNy55bLBmQb72cfNOg9Of
pajnpWKUyrzTVVtwIO34SLjcYyzA6VSN+5MgpxA1R5m8XKiPafJzOq3BzHbhWTd1AsgSY9jTHI/7
4QbzTmUkXGn1W5Dk9Qa6d9Ye+DzDknd9ubOA3J24eTnUYzvcujW8BdTIpkD71a84jIoILx0vUT4H
M5W1ZyCopDtWD7AgYZ9XmKziE4T5d3MXizecMGxhbc2NCw3W7u7tltGIvD87TczM6ZI7dD8Jx5Sl
RsHX99URSvGadgMVXHDBTKiNULec/1ik2foKSt/Ge8ftom3Y+MC4WZoIiXkVyHqT/jTl6HcH0mHd
TtxvyhYsnGRjBtuVCIANHeEds7ydDmMQh3Kwx0PtuRpiO8KDVpH+GEEmYDuWURY8ZAmwnZdha8AL
jAfGTxcNgeHYk+kZREfqBICag423dtbYEtHdtUclIBws1cELgt/JhANYf6g4lYpYtE12dWpS+hyI
6hiOcXwlit1kG/cIN3IQtVdhJywW/YX3xiS67rittkyiDzfhkK7QRkA6Tu1+gBdyKJWDFhyMarQN
gzs5at16aWMIQv37ECyPbf9eJwdiwbPYDQQsMwRaXxMDAO43yd4EMp3xkdBuFpvnvmy63pBnotXY
Hr2rVVdLrfWHlIcySKyp63TWP09gBP/k925St9Lq1Mxd5dw8h73COikIsTLW31KO9h1wdsVuSsKy
63A9tulL6Ouy6lUXLBzyTrowk5JyDawlmx7SnW7YnPKlhHIlHa9h5URNNmzKfxL8E3SW+8VkF/81
5F+MSFLhSgZQ/qbrhWZvSfbuplZnIVfmLz+NAkl+PszGNpIp5CZ4j3sQ45MscR5wdw3/iQI30ezy
KsPXtnu6eriD/5wQvKPuHpd21HLWlbGvvtHz3Y5x0JEM+30kDtrpe/2Vstu/2xT+QBexZY4OLiy6
OJBfjN3V8Lzsp3K/c6ZTZdRoQAcK+LYJ9HOTTv/BvvlRnjQx6FwcAIyjWTwPCSJ1YOc+8B4yGntq
imPN9a5EMDBDNvQsrE/oOljOOhyd2MJiLwifch+snl37uXR1cd6EncG98fOwgI/3LVQVV6DgkWFE
YluPdgQ7q1hqskz28T3cU8VY2dJO0361hI7HWpT0argObZNsDAgaim8rL3pd/OyhjvIrfQsUNe0O
H0BNJs3IW/dP57seokMsA6b5E9exBEHALrW/+XM1dc4d9iCXDmza1eIOvYweikuC0yQRUoiGPnEM
77BkqLkmRfVFukhsI6ugnPvkwzzGEVAmIuyC45stAU4ULPFiABVOMaFjdRYuPsfIgChz79FRgqtz
CqhNQuG1UPYWVtGkTuD03stjEMH+qCNvv6VvWP7v+Obuqts2QMZzX7/isV6+t/RyLmzpMMswdZGU
lEod2vIxC2VF90djU9haqLR53Wkurt+AmUG44NEyfQxRukrTYW8d8QiPf1kw+mzCTuE+WSIPuApy
17LanW3X3SOnbw/O3AeCQmugkQXLBI2o+Dh2d5nNk3KpSQTEhkZPp4ltd78LZhfOOGcSkS5XQZT9
Vpl59AGZqln1VPU+fRqpNZqR6EuLYYn7w9uB23ZsU79oe5UqM03h+HyuSTHeIF0+k4lPBISaE/tI
PhipWRRQ8VGQd8Aqym+uPhmSBFCxe7cl5PfJ4fnkKJYcTXY9rjWDtKi0PH5dpvvMGBxld7RZXTOP
NPjUnKG6kXbPXf/lyzzpG4H/A9VrxTPHHA2oelJuMBDyeUIe8yR9U+eVYzfKBuB8U69e4WKKY0gP
qUBfxWMTGh3WLt5Aqx8LWvH5PRPPfxWx6SNgNmWFy6FBtWjvboYzuO4GycDdRJIXp24l1BXAAUBv
Pkkw2+Aa5TGm0Ewx/ugI0O/kIZFpqX354LjhpWIyJsff2CGWVKJ0mn51YrssbvN1xiWCt5ENDQdn
UbQyq3s6glVhhUFtxB4v6YHy89JSlm2aOFBo0Sc4THYO23FyXZ+Sypsle/RS685Y0i+SH/8SwWke
DKHMiGT/U0md1nkgtetBGRiwJHpuMbbZcfgyr/hRenLaC519K/3DqKn3iRys+mmDvVUUMJQbKpah
9AtWUq+137qfZgYKKY5jSmMLrgcYfOsFLVvmKOK5IwBXm+ze+kpT7ZzVOMXq2JvwTb1gYsOoKXtP
wAEhCoVCaTcptqXpQVexIVYPts6QJM8qMmvL8kzchw5vjXirUSaEgJ8xagZgqTkyMYpv5/iryb7A
Z53zyWFTzW/PFINouhRgsMV6UK8kJ/qfIY9X0oHbEqbZURxdh4fqGRtoZUfT64jabSViKfvXq7pz
DddHTyIZMeARuhKO0tYU+Tc29SBvP7zNQ+VIlBczE/i9rgUoQbMXzOci7GzlfJN1LUNPMlQkSAsX
BEBfrbO20/d9MVpMxFBjQGVqRu0802Hsvzju6iKdxVot+FDLauxIRmd+FawffOau/+DGqeW6bEBK
MInXVQ0jvUd9EunsGnN8IIej/NV3kX8KKVkXxebJ18xNTlKxN42Ie5imC5Bcm7cThZj5rZZ8UUmU
BQ0ORxaQ+NJzFY3yrIPwaVcAqiU54pusoLwRP4SOKuwPMlT4HHRNqAmaZB1/2d4xqX5XQppPSarR
1hx/YvKmjGI8uLWp3Uj8Ozht6ro0t4W34U4CMRqPGCiufd22dRCkWXfCJrzzm2h2CFk1s+zvRlgn
PPx4trIYrD7pfKAvqKSea2/WQ3zbRok/l/kq7cmKm1QhQ0JeM85hL3DWjpOQz/QB4Do4MuMKZw6Q
fy6aQAd9jUEUCT5CMJYsbOdLuD62SUrQdEqwceB6HvyIPhGY28nLTnWNrcI8EnKIg9qxvdBIAiKR
SrCPXCsDhPcNpfapBsAq2nx+pOmf8otA+hdH7bQ4xdh/07VrEBTgE0STPAj5kUkluocjzyfjB7ul
6/jtr2y4L6YC6dBh+Hn+4fT5NlT811bCAtUWkMVIfLwLbt+3/W8PlRhEOK8cOfiBy7p1N06TRZDA
9vM4cSDRo7yzqvDYPqHDJyIp4vK9ZBQsEGlDuC+y2UGJPP7VAHEAJnonyql5Vl0PGhz/Vz9AvcBz
3LJQ7/fiss5gqOGFQIftMykx/9+mBEKzcn+bW+ODKWSsr1d4GL0cb09qyAJYIHsgdA5ND/HisA/u
lB9PRox7AO+uww2bJObDTriEva4NrGwKzzTCvZZujfJn/er8kkORo7fO/F4DDviLvVCnRoM/naHp
d346qTDRmNWLxm531xjOUkRBHh5vP2eaFUYT5nwzaGu0//0n7O0Yc4MBU2W3qdeytlIlcWiFsPAQ
1XnIGooetXazUuQJ/SGyrL2x+G+UXQvMgn352IpP5VuNfCDnwcJWvDB+FuFkaUFP30wCvTDWWiKh
ooM7O/ztQ0ETR/xTXrh1b5B+Bp0MPmG+kxCq5TCdzhPgw3KVCzZsIYVFOeG0M8DVPlvaInrsAEy/
XFbZp+6XSL5Y3dyCjvR67D/kVC0FRwnZnIS092VX4CafG1j5c6DIjItnY4hAybJ4c9O/8qEtlqi5
q947arHWgThmrEHpqk0CnGHDbVQ4YxK6g8L+6VDRgw4AIcYf8h8Q4toCYWp4EL9/t2A+mJtrNVAv
mBb2t/dn5fP7NBxFnCORQQ+ptbui3C7k4BBUBl+6cuPcbCG9t2j0YWa+1tsZ/vV81gZ+ihTTBXZG
xl75QgjnLL0/Cmvsje2ZGgVixfvlhBNXWiGQXqAGQpfGMV5oSwvhd0VqAz4d3+aVDmha8Cuaw6fs
NQ33Ul0dExZC3I0DDnmSdg8RwerC65AawO1nb3GZAkCbBl58lIiMUi7RBCukXwyy1pJ0A895fxRQ
rIm+oZ1rR/qe6Wlwk21EiKdTqXHxhzjaw6UXxbPsiT2xRs27oKrW420mStQdwY0SbecNURrlxlXo
9p8TzaYGpCV9CKnOO+fViCRH6vWniLh8lGSQrDQ961RgV1VtlBCYBfbMLCE9cPDRc29Asf9Pe/9T
CLnGCs7QnVA/4kyoec7BDagy7iVDu8AAVaZsrU1yCwiY1IKnl1zo7uTAqmQIG1FFQu1ULaxgwav3
qzXEEn5NAzAYlwtQN1WbW+lB9Oc0wAvTcLb8s959tJGgF8S0zyWfSVFEcUZgfJm6K8ZRFkA48Ssg
HM0GGv0NdCYI7P8uojKzvZpRpH0rAe1h2QlngNp5bZDhRkyS93Ae2/3KDlMiHpaVUtgGZPeA0Zj9
leqEZtSuCMhW2b36Va3yXvNi4yX8bX/YiDruTKKxJhJiIbx6Mg8tfCUVWDi0nZMZ8s8v67NpneAc
6SrxYbQUQGZXJJSFCXpjPfYhgW/0rkIXADjuoQd3Erqr9k2RiWVf9eiJZx0UBZcI/qmb9hT6uOYX
Tt9wOhs4h27298FGd5OSkjhzte9BhAfhVXOQ2+hqwgiLIM9yPSFlTyqDQqbGcZguM5h3bb1XqR+E
3Y+ajx6y8RnGhAhaok0krMhuKgcVms9x9abyczt7g+aYJRFuZ70DGSAavPdn1rxOulaNs8cTifc0
siuTNcHEMIlSW3ZiHX6gUEjj3qVjDQ79uvnLzmUUvC1bE3JIkr2YD6XekRnfa2n26yq/VvdC4jww
O4pg5wFWxQGdnWEWhWyebEKsK5NKrubd2g379SOuPCOHSSVeLGNzusNFPC2SzjhyTIFYoyZPtGz3
hFLWMtx6sXRPC9x6EhIwvRik9lwK0iR+NRC4JtAo9cVZBTz7GXuISHj/Z/1qwm/qc3J8Pf7E7oXd
kl3ygih0Q7UzUfzh7o4rRrSH8ng956cjnXYABElWCgr5qFxHiUFaQdEm63oeqwNKbJ7y2XnGGrd+
xjtKdtBvmGZTILudCU3YO0/nHYml/8h8QFyHE0zIA7lF5dqRpen9ZaWzLgwFWDwBKUVqXdoqqgU9
Eiwy4zXOps8ztYLb7QjoRi6ODew4WKnRKJnrq4/+Txi7ekZ6PdUGHA+KAVtYqPni2poydKBfORnl
vqjsR6E/IQ3JLtHWCvjkO8oEY4MwKgmahpMv99mYzDE4VqFE7nCEe3HzHbhibaJXzabEwxjzl78T
FeVXWGY4mUYcV8HU6UTH/76lOIHATLsF1xlAkMq/GFjzg0JLXt3TFAD0sopGA2EAAbA6DdzTOHCo
J3MJiOIZCpOq0WqX/D9DV5sumKyvWjj7Tx6zIa5ck6R3ZtEy1Xhm8Z9ljgZDkFRYgxqembstj29a
9hBMM5Ve6EbWZzSs2eF21DshCsgSWDvJzQLiXw9iWeu3TejIp0Jnu+srYqVpVv+Wws4qFnnzD7uX
Ygzr3RD8ob3aN94DnONVuxAFo4W1o8cFtO3ooC9hof4r01CYhtmCE7Azn2oOf053Zj09OqswgYb5
5PbIBMEqr41eX8Vx6MfRC1iIzLyeMlOJ132XHUmbeEPXSo2xI4cTHc7hvsa3doPqzMZgqCZj10Jx
TJleQsK1WORTyB9IWD1O/ytMUfLfO0gZBGMmixYhUSh0wRU0G6/WYVRpGoHfTabxKerPmB+NLS2d
2Qp4pN4Nfp4TCLQ5andxnc5jndvJgX/XTAFOBBvEVn4F9tMq7kkp6PbgE/vC5bOGBMKORjf5SpkN
An9xkRP9wWJQQwImreo3HwHbAuflepAQybpnaaxy5ez/xE935KZ7pRU/BAI9s4uUIjsgx0BXCYpn
TnWwPhVhlH5BhzuhQ34izv4onQ8OYmSOMiu6mKhMDWVo2XzrCK+YbvTJ8oSM6DJgRJfLp6SZVq5R
76w0fJZoBAZeplspRozbGPgftvwVs0uiGVDVPvwqZQRiOaOo/DgkYJTR+jCdEgNC4rQOOWKMmdd5
nSw9Tzwe+htVZMBtuPZ+4JjAjWY+YvMos2xAH4xIhG2oW1Xcwwgqzc8Af3t8psORthH7+clBlgB9
LfaA9LFiwahqTTLNjhCFUCgSJaf2fXBjXfXr0NFOHkpwkRn9lBl/BCqx7XFX3cskSo4fBR9jYOY1
tPIjE8B1oVUuR1ubg61mMr51Yz2mUYDv4MUJIm+tfNN8DjDMkR7tgYbhdUnnqVVjey9qNxC4rqfV
IE1tcyEBvYuoK6AQ+wAWaFqnrXWALKN7ldE3UrZ6fqRrcl5KGF0aWwjacd1lv7O5iQZ8RH2ZtF+m
XVUddiwoGLOo4vZ0mZ/4RVf672v23HA/C0GAS83YzY1YW4WA3StTVGvRZ4S/svV3u1Q32pW61PJU
rC5uY0GfxWJzV/QX5NXAsnMRfBnB4M4MH6JTM3riS97MJykwY1oupl6LtIvMfabO+1CEYIwP3FKn
eczxM1FVHPKmeC11owj0rpTjHIXmUy448NiqMvObeHSv6tIfpmGTXo87N1FPvXq9JcHSQj3G5C5n
2BsCI7AUz8eyzdf8Qag1aJy9oPPkCAOmUeQnPD157t1oXt2s0VJVBZek9W6lTlImAYAFQkjxvySZ
GyWRrLNE/0PpOiEyZ23mJfvFzTnQDWrA1B2U015tBYbzUEXi4RnJhlQVWqqJJVXx4JO8GKmsExp+
YhTPwmg19e0yeX4Jd9qiSYcCCfNJ/KUBRtUIfvb/kWzXpyrHVfsbZHOXuhP4t4WIGntJDs0rddNF
YF6YvRv4zmYm4x6ukIZs6Rus5CkOJoOzj3I2GltXIqtIYugaan+0nctc3CB9ys0Qv3tjBNtMKnXS
k6SWkgNwAlxToiuDb+DpCVZSPRXDfT/TCaHHph4cY+IjcAR0++gbykhWkUcTC6Jdz+nx1sBMMANZ
/6tGLxRs1ohiitKEHwBE4g3jLIhVg8Cc3l7MGLPMfboa6apEJh2798L5SbGKOfCC7dL/NwDEVETQ
9D2Vr+iLMLxA8ktbAlbdjWVgxUjgY2WJxaCk7+qYlMDGD4Z4HouXNaJNRyQtDKPI6badbe6VXlv6
IkyJoGsEzarBehUwbUOxLTtkhY7wyh2p34VoM5g+R+YGv98po5XjZfhrjSXOBaJWhZ0g8CUVZMHb
kvpg3UOOIudzszDUBm5HFz4pBBDxEufTOMJoZv+KodAxiL0ftYYCb2vi48sJTmtxHHIYCEOPjd4X
/C4IMeX16SsFpZBALQdAeL4YC2T8lVPkywgVxWFeV1bxlhW1N/xdRruB51LL2nuDx2MnxRWNSQ8J
Vp3PSyZgI7OYDhwuCbeieqoW5N64DGuOkqwAHuF3NCZvPW5CumkrwkeP3M1Im6dA9M4ci7rb5mIf
+ejTH613p+JHgZtfW2eDRdwG8qwc4vyOBJtylEAGlw4qigUbHQdf9H9zNZu1WRoJuKxRgajTWB7u
gaDgtOVDEtaPhE4AghsJ3AL8dsfx3flvTk07k6EyYLuSt+GcLmtusr5hJ4jJ9h3TB+O6hLvyqlXm
FZzT0JP1y2gugizsQp1P6nlO3RWHPJVOlUvsIRbV9h8UaqqNiuAwLNUrOhgJPhsoBo6Usq9VpEo9
2BLxaBDL/Ot3XlZMLQUukuB98XkGLGNvAOPhno6fuxZOM5PL+uNUfmR0fF5MqJtvLH+QcZVp102A
upUOChvuC644Cr4C2jTGH76EMhYxmRlCJUSRRf0kVPlX3W/ru7IJp8DBTNlu3OXzZOziJbET8H/M
zJk2DmfxP67Z7+B/CU/yTBQrzfWathH6T2LRxbO3Hg56a4cd9o15icUTX2Wp/t0oR7omZQcxixcj
MJ8tq18P2BPp2dDskywknPpz57iptXuyb3qXFK4+HS5Pl4FS2C+alqVVFNeOYBWrZdAPkTviWFns
/oM+lR+NH9Ync8Hy/qF58GSoJl3k7XmDNMIhl9kxsfl/Sic4wbvhN85/FVTBKF1sxWBucFbjPR6T
q5jnBXAttxipK73kOviKXoV82jzVc4GplwqOBydJVzGim8Ob1b69OfcEacDxFVRAuBrByC0M94xq
N6iI7FTS0ISNRayt0maR+8KecWWYU3wZgRGi6foAeWUxeDZPwO8vkwS/jRVL6YA3kNxQZtywUF10
D1u56KFdxyWqEO94BEdykfSGAm/aUGfRJHC/3aEsiJ80ompkYud/lhpOYZPYpUGRQKuSde9rWeVt
hTO0AMRMck0AQBlHxUKchZXAywrVL6HAU5aTEZV6YvhDt02X1SMxSvYnA3IEBpDsau3hrXtGINYy
q8pGLgCuOgX9u2zFnyZRPBEsRv96aUYTSSILciMimciqjm3/g1LqcXSwKILlIzhBZIQgBciqEgMB
X51aRVeZXxke7DsabKyssubJSSnfC/ZodDF3aSFquevSMh/6weNbpPInCdxIGZOgjBik45kN6m7x
qE2IMcGRnFotdzYOCTjGTW+BxazdKyH34xTveHRou5VCSPlDWCOMLAcHhr4swFzKawinDoyQtmrx
iYvLEj3X+m9dkVt0CMXwxvQlnmX6OvldGDAse7YuNwUt6XRsXrVEsGET6XjDjM9Trhrhnbzm9SyM
SVj1J6Mos1UnyljKwRcmSmqU6UlRJGfzRsZuqz4JUalhjTVy3vsjD/ZLwOlhVWtrHAan9oIvcZh0
h2S/WotRXxIQrjuw90rL/DhpOUGAxuhvSnoC8GH7zgFrlG8j203bI1Ioy9JX+kd+qqQLMbylW3eV
7v+QUSe19WL9d/w+/n0KYvDIX/PCAn1S2tUUqab1iB+w6OZfj2FgNEVq65p0YOJdrXCDq9oOVp91
XGHiMHnnHnDkzAmS76vIlvVC1kjd89uZnbSp2DZyR2SlCQze5PLkzrfSiXSvb1DLgOFUVYLaBZ28
7hF3NQHnjlMJEocOh6mR+Mv5l0dwCR31vCmi2LTkmZnh9xOUYIOyshZIv8qE5a+1wx2APmDT/Y35
PHggzwOHPod6DFFAkFdc+a77RZ4rv9PFNwwuR0dTkJP1HLRjzAuIGGOWgnvdLdCFF6HNsjUnSwa+
ERVPf+D3Qk5sunPTWStAKKpiavxPJ1j97fbywpvY/770EdKCoz5Unf5GsZnQcImWmlJ+venCnJaZ
p/Dmwc/ZMEkwhinVHktI0X2IzcbNkdetZz+DlXqsJKdYZRF4ipOHu14yreI1kp6fQuX4Z5ubMb6J
i8usfy9hJbBz6pHfiRsTPnKBPvJIDFV45K4EM2QBlVrnf23ScRBwy9YcI1SK3h35htxPBCrpKmEl
upajAUDcb1IDuYNqUqmoyB+3x+KY6NGmwyRSOlngbxpWg/THFYy2QaU2afuHlCHYoNn+Y3doDNSF
zmbkPmpPRRmPANDC8q6NLPdhGAudodTKp0naMeoaJJgZZXNt+W1VuXX4u7BYlbKiz0xn88ks8CZz
/kSMRtrFRW/OaEe9sdU9RT/n3ZZNktmJzs6vuFBeB772nEcnUdg4qtKirhHZKX3wbAJwqUXS553V
rc9MsZkQ1zeVTDEXDLPAvz7PP2n/2hsuqb163xO3pddYfyHP0eil+jqXJFkJ1TlVRWhRIXvUfQS3
zVfg7AH1DOAv9gQWNJCl1zO7VuG83EyOKmtNEv9eloT6x4TRNqRe3wfRN4M+TZcEDDwMrzSYl9Bo
M/gNRRyZUY3KhNg0+QYxkvlHDgVOwXUizBx3jXad96gHnQiyZstymMNncnSJSyPWes0ZLke1oHHR
1TZbA/a9kdp8+6FaUZFihW2vEzg/PJk1dhRVnIcbA19FEr3hTWtrpOkaZwyg6yj+nNd+xQIYUmt0
agsVBkN6CMgOQqz3bob7DEXQ6UUpP65hsqMmCJMYIrRRieyFmgVWZGRjZNGS8NcakeS2oQbYgGjM
93CFZLui5kJWqRPCYTsSbk77bDaADIq+y14qORbF4DwqVQB2IUEN5l7r+wcyo6C9bEbQkbnMm6OX
Q3hc2zLvmv6rRwH/lAvfs/zPQiPxmIw3AZ/Z1NuSTJ4///6gzc4DPlnr2BdRfV+tNVgnshjScia1
b1XBm+sT4PDx+GzHjAbIUjY+P1YlolAcKJlb96xo+WeEd7mffa5nzaOb3/CcW6uoC92WmgLvcfGl
BP3OHPF1Y6h8f4pOSPO7QleFCSZGHGTKXK8tCuRDKqcdvm0WpEkpIdv1gBapwoF41UJIU8NDfd+V
Nz4UjVld6gTLiorUvo5i5ey3OGRBHMHXbCA5VImlXD4bcxfkUsGlD5ePqJ5cmmE4MH+ZiskLor8Z
794JRxC3M1IVSik1R8u+MhJ/BqgaKSiCh4lNpeGEUedRrv+/Lcx5z/KpD3o8C8KIKPM0ryLkL4+0
cYVPxJ0Bv45g7JL8FtH0i6Zh2sNOJD/UbnHbZJudoxTEg3vRTqs4SlNk4YjsPG0c2IYKghACVrlD
VQ5Oka0pbVYMqRQjWIeXx5rBw/APnwm/WiEwa8lvoreJNyucqtsHfFlzdDy5+ex2cauRqG/fi4uq
T5PM2TWYaz7BQiWL2+aW5Y2YzqrtPR+Q+C9qFJ3J4U1dkSEqWKFymT1U5hB+O8ma9A11X3KI1BdY
VNmpgUVU7O/q/YTVbLIgt2OlBytQ1rCeJNOI+YNioc3q9aNFtX/JtPa1XQCBzMq1di7N7f8VYCEz
XqXLFcn7DLLwiTbcktyF03wSVrcRszp3XSi0tZyxvqDTPaa9yMKmxtmxjiLvZhYKQi9Z1JYGsCS0
N5UA+soleF2yLzJ3bNrmDFgsN2tKsxent0OL1EBtScRIgeLGcvqwfsk5mtZwYFYyoKbLJiohc21k
w6NZvYY8/2kV6QI4LPD2lkDRLYiTqtK/cFvYXMDtcpEOX/VeYlmEKssC96juCrWc4pu3Rnl/rRH8
FvaVlQmJQgTAzo2CKV1Ke9eC7m+K3weJM5zslu8QkTE6WBLJtpdUGrt1K6VD0CXn5YahHGqPkjK6
4Vme7394/6bpny9jLW1BfRkDYZqNz/da5JYLFjvrNlNCrFWn1Deq27iwbmnzVl2n+2hBvgcaQYje
Hn7zCij9kc4y1Xgr4bFIGjRFbbK33pOfA+CIFUdKK1rlTtW/qPRRuXZRsLiMoxOsvaKFXGCvmiRy
yVRnQPMpyKMQ4/NFqcVTP1gW5PrZGF/VGPzJFFhnKiUHP0kBYmpM+RoX76jTw23YAfAPeKs30iie
oXu646MwDwnnrYLhFnt8dtoU8B32S9l7mkKmqvMLstFZ3filQICNWD76v1Omg5q5eSaf56kcbwet
55CO5qX/5o3ATNY82rToqBDQX7Qudk/nKkzK2cK2y8jyqzi3gmWFEULGPFvIjbZgQe+3Cav3lvQP
MFhX71lz8NpUa/ZyGO/hB/QbjhVyKlIsOzt059qtO0Jo6NDAv/5pGFonDOO5lwIPPd8v//trenQJ
gj8RRC4TFIfak882nLb+lQD1aGUA5cQBOsnA+zd4Xxa7CLgdK718Jk4bj7g4GC/XsZxIG2G5duKY
WNtix19OaVA9fUvvSdSEnf4/Wg0kPqt0dt5ToniTYPq+6kIJvU4amLjWlVXH3CfNM0x74YaUU2X3
Dh4g/9oMsHGnRdV73TSrmadaGNrY68zTiONWLpd0+HSIRQeYZf147JbhOeuaexzMC2AGj21PXHNy
4pMbMNHfgDff+P1ZCy95ImOqYF0DqcE9inOgWS7lPfO73EVIYiz0ObWNUHzW4+jLHPT1JieYLct0
DG6FbP/T1ZjE6COv2JeAwzqBxOMywN6UmB9AcMUWHYR134aHiqDxFAmHT/QsqmBkM+vdrl+pSXzs
G4QTyx1dkF6iLKvGGnSWfrceY90zEgk+Wb4+dm5w9JZs4Ba2hXrNhpxrju0IGfapXlQcdMoqx481
lWd6ZQSEy3ZzvUgLqFWcmpFvaZMavRNH2yhCqgFx1FN4Zgx0rgCajT/DKUDSuopqrVoaWz4fnFdh
jALomz2dLTeOJzjW9uNLdmnFOxc/SDNvFmCBaZOncxFMLZVsw7Uf66ZjX1tNs0JiMhheSysefhma
LGpvitm57QZ9zfOA4jBHLDD9UUHeqSJQnJa6/gsrT/vibchRDqsz4koy56C3/5ZdrfDlZFCXe+3y
YzIdL7h1h3POMFT9t7kKcFxBmOO1JIhkTIYKLeRELX8lJjuxku3neqrzWiSu+kVxrW2Z9JeXtYm1
cT2A68nqKZCRabmXABRiMIrTLw0OwoIb8NA9Pda5QUYZOD2KRxetKsow4SUZI1iZfxaBVz1eyt95
fRdfeZ+rX39u3noUKLru3lv4Tl7Ig/b6PUS5yIVXFFqy5tC5adYaW1qCJwINzXTnSlpZF7hH6T5B
K/ZuB939eHX7UpRfX1NV8iCauvu55FmOVcrWcz96YHPISAuP2tvN46hFjymEkmyvtoE4qUp/IUA9
58Stzq3XCfs3nja5ZVpP5tQHyLYJGXHN2GOrQzMBhE8OJ+F0q9fj464US3i37usNSgHNOJynwt+S
NUNCZbFPqDB+Xu+/hKMFTVUeoxU+RIcWPX7JISz6R6Jn6ymA2Nm7fwg7RQKMVsRPZUu2bsBxJEXR
zqxc+Pu1o5LaJW0AEle146F2tNzIR+tik0OKZH6CMcdrwO1tP1dtDX1vnXfkYK/5HI9+kKogej/0
WrQbCydv+gdIb2dA9F8Q5zjnd5cfyKL6ib62HaOs+xCdNA/nYzDl2xeKwShqHw9+g/1w0yB55nxr
7NsdqxERDR7D8WeoqAXXiDpbVl3O7FC4SG/ggeXwHY3yQHNF5+DZiqJjqcANDNI7EE6+hLd35DaU
nE4wo//Grb4g4vPppOh9088mQPaJh6f/Sk1kvfYy6ClxdADZ/tnwIOb85K9hoHNxK0mRYT/f2uEH
LU8fL4WvJiQ6eJR/j8jyTarSiK2CWMciP9W4sBZrjMZHabFUauRYB4FECrNkPNIFH3n+Hskce4E9
u/tIHkqQ0mGm1ZhxxSfDt84/w6/NPz/BBOuhPRBbJx8z232WwQnT/wf7PzuuxHwIsQsl8YVysfvT
khztcLyDr7TkrGomv4pFFgHE2Dq7xZimAabs1ABKWlM7WjINwnog423fFuGaTC9F47WqlNSWr9Th
ffV9baiZzA3F8mWVTUPIXmEKicbNdc2O/ruWPGw+ofMZE2QQJWpRYXlzs2EJI7R5ywaOkeJb4Q6K
y/Erfg9tT9EiW51/rdRUWIgdnwf5T3JRTxYcZfdiMfk+NyjFrpwV5hFLEd48R5g65ox0iW49fDWV
vmIT7dXMVoJSSPTbJHjzAJrpR+B9YZvd+0URrR5QavdHRSrFI9sx3+c14UVdEeNfF73fkJcNgRYP
bMAoa5DRFHLyrxfInhmKSKdKZh5tpswxZFpVtoUYrwL7YTyhyrHJShjpOaVYdwC2vIn/GRAgZjXO
I4jd3orJSiQ2Zty5ML18Hn7OoVVBLALNpM1XcYQzsVRE971RQULwMPw49TkHaf+4wk1dDBY5qV2/
XH+whMarnwGGNJr+opy82Z6X5M3TH6x9TD/GRPzzQe/4WavXUgYGct9GGRc+x1/Cx7RXU4K7hlsi
UaEaCXDf6pqDp1Vyd+aAD1Fu5S0/FR0Pf6p4D7FyFy+A21H6KMa9+Ag7Uk5vLDn2SxaRUV8wFmvB
PLYtryVg6O7AjTF67VXDy5udMBTw69P/fhmCjp7xbjkiinSh54ZvpspSRjDjqB+iTH0aCw03pVXf
NmoG6YeuaMl7g+nKLuGONq9ZWmjgjuWDWJGVzWuAa3dsUEOc3XZNWtgSBytmL+eQi2bM1PLO/EWe
ESpZJnoyyBfm63mhBn4gP/jiaMy+26Ic/09uNKWul5hgEg7599o7i0+zmBnEWRRzTotQ8iWOicsV
0vzV/F8fW3bJjOltCq6FvVU460siBK2v1ucLLumM/dQl9yAlBFm6P3v3sEjbKLTc6zV7StVJZ8NR
c7yHj+HbUeSrOoPDBJfoKz3B+IRecNAwcGgQXCxUFqabjd3jhjonM6Bj/i9rqKVMX9WgJuPeebom
y/mSLAercn3Otp3mZeoOj2gxppgdC5saW0BtqEB1Tg0Hy0yVPps3XnO5Eq4ELOZ16F1maV5h3fdz
TJNwr8kh21G4QzcsS0dV8cNg+207zsS07XoaV+DlUZ4AFEhEeedtmEIEc1z8GtNxfclMXmcVAPQO
FSfK5D2o1Rxd7avJBaq9vThubwFq1BzDrGtzlsLqBPPTx6lMgvt606SZPgAAen+In9tM9YOZHL9I
eMCW6jaqEtgq8VZ1659YSSCacpS1FdNLMrwqT4o/Y5HJKHEntMX6Cuo4AnYzqOiZPeXLOnKChcwJ
vXlmyR+XaWmb+Q5qqCv0wcgbVY6Yq+otmwgniB1IMTUqEarQuis9e58feS8nu+S0HBX3OeqMAPl5
P7N/588LkZWKkMMlMKxQ6QxIETF+Q4BHlxNSBcZX3cwZCNCQwgLELOPJoGZGRnpE8F6XhbmDf09M
42RtSFu7FBMk4uYkASEvEe2zqJ31CEiBfBmr4Z/m6C6MDq8ahRjk16wtfdNvkHkl1Ay8GoJK+be/
odS1dHb8nKCLGzo+Qaa3Y9+SPUgKNJEqS1POaxsyflZXjUe4++0T5VAlXdms2bUuf8Bq07zJc5lN
+cyzOLET2GU3XlmAPGjFvIuw5VcvS985vWWaqClJU9tFPqZ3Zc3CZRKMaHhLQOnb9BJGyKiqUPBW
d+82TjywEtEUDt89Iz1O+5xkvGLobmfydKkRFp6qOU4WuinRZ5+eUBurKHnLqQjJ+zK6J99zPXgY
N7d3KAPrtdrTiefxMR5Btu3am/0axwgoFsMDjGV8p25efZaTFNwlPJGWidzOl5ZrKjTnF3LpPxD5
zBLRgOkRz3Yo7cfnpBW5tvljEIhE4AJyktWc/tesBfWcl6DOTtYn+eGjdIoWAYN/RvQ8tV4/apeH
7Dsd1A2i9YwfdfBJurBSU56ewuyVx0BvBiEvcFo7Zsn62d6wrmCYotayD+pTUkubn5dsqQ/7yS5z
foRHLbd4D9SwBcwQGJS6QpCFkvibqOa+nWRKtJfTPNzD9UVK2RSmKyeGc4dtLRolWxntx+uPPNFy
Mnnlui7ZzC7uX1OUBKZ7sj8P/OE5RnTitFVozxSZ5q5tLZMtWe3/fpc/tsaLElUh7YbEzDL2eJkr
Ce0DmR1jwclvzZoLrXo8AlWdeJbVpGTHWysF/Y/CrwvaUBQzXKiTfVZjVHp3TCiyYNUvNs/+wBqv
0DjvmE7r64mxv3JLz/WtfvYVb03OBf2s+r2uIAzMb7RQAwLtfK218X/V5ruLzPXGMmcyvwfoeMBd
Meyorxbyn8qWS2fJ2Tztor4dsGlQ13GdkM56NirAjaqhAKVj2Cvfh9IYPoberERfwB59vlkxwobG
bkCNPCYzLyWD0OGoiWPszGLeZdwOjxbw
`pragma protect end_protected


endmodule
