`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
iusoVxay1geNO/cptBl91PSzO1ZBrPNdBTsITWoL6/G7S1hGnAkqIsC2eKWvJUOEoN9PztrRj5j4
nkxFL+oOao92bXOzzxDQm/vfwNZsmDUJkoSa4Ytzbtw3CC8hxAcYgz3QLAHEpvx6DoimV8jbBBk4
W9VNcKto9NKjt6zcaOud2ER0SiXVCujRtVplZy/huN0WvpFBG0CaUW59Ba4X79onr/4U1yrP+j/w
lP7oGtds4RvMQgk0zw0cKGwz3Si7swbJESlma2Jez3SVgYEcXuZYYYtD6wOXzPOx3vvzHeOnnqWD
NndtGAHCs4esgYF6dDlVGbdpGtKAdNYnfxoPXA==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
oT9QJJQqRWGoLobCMzKfgCz7BH3SD1mZ+kTg0VtosGQsfEm8/ZwkcxuwdFqU9j0YM/DZiFHQBCuW
DTq1pbjFo7P+3ioXEKn/X0fCBBCAr0yd5ySVUMqYIl4yGvJybRY4mWgk9Vq/XMrJUvxUKASe0+ip
kxQUUABkd7LPx7k3uKc=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
T7xbJLlEvHo6/wJ6lvoP1bz8Jgb2S0WErwhThpJUvPgQJwbC3+rbmMW7F7gVxhH4pJ+XziSWISgL
L7g3+G5809SKwBDyVYbeXTaFSadO3kp1v0w2w5bQXUT6udn5bTTB7IJgzxD69MYaY21JRcpT9Fl8
xemwWua0Y2cShuRIlI8=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 135648)
`pragma protect data_block
GZcnHV/b/t+uWBM2Gs370IMe0CgRWBvevQHI/Drnr6XPQofLZAPQfp0YWDh4ek29QJmwUMQYjLII
j+SVpmzMrKDs5ry0Pc4ewbkIiWwxyqByg/32QcYWVHRwKSJE+s+e9vqf/9QxKsmCv/F/fW4LneKL
7ARp4/LfeJxsJNdEpTrFAk2bXLrWdABISivMcoWJfnDX2kcC413uRpfJwkMHr6CpEOu5WRJBK9ja
6gCGV38QP6i/sGYbA6YeAxPfH7PVV7a8TqJoOrsLkgY5tFgo7lQ4lKYyarWmNi7EUsm1/qb8b++P
4Q2IoF/nfrp3V4zDU417dW0e+II+mXY6RDzNr4B2LgZ8wY8UBXDhbZxxHP1I0o19AFXqj9d2yErz
kBIhRLUsY1REpEeA1VOXLrg6v1QYFL3ISsW7ucuDvzySzRlh2fu6T3YUVxrf0vXdpKkgVwfD29S4
mseurGoA97aQxBLgvJ+ONXFJs2aeU9vubuRM7U3pwIlTWBxq1QoQiUaeDpliuVUS6UznsvSX+GKe
xS5YIbSCuVvOxQm0Rjf+i4xM5ho2XfBTfHmbEG602I4xYT4iKattuVLUSUrzrBirGcUKmjL5KEfC
iEgsn2Ppueu0/TyAcE6jCveQVlatEpPByz0DPI7Svvw6uEZyuBbZGxOg3Ht2t9IMSH+8Uj11ENFH
XzbmFnqsz9Er7oaKA1/mJQ1wJhUWKyP5zQHcvk4uPyLcXNvGpT49aPXEb7GfD33SsVaKvC6BXMTS
8wOuHYLD/68lNxp+SXiucuTthnyNEK4rky64hi0Sl4TXs82FsNy9HoS1jikYmeLKwb8N0Le+wtJK
PZ+1NYeL+W5OH+XzJ6nVM14a2kra2Nju0SlcLVyCTQKmD714UshrF2oWMJtXqCJV1CRUylDq9JXC
o5bJI/IKQm5UFs/HBFD6DLwiyeueDkHEUpFJCWS6GK0gy5ELY7qbLLLjTIId8gH0pKgKMo6fklKC
2zoRvjkM+kF32c5jAER05I9ZmAZ6dT9ULQnv2w/U2TOWBad+GMy9dsFP/Y5BLyWLAygLgFCSq/Wh
US+0u8lTSwTiyj70/9wB65OBvPW+kWZOF25/UawPtZapvy7niWh6i/nYhovr51xyuiQy3/Ggr9Q3
+MgVM2Zvm/xsKYi9P700OMqkAzxNLIV5toRDpxrAJApy+7oqKHcKeF2YPwVNsoHTwf7bn9m5ntFY
Wlpde0zcFHRSGU1PIQE4mMf2J3FUBYm9QaguDQhnUAfq+b9j84HVWfxPlKGOWOhvmtWrJ8j0WSIc
MTiAAhtYGXNuPzBoxBvgH9AEHKtUU4xAlvtqttd+F0JLRw+TWXMbDgKoS7NAEP+Klr7wkiB7FaTp
clIznD/ZLP2UIYvSWRzC1odH96z7VCFw5FxVeN1u/Qryis67riTEXrjm9vGNew3RpXf5EUURSEWJ
hKwL+aq+5K2qhgeesS5Xk1fjxgNE+RZiMNux0Txi7GRl9z1H2Mf8NyPyKTXysHM+ahibErNVGHn7
OECxkfbGUZxIlbhQpKbQPaOYTp9+UWCpXGdl6Hg3sQYXUIo8pu7tSFk2aMRaO/MzfubwJdT+Ml4S
BxddeLPZ+pOBWij427AQw9LTfVAVs/ykJqqwZU4F0gX2cm85LdX7yVEubE/avyBBTv3KqkFR+7B1
HOYl+7QWAnkR7dlC/e0Yv1r43I1E4qVQlAbf7K4fOgKGY4X9hQgbAZEISu5zopnymwbgLAwsfLN2
lrGSl5zOMB/PyaRt+F9DwIjBVWG4QN9RqqlB2gksRuf48FEydSXqKRzjysmvNVP1n2aaKWp/x9+J
vsbmXXGoaKlFGSjjti58mOAvN6zdluJLFwrUaGDJfYM5yBDJCNDdeX2vW9TaoTM3e/v3tMN5wqc/
dLTHnZnvwgB8wYSUjS5JM/awh50AM7Ni+NE/8MdpC43loYJgMDigkT2BZAj64PXdDeHe4fvAOzqu
/Ie7gP9w9+/7Cbz42q4bunqz6IRTM/wdqRTOmC94okxRxrlJ1+Erw9xdRPB8pV+asJ7SASGtDzie
IA8Nb3P7xGsQ06clEfUSvwIQ5deE57CsS8InqUnBYCbfa01dPFKP8qxN2WtEoAaXG9/cCnbYVIPZ
BmYB2mljDTGaLaeBDvmgJpaYAArNdsN1dmKjHDKGzlTx2awbjOepbvjUILrWGeaJdkuGtucrUngN
2Yf7LGNe9/bO0ixYv5T2ZPmdEVND78eUE/RAPs6rQcfd+PKhOEspbvhW7dAGkMI9KBz+2gCXVsqy
qbRteeQJQsMlmnYTXSV4o8mub2fIs3xiRIF/Wrn6eO4KW2UJYuHEDA1gc4n0HK/2FY193iUlWH6w
SsrHqCjvdqwrBn2u57JxjvT6jFpqgBiGvIVzEgyQKpCcVjRnzpRGxx7YOivG79Wbg+8Ouq31OHdw
Nz3WTGRKvLnthxbS7CxNyS5vBYDF9fYcRLWcwZHALGNDx+DWcz+57UI3y6tfEFZuhyA7YmG93AcD
JgLj7FFjxgDksUmmjcrxz3obP5TvzdgzYFgNvR4npNidRE6BF1xOCeroAiHR6V0LaqLKkeH0dmtz
jBpIph/COEsH2pqncJj6xRB9V253/so4P6U8nq+zfmjz+6jECp3TLCcL7lJpxgs+foTakreei3iS
OxC3FqopzwIPRzuP1IoHg43lt1EfWXgYP8m3hXGMhaXY3w7Ch/KTEk1spBULRLgROb9DtxCzsbXn
ezm/TcordZyorVgeXbk8VCzVoyhTVE5wwqNAILK4Ekkar7YIdxGMOtMrQf4+vzwABNQC1tXXNddn
nxvfXzz8xdLAv8eMe6kzXAtY9zmdTFfKgjg1bnAFzm2lcxFadAGEB+OXUr0NA5SvTWgRFCGQO2ey
0JKjDtT/UEi6MTTUzRaImvUDnhqPr1zjUumrhlQfyuFFS6SSZUbKS83UnXcCf0j6JXl9lrJxoaZ6
dijlZRJqu5PzxrMsEu9Za8gPhocSJCszHWO1luy2RghsaVVugwsUMm5JYzq8GS4pDtoPj5SkDlSr
HPgoc2X6FpZAVBh7LJO3Zv+y/8pjiFByVnJRUoV6gITdJfu5Fe/xDh6RZHnLLzxGm0/rOIqMfdjt
qgdvKIbUprcGNCxdTUF2pi/d5Ilmaoy8bM0rh1tYkZN7LSam/PALjrrEI44dLMyAhxaUzmtTIRtp
AdTwHs3bz9cg3iFqATZ33vPj0JwkCTnFJktFr0INRHuXQQbDU3LD2344BDXm4272rUj/kW0PioES
DmLrYcP14DbK9HeI0dT/XDE8cd0bjzO5IYpyxoi8eCuR0ovZS8h3fK+xyHJHGMlGoWe7i7dg89YP
rzXjmjHQMhykEA0aOp3NChewG+B0Xz5xJe0FEYps1k4p2oTYTtA2VMDETSuKL/lkbacg83bAcEY+
VmVe2l4qiJOm5r4iAAiTtT00DKUauAYCeeSdFMVehTkGkIkIaPajJT17DZsDhTTNN9XNL9SmlRSi
umfUhdQl3Plbizzaf1QE5ShHIBC64oYWn+AW/mfi01AqryBlks7EZdSukSbGsEpf62A+nBYosCqK
2hps0BjsCsnGbl3U4QMR7ZOjPrsRjF1Rv+4w1uEpN9lvwyrKPTpHZGqwA608iUTKggydXfGfoIRo
U/1V6SD+js3K0F2fUp/SHClBcSRVBaALJl/LFTLr2IL5Fuh0gzIKy8u3PAE2GOCrv++ur7AsUpzM
jogZXW/5kzDwCwGafTFaQmpMwZ7XWYlRNxBs4zqQ8SDdomyb6HpubLvFWhD+3q84G9Xyer+1IJZj
z5e7TFF55DWvEkjrnPgUeAhe9TxQifcfhOcSXJZhrYnPoJ/fHU9cac92JBpk6HbFpyrJxXbACdMU
zY3oGPtaoB+oQ5ih8hP0wo5HyQpm1wYmO/xuNWe6N/5fn71m12inn7XOU03R4dJ5dRoXc6y6e4Ci
Bl4oqJM6tGvCahGHH7Amfuv/jia/gPCbdCcdEIU6LQCvyu9luTmnZB5VBxlpwndd2aU06aFxmJLe
TAWWlAMZEULX31+1+kjmQ6h3MEuJf6utkWsZmSrjr0Uhxll8J9TBV/ltd/+zOzgPfapdORC7Qgvs
M2Y7AkR8z/blMHVQJiikmhQfN8E/W0ce34qtYe4zZmsgkZ8gfTu6splCFxnMOZRrPO+ZWS5gyh4V
1E/ZUZCZBeQAym+e794f0UPQs+AiuC5Uo4YGkP87ymvDRBnbCb7H4MtPqDoSosoSyKWsXKarKrCx
wLFJ9LDB0gJiKgpOx8pdSN041Fp1x7Pm8TZFRjVG6gWcQF1qNg7MwGIl5m/1iKf5I/zbXy9fAe6X
3NepJJRv0LIRl12Zs/g+uOPgtARpmMfOX1c+GbUYLurf7VRKRVPxiq10jT3SfkFEdAfoN2nYXlIh
a4J/A+6DURT0gfWrtto7dEINbNZ3TB8tDFDuwoln3D53xy4CwbtRFg9kfwy6St2uT0BFKyY7OTtw
Js690/low9amWLSdRp6bLzZVBjYGQeyLj+EoAxVnsDHPwMOCU4OHrB3Q+HdV7Cve3b/FfztHcewQ
/ZpRRnjwp8INSumxWl1XuGZkBsP+ZTb7r2aZSeEXmeyGkDLEKVCTLnuht0dE9IxEXVHYWPLPFCM2
kR9dllsSSxTDFyUqgigI+1WhfwEqNBLJxYRiWSP4mxTNU26gQDV9Cype09LjZMNwJVEs6mxBwk5f
nhSjENVneaiSy7lXZCuHPqlHEDX5Z/lKNI0+wZsnu8wU6RkKdFcvpSa0viprCod8L3LyLML1zJ2i
p5W+ogbZknXLo3UPRB91OQSt2VIeOhaP6tozYEdeccBcnv5ACYZSGT9ABOF1lebAoVuDyTSZ6NaC
JuaE84jOBEQrIVxSIu7j6ok3geWjnf3yrTl98pc09v+gYxAyiyDzRxzND7TnGJ7DDgOIQZrddS0L
sErXh6kqjCFx+FHmRDGjQ64wVPqQoWrdp26o3v9NHZy/9piCOHeDImKr0nv0GLyi0sjPYUh5WX41
GvqeD/nYab/Ulyufdw9CgsKr/gEC+6UgWI0/NmYaCux33Ctj1bPWhTjwDoGSYHYOtfi5PEJQ2Fwj
Yob3eyTppDCpg2bZpaoDhXN+hTUF5LTRF0trbL5B5biJVOCOQTTB1rrHcHdjyUIRnkUCvUt3kN2u
qQ+otL00Sx+EN2U5WsfonOmQv7YImSU6WcylU4A344o+nELz42cVHj7ZDSytCWeqM9DHtbRZhecG
k8QsyZwFP8G5gSm3KuiVOjIMnxehUJUSt5NOSljsIuvvW73tDZHdGAlo/BptO1adGI6jq9+yMmdH
qsI4EemuWs2+cIq9AuctRGsuUpWsdb6odrQ/R7zQMKtcSGzNyQKlr4W3bupvxemZDQtnr8/DqdRA
gfEGLhtJ6KTKE4+71KJFAsW/Mt1j4iYz3cGV3woaj3n0/HPekd0LcNvQri+qA5Fl55WdixnnIfKd
6NNk/OYcgpAPyf0JT4keWaFaCcjcQzNZOImjnpKCbfQNrpA++4loP9TF71WOlp6XJADvIwwx3K+0
QjPVypzoUXzVk9c1wEmeGjc5gH7NdSQXUu2AwailpAtrPMOR5t3z39A36LSewQxNP6zfjZ9uxcsP
Ikj4fkl8acZMPncLS/1m3AzG4WfZSFWB22PNIk1dBte+qj3jAPH6/OA2k8Z1458Rs5JK5GOvHo1y
bklxz4zXiFnW2AT9oMd4tCCsxbS3wcn8omfc76LWiJlJAEpW3oUSuX9Fki8VtbJtlarg2UM67D9K
xoqRmRUQDhHx7KD+rVJB5gZlwbpzPTi3Tew6IStMBI4JBZhfxcqrmB72jg2pvRxMf5giNXEb50tV
iTtw+fVbK9v/4lCARjF6FApRVJe6cNRNyfFxJjavA3gF4fnWJQ9vywk+6D11R4gwGujdXK6cmErh
8sl1AkfITiTCQpm/AV4/4vggCDsyifishpi1NPYcMOjgJbUL9LOhpyznsxcAxswa9LuW+I8XmVkq
y+Aukt0HRgImtbSqvz4yn9cPqEGxY4X60w8SkCzWqhiTdYTR8OqJSAsUfFyG7ryTlTq4ysU1NYZP
3ptZkLixy31LmPcNflMUfdTY/170mspiJN14S+X5B/FPgQBDONnYwEhgx7trVA7EamPQEN86+/U8
PRYp/BdwxuVwe6Qcc0ysUC90BEo85QzRCd33cEYUvfrt4dIV6+i4KO/kZ/bcUBJSYiTKmw9kHMx4
UzOvQR+hSCDK2uFG1/nzmmYpgHQGgSIkMIKpOvldcHTPeYMuLw5mNbhXKeLpS1hKDThPf5qG+f80
FdaCXBQI0iJjxQzZct4sN4I5enzCSVMTqDsnjsGGSe/3mrnrEEFyJJMGgVLtFgF+tl/AOHG4dlDM
GkIvjXklj1kYSy+4zJ6n2iGEx6ZSkeXV2RR9MVsBa0kEK+ArJrdPLaIfmGIoKEqkxwSGvnQ/8uGF
QfSXtDDD7SPp40Tkq5fSwglT+zcsiLGxg3lXwCHEKw+EUgpfR2IE4x4kYi8RsI7+Xrd6Kx9FslKT
5djpCPusLrHrvp8t9cYCSoTZiTKxoIuuzHfJEdoG+S2ie5jboxDxzPzFt9Ms8Zl+RSoDUOxM/hbu
H+mrxrH5GOpMbONPJ3ldQkjqzBKyM6qfMd2CCxiU6qxZSJOsxFJ+4MauEoShOTC8O+4fLdzrAbiG
fgfEbArojRB7x1Rako2nhX0kcMF5FHe0yk+cmD5xdqMvcSbfFgUckkC9m3+M5kfwysclcN1WVayY
BypPqhDZOSbvGijKURXlowN2jUX/hYQaCMhdeJq10h+Ea7BJ1OKaEeq8Fexb78/rjcDdEgwGbKT9
k4noAjCmIoSr+SIEPXjJsCXiT1NpwNOE8i5eSQbjc2gS0nKelzjhEDaGX06JCsqGx5vVT/DDIYlP
DDBrZHSkFMyJxQstG/Bj5tPs8HxAdMxcZGrwpTRsGCivgkN81HXaIw9QCBU1L4qMBSu2bt4sBBsP
1bhqKcgOmeunEKhjSaR51T0CnLiYhHk4Ri2QTnISCUTxS2YKGM88Z09F7PVrNsqqmhrue1DMsnf0
WEhxWaNrqqfzAy78+nkmrsTe1AfnOMqOMwxEA2URq86X5lVc20z+Fe/Lc6TigIIBH4TI2OHMbcRe
lWRhFm0VR95BlozYzCbztoa6Qt06uRG7ZIYcScsPT8RpqpKxvwIY1ADKCGwKqsKkIB2orqsPZYld
mSLc+DLghlxlDSbV0hWaU5FzKOYfm8OqGuBDZMLLd26CBaTRog6rXyKJppu2FwhdaUc/tQOVi06v
bnO2imVGNith93A37sj5rYEprK/GY5covNIaGJQqKMlI0X1vIOqKp5Ookmu4/aXjpAW3/S+iRN7z
ivFnLhE1N1Vdq73Lf9qLdE4XEGv9COaQJ7zu8w/udocMdo1yvDnxZexhT8S/hizykD8KkCfy0P0p
Vcil8UtDpuBgWSFBwCGxvL39QqT6jBhy+X+ikWLiDusbsPZaE+Wkl890U5T9Op2Jx4/AsKtLAIi4
O+qYoBlmjuDNHBn/8B1UcTidvhsg4/5gK6o5F3fYG7sXsB+ZxMFEjgCeIBTCJBi+FURFIF+SNLMt
/zaJA0vmUJDcN0udOmH4UrfDQ5pYwkH8NeTqpPP3eYb0l2X0FcqN2UzVbTH3RIDNqg3qMUFLABRs
0fnomS37QMxEN31GNs4OtUtVg8cqALNbGaq5Erd8qkHYdjCAQILzlH9NWl2PBR8bIrhClb3HINcX
LqUq3tV8aG+yVTKnnvEW+PcGB0o1VYZLRBn8EbSg3e3pPxjoPoGMcKobqDkI75S/0/vROsMEv5zl
AYldG4MfOoHAMNLs2yQO/o+DdFw39oTDNWFmc+D/n5fpFEfNeVaDijUQsHrONZvDyHmSsM1cMaRf
nTsrKQMxLX5NM6XtktUwnbOp8kfJImN6rWCSor9Xy+XACqJlxMZbH6erFORtqTYW6L3KLxvNIepb
OWpKsbm1opGK7aXOOSLiXQ/nAi2bN78JEokzBubwYcrXxvp74BQaJIURb86FHvhtdy+DeqZL9ric
y2kECAX75SQbFDCcns1u66vKWbYce407prEKWqbTZlEJxO7Iyg+jWiXIdCI5ZksbAHacpOTUQ74o
Tw8JLjC5jKC6HO105gnbRlFHuWf7E4msmDxeZAVog1aVoWP4qGzUso3kXtmGpgUpYub0ZOWD2fxt
Nb5h9HI5BMNl4+DplNbFTQVbovStXPjpxXJJC543mluyuQhYihYWH5zjqcs7wT6qwsqr8e7PizqL
3kqO20EGatatDtOLe4hmIw7jetK1ruD0pt/fFiJjapXXYbFNYaDO4maQ9FphFN9Is/ubpwzSTljS
mFEYPY05BfcG+DZMh9NHysqJMLwfQ2/F5isWqMYtykae6LRNYBnYRykr+qo6N9ZfU8X2G/8hvGkv
ArtN5KTsGMG3pjKq4zA/Ly9M69ZmyuH/EcYjIiYS3wWSgoEwiWRtO8VmPhnN74TsyX6k4pamKu8G
dyUQrQ3tA8KIb09leLTToBxNrVwPPnykR0rJJGYMI5X+2vNW9hxPPIFL7oLmxEJYeMUN0gqsLaN4
eLN7MHFuv6v/Qs3/Tc38j+BrB1OkaNvPN2VCEyUPAbMh+sfnCcPh/SOtcCTrW8iPtKMQlOZ0a7Hc
UN0LOlQ82JUDXOCyPxJ5IOuYYz5QFNMEQdvJewFGdogZXR2CZA+pVosQzEICAqOE4ODhjWitOVOT
pNPA3DMiY5psN9Sxdw+MHQM0d9YT2AcqPF39VoJlcC2HfA828Wuzn4a2kWatRDaEzGKwxZBfZi1j
gCuboL4UKb2qXYP2Rg8ZMAeP67qVMhz3qhPwlpPxGeMgXFECMrvZYOpfLiSTxiNHU/xKn9/Vywp7
QIxqq97OXWyL54xysgJBGltcLIZ3CSzoLsZb2jMZtUG8nlv8bIczswjyQX/kHkx7KCXWSSO7OqDK
RBuJluALZ8gXYvv519IQSR1aBWLyiuricEbnJx7wUGPMQFScHL7ds+/gVj7KEHW1GCZr7BrbHmrl
yAUd+EZWYZiRphJm9SPngisKrMc3l9+zZuul2XSBkle9Z8PFnQA2d8cmdDZ9nAadPlBO50kI2Dmm
pGi8HzpGusXgAS2cym2cfimqSwpqH25T4AuRTO426f7jFu1IM1eX2GN+0fTFH8ow9u/0V526Abs5
wci7g09rcTJodtVrW2FP97ME36zqOhKbJrbeRjOFjTcDYzs6MLEeZHkJTpWTmffAL33ysd+RTzsV
GwioOZ72O34fBDzftV+zAf4xrZHu/7q4WmFdF40krQPmdZQI76gwXqJQbWze9OMvQRINrEVsnoAQ
b6ihoazgEZ3N2CDKTtb56m1v0mwBl+RvW91wbFgKuSi7oocmK6mhcozWSxPivYS3Aw0jyAApgrsV
39CdwlPSx8erV501bA1f3dHb4GAwqkn86w0Nz6ZE01jUpw1di3dO//8/4gs6gbv+/AoWegjomQaw
jUEvL/IrKLbj/Q1inl049U64z/ZKP7scob2xLxWY7WwfzkM3tNJMT5XHOhA2S0CRV5Hm7suZio1z
uSmJht1PUrbiH1p8eT3yI2I/DNGIEq/ZrgkPl18rRO4/4FwIu2qVWFdr65OqrGfNTpnlTWi3dlrt
WaEJnVIWdMrrlxGDx9unGliDERf4caIn633UfJpPSAi3K9gpnAuYew01lg/rgu8FuF3BEfqYD8GF
+5fzi+qj5CT07l5Y+fw8IfeNVyXiDRRgu6jjJpFY11oi1OBedbF3mdv9JjZs+HnnDsSaLpLUHoI7
Dmw7gDVLQRNo+JZ+ndUuGkYbHa98mz8mAdy+yUpTxU0DkTSvLfB7hFXk9hPqEbtsAHDfb0Gijc7V
iw2Dc0WmKOBxcfzyc+23qdkOW9lRXuLcEckKEYbGv+s1pl1W8Xa7PIuhNWb6GkQg7bp8hMO+oopd
9u0O0JIaaNn8uzDyP0HtwJiJMYl56RG/OrGCwkVdYy0WnA3N1HpqUHyJ60xU6ktafAkBtmQH6SRl
pesSuxWjqNjfj0Zxrn3vk0sKJLa2Qcks92gcLFoqdmdNj6TxJnu030OjJJLtDmfqxTAkZj71msZG
mwXfDhrywF6RCc9K8nDXcV3uv8QEeX5Ze61B86xcnCuNDfsAWWtPaXAVVlTONADeh0FvPefM98Oi
7a7gqeOh7UC3yjjnqh5Mzn2WQ8Q3+mMZo07X6rBH682cuZcubTeO6mAK5HR+17Dv0IvOfA7qJy4s
ge3gKA/sTWw2haycP4SsV+RIhLgX8EcJv/a3kB+xpFU58yeISDAuuKoKp7LnaccBjQUEfwKVNm7y
xFe1APmI1JmeH+2BWMOsymfqbQ7Y1h2Bdsze8KpISr7yY0Y7r1m132/zcwEoMfmr7Fbc42EuonG5
Lb2Qe1du6L7MLWI7FHaI7tP3Ok3yTcr3ZVLMDpiHr40Z6QWzh+aLh9bjqLCVZXQmBzmGmco5PLlL
Dw1IpJUEjDW/Mv8e1GTqahF+xFwgL4d2oE1e6NEV8T5zvSCTac5ODCZ6PaIe2MLN2pdxnUFJGDqi
EFGyDddrn3dzaFqIbhc8rMcCAqnStpO+x1ZpbxcuAsJkqdaOSF+D9zm9CT+q9z3oWOc5SCN9zhGF
o72gYBSnYIUUoiSh2UUq0Mb6vxEZHFmj8oRRyGUsSivvGYITMmhNKjChcNmpDcxhZZvB8VHZUlB3
RBE24kWusjvbYkra8zOvuMPizSfTf9WE8DXyjXIGMOsvrn1/AUqDEiHMt6Tctmsl5wFMMtzlD6NL
Aq78SitEqRloD+1JCFzInMpbD7hHNhwar4rHY0a6t08kddNGaDvLQPruGspvBw3A66DLoHVqf+8K
RYaGms/7N0smgrZ1W8S8CNCLimYZrDhnQy1ctEMlJJZava69qT7B0/DyBP4wk/7H73qEzBDbBBrd
wV1jd1iN1rqAyr21vrv9bE01IU8ygIPpYVhJZqZSuKuCYEE24RajSHRi77sEdd9vrS+lXgFbIzdm
cr/NKntyAcA7hMx+868lctMFk1F/OimuaDRW+6xJVu8+h9RWGiT6ERqSeJ9C+dI7/AVkTUWdEdaN
s8dXwYj3X/kz+v0V9TCIDTYWro74oRYd7tHEb/ca0Q0u1GoGRTLB0smkAeNsNgdvL8p1CtxBpfUo
W1eNrwmYih5BflmopbGnHz/kukKnbekxm2sbjk5xWVtuDlF0FLjdcYrY5hXec6ZfCKAQSzaSovWo
jaXPxxBE18oeCXk2yet6EeTow25V1Mx6LlnWaIuvTEwEbSB3e5wik4/lhD0mnqLoEKl5JPPQzogu
D3K8jkTCY2zCVYYsNEmee0w3RwDa6keHZaFUtJ4UUe5uJuB3WCY95r7bwfQZgpuaWs3yDxRJvZ2H
Yd8nhoOQcQRjPvuSvmS5j3HUycgz2lBH+NbVFm8I7UW0BqQVYc/GnEBFDlWZnK6EoY11B6ClPlYz
1cLt3mzIP1zn9IpYhhBjc9DMhNCC9nIC7YiAANpXdquCChgEaH+UkuTi/Fm8wHjP5N2cVVmxV++f
m0cCsAZHggKMmpP6xqKfBKUOrNN1sdFr59lCefML7wv1jwWxVWhTYhv4xFetvSpwStyUeUxaKvIN
fjSv6j06r6fkPrGR2Fg1qYrqzvfdPOnPIH9FG9QczNMK08ZoQFmVgyQwsMuidRByEH/K0arZUGh3
XLkzolEAKtHGCWNUx2WJfAfBHV6NinpG1QWikjEPV7T99WzraTsRV2OrJaMfc+sRs1Fily2+h9KY
78eaQWL0+aQutnl4/fL0FKuLNNu7lceTRia9WxkhxetDslwABttuDgZ4MzeihtJbc55DGINkWdXv
WenGgpKS+BUGtAcyYFwxwi14AhUPe8ZLJAZck9OsIO1scf7Nfgr1cjXWOEu/XxiZs6tR3baAlMEL
iKKvdLH76+Jh7d/E9jrcIuj1IMzoL40UwtWtxTMm9AXZmDzaN9GdrFgVZ3ETyhQmCjO88Fr/RHjA
YvJN36T4ztHeTdNx6xDLKNrxWrxWS5wYVICyo8+IQ71oBPNWZHU8a1kcR4U7eCQdgTyTVekqKPj7
Qq6CQh3TVrLH+NmKo4DrosWqj7OOBnEIEK3/5ZcqhqdO9yK7At4EFzbabSjC72ScaRUT2BWZO4V0
/T+id3aaKPbGZIL778BUV3FkBnQCowXaTidTIZDz3UwjczEd4980id0XKcWZZeGymmsQnaEpT1QI
i+Ysu84i46at1jbD2oOy5s3ykvo7HOUTCNh+Sy8bf0Tr3vk3kUl3clbFz0cwXL+ca3zq3x8gcd1T
UuhC1gu/ZhK9VQTmvwXHAbrI06cdj/yr/U0YazzQU9YXPbFdqS0je1Mw9UPkCtl1h6hTL9ZhYN33
VscnjQxiJD+qLThDh8wY7GNaKGVLwzvo6gJW0eG2a/ZBpYKR/Y8+1yVkrvGAHPScfsdv9hP5fPiv
qC1E1dagI2EbqxoZOtrCEVKyW4FYk7LOKf/U2gZD/6ws/VKGkll7hT7VhOaivt6EkZGv4kOXRJ/B
YEkzG8A64CtXiPlGFagJdg+S0Atl/ZaWnId2Nmd76Tn0COw3jGoxHyS3yqoduVRmhXFw8i/A1r2Q
HfPtfHh2+knO9K76oli+H0MH4zQK1SrRIMMOyHYsGipCy0lm0cLB0NNA9HNwa7wpt6JhlsZZu/kw
061x6WGQ0elhqcevP8EMyZS6Tu2NLyAsWT+8jmx8EMPgmKvPmNKDh86E5uvFpV8XovyZSCI0TMU+
IQDeC1tJag9nCZx2hQQxKqD/KD+itumVINSGXHKJ5mNVRVcVrG2CfR2isBju8grFFfc7K5OMguiJ
J4lgc4PQi7Mmhkg2UjK1d3wnw7NF0JGJSZ4hke+mFpEzowvNZvq7JmyTITscsDm+/qADenzcNqZj
u5TUiYnQZI980tiWa/ycQoCB1LkYzVviuj9+pADBTzjwv1PW/E3rrxRLmYwg90dN2UZMfMxmQ+vF
5/yt2R3pPDrNreezcfJSgrCHtRt4jNPePSQN3L8s8r33TOfsvlGkv3BdJwfV/XUrzakZDupSicrg
T6Cia/ZSl2uonnPYJk8jRnv+FUE3joZ38bqooU9ogyaCye0gAO3L3vNEUGAkgM19wRl44IobzxjS
f8Yh1G/UYk3sQ0XhpMGyq5bDzsY/DsSSeX1nap3GfRtCGqhpbpuPp3SWgwkqG1NjI4Mn9Wma2PGw
WPv3wgOALrops0Ux+BPqolduTs+wSvTpEG1ZMv2E7YHU3E4bUjfWQrHeTvkZEer3VFHNIOMs2fdh
6BfbJBAKpnak7vdhO7QDze0o5l4YewkmM0FCw1fJ0PEPk3C4OKRHXcywO5dGOZQkpsacn+8W8WaJ
QIkfqvNLUDoSgp36Li37Z0w8gQQpwYkPtj31etNbCPyK5iAMSODHY4DSSeZzJTwyzxrr8U7Vra4i
8vXE0duooFO6cKykYwZqjNf/HIBK8RIpmFZscBYpEjpTsM+SKdOPb3f37uud1VKVyeu03bcIAVBA
5jLXsFt/lR8KbloVzXQD7TUj7VzyLiCXqLD0gEAfjWOLf5CdYk7Z/EpGRjToSxsStm7Hp/u/UJFg
Q0mQzsKSBzECYm2DQJxOkWdmh0dADvWcUfaXu6f5LROaf5ChsWqphlOcEtGOn8G0mPZ78L6WSnYV
pmDkagEWRk8QgNYztxnMTnq7P86mMM48DyztPMo/kZbV4h3kanoXyEPlvKN6U+DPeGm4JklSd8gL
cUQvvsaM65F32Vf3zvG5Avg5fzLw5QeuYZjvyLec5p2FhDOsDdFvo2un16hT6w/CZCe54xJmK5oc
XyTfwmVRloLte8uxh8axOyX+KQQ7Siygrryre451DWHJX4mXdxYf1ZeAl7CAmio2SEqV+fB33QYA
psXexQDkSqcZCsnDnPtvXjazbdZcuuKvUmFZRxbMLrBTpIyKZh6EU04iN0EluvnH3RiMg0HoHpwX
gdbXoHWsupLls6ptX2Xi+ueYjV0XYsOlATY+ckzmiRrHolPn9VfKWrX0CCjrk9zaKwgyrso8bEVR
8YG6zjs2i+Xdem23H0I49qdxKPeaCYxq4C/jHs9XZsvnzogmf15ttBZbr8qmhqj9ghtqddq26TaJ
Ib0eDx0ZoCyDF+zRQp9dDUueDsayLP5WAyks3LdaEuhXTt2rgi1sMl/FyZUIpkSzDZyQlj8pczqU
hCMh8to3ras178zOVlnnFELWcm7V3mFi1v+5ok7Nkytf91JN9N4/yvkZlLDPrqDe8zoIzeaoaq2B
bw+SAuGGOWeco8ULGRo3vsvGVzVr3HRclhNCT604O0/Wcjc0Fll7zeojioUXoNlxS2JmBrJsOAJi
/WZ3befJLKYJo4VEDz6f/NJ/PY2WEeTbbwLj97ZAx+sKqEjOLuFv7DfJQ96zqOcFMBSW4Xis13Q0
VltfdDCgLgnCEoy8enunXLDwQWTGY+OOfKvXr0EIL1fJob/7s+xBXyCJy1PyqdrOios04OtnAwzt
oOgTbtvFoM3DdAJkI2iAn3Nj9uohQ0aWg5ixpXzZgijsfhhz9VJBC/34fqlzOkRVoUOPRw5K80db
pMODV5sX+QYGKAwSVNT7AarDEeMkWTkk+PnQKb6HaCAe1pqvJqxFxL/5euBy6qR7CtDDBTcAEA/B
cSKgMYnIeitQ8yI+Do8KcGMOqPzgTVhlBleJmwqMVa3lQ6CXo/hdv1lCMcNwXg8G2HTFhnKfDGIT
Ftd/W3Ip9AGotiiGYz146PXT5Kf1oo9Hes6iX+k2jI/5979ZXym5aPsqQxG0RIP38Abirm4SUZqz
XCF9ZpBBqp6F5y+fwc3fl50y0X1iMCkopXS/M7suZWyLgJUdXjdnxILADSswbZNGzcYaJHQWVdFy
7ylybkk4fLi1dJ5UAzugltchE5d2js/G9u3rQJjd7oWZ1/Xuak6RbEyCy2K0uvDWiqxJt7zRQIq7
KA3LrLozPFySrTf898XhxJ81BZAxbWx6A17IZfsYRdNoklUHaP1eemMkl/ND8GvZqrilB2NEjJtv
mIKX+QBBPy0qXLofNcHqwUGCAA2oeuBr5ZKzQ1hmTpHcZNyc9wZ9v39Bm9FACHU/EaqFtTKug/FR
x+pb2OLeKUk/2+2AHaEE/ulvQ51sCxJ/OH+bNrbIk/SyopMu/Ni1SNog3qCYo/ugB4aAQV5bwjID
ETD9kLUeVkJtZCg5BcLlvaa/BKCpl8hhwu1nnV5RH+uHLO+LwBUAoDEdftDRUXAWhTGBwrgqDaF1
n2tjZseqyEFOlYRaYbMZB6gIAnVjXsTYdVXWcJNfHTf+ML+lx+kSs0bggHCxPzqUX0OhORrQDNb/
zTOauSYkSrzeTckWyfdKvHPwyUsd2b7ETocmLA+yaFgjDnSN97S+DuEkmqaS+InaYUoiAuFuE0XG
hxoGnq2EtsE3kiqtRejjJq7V4Kea4tcCTdqXLPMBWt+q+li3Fl2gCMSnL4q3mOR2YfRGHnh7ahIa
hxqm0vlhSxn3aDJQKOQ945t4bdvox1lc59p1Yy6Qs+WJNCC8kp2BIqSkhOhQi32oTexCul8tquc4
9Rqiica4Iw89iJ8dyhGhfPSbebtL0K9M47j1CAEeIS/4EC2V/csdbfKhPq1z3aVZDiY7u9wHfaEw
a4gBoMyx2exoKHPw0Mqj+ojQLnRbOitoLOGY/YVKwcmfF9riCt+CooaRqcj1bOLSdIgW2xGTsXYs
QQPP8qataQH0b1EdV8XVD0jE3il7W7plIsH+oi9WXpldPTN+PkqDPN7B2VftL0TXBnfh3qtPAR2u
irjZV027dLehtqWRWZ/uKvn2bNxOzE432lk+bWobVOXP7aJgVjtXNZlkRwsTjw6GZz++CQokDLaS
7a6Kaln94oIFrFLBvRbzPI88uxtiHHc5seuCWiO7rNE/raboclARQx0tukaWwX2Qo6fcLCSHIF7Z
RJ/iI4s99X25fOvKi8Mc5F6MT9Euf8l91+/o9vbv3wzClcq9LSWsAC3cnNPcZVg0rqJGvX1JOSt6
y1WcZqVTwL9KBzSSy7uowU1A6172vTd9h44DA4NNsqBSpcnA2DabtsPaUQfaXn50T1ZxKkZJPv+b
vkZW3dvtGkJ2ok6h/UD9XMeir71MCF3hNMzkP/0WIxwfV/nK+QtO9prwTjREvgdunBDYbd4dvyFo
c5dbpaG5SwbjrC0XjmK59pp4XF4LI46tlwdvt3S1raRTgsYcyDPCuj5k7MeayWtmPzTfytwiCGos
G0w+TOhDCCXsyxXO+GmQDsB2SpmBrp7rUM9+Y+ng21jyB3qj+TuULAOKRT+lznC4qJZT8ueW21FQ
ofGSAZf7mhJKGvIHFl7+RjwEwT+RFSZs/nZmkyl0rB8cYqrbhXqP3H9KaqFl2pTdu9wFOK3++0Kj
ezrDiUnzGkTSKXNuSxH+T+mXxE4536iJzapD8V5C9csOUQeOaPvvlG8zBxoku4mGomMWQMHa6+2X
nLKeH2tttXvEu9aQiJquXSsgMsTijlVAsQOAh6OHubjSsFneEUTAICxawudG7iYIWdbyZA8QdTnD
mdEG0bbEux1preFZObYgWEr6ddKkr31KfODj4AnmeOON3X4w7hHgUHqDUItragpBn4hJZ5WuFcaa
xhQ7OVLldc3Ohi06Mvz91hP7csbSWA88C01WLK7Em1/Ppt8azhjHE4e1/kBD2E3Fr0deUAdlW7I7
odqab+9UQixjhETJC0kO7smIuVPbXuXMEoANt9gnpeU4rIl9/H8CBVOOwETVOrkrTvWz7t8hpSKd
+bngdwvY1nrWGLiJQulknHnnWjnsEz8XUpogxLqvYv1OPfhM1jVgHe9AdAMmENQdFu6ZenrNLNVS
F9XM7PQU4kzikcaPAu9EoyNTAJag3RqXgkHduiTW69Hb76lMl0nd257FB6YocOqkA3AdITP6KYdF
bgGcyZO659uSmI+n6zzxd+zk7tRPY4pywlzw+1RDaaW394Svthme5rKf2P2QG0YXgbTUL/3yMPLQ
aj2sS7fXpScV2KyVbmOYc5889rk///IcvFBV1XpGxI47GJdP42IRUH7VwPOr9potzQEjaAYquxdt
Gymo++r6Dvas1WsE4IPwwYWH7oJ/NIroOnYMvTmtK67zn12vetjeJgurE8t/zepKrDMTp5I5s4K1
zz9xkaonnVBFRcwb596mHO66VqpYJV8Xe/00OXmNDL/V3123057yha9UYnqjtr1EaeAbCUD+G+5x
N3Q0CjCbMCtk3P/3fXbUaeQmXvWpYKN+8WZspmQkQbPrenmAglDnsIbInDB5GJD9Atl9umBM/0Kq
OQpVUzWFaC6mpxQgbJ43r8ouVc6TDZcRrsCzxsywFfh6cwfRzFvBGKvyGkqzwWYdoUCfJF8s6yBw
bxzaAacHFHcAQGTkl+hPI+hu3R95kV/Myl4Wlissfg0vLgwGfl3HybdmMHeYDXzD57svEZICo046
Y71juyRKXM37wdlS3vXgAQ+OBAtpGp/hjXy+S/s/aaSut4zgHXldZdfbKmFB4dhC3KkEbiKGWVCO
h/eA+bhWhkYJKAG2WKy0BaIbds0HyuMGuEoUzY2f9pLFaxdqz0n3+zeQx+n7KodjHUy2hghfaUml
dPgaO2Rx9/jPOljPt1Bvt/bhUvNhHY378jI1b0R+nXhN2aJQA/ZESxZ5OLFvO9KXZj36PAGDeFAG
lXsC5cUulIMONAWmS3nzUaPjvUVGm+4yDn8HxL7+LjD0Xx0c+hkYM08H225AajFd0mVoIbta3PSD
0W7HkHvEDcT59Cmj25ohjPdQI3xGMlcW4D5fFlqlr2P5dBGWrqckSRbT/P9IaMN+e8fwmICWqD2m
FvlnSeGpM1O7Tva+lvI5Cw8J5dJ+GBbUydkDdjOrT3OdHaK+QkCnXG4C40HcQnqn/wT9ywuwlWUy
rDMIc87nyjTeoOCNKifs/G9P4Inm0dQkKCftDq3EgqVeXbtGrlWNLhCjVlcPUarKELcGZZDIt+LP
dM/1oNiXgp9LGlxEWltQFCCjFmjgBXuSifahSnFNuOu92uYar0LOcwZri4nH874r8geOp6yq50tZ
EDgf5LTxdbPhBViWs2TQtsyqBumyIvBt9lzyZabLqP449gt/K0aGzMdIRfMLrTKo8/AD0V4ontbs
sB+zK7i+xiZ+EnfHz2bfzVMMIv4EduzN6FCP4nxoHT48BkRjZqhwdObpQQ8x37q6ybHw057PpxQT
FiaElELG1S3nY7tmp/3TWJpfBxK7GPo2tw0J6hlk76L+OAI6Df0K0o7wASXV6Toz/Zqn+MyAXAZe
XmxlE19xOkuF6SsKmRQZyUMQU+nFhoV4UJU+91GJ4dMbDnKBYAQEeDKpG2fNxr4VFZXITTRZPvlG
AUqPQvZST5PLbM0rPkmI/ZhKkMFv++trmVwQ+pvy+z6BIM2A3Q3nX8hRzmj5ifz3YGTJECXVCr9U
tVqtaj/hb/eZ8uAhSI2KR1fGWLR+4OWmpqTeyWuUhCRfDVAHbZENhqAADZDLYKqODcl3/I9UpuiK
PXH5yIIJG3oFw8AeM+SaLvby38h+oxuWKS1rKXc2kxDClGVTHA9HgJE4HwapdbuvKDG0NWTAzyck
137fpq87uVyR2vHRnEjMYHVuCvlZVXOBCHrCC3je5JyweELnjoKe9hvzuJvedaIyFhJdHzudKTrH
oDqhC6/uN7Yk/O7ft9wpAfKPNBkvz02aj+LcjBgGiPokAZjMU9LnZlHcWq9KwBQ/ZzgVHBJoBJM9
RBI5itKsCnVKuWGdEJxaNRh9QM6sCOrxtjYFuuAFPRzkd0ccl18O8GlJ/Qr0ak1MFMqYNGbhl4QI
pq0nuyOh0rSKoLbB21ohtAuqrFKvoe62zAGAmY9IvIt6GXfyF1SUhPDL8Arv+R+nivYlAV9b/U9+
t/c6YfwKlMBWOhuHNLVE8VFuIDbdmt6fxhaJZLcHuFEUqooJJwXnz+EnmBTRm84oRdCEXCGa5Pik
edY1ulAKW7YO23c/PM407/xiSPTKSanRrohiP7epykX7WJd7cynbL29chIKwbXDWFw0Otv291WVA
oXVgwuqStaZacoM3N0ngXELrosc+Mtuj4hdhaeRiggBdtZzei6a/j0BHQVeNaazUSzW884x2wEjt
thU3vJaGnGgg2E8aUVIHQOnh1gySKBYHnVedoHQrz8hPeXULkKJ2KE6v8iFLtbVYchO+laChQt5z
I6l60XUTYDkWtIj7e1q/w7sSIyoU2Pjg9yMO/MdnT6ZO/iK8BRwb/iOm+rD0zlalzEpp+ftpuxmg
wjFhfyB6fuwZk1OrjubJGQ1wxRgWj4spHFmcKJR7NVybppgRfHAOlsWVLmB1HgJmy7ZKNDnrlHty
pEqplI4NA5ls/Sc16ZqLJMzxmloxwKXhBg55LErmeb2bJ41S7LVheBrYSIFNA/LhcJq2gZ/ahtXm
wk2q6nXPRqos74VP/1QwGxwUtqAfv33eKvGL4UxOw7/A/8Higo88wp0dG/v4WHx5WB3QPv1/0Lrx
XcC1aVbCKiInnL62XSJyKoVEnbHOiknsUn40d43behgMG0uRFZqdIui+4K3UWvsZQJAwFfpZLwoW
qiPp70hrCdkW6vb5L0m6/2IIMhhtBMgOQt79ReIUA+rnfDItuP39hUpB1TXbNoTFDka2mAk4a7Q9
Fwg2FsBOEIccyGynCRX534saR6NLGg07dCqB5mrZbwow2X+uS3Bm42sZdW4RzbtOpatFcNBkyajh
obrn6D3sNxr8lLRowwlxO28tRgu3okyDh8yj5417XtdlEULkMocNynyluyhqQPnMHkkOzNJX+IsT
LkCNqPWzQnA1VGygmTDvmPjBlkYMgIRGV85KiCLT4CNXhqABsup11jcy+ykZd9HMtzGBOVnlKZMJ
289voIqzaVVOCCmLkntds6PZEQTZRKMJLJEShVtC7lGsrfrtVn/C+4PsFw9x/R2DfEQ/Jlaw61w0
hSN0w++OqXz7C0jj5A7mtoGjK7f962e8HHrHU9qby2mTxLIyz5krWCc0v9c0X+AFKwhvoGuVOLbs
mnYrU1jbtuUpUEUxI/VDTvhkfYYQDKIokqQ1t6d/LoaJRMOJapTQ/epVCPLuPdeWwMVw7j60mbDv
n8SIsRbVafVABgLSr7oD5a9OwzlbV0DK87eXh993ahKnEMNwmcYrHeOB9vXpNnJs578YWas5fw5p
6ik8EO5FIeWbPLGo+fnFzUvrQAGVjpyQf5iogOr5pD0aBunMSyS6/NWajCCu37UKeEbGFFOiqRu5
tZ4l1qnQPTXZMzq/mviIbtJogTdHmrl1vjduj7OoXlt7P+3BDDvyrONQ03z12YBGol7gMnNpNqeb
5BRc1s97GKyNVHtAiebsFyWuXP+lTvoXvPeGYPjWhLExEO4YyOxdJRmONsA/j1SPFw8RxOqiCaIh
5t7VN+iiZePuVmrbh5AzUWl/zuaXlLz2jJ1gDjp9f95Z7DaumGik3eIDGCMJKqLef9eYjoa+ZbL8
6sNZhxJoqz0jq4ztXfoJSQoT7iBEGJYvWC3PUNl5msjlIfaOCw+IvSAwjDX44AI3PxpPGiZBKZpp
E0RMEJRg6QI5Sy2ZPprqAVm8pG90P/GP8nfC/varGiAQm0WK6+wVZvZ1nrayLZi7NXQchlDt+UuO
dDn4rhQX2CgcFfgN2d+WNmYfHVZ5OpsKK2gQ2fUndaK6XXJtTGdhPtyx9Xbw5MpVrRnZtawHI5nt
DZ7uXArK3cGap59M1r4wNosBrF4i7n/tz5aKnjHTgOfTEnsDqD+xGNaOCLhCgMFW/zykn1tSMUyg
v8WSLQK3zajmRNBgNCZNXlip+9qy/zErILRTPNKKL/hcFZ/37rHTXfud3taK5rybBOj6EKGHeAVp
3bMWKxAx0hhLhHQgETdOhtWRkfIQDPhniMs2wqXuKkrcyOU0nQ+hDVpCezzXYeLoT1gjFu41Xz1L
WH+4PLqwlvU00Zghzo3OoGl9sd1urwQ00ZLBgmOYuVvbrYVsiI4nwna9Pbzh5sE2p3q3DGfpFwmn
rSYXR5O89XKZ8BS/Bmv8VQnx6cFWNz6e1ZpwxR/VWmv6RWVKKMTQ7MiN/EgJdLi2aCZAsqvoGWUi
ZP/WLIe5PczQWEkIxaU/aeAIRIXP3rEq3SeJVUphpYsA+8Pjz/mgxTaPcBRrBDOehjwWtqpDlJgN
FoQ1M4ocr5hvGPuw4wRw9lh1SGRMjf4snCd6S7uIHfGfh81ClV9hJMVgkNMd2hJXfqUVmCaYnPC9
vqhuUBQrv7/OCIXbw1sH6kpV7VM1K4FO6z41cBeuPCKY2/Sh5BSnh81Masj7/xbC34F9iSBg3WC/
jgFO5Vatcktnu+AMi7rC6wPUaeE38PRxJbzoYGPXG9adX09FnkIU81e8y23p7H86HaT1l4u0evGF
A8PsFeRa9EgYAX1h8t+jnDAqrmU88x6oZDvi7GS7F6OloyWo6ZiCYXt6raiNoqm+8SnyB4zXjUs2
1mWyjf11cuq+7BeYRjjuIHN7zyXOwqEKWLNCzlfotWfeL7c4E3g+CxdL7GAH93IRdagfYqIT0UTZ
YKPyV44cBXS2+U4m6kA5+r2OFdBvB3h6mdCMXgcmP+abXqYFt+SQCyCUoBv6rqfRkODr1/tzX+HQ
t9ChhHB9WT4k0p2/xxA32LQmlDSCJUPTjJxo5X152MxAN/wtcoolypfH7yi+yn5hsexUmDy7e4ns
Dr9cwujhcOtNZlTRQQHYwGb5evU1r7Hhag1cldmtHHTsp3QbtXa9Hedx4XY36n6nS0cyWCOyslSP
reZ/kP8yZr+VQ+XHp7lcCSBz3sR2nsTQr6qMoQ1JBnGSP40Ed+/Nncx0d7/B36Vp/vyzPlkemAxY
CbM4apVQhC3fCpC3g1oPPewFydwAu3SXDJp/GXm7L5XFv3kRzxSfXlvaATktH9VPtq9hUKcI9mgc
uCBPGFqUZO96ppdxRv78ndDvSzqbbrtwWNfoLt6swhVT6TC5Vqrn3LNbHmbAVo+9q2HDEYWuvj4x
sdi1je8bB6H9EOubsbm8+LMswU9FVZQ4l5f4CDPQbBZNUohiCu2LIdZ9VZ+6ZkuZGWmEGzW9wwNQ
tH68xGLhzFaLQOYIZhEdlhe0n25O3HJTqWYoj3ywdozdX952VVvJP2gmeD0TI6qwQdADdDNx0WuR
2f7UGAWwRPjv6vK3demuqs2flSg8VC14a608EAk7x7w6su84QT0OCLnxu8kZbMJvHNK6jiHsz6fJ
p/CpnbfJBXSQGaWxEyfatS4xZb95yjcrgdvuXjpb0v4OJ2O+tvNzFVWkGFLgzLIOOXm5O5mmgBAn
UYKyi0JPTUUVdO/g6SMxe+tc3BbaPw1x1Wrz9X8rhKLi2kefzdBfo/ki+f4hPMYMamG9Zat2tZna
0gLdJ5CGCxTaPTBw8ecy/cNNXU/WHhyjYIqYA177EIVCAjHAhchJ8DpKjLFj3EzI2jj7YC+qpgi9
e8ogtKgn3dhv0tkEar5jfG1us3Am8b7+NMHXurW60WPNvG6/+m2hQfU+1pRnZhEQWg4F8DTlsJ9z
+SklQ0C8eF7/XvwThMd2ec09GdrLSRO3vyH/KfkNy+oerAzeDz+VeX1zbOlByAntefXdCpCfNYnt
c63SekVC/b8+JBCe/35klBbnx7TziU5Fpf053Yl2tnlBAr8UwmrWuEw48otS+yuZyvNsgulXnOGz
2aaWwlzYLJR2GvuIFzAViXINYVnugdH6d0z6UBOIPUJqaXvHP+seiMw270aqEcjqENdzk4sIe6TR
Mu2RC3Z4GpeimnCGeTQMADBnoOw3QEBiXQAEQbVvwivRNGRUOS/0h984FEY3vcYpHj0dr6aZp/Rc
M0qkHxlpz/jelDEYIzgcG/T1Zayyotwf4GgKwlYgpdP5M7EvL49RLYiEuF/jHh6XSpcoNZI5iaPk
8Z4VTxA4toMahPKz3HvFeHkLsUDQfoNP4GhiPSZB4u0xdqD3PT0n2tsolACV3w3dW4EJncYkDAFn
rP8tT5rfEKxBlEogZUEX4p6UXquYP5FBBwWFwFRRIiSovbEOUkW2o5tb1ltqNcO/vJvbsMbRUBFQ
UTsxaZmEtwRqN2BRrzFA8UbWWguU4R7z9cXncks1a/PmwkLfiED1FAI/e+FQFrVk/iHlZFmX6H68
EzvW2j5yZ4Gmr0ufHqFTPnDjENF3bgLSzMk9bL9NSwnBDnvG6oz5VE5pTUYpa7RUHKdwUNKxDARG
v8+GIqJQQwyoogNEcUEX7wTWpNpkuEDRIx7ftWOk7YdYCc9WnIg6uwdvPR7TXU55vyf10NpWvoeg
b6voTaaGYnlm7yYeaKh35vbiCSR4XNIMONgUyVwEeOegn2eXVSWpVM6lRAPdjnpxr5I4Gi8WscYn
EoC+K2JaZbz8vp1N1G1VpjScpPptgI4SAbVgyOq5jehiTyyTDBwhX9iettreF/S5sgVa0dbQsn6i
b1d2aYyWwFKwmGHYofrFCwteOy5EiyFN/ldyk/8bE5nNK9m/KS1Cc3up18ICPlIfjiWivi7wDS/9
+KUi7J/IHQAdtPO/lFrXfegh6XuT1zNy+k7JTWkzYlvsQrNlp+FMmd/eu8Y1i1qPrC5V/b/Ooveb
uNN3csrn0XotZFZ3kPjzKqVfIvTWWHvRH5Ug0l3oniwjjinaRQ//agY2uB+tx4ln13rD01TeXE+d
JYswo56TCDKM5GKJbl0WNulNESQolhrsizj2GT/kuIzZyXIYbKNY8R7iFkJcog7LjJZBr6V/u9FU
sASyME9HVaYsGV3dBzuM/pIQx31r3g0w21sKmivLXZ6V7BWc2xBm4M4U/q9lwdi9CYB5QgfHujvr
Px935XJvupKzFKlTfZDPlxuFVxqA0lrvlcFRbd7IBbDi7a0Ozb4VCrN4YW5M4nV/Rx8/ST7wCvjL
LYWdEu5IIBnAlv/C5VEPNVmDMXQbvaFWnD0S+ZjWTym2KhadGGOw8sb7cxCVp0OjXMYQSzNW7Y+d
OIkemxhAO6t6geHC8acdmg7Y5y62JOviOhfgovKGMs3VDjQ3f6byUIi0q647NOHtCAv70raLvYHr
JGB73OqFMqAMtIvYV+6x97eOqHEwxiVZFH7YtcsbfMWGBXoPZ9wPRUXqwGcPa6RHhqzO/ld4qgLd
JhS/LEVUbGqymVcJ5lpaBrkag4EcWCRpcB4z6UrhGC+wT7dkwjVr9K6NEmlHzcmZ84b7z1is18mO
WijdprHI+fjKzWB/dxpscSuqq0s52oaBHQhpx+KxhvQxlvG1PzD9WoNHh8TTMMzoqwES0B2FFxSV
daa4qBfeghBKMOMfZL+8wekW5vGTaS2bY5irJqMRk6ymwfVl27715sl3S29+zAume86tUKcDZ9Sf
EimHsb3+V1Z+J1ThTbg9Xblhmzqcukar6HYKGTYk+oDOMf6+hVUW8jaJTTuEa0uYIjL6nUOsFL/2
5nwBXWV0NXSx/HjGhYJNJcW0eho7dYEmuJ+O55EFVYA+kaU8bKxj4Pfm4XxfyB9zS8M1R2daTIE4
xPZe8EmW6m0cdtaGDd9DAg7lvApWh4VWYTG/pvYnZjsB67Eh8LORwKRgFzu3bOQ0Qu/goyEWmp7C
6McdGULD3v1YOJyOHbsKHC8gtau5LE808qpAbk+nAMCVU7ttwRiiQMOrVUlhZi4YvmPGCsiqGcPS
uAiGvyLKsRFeopjv7dVn4xw+VKNZBNLO8j/TVPR/NuKNBD5U62LY6JNtO9VcW533b5eMubOm7MNV
cIIVKyTb0TZBnwiTCeIStrSSbAcfzjjbIbmaWS9Kzy6bvCq9BZHS4San8V0Ex7mIdehGrp+vueLk
l66w3ShMddWuPVCyPVy2fvnOq/8jfh6G15Lyls+5DiDTT16U1urAuqGsoCLF0NnxiF+IFxLcLCUi
G36t5jVaykhXohgw/AJ6nlQxsijRzMVYZYi3tuHwTmu69HYBPjRMouBaExe1m1iI9CStmgke9S5d
jyodTvcKooBjm9UogkWABc74nU85RKURy4bLWS9Yhqbqd/5KqmvxMjb9N2p6lu31K26dXucLf/yI
GNonlsAJvpvtlQBOeTWSbsbt5/YYrs5Qtd9Kqg22UGkgoYIiuqr3GXRZDRGr5llFXJAnVagZ/11b
85YJZ/RhDAmmRlYLtXWDj+tLxS25NwXOTOGBvulVnUX1dkbtR4o3mwVn/suOzaPq/c55wJqv+jAQ
Uy4g4LvFVv/qpA909Qjz0Ym7qsUJT4rLoq4epvgRrcfeYxhZeaYse1/FQJGihePu5uvwHehHRidI
KFybEqN/tJktTVkHlcz3cyxe+TS/vE0ayl8FfHJD9rC+5LDvOSt0tQo1q9u74cfB1vzESCMG5CNV
IsddQYOjwST4MttaFkxUVL1wkGMdXHvUeDvxpBcnF1OWft5/pY83JMDAM8iXcxY7/YR73c/V6mnK
hQK6cIBWebGLn5PwYmlVee4vzW3Ie5srnKSHOdjZALXPGMuCkJvrT28iG/XMNglqmvtzWgKujOmQ
cTOqTAtEal+eI3wYZ1/1XYVrwb7A2FyCZhsfliRrEZO5jhZd3db+2MWLkxcVwEyoS+RCrbOxXhWg
ZCf+GWp/zlV1Pb0asHuIKkSEm6a4G15WaYjfTKC4H/NkoCFVjQ+3AnYWughyf6KFBaA7eni79jn6
bmoaaLp8gDSevi2oONkMoN1QRtj55eapsfhV7Mgn0yjU4ZA1bYnEd9hBmXtOLpY8URPgteL5xLdp
B/asfTBkzih9XW5Wo0zHrTlWvZNizGpuz5ouqxDdmiL/sQegK+zcInWCxTqT95wYkAE6xoNlMi0S
EV97U56H7ndnQDzrLXTfH5JMlJMD3ee2Pa+DzUoLYGYlMsWp/5bR7YJMmzV5QvGgNXsezMKLH4e+
scrcadeCtFFKZ0UNFpwiiUkqyI7JgdRbOgLTAPLcFvavz9AU2EsnYa7rYa8gVftSQhXFbonmabuV
Yry/BfHue65irTd9SqTIG0WFqh13OasXrBQm833S+Kx8V5a6q/y7IE28TRJhRGcicmIKmA4g52+b
fNGEWOk5urY1yX0F+NkHZxYFg2e1eZctuqpQE9GDJK2+wyiKiGu//RspejsS8mlmhPew2m9osfM6
9zrkMgg3X3nCoxcpqNJ0qlR5RVMnF9NUp5GU+90JgcjtxagyIBu8A0Wxf8P4L9r8rhCVUjl6ezuh
qu3R4/wUPC6lsvWEn4IKI1xRzUXQVuSPlT2TGhkyVaTmailKB2PcrFsnEOv79bnvzp1NjzajuNic
JBcSey2ubZut9gDW1HQQayJia4eCx9Aq8xU2pYCgPaN5wnDH7H2Tl/CdILu3RH7ul84jeXIkiqt2
oCO7px3ioN87AIM3+1N7Cj01UhPXu3PocF0DbhKOabcJn2bvnvk1ZeIRpp7gWArjOo3G6SK8DieV
/3LvsYRPF7wS2g/24guuN+8O//QDvSrrpuPgPy0XBYc5p+b5v6KSgg7A1L9KZwRpyFZ+stPc3tEe
Pmgn3nBNFiKs7NhhdQvCaol6KbtD/5+lUuLesTmwt8Z2SnDLazmQDwLiQltaNp/whCIEWZFL7zkv
51BK4y35Y8XVVkBm7OAPAlD1+BLqlJ604CynYjaFRoxs7XDiXQNDqCGifjLALc9p9mJU0IAeahz0
xK+zf6+yGkNyyXGM+k+xbbFd5tS8twjdgbUIQUoywOQ3rYs5hhnUA8JW4RZGH/WyPUzQFKpD801X
xwHg898JdUBzJDxB7dLfg6fwljp1mftlRvkWUfkujM6qLK33CJwPyT1jSfey3gsMPHqCyiLwk8ZW
UArfSNoyQ9v52PkVy999GLYB9siuiMpnQaoiUDNKX2rgz/OLMTi9y/M4Lbgw/Ig/mUtm6q+bh3tT
yIXXxuBwiaLvg9MsCbkQU2Ss76/0wXccPzmfkR22Ago7kz9pg4Kc7WtF6ja+Zq/JAYQA9WfSLUSd
s6+NHkvOLKLPIpKRvLztjVdAB8Qfs+JS+XV1pXyqMvwdRv0SGbWh+dE5QFRhBmDKEItq+69uWVSQ
JWgawtxZEA4EsEZU5x/315pmtUymR5X9GkS1CM2IAeSqwSEA8dO7iKxeL3z0Ly/h1flJkL92jUA6
GlYJ/hEIRzy5GwWkoY/3Wxr5swIv2QVdh8Q+wuw5Z4WABDV5IXDERt71HGkGKdNQXsbzN3Vdj/oX
ETBP6NMJ472trrzEUDJCYQAfimxRuyS1l6g9exBKzBgZCBNYgdnaK5NXA55xmRRZRr5pKENQ9HUc
U8I0ephRQnvL2W4aDaAcPBaxovc0AL/6Rcv2UenfBfhDOhaM52FFFctCgkad0B9urxNGFZ4o4khN
3kuM+sxzPgCPKt4l5olUg7QM1LTQBuO4eVPLXF/MG2yF5N8IZiigc6O/Bs3aWZun1RUaz/xAZfmR
rUcWu5s/w5i+4cdPKeqc2v7BXQF4SPBUMIQ4+FXpAvpn06aTa4zGUs6ooe4H9VGEzI+C/m9cQMNz
UEwjpp/iyzVs8CTtWNuCXInulebZs1u08rJbFv+zwpNFeDn15JZggntKoWzJ0jyWWbset4hz4Pm0
1KK1faqWOECm5PraCn3LV9wTxWXqMvYmmtwnfgisPcNHzsyfIrbEcImN7WpEXIBnkel8faFlWfU8
zj6QsTOBZf/XXAWOVSzdOV+bCP+DAegKX0dyH+vwjVze1NpnHatYzZy1PH0QA2UsOMCbk1EQUbpk
DvUV2aG9xCdg+WKQ8BvVhKEqsldJYFphzm34tJbuo/v64IvyapbCF7up5QrSJpwEiy/0YxItmy9I
LW/IW7ht+xHTnbPys2jKskToOYl7P0hxfI6c99Vr/OR9S1EKs0wM94dv77dhQNfzA0tG5PMuA8Fr
0Lk2hxTINMoH0Iw/phS5KNcBjHsPosIXNxcU1cW5GG9QoOqYdPnXZWxT4pzOSaV9BERfSjdxywF2
yB5pYHr3xloZjd1JULRwvvgsO9tyPBo8gUAcxVU7y0G9/N2weNhezK6coi3hXlxLfAPT/ON1YoBp
XYMAGcquvGPXr5I49l1M4aWpCkKAQElh+4DgEpsV52PrZz3PLNs/ySMS1BPc2YYmKiQ/WoH2jr0F
6srUoCGH78puuSLw2q9PZmhwEFCgPlJvMT8N5Oog7Q17qY8HXSsL4DlxYxKV/FM7d3IvzDEzI5Up
LWimJk7pbo64DNoFgOpCNrdnfsLYYdgPytjiq8SoRZcosN6Tx3QI/oRGELFHfr2Q7i/2kSjw7K+p
4nydfQ42aSbDBBS0aaxXUaySkrK/kTaTbnWgr6fGxc1muTHxLzJbJaUgftMCiftyajTgerKOjbek
akhr0eumzVikHYxgdxekjYQ/R1exwHf1/vu4w4BVB3pWih46mCyS+S4Po4eqU2tXWAIirir9DOYI
idXA6THKUR49Nm4G7PwG1Bq98+1MWxBT1lO52xDLwxCrqTeuX/AZdLSB7vNk9blAMaaGdgwiaCrY
yMDxegJpc/6C0aaZfLj7ZCX6GB6eRjPWIQMCF8dciWL1nJVz3yvW68rw75RaFXPe9Z9jNSnpBYQt
7+bSwWTZldNpZmziqCWaTvhPbgWh1YM0W1lv8qlJrkehCF45Zze6UB7ulW20Vdrhz89G0Ok5tHSF
HWBZKjxMZt/RvjZFbjKtMdnhic/9N7Yh6KapVxqGyWJrNRXh8hLbs6NsA3X/W6jPdqNbYHBh/sIG
wlb1yS4V19IoXfaZlCnlmbWE6rNipj90FakJkdumpqpaaTvgSluMGhm4mtD5wh0g5cR7Bf1QwLGo
yltbVkkgFvp/x92IeW9WBnd2SS15vlSSFEdb/eHbYoO9JlGR0gWBNJUE8rFe3ebmbpuP3buosMFO
DcwEPARJ2UjzEcW9SmgBGC50s9142duvk7rtBfkmJZKDsC92m/X5xULJDnFyC7rDQ2o+04lZAnF3
7F87+i2cgnT8Gj6vL1m2b/sz+cTl0WxZGQjA9wR2b7W0tTujPaatmGBWllDp7LSHEHuB8cYbOYS2
bA6+GswfMl47qWHaD4d/roTYr51ipZBq0llWmmw2uVOiP8dp26LKCXVtGDBezTWLoYd3uS2rVkwp
AcK7JgY1WhIszqGt4IxuIFH56G0dY7jiTPaOqGiDaOb4k3cRGdoFUVkD5q0FsX3EAroDmt1Ln8bX
2zQd6i7pQMvMJGqPhcH91BMU+motDTx7tMlVrauKK8pNpAr0Oh4Y0uCM5lu7exWy+Lp36YpHKivR
LJRaahbH4vfzbe9hfjWPMsP11xfxJGN/x35L3tJLvKJmcGQRvtKoZtExc7Tbc7lbsooP0HO54AAA
1WCe1KgFj3KymQOFVzs0V3upV5rnVb7enSy6OPRHHoYIkLiCkGneIlyaWwht9h99J2kfcX36uTPZ
euwk+HmBK9usEaaWRW0PbxKAYko3dAScxufExH4cY+gEpJu0HlNnjGakIdvivguWmz28//Evb7YC
RpggpajYx13wdDpqWmwo8EQZQ2rjBPIUrxfVe/pT+Cleai0PiIVoBSiVQt1t1mvcU1M8V6o51plr
TRDilERyIFbWo8iMt4z83jAoJJaX/jkemAYmNV+ABTvwhLr7r1JOhdCEaVfMYSJm+7w0V27ZsHaW
CD4tpZd2BuC6SbBOfPk0TEyT85yevvEpW3D/I19PzNdt9+dLr+h5koIwy6x7g+uL/jOZM8ylCBR0
OmOCuOrypvGZxkhRyL46WUPTbM4GZXJzhmHoLTAx6rEYJZLe+zwzSWpMNVQdh5ii4PbaSwG3JUkw
a7fBnWuDZntFzRHZKfWhj+MP89vb9Ed69UR2lgh+oMETojqnq83P1ZnXt8pQv0eC1nGgFVTj0cO2
Iaz5qQvWNzJRUHaHJRGPeH/LcSF0yEkm7UK72fGVwU9ul1eu7cFz5QBIBR1MCVSYmRpcZgcMC7mA
dJ8qysqYD3RRy2tFH0UYc8wBnOc/Oa00a4V90h7L5KRIjbQezLvlORsw/nkDcDUrY6W8fOzSNibW
xXvhtFjqOxJztH0hrlIaDumEIPsfmK6tvs2jogyx/I3J9WOSXU8ShemAdHCcchRNY2n+UqnMfV2i
jhRKznvScDSPtmPUpuZaJ/Ru9T9qJ+hyv7S0ruu3w0EnFClZSjjt7MZH1Z1ge0CY9dZ77pOYFA0k
W3O4MkIA1DhO3i+GrnIpYWL1/f8uLJUDPhOBiCjqyx6F+qwlBssFFVIXpqeXm+N4v5wQ9hJ/Rq0v
cTz0zicWQHjDHGlHoDyP9gGRZjUf5PDl0Ij/1crogjrsxeehT4OmX7cddKNJs9dFEEW3Q7OOrKw4
XFR7MP7IL/Xm65GXfA7wwhGpYNCsHB8Y2yw9Q0HfvFllVpxX7uRCRDZ6JCWq2pCDA/gsAyZF7p+D
jG4MYMGbhZqcfPE6h7b55KuD02bD51PUBut5vCxvmHsmLD+5GM+HB0WKA1XNozDbmyhbKunBcx6j
Id1QV2e14ZA8aCRuEZOeBrQ8sJUhXB6+0/1h1BIUULc3Jfu0YhkupJIu39KrlizUP98iK0np6cKM
YPjVBISSrSCjJMGN67irPDk07yWhvlnPpkQW40lyFt5lOGSmne3QoXYeF2/t6Tg+OG+8TwruQVch
d92U6KGy/RvaNEZfbtVCuNwL2WMhFUMYvC0e/kw/d0YMdEVDm7eNP0edWWwRCKzSUzird6X7D+Ab
ZWQZqtL0AAYR+TpbYZ4uo1JLb0/JlCDFBLmKzcvfr5ajZM1pKidTGd7zzkQIXJTiy1zL51Fa/tpZ
+MfIHQzxQovHPY+2g7iwGYK+hSyNBa5CJ8SyDWjSrhZAwiUwGA7SGnHKv7Hxr8IW0oxuAbKYv599
/BBY4IRUhKSbq3k+14ysEYXWTlE4ngCaY1bceLcm4VjyiP5Cy6NfCwMKGzzeLwKIqgZOrrHgpQY2
yCYXyhqXRWJr0u2xM7TfKmbclYSXsF6oyUbD/ue2q5O+EuWAekYEcnX6321bQfGl/gFEreBKN1Ap
VOGSA3J0JwECs19/WYpbdIepQ7gbpZhJA29IlwtPsX33a/5rURqUT2yLZOzN19F13qebCO8XJ1Ts
dsGm41LdyUFlzG6nshkOldahNoka0L8mr5U2yeYUZOmcso6b1+d+4GysfPVciVxU4DQ80TwEWMOJ
CH6SQmkbK9iMbCzVVo3XuiYPsRiYnzTCHfBjZwCaOBo+a94u9h1eHzskZBFjM2wHB3GhwHaIblvh
uztLoT/OFtZZo3Erho2NQ73WealwueVDSYpN+BkoR1En8bcOxy7VrBfN8cKJvwHQh1JBdRzoW+UX
pSXPsPutac8XuXCEIXmmDhOYiLH/9VdZ1ymwIk5uh54E4bTM2GWNypik7e21tlbVehYtTMInfybI
e8mmAO6SMpspj9nkOgIhzH0sLJoa2UI1kZwyVKMSG9gccDmCzAMe/SYd0JXLBVMZ3Op4isFpy1GS
MD9xQOr8TzpYyKU/5BbcEA2X2HhQewjzgj1FBbAx6Moj4V5jamrjZ3lwwA/6c8Yn6RMHuk8szqfP
iWe8ZW2UzdFJBt9P4obMuizcWI4msvhuyd6Jv03LtzXSF4HLWWGgdZJqWUzyZh+nz2q3Yz4MlpgU
khUUECdveQF/MxohwyKmyx+UJPzoaTOb52OMe6tcvcd2DkJB+NHvPCvwaCTnGNCU9AiGJH27ushX
dk2/LPDjU3CCF8mQwvfILOPl11cf7nZ7imsygPnrAnKCRlhQmzJFz96A5aU8uUkTYCkleok1uweQ
T5ZAAefMBTUQaDaAo14kRyy7tgWOa9a3qA4Xc/JPEQyftYd8CdKN6gZgxsNBshMsqIl6yxyc3JAX
eAlGfezI52aqnM2NerJrKDk5yz7vo53UqUFORhwECEpfKlOJ82N0a2TbzYsnVpSASC46TAFfDRQ+
iWEr0W5huZYibwYAJfITQ++xCmaVMzZ7zqioWo1v51UMOQ3nscc6J/N5HC4Jawvdu7FuU2CTQ+9a
lWvstazQUZBSoXOUH2npH4x9uGUVV/ycjUSt+61XgGwmXp3pNLvb66+y8iguMbI309S898FNoPSg
r05or/ig3cyHHYRimkO5ScNc1egLkVqz6t1wBHKVb8Filp+lLEZ1Whw0IEiKZ7mhXxssEBv8IUW3
ulI+rlPysQrDxZ2vwLUQUhdyvpZfijaqU/zqJOVyAydCoj2uojXMBRrxp4yC3dw0QFSJLL6f2lze
si/thlMidyO9Yb3kJcgGcqGUoQ+271rHUhDpRknbqNZGpctjSMFl1iFumLa0kACHFY29klUMwqE6
RcDEd2gIMw4yMaZ9117Qhj396gEOwZktOcIU25QTBZtKTynXUbvhw3fAXiT6MGmKZVuaWgL18Gz3
6NtpcebvT5/8CE9Dm0IJHaKLbvdn6+67aoPKf9AEOgV0QFOohiwcYb66VllnDUHXF2rPWqk5wbRD
KRftdsOOfVFGgui54xrMErGZApGBJvnRlsYh+F1G/EH2DGl4hAed4BG2dzxW6FtAUBDWOX809ZX2
aJ/KOtMFvGTGzJEMelmuUxw57OHy6rrJWHL1bEpvYeA724yPYVzTIPoSsTdA+6/xTCqON5GP3GT8
YLwnQwu/6le/XLevXzG/Hqis4SZtBLzCeDmhIKtUemjPq6F+0CadGaDrDd/uAt8XNLqoINJ9bZ81
0iN8sHkHe7CDIMA1EeS+XXRK3wBZ409UMsjQIEmuhjGlZJniMHVmb4glSlsMmmY6TTSlwT148Y8m
hblF/XtU4UHmxiki12qT/xdCktj2qCbIOyoHc1Qa6zY66hVLb8q8PakbNpcgwgrji6eEcwl5t5el
qXM5Z8GAXb9vTf7h8/7zqB+RVhPurAVZnokxOXIl7Hg2ONp366SRH4Y2PZ3j2v5R3OcuVfJRfK49
4XdASPIsKVP9YBr+aXNtd1LYTQIIscnofUDPPtZ1PdQgRkvuoTUx22PWdOo+xQdMoIPIkDoMTzsM
jEfOTO+0mk8F6jufHMpLq5SsVD4+XY7sng1Eop8pVMbIV1PFOyMTMgv60RgPwtPlWeJpiV/cudHC
eeIJ6CGJYUA2LXsyE0KO6FnfxlZiK+sLwYAgVsY9ZdreeGW98uQFXt1ZLhyzQIWHm4LebsLN+13z
zF0lCPA1mjh8vWJQNJmkHt6ymf6HRpLhoZCV32WeObKqiIw5HB6b/3WHt0+r61Yb+8icNNisbVTZ
XQhAhAog5l9dZDyFhmrOOu/wVyXfxKGF9DSPH+YoKcCHvy58a0riDQ87aPu4Mmyz9fk6UKRbIRX2
EbgTOqljP5BA+/TwgLzMfJEyhxNVMvov1XK+SZunYz6Wl2TBBf+//bulXDniNuqih9OsJ+CkPmvD
z/UedY4qU4AP6PUV5mgKMpO22mFl0hfHeziInVVAxIb3IRslRFRUwhf30phsprvGa0RMiE/Mjp/U
yLo2lDVut4+bNzpb2A0ObPCfUzUSF74sHsN7mumb96O6jRLHT/21T7xMQYpcisgcGTg038Nb87Lj
LMA6BqYANX2RnAm4N4Q2gHEf/4wNgT+gkX0e61/JeRmBtT/Foh5yUYP1GJreNgEoSmw0coVXWL3D
VhLuSy9Q+qcdCacO+qhx5NotGjT8qrgtXnA7sDJGWVT47sbGpD9hrNVfpyX87sZeQiptywej3ez+
rlXCbflhXxq8tSXOErXNwKi5Sik1UAy5QQusNfblFH6HkEdqqh9o3whtb0VCeCB5K4u9TEo5kVhF
SCTfNSH2m4BGYNRgeNgr9Hy2wfoBnD9w7HyKCF3kVuHQARyOAKYGdPv6EhHlUdfxebw2x/AKz42u
F+5zkc2t2y3L46HPTwPu4+tvGk8u1ff17cR1v55R8+SsVjs0Lq7rR94oeH1NQVJVY5JiC16OaC+r
P5GANFo9et44VPD8zHsqH0IzjtVOvnit0IHNHms0v2avXI1HNiJxd5Vca5fIkzzhyOD/kPdhOi/6
hfbroc7JOEKkq5kN1StkWaacVArUi3AQvWTvcTlpjBDAHigzJ7K/GuqpkszoCHav6jMxzx/Ti4zU
GNlkeag+cDO8w4g7uCQ0ZgMXSAsV4FWHDTHM2Sy5nSQftPP9E6bITD62yvjSJeAIV9vBDDNc9cDz
OfnaScgVjcLjDngXwi4am5U2EYfy4/MQnLm7R1GTTtHiSnJdUeaA0lHVpg0iAzILllQlNzPn5b1x
0GBj1FrN+UHp3ulo0kGDZNv6C7Fvu7eYQSR5V0HmHHRCvRFBqtVxlBtWslv5DnElCFuCR6xe0fiG
J+M3oqi38VQxXY9jrIxt7EBf8fZODUM2Xs/3kfMSo76PDNbnqGik9qoo+Q1Fevo0ivSv7XNiq5nK
YvdTr5StP2BHVjYTfCvuSS4dMRFeZHjE9gTTk2kRqw5Px/4B3AMoMCGVmyhjGmswEZ9mrHGxIMb4
WrhOSpfB2Gvqg8hxfFLW9wDTklNTMrIbgkZfM0H42gETHFwJnPhOaY7/EB2iN85R2vMG6TzXXEZl
JQ71fAPTzgMKV2ayKvKpoYTWlZLjl/eCGI+fzzelPglRqHAavbM6hNPv7myqjZOapeFgyRYNjz+I
M4m1AfXdkm6o9ayx/vFAcx84ax6a/NI3saBQ0OHBi7jwRh11m6cOD2QJxSbvjyycgQZnQJD3/0pf
IL/KIqXir0GxLktALGwh6rrdcKt23v7ng8ZoazFoty0bWKnQW7hDUWoOHyluCZqpZLQo/qwezUeW
EszDGLrOTRdxvUfvYlHQr2fvfVbB4+HyX8xOM95MyUi+PZEDDAUsjF1ZPYcYzjXT53XPo+BFW6Ls
cgB/0KOlXaDisbpsvk4uUbmquPIfMfPmwa6KBo/poMZhC2la/JdZe9I0GV9CiU/kHkGpinetCY01
1Y8jzVRnj7BURj3QQk3Bp/D10EV9J8hWwu5CQy/y+TymY5NJeCN4/2FlQ3JL2vsLR1cd3fbt5amv
gS4wk0ZtUhP6ZwK3Whh9iLKWvvqDW00Sr9MljtV56AOulkOSbxrEWF8mPjjTYS6rvMRaFwmcvdLp
yOgyyNlz2FPXrpcrPEW+41MULOwCXN02qM6ZVTv2V7e6zRZnIKbg3Po777iEQJpGMYDLtEtLT7RJ
5IqIpxf1irhkiwflajfCH5HYOJKOQwP+iF1/HQAVAGSCNvcsUTZjNC9fgRe+Ziwb3aqwSHauyRAD
99WfKaPbeip3qJ45te1zZV8BPlC5xQpF2fM8KD6iyqUTIya9NKomN+Ub2EL6D1AgGFV8XJiBO4gp
iEBqBaDPiFtBPQ2HARKSTaicfaRC/87tw1wGv9/XaPPW5vWSUnYeBanxjHFuACpfKRmasaZEB/dm
T2nUb4Q5+WOp8MyMG8b5pKlfFxG/mJm+8O4SzEk/rOIb8RK1KWL9CUKPw3LCAcML9AfTTGzbRHhj
CiMh6ipd+B0PGiBP5DksQPCQ9dgSCjKUy9yr+Yeen9jeHJssFln22LFVCfmfKJZAy/DqnI7GaCwG
pqk1auS4I2ipmbKPojfg10E1AvDF5vggpnxyRyQxe5OIXp/67IO5a0r+Iz/zfEj5ub7oHNzAXQJt
bUntBJvFtHY3wZKGkbiYdisZIP4sPUyPACm/xn7hcBJB2V1XNiw9yXp69Aotbm4VwJDDk19SIS/J
Nb6k/HITLOVvrwLZRjFjMV8ODgd/HUhPEA4e2RgPVH3CLz8rQ3LUwQ4DWIIDjbc9Fc9HTM4FPzTn
MYvdAWCSgkd2o0c0Z8r6e8+toetScbuR65P6joVhKS3AYpFKNiOusZgekkrbS89M4yaIovr6+zh8
BTdvlWHyjOtcMFhdEdQghVsACWtShlbgxeXjej4aRVAuohLobA0i0TGWhwPNWfmbvlomt0Oo1VM+
OVAYhgWTR0XLuYyGgQdagHmV172ELaocN7Bnoq2DO4uy+m3cfiQ5BGik+rw6m+crsDBlr3Sq+AFS
KArnM1n6vlped8rLsQldSym4DKul8VWozjmVjJw2I+BsXd+FX0O6Ibu+bEtHG96k32wC/z6BKOrf
oALOHA3uOAixZyDAcjrFb8lEfVX/ajnigrhV+/J8po5zubzE1LphXZISKI6G3VfMJvrVL/DYITCz
AJV8JjdD6k7rYsHhAb5K5dDvLkXxlRLN7taCMv+yV0m9VXDCjfdmTyv45HlixkU/0bsjdaldVdQ9
5Do+VwcWQTNToByZye82BhgYSDTfQQNgHBq61H8PGJgFKIYE0JmSdV00T+/3CSUsWI4p7jYmwhSs
57mGyFr3+O+NnqnqNf/v+Xfp95tNCz1pogYYN/Af3fNGwJCVKVxCzUExnkNRw0oAHpQhjxgkCtSo
7F9mBKRi5NaqS6K8uIuEnpTnuqbTAfQmXHlK0BbEAEO3OFaJb2P28bQlk3qSdHhAvXqBN3ltsr8O
DUp9r3KtFQyHOv6/MempDYJT/AH4AzBpR83bzJxGN9k35pdYh/3UdjSEYvK+G5YI3VZYWQw5ez1C
PK3ADCRlg24KQd9PDoKAXm1xMufT+auq3pZFP7P49i3NPN0AIzPW1LLaD+fmea5E+qsWegZs59sj
pEbHaHHOaNaa3d8PZS+YrwglrYJX2SJTpunsVWRZQXBFbTKOTrtMcGDAY9zyfhhku9ph/pR3ME3s
GC8X8puj4yFIvM0OhANdhXqCjtSelpCyaXkGRUwyWgZ0zDhHWdNNGXZ1OAqMulYyuT9mknwvyitn
PeFdZ4Fvps4LLTerujDEX9PdDZNXCN32cDSHWBukPrZQYSnox3Sa72ZZ0NfEdScvu+Xg+TgLQ+BN
ht9KH5Aa+07MDXlxXTwuyH33DH6spX8trz6LTajs0P1L6tXG6cu+ULv0NOD7x+dpjidmwFammZZ7
4U9kWmgRgTVi/35nPBUy0m9rLmCW1HEfgim1O4Exhwh5HNLvbFTN9rk2DdhgLSjbmxyD1D797yhJ
/MsIIk1IFUrjfUtZ5fCCg1uMAIbzP7sxseERscYa1MwFezFQm/YJZzIL+/lOvwud4EvncC/2is4C
CNbBa3snmJ42RbqTBi2wQhtaZIPxFyVT7MqvHOV9wG5CCg+uD3TNDCxqkmdSO/rzUp3K+3ZbfgmP
VHB07sh5CiySvZ41d1qWZ1uXCpFgEu3hYnBkdrUiml1sqKN48AImlw616cGPhHcmzXl+5rBjuNB4
bv0czmebtgVqjRmV2NITzBvb2P6eGtU24WncM1JgoznT0r2i14UYmISO4pEQ/fGJ2qhmggG11NcQ
Ni0iOuokELidt4q64IC6/Jfsk0K5X08GbJy7Nh48XcF17J9PUuB1BMGOyl15jaC8iRSquzWIxlvM
AijojExBmQtTYFG1jR8RqthHjokRVkLcBbJc91/S7Leje3Ft/xBYfitzHsx0w2vV0dOmo3HmTl9L
K5Ui4UlMyaH4Or5NWvaWnh4FbBCvFQnyc8Y1Sdo4Cc0tL2EZvHul5tf0AyPRcbQgPLw+c/BW68lD
cN5rZT/vZLrQ2rxCBlUUSNGAEQ8ZBvbUeT+Hwrvxumicx4ztncnjY6FAFSJwKwcSatD1riLpmqM/
/nsv0UFs+q9WRo85gk3OS8DYOS5JJvx7JG9OYrkyWpA8JuLapfPg8ST9zdZn/AecfEgt3NixzsE7
OHwbewKjDKe6+MHLBw68efEZgIRPxjEc9Zh3zCQiK3BMXQVtGMZkAUX0lJ1lH3aB5AoYH6xpcDmg
5Zhcz0tZsBqfM9KjQrHVDeVBD2LvXWkl1/QHJFpehsg2Cn3ab99kSBDlPKax/LRYzbK+ixiXGJlT
qrIHR7RnMzwozVECB8B3YDicy0AhO47VeKQusxH92UnI4SchoII0BPvNRu9J27iIyvqr8epO7Mov
FAOONeGfD/pEgmwCc+uWviKV42k5RdGqRfQV7Y5QYdyBlA8Vvia+IIecl7VYYvs2iMHF1wI+JE5k
d7CpuQiGxtU1WDWo3zxEjdx/dE7RtCOL6GRg/MwNSxV+TjwFrKT7XuKBFCytLzhhctxRkxA3B5th
L4ISRmEoty1YnRs11Gzib4NI/YPVahctdnNr8xethX1Z9AVqU9Vx+1VSM947cZXYLMutY4hWs04g
RoARswyhnz0HZJSx5WJ5u71yz4DZROOa29JOMgCihN45YOlho6fFCa7h55VIV672JLuvXTW0E2k5
bs9xTVi/TWj8TWK5f0DJQXFKfAG7OomS0Sv/Dxcn54winEAI59fnbO4d+slh+cpTJ/6CJig91VIG
avR+lbpnGR2dMr7tx0FigtPAGW/pfYIT0Dyc3ODvJaAbKJrj99TOu0TOqKt8rvMm0qnNDWxsGWHb
of2IWXx7URI4vzgr67jk+qc5piqUQHHaQW6R4Ku+ozEvbgmHZYmGNRTkcs3VF9BWXDbilv0aKvrs
vz2IRgdGJrOf2GyrYyOlkdqj6XZ25Yixmj0ejT6B0FcfQI39HscRH055TVPA9C6+ukHCpcWK6vUQ
acqqrCdCzmslOA89U/GjLz1vmNm9JFCunLe4fy2Myvt5+L0eePV46wHyY2EsBXvFwO6s/x7FayJC
FlIRLk7H7B4n4IbG7SPRDBzMSFukvWaMW0KqOUnmORogdq+0g+s5LIe1JxrH7KrLQk/8bJiH51N9
eIRunym1AvuT3V/GmLkcA2MRcYalDDYe1FTlKLcFjq/VC8AqFC5xNcRE8FxA7nvKYHRMr02fT70X
GY2zaGM2iz11FGdCQjf0XPUOHI1blOqHH3DY5/j41E6Ox015uJXMdL6n7C8vc8+gk70HO/v+16q9
LY11Rfu8p8JqIinoqboJHsTtsBS7bOW/EUlUqVVzs1t+JdwfhctCOZ3IlmaqC653uS9/1GzqO2oE
LS9c8gdDRAcrJhlmFeYzTJGmjMM0I0KF0jYBliJnf5LVEWxEPOsdjJxOOpj31cwh/ttCFe5cSxp7
dO5bxjwFUu46dzsGC2WO7rQY896JDCBBAeF6sXUWQZ1VngJwSGinNqGB9LhWEExNY4jntqQxGYZ6
MyTxhcTrY9v7F3bZXheBe7QDctihExtPIjlNAkXepa+L8MPkgHBWPd/vWazYRqqpNUMvL/Rd1oN9
C33QLoqW3D7tpRE7fIpKKItIKlWfGjmrRbJmx18+KiUKNbOp7hggIuLol3O40JSTPCoXZap8XcX8
SArc6DhkmUelHov9ZrSUt2gyczZGWPuJlbZJRgBXf2nUXvxSatylteDO2/sHbujUiAHjbM2huOW5
d3JtMMUip/GNys4LHLShcg6ssZ/zWDOhG5MCmjcZRanLFiJK3nLABNRtlPlRq3VeV4J6Ja/KOVSM
OWpsR4Bs4HSJ2RcLGmH3nlw3XLKZ2yvbtnZ4HavWJ48mwwJksrRvJnP+82DQ4bQpNOwcL6IYuRi6
D4p4DYqk8qT981uLepIvmFMN8xVVNUjc5YWyV6Dbb3oob4v4nglDTTAM2LSMyQQpozu22Lqbb9GI
Xu7QIeZR3A79y0FCFhGTs/nmOdSskg5BswIPzxiwW0YDZyZNNs/+akwlvR04nLA1r7/w1EKomRzY
N9W/gKb653Y6LlzG8Wf+KwLkyWGNrHCLZQsNsuSv8Y9EpdU8lU8mZCEUcEqw2L8R3DyB5I06Gngi
16dQNeLJfJ6Ubp1vvq3eBYVWOoreUzERBQFDBHXjAIpfGcdQEl49hSuYDN7kHGC2+Jf/qpmvN0JR
91jqHwX3elbJqUBIcgmJsCjc1TTAQ+M0yYTZ0sbnynuNAKfNyZayulxljRq+w07Nd8qwOAhYqfuJ
rmrQvtYYdyhHZ1JZNusZeFlCAEhSqjfDfYxBa5nKo1jQ0Rn8PB1D9YXisNYtx3xFrRiJjtDRROgP
U54ecp8Qlgg7s05CTxHyQYMMiKh7pQLHSWfm2rF6pnvKNZdq0MhDG1hZKxIZTbqNSGNxTh0YKyaJ
gST82uMq3CGrpePwdv2068q+XHtAOKEiIw5Zxz8MYXIH3eMrcMqvTc4ceUmFkQwH4FKgqKzm/cy3
UCEm/ckfFCnq/CXvGkU3w/3U7jsWjmObI81k9c4ldRNl902XFHG52vyq2U5YJjnn5ctT4ZTxk4S2
jh5otIbR/FwPHM8r50Q83ekiEAKG5aVyPtuTtwMif60mgcVpyFJftOw4c25MJzBuH5QO+1ppLtbn
LyMJ1F4JQBU2CPT/t0v1U6IpnJUOCg2eRllz2hpSktdBIeRCBsjLdbm7+JZqOeF+h9SGl++i+a01
PnOrfnBs+tJgE+SWCnLwcwxWXtB1OZ5yn5aSmPgToH4OABDHQMTr5xiBM+YrN6B87gOK4430sELD
7ayi+a/7h88F6uVo/DJ3yK3xuPtsPGGqMykaF6vL8xzr5DDhBE4sLXsnQjYTRvphDQmDh0Fqkxy9
/bSjpTAzkSTmRFAxI+8fHFa0gYSsMGxclL8TM+yNCk21Td51qwhi4jKbuGzwi3sivB7Wjmyvp1M2
1u4ARhYNzMqOwpNcE9d5nXdhuYJj099jaGhP8Kpf6Iej5XEU7PUE0sXodFX9rZOlZU+Df/7jZLg6
dBYrjr0tRtdEoLieR+jQ7KmxHDM0UIwHdsYPXo52vh0YTQNQXZO8tu+3nRGHv38wts6Sm/3TAIV4
xU+f5odbJILLuS/jf1Kut/Lk+erYzjByxSJvCgBf1aeW+r6722iISriMWbAYyRoJg8yomtMxhtXC
yyFMwtCZPZwwPysPSEZVglUqLKSBp9Y27V0JlWDSrAgrJ3ZM3UdsYvQP4zzl2sjeBCduJju2OndJ
Ogbgwjf87+cCk8jqvWyQJsSly68PQUZPwQnIJD9OeCRZYMc1aja/gaKtmYjpRuDQOq0DmDxUYQAx
lV2W5MK2VyuhlMnppPpPg+3XD0J/Av/WOo4Kqror7kAoUo/JjefF8uRqnwdP4fACsXDEHlD2+jro
Domc6UQNywGdNGjgb2Vya0MjDVqonuyj3NNaEZZw25UnWWCEfWbHfjweZkTIXNpTC2qbOvtfb4u0
7UA8AbjDRKsp8KMMTPQrYYQDeDotsQzVk40bgGuoeT9BoRGtnX+X5R8on+9zgWUE6HJepJXrUp9X
O+m107w6KaxGQBedcpG84Tvp9mIE4yfa7OH34jkF9AsFAwEGI5q0Ze8x9LpGMdPiwMABJzShmNOv
d4NCWDMg2CPFQQkTrIuAU6Smmz3kXSyuDpL6EHETL0+5bd4l7Pc3qpy8z+++a9SnOQLjCHDNO/rq
xaE2UGemF6f81MwqHTT/J3ALvcy5c85hDTh+GYcYDw9p7jnQmPYVkquVzVf2BSy80RwNCssUVbTf
unwQhnGxCSm45slumqWsmsdDAK1hjdlQdIqr1G5yDCBOn+pzVsV4112WMjh2HkbYxRskvPPd57wv
GXeW3adxoJwmZQYGx6HArPCsvv6n1sEihaVHjFRP4URYiKzAthMo3ofTn1tYcn9n8GfFedfGceWM
c4HWwqLR2lTNlrK1AKaJjnkN7IhNHqTI3KJf0kGtj/IWHwmJ+vRZ+jMyCKXyOYRnOPcW8UqlfBFq
WguAieHWFC1sq/AAN1nbMC6YIEICZmt4HHVjda2NqF6L9wSZ9z/cuJhIBsljr6E8P42r6/yU9kxS
SE/+fnubZfMnjFC6bYj6pViyQcd7J3BhzMd2nKyuMVgOD5U4acc4ro51pmksBWU8Id6/ybzN9f8P
MWvasmMqKu/6Bg+GPzpw+zTTzglM9TBU3ysRXEF3J+Yr17WoVPcSTGbu/kcAB5qVOpUO5GGUH5+W
jmxTq9ItMrg/LeiSByK3nP/5Ro6ZI2uT+hpCGWxZG4Y6SwTv9WXggvLNT+et44W+99E0tEQPwYee
TW+ECB1tF7B7tXYI8TsLoAN8fADt9DZ//CtE0eWF2NJ0hLVD12YwDHrfrWGJXKrq0A539O4rbIWy
B7oivY3IzcOqfwCeLFghkgHdOK2aGhn2V+CEMilsySrMj3aD7FZDH9e4Z/w8Gg8srJdRGA8VELth
dfj6/cqW6Ev9S64jQF4Bm23cs2xpRuoIf7vHQJg2UYHdKnVnO3rbGWcruur6ebo3pIHVTDN4eLxP
B0iiTXQxNBVXZ3iW7dba4P47I3/Ogyxt1y8SnYo5qnH4d84QcRn+1KigkdXOyAm0dXeYCOTTp2m1
7qwWOfn2nd8asRgHadb45HMXOZDKE8rzz3UnZyaeSyG57TDFzo5ChST9ZQLSZWEZ9MhdEvVjjywT
dkMFbGbGcU3mdiJb/uf3OPe+VzdK+BY1jSP8bv6qxWV3qny+mS5iKGJSj9iTOJult/nV+b27xN6e
LEfnMqGA+7gjm9VVPS1MjnGKsiSBe5fIvMc1ntpIXlYwZIXx7PbCXH7rk13XZVTBry7ahGYdPWCV
fLqHG90QIg9CiuQVAIS9hS3K8kieHSrrC2z9oJn3RUe6ubP8XZ3XKLSLyWbZ71ABSRm8publhjRZ
EctPL24dLjo44zynR3J7Fnq7AaTOvRENnVx7efAvheM9LK8PhyHn5zPLG8GDZV4K3TCaEKyZxeOv
wnnJOP7VF0ZUQgbDXPYDrS7RxQZqRI5mR+hHg9z6KVhX+jF7tvWnNtLts0RLPMOescslcueW4Doz
8cv/DrEPwwVft9CSQJyCFvbehPqD3rji21Eet02VyQTc6nMALoqffKRr/u4c6TEjCiZuzDMChuFx
ipcPWE7Lvom1XCpGHg3DIk2qUzeQukv7cj8k1DTupZpNCgxGLXoI4oP55scZ4qzHfad+qCxfNf3o
J8BcWpjakIirVaV8I+npGPaZeEpvj+3Qmfny9B24Wh8LqhJl0uF+oOfLXhZeHaZfW0FdrAhISSCF
pMSj31NvnXVX0ZxF0sWZPZAWW5Px/Lle6ar9kGutvIiygEsAvKzh+pm4k7HuGtWM5dCXxyuin+fh
zw08N9hZesSiKxS2IHGAeYwYqQ3H/h0slvHRRYr77ZGdSttWwNgjYXAXeN9wwwRcKS0pZLpSMUPw
iVY5VieJRmz4uLP53K2jbD2BoSeMcI2KePb/s7DdPqfHXxh7pQPXs2laTNKcTmIYCjcwgdQdWkSe
arrLsBxt/4uhy8cDZoib4cQLcMJp7lgaxzdiQtyUcLe8PqjnJzwEjD3ALhv2wnhdeaShvPV6q9R7
udju1ZnDEE1wZdeudtywxu9GsIx7rU+O3SCLBa+lmyfhApl35gtJkr7cxxS38GNNGha3iAwsvk8Y
+tQ0OWa5NfoY1e7hJKufQabr58yHPMfdHL9F9GtGi5s4nir94gNHp7AlKE375uHpRhinMQ9CLMm8
wEz43ftIO/691t6PKGSloXposHtnxDz3sPjsadJjKwNdWlzhCaCN3gVW3hXstT+PgZIRrDeaeg1/
Tt1c0C6Pq+g5CxmiZSfGKH8zX36/XqQoxG//e0eRrIU/r53QK96rJByclzO9Uvq0KKDf62ABOEkU
nYH8sZiuzqFNejNRGSoFuf/t8jMOz3s1OOW20KuFSTQmGW00HOdU/Lni5mx7qhgeeAPw1yavLDVw
YATDjDHf378ufuGWQuTG2AA/SL9uaqQAfY472rFDoDQ6Q5M0XlqkfxgCZkAdHxjoZjgj/bwz8Ae3
P0RCfUlYbKzVG0PqfSdwrR6fc1pPi9vqWKrsBJz18BMAgASrQUkqi2up8JymdzoEAypIH7Qrpj8P
KdREv0FrTWruIWkRGS9bR+Ped9tcP3xJmWsIg/14cn2R4W6bRHmCHFVEVTLRyuyCGEhngrjFWymo
kQee8aTNVKBnYMzcLsfclErYL26EXUlyGlXLPjrT86/5opwLM18ViOLMnjkDuq1ZdWRBc878/jZQ
zrT+33y8JJuzTWTdubnu6mL95OD+UQ26+ui/wsh76Yx8RnGdpEebipUaEHR5BCQASEEDHSJMg5+0
roaaERzvlyBZXISWvg985lQ2rbnZQoNjphIps2xhBNhVKtIUyDJPxX7dwMiWDx81qARbrdU7pjsB
FkfykXGOaJQfvRK0tQSFYYThxc8G+/22RJ1BYXf0Kjvgiun0UB7UVZ9HSZ2dS7RmACiwR2tokF6z
c6WTUv3oJACTSP8b5Fju54Tt/CQBAdjlM3i33SCFThYzgZmYMgZ6abnVZvWOoN26o4mZbrUVWMk0
QNjtvH3sY1dsBxOg7OIggPOlHwL5TBPIAnlGyk9uzKV/bsLZV6Z37glOA2F0LocYYbFnZvQ04D3M
9uUD1SVnh2YtKllyL41Cd0NOyDzc7IyCEmDi1GTEwVp46kbwxWPsjtcz0D4hhwezafmxMrZhfxGg
AAu4NGLvGPTotFabCjAIhPgXvHUx5ufqUq2/VYH9YTNM1DFF4iMv9XljSC+gtDgZB6bQ8Sr6PNEB
uayHv6rjxAp7oINbrMYZdXb5RHtAaxpOk8rTVhLF+caZuHX/1aePkYGhAFpEYK2ltdgUPShShJZA
QYDqAurVfpiX/IMWDnc9uKZRUSN0spCRABBdSsqZpFGgGlxFJZaEmlnECBac2YA6Lt6FZVnYCN1k
VDsVBxilF18zcFmmwtxR+ka8Y1fhqrx9Lv7k9AnNb1KWpDJgz7cbgiDQYR/YdcqDWySq6WVu4Iko
ve90NJcRpEotu3w8dOr7CdwaawcASbHSlf9FSBUVbJdpGIIr5+NS0gftSn/JAN5j7c3Vukf4/V4v
zr6HUtJH2DkEquvJ0KpTffWg0klelsUgJwLgPj3kjzm4UnZNvI0/tAS/wcALLlU75sX29uc2n6Pt
HaA586/D+MiF3VJzKtb3C1XAeRiicjf5MVUDjiFTuzuuuEpzkYJehGEi+rKkKV/O6koyuiCe5ke6
DqTPS6kNUzDHDMYCg/BOypZmq7/MdsEsNELOZSJEp+GdU0Pj1dy+Fha0++MCdNjdGnhF1Zzldsx0
OsVsohscP32eeHBZWl3Jq8y4qCngaM0ddQ0ESFsoRVQ43LaP6U+csoPqj8r3rbHQC6zGCFlyV46O
2jberd+4Ez97mrqDj3+Fnsv3mNOp7UD5jQGrk6BhiT3Ecy0axzU8CYDMikZbHCG/5X/KqJncvuvI
MIvX9VzB0oJtPDc8yHlNiYhybhVLdsUu1Qrfyj+MHbhPkTWai+dUPj0m9y9BNYsbKspHw1PrwD5S
eEcSER6krFtcg98yQbNBzTcsnbw0MI0k36uANUqJenPjIdTgyG0e4ziBgZ5ej6F+fI4QYpL4yewf
dlOyqe94bnzD8Ed++IwvLnFUJBH9EPRCbY7Gc/kIHxY3Ig16QvQWWrKtlVkoDCYp1UG5bp8U4DWx
eckQgLEGV+9dTbiPvDf3tlGOqtXnhhBQc3Re231CdAwUYiQOHwwC326pZhICtKvtBZXRzXdbP4I7
5h/tNCiDii2ZJILEf8vNiQdlbcGiv3tsUtNk+duEWCOvq5eC1zKvONdfnHXdFv/k/tRvvbq7eR7n
n4OntSppkBs1MSuw7OvLG7WWQoSNiml+43m95+/N0/dRI/nfIKbbhYrTEtu/9lANp2EutiOK9EzB
e9f4u5YGmYWrX7fY9Ukh2avYKgBaNecyVi7a2pJwTp5Dxb4KkgCsATSPeP53CoxCPiYeWi2jPgkp
BoPzG17CRBxEbvfvJI/xwqBJFtxnzyfoobelx4OjzE2oIHNUg9kVn/ymubC6EOwYjfKug+IZqHxY
DBSK80XwLaecIsviXVCffenjrXh7z7Sf7WLf9gFD+2K1E4XM+Qzy2Go0Ab9wJf06BpWNVB63nn8d
z+BVn+XpowIlP31Neg0LAxtpAl2L5ds0csYXMM+v6OKnBDa2NbcSTZWv0+56HBqo2QQGH5DaZuJf
PVRxks08hUndTdFU6g2Va6jcI9Lr3MIi2SLzfZnzrJdqcACnp+Jss/BB0tXCRlbuFq6sDXiU/2h4
ptZc+vODxUlWEYl71dmrnD/rFOnkVhISB3rkPBeFD5SVMyvG4Si1hQoBkeCxfKyTFsDemgL2CBIs
bOJOtlaUz0IaDxitJPzyMQE4mxciw1/iysaLBTma+x+pLmjXn+i3+7+eurzl4ktSNF1ZaNSXW6F9
R1P5v4eRXayu3ndRilYh8m1JxGpAY8K3DbEgrwxn5MEmURIqZap1AkejROKG+lSceaUJHoTRfHWW
Po/2j3ExzwGMeSSJrauf1BFBF1h+/uY+APjoH8Bk7wPocAgXTeIAk+AoNdNpyBjjNKBcPsFpERaS
pUAFohIGAnEoItjUYeSeO4q0VhHT/EJJdTi8vzRdP6sb7YxfcTolKHvWUl5oKXGQIi46NXTYp8pR
0tU7xJ5JQFtIhHNWDpRiwCtseHI30NHlCjYIb9zZ0QkG3uWQ8bv0kCaidlve+CtUl/2LWFwfPcus
Qaa4KrzYHYxqUCQgUw/PQcm4mWZi+jZOtMrGOm0qddbBjEuBxLJ22SUDOBEWAp9MOtgPOjIHjWWB
lv3F4YiMOa86q3sXvVj6eiHgsQVyvJSk5hLTHzjYp1hAEInyeE+DyK8rRES95xyhcw46fmVwFBZZ
XHVI2YbI3yitG9nRuU0EvQfzZKrTbC8UswPsJGe10GmPtxjZDTwRUhBvRKptCFeP+83XuvcXc3Ph
+AklorxyHXfWZhyIO4L30KXGWdfrtrXT9nZ9i4H9ptmTpmHVywnwMMzg3DtqlQqiK1qo7RlKcGih
GB9/tr195PZQhlm+q3tFhHMdeCl4+66sv5r+FEk74Wfwc2LdZjM1Hh1qd81ysqBqaXVVq5v3fwJy
0H8bRYnCpzUTgv28zkoxMuqg0vKd1vwZrdvm/OYMZmF5ntX4xAkzj1yj+6W5Xa/5gS+yfs6l47m8
aRfHWFVwaaJ4/yU52NOHU6BoBeAQun1KqM5UO+UhVqs8vBBg7TJUX4hCrH9h5TGDZSRvlHSQbEUU
W4CwlA8MssINP23yP8rpX9w7k5H7xSiZmVODY+b2I9R74yKe3z7fhdkQ7ZU09b9jLW75O48aHkci
qx84xmF8/cmUypi3te46LdlA9Lss9ISgbCQRJDb6tXSmnnYnEjNG8vnDd122QW1/py/b+h0lLBPD
f02WHaOlZl1oVU04qzH6KecvHhlKxiBf14JAYXsrsxGhj9cYxbdHpK6VFubJqRV3TX2y9zfVRJ2W
JfYQ4dLfGzyVb1u/6K/+BjDsp0RsQmA8qOKqUEQzZpjar44AlM37YRioxA/xP4L1cOjdNEfnQjIl
rbAU+Xpsot0iWU0lrT3Y5+7LLJkScacJZxewXLbgeQLS/ZigD6y90b8KUMh5QGCtuvEY72L9yoGN
NRxZznu3n5fvPSQAGYrFkG4PKWr2C6iiNu+xl6pWWQK1XZ0L1/V6YPLohpYEIvr8znfsZaiwa23A
AYgeoyyInEa4dZwGokriR8yqVRPWC59tRaXoAYMs0qJEMHl9mp2U4adOGAfjoCnSSPayTh9qeirt
L7tTqmTJKE+MBU8t0lTlyLOXtA/YbVag4aYkTmPce+81wKOm+u6pISHFIhbW5akK3c6xVPq5jALO
/WUf7vl0DiL73F/FglWzwR/0pd61Hfzwfz5kQuib2QuWUyP3lMtXgr2nsiUPH9BhJffsNDuQKPBS
oVEKP69QXtJB4gKKSUbRAWgXXaEyxSUsNfmJ1hHRBc8eiX+qP08i9Gj/6xsizwM8tKH4KWX2FzeV
PPmEnaHHXOkLJLx1nllAZbg6rlAHiHRsK3wa5Hfce1ukctcnIb4up6rnK9xgWPA9B5VkIFjbr46u
R3lZFeGKDxqr0nDgZM7acOr9Jo20xTn0kZrGfglfa4+GXcGBAgvmabOEAv/7RIkv6/NjF7xs1glK
eQLa8/augK5vCMTbenZL5w4F9FN/GiTCK8jC3XiBUoS6jqm6UefPV5x4/G7JBAXnKHrxJtYi6gpd
mvnuMWwaMZUYxdMPpEu9TrkX9Mc4hrKszQWWgkYK5hhN7c+iNM7hAmALB3nwwXE0JLpT5LgQLapc
5ztW4Enw5MXdGTtRcsuE8U4zy8Qnp43UYzYRWbmdfJ+EMgmwPncu2L567ZQMXMKn+dDwd6IULFXN
YF3Fxw9XdEHks6TdAP+8KWxZQpMWv3h7oYFskShQIzx3CxlXGG9AEZ5nHyx5lh8tX3HST77Wjid1
mMzaru7ZkkK5/sFFW+xIL1rzDST8cApN7OLPBtf2lSfGTVh0ytbNBlYwSk6at4qeNWX2T6J5wV61
O4zQFIP8VUH66W9YymTGn8S2YGmgaCNbAUA8OyuLJX0xqbpFhPagJU5lGqcmYEupX1TN9pkglF2y
ggXOvK5mg/6Wd23/vU7/JDWQ2M77qnxwrqrVDlC+PupAkK0Do+IKFczKl4ZzkzfO5K7djBinejeO
tlBBpDb9KCXvozGAz51Cs6644cuSsW75VWLMa87OvSqeuKqjqB0CMq0bhsdi7/Q4sc1H+AjTZo6R
Rzu+hchT86e8JmGgw6J7asZcokf0HE2bX5hRqEYEqnhpLC1mT+67p0sWaKTGZ5AH5uzMQuhgsMEz
fcLaPqfqLBPpXEY/FDzEnxeBuK5Pj/Bo0LdPbJfsH5t8I9wfvUQyklhgfYmTl+WlP16FPN4hgwsW
acF81O8TCHuNsXU2SYBrjfgneWlSVaQC6EZh6WwzpSexHesSp47achq9nIyNA5fDdIAtAKsyLuJW
wAhPp8jwKzDwtuh4UTWXyc+0nvYgM7S3lQxvoo9tYZjb19eVjmeaYlDjM81vuBq3GDW4hKeH50RB
KAc/FUAYPdOyd9NU/SwI8amOJsnGbBD5kzfjoNq/GRxEp+rBbfq2X6/zZZZmkuzCiLW7VpK3/Uxw
3/Qn2mSY3VCXGgORAocyIRGY9zq4N+j7z6PCuQlDyjAtkJxaTuJYKCQlprMyXcRlYPTu/osuJDkI
AFyyBtsPpuiBaYCwlL39vVjYwJFTqq/AqXfkSVOLwbo5Xogt5Zpx0KomRo7Cc3ia7jQnBnEXihVn
ySHTJLOxVEj1m9+9yHVUX3VciYyHEz9fu1wrpTZZ3+K+K5MUzGU10s6XbQy1FFvyBXCZWE5oJSB6
gGXCMPy485tRZw2KPnJeSVyILrOvRxzZW0Dv9Zg/c/E3TDiuOv+1/81fU3hyI+J8Sgoten1VQj+M
gwWwrVvh7luE5a8wHQ+NhnCwagZQZSe+wwrgipnOetp12ZKqBcXSNaRDp5jzi6FwYCGYJQ4gi3Bb
xnef/GYhbCNpo+qCe0PnQBzOc3v488cJS5Leiv4f6GD2K84Z/M3SbYg4+Ila0gyvi4zWVjXBABj0
fVaIDYJdsd0e8qxUMUHeH4qt6bwA1eqC8xmob1QCRuZx/K/dGzo4ADPMtMQybTSSyfYMVgPlKB5n
nlObpjw0c94sMd0ErJwnzPLPREnnI0q/kKPP9IbGl6rjbXH8Dc32dB5LSmxwmYrJtZPsbPfjIX8i
XU2n+efiEQZpReZrieMNStgAVhyGdapV9ieo7lD1tGAHDPWwaLsx1gf847tbAO+ng2oCS9GTau6m
JcnAsBMRDJidmqZ3f/wJwud5qcp5i+6v33r8cMiIvI2VnCbZyzECiTwGnMRI0PMYBbrC/OM8xvN3
SjcEdhnzWYqFGKgkX7DafK5yXIJ+4ZxSVyeOvpIllMVpQjIsJcgG7te0WAJqhrZW9XZ801dNIaCm
c20b1Izgexae/7ZyfrsNrsC3xnb6ngGX5qYbXFcdJ+83DEqJ7jcQ/dWqf6t+2qPyAePJATTL8egq
aAH7cr+vjuHtXOzrVHoOQg8/j62C1VfNYb8pWIn4ptIdF8BZeOfc33SQDBcDayeZUm2puB4qL97o
ABxqetlcoRFsiSDH7CO7dRKUaJyGAU726y/isPWuLF4csTjpRu+U8R7KMDDf5dU7bCLflAVu5MtR
5kGnn3MgnVRmfKfbcjJDLYVj/hTs9od7eZIruOVmZHFj65icuY6H4CdHGwdiDwb0IGQmuihkVUZk
kgg6iFqdTI6TeubJhWqxpgVSkG9tZ2FQrrYsCL4jRCk1gLSxNRPkbId4AA55EOUaBGX+8tGYqFb2
xl+MyjqvBuE+ZoIzWMjHI0YIP4+VIe0+ezxJcCCfuxvgngowJMe7ySbr4cRDeuLWH3eVvdjmRfPg
wVSLDLiV4BSC0w5wv8jrnVmi4GPUG6agBxNRskRiTjXJF1NsyxfZgM+vdD3mSNwW9AkFWa7YzNUu
lQyt+QmOgHMy1K36VkHUgYroc9Tl34OvLPGzUzd+Lp7dRgQOL+Y4HO1hLY/qGuXJMiQc04gYP6gY
VwgWSMPPniMFLCqi8oNcbhNUJfHqMfz96RP8xGnOELY+V7EYGS89J55Yzxvk246EIazZVb3q2U4d
FzeGVrjEY/oxYOkq5oMkwIvLD0p2jxh7/m85sd7jExhFYH2S/5Tj5R1MR/npFTYr5cfOgjJq9lN7
4cZYQ+OW0eYivWupplppYkQyWVLcpKJZLEpX9hTiog8Ao3KmE7Hjo1D1xIfLHjU6Zkmeujh0KzkX
qawh6qDx1k1VPubB3KRgfZSaZswMzYxmHgfMvV6Zp1GgmccSK8mVQM2U4FY5FZurvE0ONpIQyigK
UxejZGxAivoANA7m4WrkoNHzkSKJXCr5E9BIoVFDJDMBnpDUFGrXMetSkq7DgQ54GdDSssm+Jc8L
sD/Axze6iz4rOPaFDdYzYDZ4Fm7TUJXtxCAiJZNCcJvOu/JKoxJcAz3mSJNgOqMDjp81XpJIWNmB
rBAHTYXIYcssaIdonKV8O+fsuMVvdV8ypLs8Frj5oHuhP+P7ByVD6Ftn3fpG6ePrkAgqDJr1ESdY
agnpT9HO3pHzw8WL83227cqeIfvqbcBpa7mIW7l7ZeHjqEgg7seSB+LqUDG2be6UDX6ryY1E2v+0
8dhMY6mpVPTvAMWsE/dTeyKvjsjn1gJIc58/wJJfOIMxnVY2LW7Vo17aA4X1Rg9nkN9cK09BCdEL
RSQ0HspD3BBRezyzZKb4geB/7MefdMt1kwFegln5CkUPjrORmNupyy61Gs4A1kZK/U9KYLJQs0Oa
FB3jAVuK2EmAuiap0SiEM0DgeLD5LtKSKl3Hz8TGhr2TBKcNpFdWLb3UZUWK6j0bXQMaw+v92yq7
/1WhRvc6OSFFX+eW7uqTo4oN5uP7zdY027iCRftl7yROC4g/AO884815oc6PcseawLJmNHKiZKil
c1HG3/4gE9aS5WS2L5bJI5ZOM9IeBT98+37j7r8Cp3M+bMjcD2jCLvFsUNiAPjSxVNwdQU74TJbj
U3U3oCseWFe6IcQpegZlSEXe5ig2+13CoIwTz09E0ts4PfQ6+Am10l4AwSDuBHDbgbnQy4VrWtjK
4gnLmj9eRzlqVZiM+KmJkSKFyDYX56A5dAioAMfZCvLIuVu/KilGUWDp1ICf9mansxW2qUoOfFmx
rhI/Y28p2UL3K91XtSr1qgbzKqlA8ub0wVeRSqyoJwtqR+f9mxGg3xxOCQ5t2wZIk8x8tERIXwwD
kIa5rUi9+BN7pdSbfTg5yLWRvoamOMpqX/lDKHqB+brGaFeDqRjsXnKEkQZvScqYl+1RPqBI077B
7bFY51TR4GYYpPmzmiyzlA5LgT3EiLQphvs4lcEyF8Ltc+GylqGqmDdT8VD+tdY0Uxv2HKrtb9l5
kl7/RiYyoDQafwMur23X4gnHCzlUIR7ellCZT3I7oTVEHstPkfyH8M1SId9pqrb/E1gYCV2b73q3
3edtVOeBlH9SzHpaF62P0s0H+DPHarCVEe/GTHJWhy3KTfu4C4X4TTSjTu/Q5cPGqyPCwgJg7vb2
ypIY9NzTrqvd5q3V3RD2gzNMyH59Mlg+goYs6XAKRTOrjIMnFBsxzJBkB90y6bvTjSZjCkGWXCnY
RrLrsAIvWf1SL105wHeOcpIK0tq+691VTLmwK3SzAxlNnOcoHoAn8Xsc5XCiCaZOQKq1tYDp9VGB
3ONJUm31PE5CB1Dg6DKWL3tSZUcmXXQGiuRiqp5tyaoLdEf1rkFhlq4IDuE/7t/zIs8Peh9lfeLu
IgIx9uG4ZA4ftrshm/BteIHtYH8Xk4h6VkSyoZsyT30MQ0pNXF4O7x+CIxeQEVXnMGIr38UjH0r8
ocp37lrJTwIF7Ys2Ngwya862hPfXN422YmjICrVhGr8aJfQredRd8y/foyYv51tAqFx9KskNe2qf
KjYjtJmxNxVjpEUYI8UvQygpAkJpnNK0/DfJt3WhKHj5yI91zQ5YRSJIuexa/etIVQLFN9ePw4EA
+YvHfk621Pj+tqdtKMT1lgQcZsWaOCexNiAd7W2lC3GIwvuajcNjeRrgNOX85vp5RWvbjQtufYHJ
9IglQV1D9xnR1KAoJoamROMR2UouxP3NPRnaYjLdylL3jlJthSuVCGQgRgWdRz4yHx1TEd/E+wRk
53WCqVgGEXNrVqW9pCUXPXtrakQqiqaF7pahlulL2l2jxkmX7abBkFJw/55Yms6K99qqdDND5Eyr
A2mI9PTfWp1+xAATs9gFqVBNpCK4y196DQwxZqovOHr7jc/bvSLjgtAGNLZyN7Ime+dV7YQptj48
sKV0m3iFkWxslAiq2+EGM1YbXUyom/OjH0Jdtl0IiDneKS4BgwX4a66ASWZWfbF5XZhK4ie8Yq7o
66BqFnpxFOjXg/Varg/JwJR4a+ztDcukTT+Oa+m8J4UPNRsxTFU/ifpX10++Ar0F6QgBXszqk91h
KMeRsPz8Im+1RMdWHKceqfKI95HYsN0mOaz8vQ6fVcy8vJskWga+ysWL0OxtzAPTCQJzjjLbbNoA
XphbJJP5f/Tx495nJCO/vlmDN/SHHYrOuKaY4Tg7faKvEbhTP7fUuADwHgcMOZ9tbzpZdAxqKkqa
0k4MzzoZAXvWc744NahZrGTeOUgOVdsm+Kf7pA08932TSAHcYM9exDPwAz0Y2ZHRD1prVMAG1Fxf
FxK3uVqLQphZZimI2n1QMe3sRUc/Kh/TrDNwLJgjj5cu5qxj+P8kWPmCJ+lHSkBjvc/PYuTHn35A
tVPsym7D4G+/cdAnj0TDDGXzODm9rI7r/0vgj+LhCUCOr251eGESfc3uERdBda/0oPkJNvwO4pzD
9ZGevgtcDkWnOhHTrQJABXquJdouB/ffIihhPMkxa3R9ResXaBw3h6KvqdWCFhnkod4x/r6tsg+o
13aARBfEZG8B69x6LsIrx3hpRndOuHnY7uJWxVtVVT/h9VKd5/m/PxpCIAn7DS/26FyM/IhIkK7X
jbhBrC5mocP8yAdHiIY1NEHsiGXYPh2dAKB14Pdgf+ToHrqmL2/JJ1h4gyldvXqa2A5R498JiSrK
TNSUiq51YsOcewAuJKmxOHqsXZRQmdL5KDmZjw5w2XVkPt0bGow6on9vuEZtnshTsjHj2P7B1p8O
3on6ezg+uPc2+kVxrneGw66Vkm4UwrY2sLBitRwdPdQN+SszeMEO3NyL8VkOUKvTcURpJucX2s6X
PzCC9x5XjZzue7j6DZEtgn9DpgvTptyMYWFw6QgwCn+EGje1DN1uz0xXc2ysm6DfEyT3TQGVWrjS
zbmssF/C2RFz4qxAydNEyxHNu84/TE6+SbMJzQBzYdfQV/KkLaG0RWIJzwXkzloXJ4TVQkGzwbQe
fj5fadz9IUdMdJmxoRAxg2l6X1Q2V0WbTsfG4vNeyBwLEoUu/KYxZuzpMkNWeaxQIwTYWNGdZfgp
5kliL6nfa+5i6I3tOvXNrXrCAPBhrJXHJ7hP2IlVY3Cd0q36K5JrD3CGL2ro6akN77TAS4f3VyTl
VCif88GZLT/QqE6R6iXw8JoPBlmhs++Mf0EeH6p0+jgRcS6tlevrboqhKxjFrsNWg3OH8EBwPxlk
FxiBdD4RN4fRQ5pmIBHngIw2CaH8BJUeJPd5HHZnYM5TWkPuRy5zjvHRpeJANW/f23giP8jL7KVd
lM60QweyRu7exb2NGCGt0zFa7U+6Pw3m1BmADWK0ScT+FV02bLzPjdJ4sMtaIKS7ObUIxqUdCq6e
k1PlSp72VoXOuEiTqmPxdR6iJAqy6SuoFzlLNriFTlsW2haCxrbHM+JjrbV5mzLrxa8f3+lpibpU
W9I+sOQ2uYUccX82VJ/UdNlqTsnetWA2OdqzrTYpRaCYQCsohcaTeREIwVjnHiwYTWRfcWkjNpRC
zD/0lxHTzyzNiUl6SQ486di1zCW54I7gzvTpWNyf8tj9W42z3SPFroA6ZfIg7Gr6PyDfqOVdMAbl
k2EB0KHSfuTFhWioVnKX/g0cqCOGDuiWAelfK45Pork4iqO7lKFcgCJzNYc9ZQLhkraVkr39Y2aE
2zCUopZpnp7NJ4yhjLQ3fzVspMErejqUt/gsZraN2xxmfnBfOjMSJuPUn1ZxHoU6zL1piD8PJDgs
7Kca9mH7NhOvfn4mGB89F5C2owAEmhnz1lB/iMiZEAJv7BUo4EB/Cp46xNWpQO0uGrQ4eB7g8y+c
XLZ5VNWbGIa0LCjY/pUWo/+91aCKTW/SpsxT6PhXdrn8ysmHkXAV3X49UFaNtf0S5zodgwT6olTG
qZ2h33pFPAfEB7u5DJX/aoZTJfKn6V63oM/TkUC1riwl302+sMOdCr/YohmGLlBtVtEEER4of9T4
JNvqfuGvGCdBQQgRA86eWIEl0qOZm+O3u1ERZGiik1Lk6jA+8WiY0YVbrRVG/DvDG+XsZhRxSA0j
XaDbsz3vVSc/8aunYFVRLwmvmMNDVdDEQO1fCh35omE6cgwIy6/4LPRkepN6NY4bciKpDHx7cchu
IBpaVLIFrfhE4qPtZ45iEpBIGOP4jILIm+Nw530haFWheYKE1Ko/eLWmgwECYfLbQgaMNA19qvzg
1AbWEN0t1LXu/rM1kNp37/4evKrpsKNEQf+kXQmiGWOVgDHlyLUGgZ4uabRkv5/WhX5/zX7vwTJW
9/00ne19e2cdkC0YG4piNZQF4o9bHJAG1OaLHjIT4PSyNCr52sdm0AlMulErr8N3b3LLZCngY/lV
CDo/afuefCtq2P4Fqe4yRqZ0HCCzibJnwVBnt+SGjSKsQ5SyFlBOeuNv2jmmCUHH1Y/t0aYzy+dc
68xZ+Fcnu1XoW6myUuT0hqyFAVfnGiYdKeEk7vFfoWW4RXft+o5SMsLv8wwoN5zfQUavp6+hOf9d
AxNfU0IGpRjgztmXz8pdYRHLAqrErvyTPmHyz/f9wYA4UsYLXGJ2dZMaD9h7xLJniyz85gWF3cIU
thoGCdC8ZRWvAm01rRb25AKq2n/sztO1VKGzHZXZMZEdhqYecvtYWT8CTkxK4mo71VkZPtd7JQ1W
lw/XofsdHxNGMI6jXCQxIVRNV7GtLCDVM+ifCPh1eUKJYC14k3DWrZrnEuzyf8pr+cHnqzdfd1yi
2cK57P5KRyKtRxADIuYgsrFJSysY0901A9nWXZPge/bZ3z5iDV1HABxy2uWCYn0xHtD5/xETR6Ye
wTGmH8d3I1Y/FkF+jBGxaKZ5xGliJ8mp7Ds5ory2uVnD8EOHPjMvMaHT4NsLldkNhuJkRrCAbgNq
9TpkBtTZeA4KT3xf7z5gtVH6pRz7Moyaq+ESQAVDsUN7z0Ct4fHu5d2mwr7UbGgO8Y3Q7zGb1JPU
n2dQilOckFa3vGPUSv537+LzSqWK9EpZr52h5QHEQPSsOC2S6hxPrWzYvA1LI+mrKO68rjhvCpwk
OdjGrOmXUIt8nOGT2sPqI6PMTm6Xe1FAZcW6edyQUUNG0kYFl9WDjsHrePSCm+jLGKTQTOjp3nCI
d5NQKcDLRIFY1mvyr6dJ4oq8RgB1yzleM26AxxjAsL5/UXXm2P6zw9xEy27a1NRDrcEJ71h7cN1f
VmL5iavKej5VEsC15wZX2UwNwHO0RrWr7Jzdx4Xt9Rp38EH9Jic9jJUGK6kwts5AOKMUcRX87q5+
K5MNfioe1oZBg11PhM/MQn7T8viScBUx73N9cuwa4xCwPvhgoRa2F+epTc4uZC6Cvjr19EKcdvob
p33mURXuQjtpBhvN11B61cLzXe6p/iLwzU8Uj+qXDorbJwGbBen2sqTdt++QK3gTxxBwMsQ45Z2+
QDcW3kDdbx/mxfarvwlWN4yYmKh+F+VsO1DpwbBCYZDiwZtG5jaizS2+Ik6jc8hYSKPJ07XIP7ZJ
IzXo7oeU0r/3DKMJOlL0Rc8PgVTKJpPevOvxu+MQBY7Mh+ZVFxOFiyIvERMUNvtSSfFVcExgxFo2
JHITOzE/L3kb/nKpUlYSkSVCLFhYTHs9ZZKi0ZOEDkvRBwU1CrK1b8dDohzo0GTnIKrqahLuMStO
Se6WAKKaBS/n59EuKWPTXd+mpTBg7v8XeQJnelUyZeNr51XdLPcKhsvemyasJY3K+vv8dEPeXbzQ
SLsJNFhELsswfaOUwO7E9kP4SQqUwwa0S4Ur5eliS0ite/LLHNji4Yoy6uMVht5qvFsOax4fR3Ol
+n+f92dzkGKiU+hBZuZfBLwrZ/y3Br7FWzt8V6Ji+mO223dkpN0oNcfMOvryKtIOVrhw3IAKmen6
uqSvxa3rQe4B/XJPpp4yMOgrFMqMy3H2pMmeUohFTi51rqmzApqfLfx0KNFjIX65k5IFvV7QkP8C
ft+YsQJ5uNMh+smJa98van3Kqltht/qbFGK+RPFtl1U2nruiQiX3PVKrTEbxrE5gpBD9b2tltU91
A51hzvx182tBj3uHw8r9j5L8fz89ctZYgQM/jpAvw4H6VLNSeJRTDO9Vo0IZeqrBjm1BthoC97Ut
orB+hzTinNJYWPyl0aOsPXGJLIjVRofa4DLXaZc2jkFR71t4cJw6HvRu9RS/ABCow8XCYhEteMKN
BfBsXUJpFjSdd7yJT3tP6PMzi13r/aHxya8VM5GVuQAmdbmQTFpQwdsfDGcPBqXGTPL07EsulhIO
MLAmg0i29y9LWqimuO8nKyjR8QLkJmWuKzpWGgMMM3bjrWnegWYSDHd25fAEXp/+vuSc5wEv3AW4
olCI1WQ509QHoFtHnZh01hRG1ugLOkxe0RiB0Flckq9hH3PjBRF4azouO2EbZMlh6DGLTAcIIs/a
s1+F8+ho2Yylbv+enenaM0VMW+4vS8PPDP9oSg8OWP7APC4R6daYULY4xhDGqDzmZAcrR92XbsPj
VWvf+Kq9G0sNkH02o0U8pcpiov1xYw2yJF5R6bK1nVgglbo5JpygORJyWeic5XjVvEkFD8elaUs9
KdUwegGadAkzzIFJbZ0pdOFpC0Bg/kFOlbCQuvaM+A7TVsa1mCr6opANcdqzfsabzw7wQ/783fQo
jpMjQJEoARBWxlWGxMuy5aaXiuST1NujFbvOdCn1JQnBC64fWHCEmT24Y9CdoEgcc7C41qwSjfHl
x8aIai/SnhNX/m69i7mD3mI6b5RtJ1/ZU9GXEJymAnP/VvEOa7x1gxfB2zPswF9PI+3srMdF+Zfl
4f4AGtrnu6bP3BtQfqMS/L7Xtoj2XcV4AcS6A+h+3XD8/fLpjcaOG0NZFbU4cOAha9CCdQ2K57X1
abeBfSo+EV/GjFyuvhS2T8clPYPfhxCmvkG8hPD6Gksg3N9SyOeaZ3xwRIOBZNLuJDBIZVfUL8Ll
lfD8yMN+pz5MjCXfi8bogn8nVmjs0fdDKV8/f75cYd/HOG9hs/Ro0/1/ETk4Dgs2kHM0JPS5PIti
Rvpp9bsTMXTmP4YdX5DHXIQhjllMoa3XBzH4/nRd286JbpIQr7Yt0cZzCNJQik8LuaKZ7fAtzE+X
4rEW0a0N5vEmn21HBq7UZRMvIUJMXQXWauyJlhCOH7/d5f7D5jYzUiUUiGA07o4sB1OuLn0pCd3Y
OK4dva8fqvUmR3ZoBRb0Xg2LbSnzTjbH9jntUcQNeN7bITZLjmCoWE5DiCZCFt0jOvQHqm1G4CjA
Py3XECjJhpxV3gZETnBitU3o+PymRMKnx1FFTrcfypudwJEOMXp9IlFv3gKW1Ex+p7M6FkBfqtNc
FraokqHzC6I7Qe0iXr9L96l3KJLRyPh6/OBXrVs02C9M3+VVmNUrYgsyTB/5gaO1nw521ln7orjf
UeqprILUqonMbyuEVPnDvpumY9ymTqlfD7oNH9axEhCXTm7x/ih58tVqzSMKGuWf911kVCnkMYNa
7Fg5NA/TWHzJhvqXckK9SIAmILd9p8dJ2bubLDuCcVEvx7PV5KUQ2TjGWcg/wCThm1eSbqGspaNO
Eukc5yZ0EVYt1qsz8lqfgbtWdUUlX7ZrTzIGuzzKk9vDj1itY6XS8AIFDhYe9hrRGeCQCD8TcwAo
Ir9QKDfc3g5uM2tC+8Gr/2ycPb6F1s02JATzJFWEoMolcTVqJxWJ3wzrWv5AVAnOOfUZmnFPBXI7
zNv5Yij69Wn86FsHZjJLhkiiV1yuDGhxyz2Ari/lMt3sJuQKfUAjVMPdzp5SLxoRSAMWjJWSjSL9
i4j9PgmW+BxwdUOD0uqW/SgL7XeEWxLRWbG2klTYtkRNl54odvDkPRT5jpDuRIBMzR9vjB9hjjWg
vRD3RGToGg6TCIhYkLkaHkSeva0gANcYmiCftXWg8odR3oh4Hth6EXkI1hHBXMFGkZUXHGnnxaSg
bsF4V2gqTNp1hPnGw9vEbKCY8IKn993f9Ze2Xdu0yfUn7np1gVbRUu5cjDOLdeQsncLhMI1iCqW3
+lbp+Ols/1w2J/IdX2JDc0TXkfDghbvXuADsY+FBQ4X67+Hcgeoqa/OMZjJFHJk7qTo4qawh5ZUU
PAhcEgen+3aemJAHGcB0c5/rMPCG1NSrlAGf2OnqD6iEkcevMy+EN6feuPm4AAUsTVpby3ksms9x
X6RAqCKJ4W+NZv/2WGDQKPZNTy8i7pkCcltku+6xytGmR87ccDBSLi1bdwVVLyJSeWccdCqT4VSw
KeNQqyOLUF1Hal1076NcubBD9mIemHnrc/0FeQ2gvcIQP1GtI74y5wRBd0h6V6B7Xy8p8z3mB8NH
nB4fRtzzGBgvU2eZfIBQOxHy/D416D4ZFRztTBqnDxNIJfYxexS25kQ0cgbFbD9mVCwrneqOjGTV
OJIC577iBJyb7x2o8zxi1NvfwDFIxdD28qrx9UCUcUnofaUMoKcCIiclaq8ilGz1I8BLw+XGaSKk
FGYFOR8r6Xe4u3gVsXyrmBo9UIGEODDFOlQYfLDj7MmfDVtYeUaJhVre77u8kFdUUndU/4U/frhZ
I7+fKewLWuJJCDbthsCX1paaRuS+AD3ew/EuNEv+XlkpqErExE4YbnxU/SIC9SxXTN0V3C7+/iiQ
6sSypw1DqfaMtAwDgq+PTfBlhpGNWxmKJA81CPPIByTCTGSGTzobwIEjvwiHU8lltJv/K1uzwMrH
CLnvEdBNwOcoqoigI4fNKUdPNtJobY1bOjZidAjN8DqkGqzF6VjVg4pPH/mNxQMI+KNXV6xXm8cw
XpiGmZRJZHo4i7o9Z755X0FP42yTg6ZNs1BwvHaSLrs9JQiIBsvEGTLIN5WiNiXO3xNSDCezSe1M
ObgzxseFOvY3fi01UXOW1SkAxOYSv21QTsq5I4XzRFFVH1Mtyj2K0TacaxSEav+zGfs1oVFGjldY
wwSb/dc2e9Qx4E06M30wdG4SmfhYtY230qR1+tCrguaPqamp0MfwfocfZYwFLzGs21uNYYfTedTF
RXO06ufd1oejjTdbqw0PmsXo289cQaA9i6PujCic6vCkqTQR79So4ZoPZvonBPAU8lVh+NlFdFPC
acmZqL59fKryZhRHJcRMt+jyWXRNwson69VA3rMRPaV05qYnrbDrs5M6VkUUx6WOGiuaZ2wTI/IU
DmxfgaxoDZMq7qxBg6VaJqUfgXR+5jS5v+HJdetCD/f2HmUQ22drPTOji+Rv1q6HFnxDDtsXLkUW
XJ/PNUhnqXH4CBE030mil0dDDlKagrGLG3jDzX3WR2K/fskdkMl4OpbC6h8+n9jLE90/bBHiQMY8
WjSUsFGGHo11yJZW5SWjMWwD2RCrgjk3vytpTLf0HtanJu8nhx88FQj1qYG0vVAptuSWpnPUUSK4
ieTG9Tt387pl2Cz45Rd0AX6g4G0HukRmRrUoVhWdVi0OReyznd4HsK6tbSG6JJyNGOES7ewEs1Zz
Mo1pkEJPMD4bDhUSEaTxf6pVVOPxfkbt2YmmuzYwCMQcYJ6vCl1OsQt1OWzw3Tu2Dd7yGXTFDDx6
qok4MDNq8ghB35q8KLEcWqzbC15gZuM9rRp64K+nQq16GVbujb9ZCDudNBCKzLZ1YmqdvLRiED2G
I/kO1UNCzsp4VvXX0kIHJa7PWEMq9XK1me0EEy/89fmwE7mmtRjbndyXGKyBRhQdKmTpeAnKikKp
wJUKAjKZWIKJSoSTwVjAM5OlzevTX7qCeT7xTKBJUJ+52SAR6gnwGZFkm96zksb0cALKskBTRQHZ
WwY9M/fCe39Uhzc72ID62suWtRiIUfsJZtYwvluHUooVASaxPfTP+iIZTpIMQwes5GJmECbwXX5k
XvIfa34tyHiY+32b8BeM8TqyGozkvc2cf4JP+Jai4gnRImb2Syi1MSlKzN19HdlAt470OpFBsSnC
UN6FbbZpuuuM5rEhVqeFMut7UOXTmNh9zx/lnip7VBVH+GWNR4fpsm16gYHM/VtERdOHTJLDyRDn
6HFF4FxxTdq/3Wd7VNrYi53OGpRJ5s0kczDHTPZr0pXJjpm/Np5frRYSfQ5P9cg4FtDmxQyCtTwI
s2vAMozMG+63F/wbDD5XcN+1OzwtCtjLlQyZAYiXUgj8dYV1V2r4j7+pg+W1HXJcFgSSUceb18Vg
CAYwZTyHyf5h7mts6gKYpVnTdyh6n5h0Q/mOtloVU2yyJ6W/5JtH3gfpQKZKNnuqbIfpRGrAOxQ9
5k5FCfZIslSvshbNjvUFMplR8Y0Vf5Z7K5kvaAJ6FqT4F+hzA2UgzaZWSonDbT/5hhwsqdJJz4X/
1Je4ZlGwMWbn28YtDODdCV5bK/2W5r8kMC7viyV6cILem5tiKeI8OecuQsrInXN1tlaaM4847Qo0
wY9l5Y3Yf4/WiFjoXbaamEUV8xokC6uHqOVqFga2QeGqRww9jyx/iy4qY9zYGU4cNj1xAzR59HuB
ZziI1aaFq6Hz+c0TNNF5lhVoamTQJMNVwch1a0+8nbnGr94GQodL2kbAqEkYcsPBFdt3E4gK3acY
fxbBN+gvK8Dfb25eZqnP4MwGIP2oRZtLta3h6ae2KAiZhQSYinO8dk6kaZo/mg7FGhwnRpFyQ7C5
fMb2NEzHliGLK9vDbn9FBmjRH/AB6jXwKgK6KqZnpvsxb0iytv++heYwYQ8NfSdBBbDAYxOvStQ4
LPMmRpiVuwb8D72AiWhaPrME3BGysq9p6vw+b5RURSDLrzmxyem+gMfAcVXGiFyZbgSIp88HUW/X
JXd7cvMgRjg5mftnN+9zN+UD3pRiC8HoxKdpYtWgZj2tgSpCHz/NpORx8yweQoc/jj6oGldCrgNm
SFsBsB9upvYu++sbGaS8ZAJIWqgVrS4/jJU8b0GdsIwaqqt3y/rLIrsniBl10ndkfw+LyeVQva7O
q388AWLsbbMPdnEPm4JnQICEulBLqtoimPZ21yHf/W3t6GisFToQDPgHUozj0H8KoSYYFB4kSiiZ
D6ns6zoYNZ/4NEsEQiVYyMuIcynuSrKBij8LU1y3GiyXR+lAhnjWqo7lIW/mdYXnbyet6BbBaMT1
ttnlVFtBkivuNekITc0ph31UlR9qjhEl5kYkL/iewVnk8FNVGp3KWkRNGVGsQ2k//vXO1kJAk9cY
JLZxLJxwxnFGjjOba5OH0mox+f4BPCCbtdixhMFOCaUVY9vqTRsgT3f4YQXsYoqTuWUXfl30q7aP
AEFiFHQYaMRwP0bIkxHD9X7eWxbQ0JgD8VJy/3k7+4jzLfdRMa3ieJb3HqDn+akvdFqWUp0SUuc6
TJoMVTVUigIACu0fyo9n+o4JiOUKYuoMqrzhj07Uxe+ffChqaKl+VXhd4N3c9vtFXKWGmP9BcWd6
h9Y71OozC6SCQR1hR4c4MqLIvo/L8Kjwc4VHjUIW9nLvLOZW8L/V0clweRBofgoweUymL0UJ+Gnl
MYPPTZtn1t9zOMiFS8wDsoQJ8Adwp4SqZalv1PZAr+MUPo8tBc7dtkYtmOXIHY1A82mYlN7tp3m5
ujf4jQmgKqnjDILOESSRqaLlO7RD/LZNN41gZs1zdSr0Pdl/QZM15+eeERd+XkxMsW06B1hhay5W
rJ04A6X75Gj+8Vni7u2a5cmmJ4Vwko2M5TIGNYsVqRtraoYD1p3cOUUN7MhZ4Mn2lUhABf9JGdgU
CT8QukCShIH5QsBQdzNebalT2z9k9YlIKawkF2r/RClTUmlohMB2OXObVg1IU6e1z1gApuseHEoa
+QsF7NdPiA6aFuoxOKBSvXfE1L6qBQGymYEv5i7rZSltIIL9eeT4QlPi5UDIM2fbuZPsqKx2gqZX
rag8EUsuavtiRFMfUnWJXDotKdudM4OYmVgYIgsqh/PmaN3oOXUsHQtm612A3+ElrabcRTjW8Z17
FuOFlor+tSM+arQkN/4rpycjj7pBtqNDvDRNf/pkMr25arDPratVrvcUhgA2+GDBZPNzyrRZb2DC
3/pMNoXiSQhr5wTc8xQLnuqdCGwMoh8DfD11FfE0FZnlRql33qpuVSIEc3trYH8IoIe+BXXvLju9
O65//1uSZlT0AYyw6hHhxa+8VuBmO0/IGAz10i8xlJ9kxLHOBf5AYvd5FI4sldWHv4SZxGLUMIrj
UfWJEvemwzpbiduHWTvJgzeZEAUsEo34stUemp29/WTh7PlD3AR7HN9JlHr1ZAJwkR+Gb0O9CwmQ
MXlVUfk/IHLbfCPDWA9Pb1WCZ1uPxVmzpMTLm0i0dedhAc6cJ7O6xTkQiY2BfsP8nFprxQjxfXgE
gznHEtwrCTyg6QTrJeDoeWTqyvv/P/ncJ/OIPUzJP9Z7GFSc3HWaSZjoTLUhp3FMm3KYAGcXiJAv
uGA6NvZtZIJUVb9U5BY7YkqiOhBtbGO6nMiSveW9T1xo7Cxf9KEonmulZkqo1S4O0QQbrXHXeN9O
m4QgUV1lm+P2Tge1zc6pHm0WMaJi+6wIibmWeB8CqQifHe3dTxYfIMfMC/eKeBrr9TiWprK4wP9f
A4buG6/3hTYoQIJ3cAllWLFaNsUibbKaZe3LQnzDLEWx2H/njLKRsJlNJnYe9JL5h63rxlRwmQex
M4BdXQwJ6SFciKCV9vl9uoJkSeDj0EJJxlJE5sMWeio+VjsgrilGsT29ydsFRzaTLbNlIs7skvUr
Mf+PlKdFwPVHaZz3651ax9YxTVmAwoOofeHV4Jt04VzBbYtdlB7Ty/kzZ2mVtQ7QsQO05ExmbA6P
WrrKWoftICdcfOhy33kQh0jHcczzaRZw8LjDTw6y2VppCfg6Sjx+xzJrEezV4+ubL6I/dnunqcuY
Q003vWJ+4s1GZbcTQlR7bjxAizYs0bqKoSvwF8XoYOXW4Xnneniai1RHDWcog6Ilu26T+1RwcrSm
896IETHSo8zbOuLRdOJx9k8IKtnjzc9eiMXy1kZP2SL/qLhracochYl0iwYOmH3vriQarWh8+7rP
mZWtnRzQPaoH5LMa1kw2RzL5iGyIi7bN0d3bxHtI2EKGG1rSkIsDABxOxV/Fz2gv1ekKZjitunz6
GW/ihg1w2sR38fy1EQk/+035gfF9t1Xx4MDUUv19bhIinooryTjioaUq0uugTQhx1ZDORHeDwBH7
k+da7LxHfQC3V0I/vwHwuV/Ba3pNkXD5PC9rH7koKrfPgLlJ0C/aL8dGKTjP9tcDO5lAlW5HXNjH
f/khfDpCH4EdE6bRFrtHcyyr/uH6tDzzAfSyXvCiA3pxz/hr35ySDO619ERyemnDIYUKNxd4recN
ZfUQWBYLOkA6hlCbu8DcxFXh6pJeCzEDUh4NA+szkgMx3M4C4ubkJFoD9l3Y3s/ZIiF141Bxdfdg
fdvJNDXo9kJsUSUpx05dQ9llHDOOJ4ZfjrWet4vW8YYWy52dG+THWGyjaeVuhGcmK3cdH2pdnUtf
bDDdBLGBTRULnXtPaQUGez7shsoTXB1MuW7fjbUH9YBzHVSrHN5DduLiwIYkkFK4zYW4h+P0OKxB
rsuZwALnfjt0mGMqhzMEMsnj9D6lw++RZwvKo74ehXz02BjwVoLYHcGTa7g7PMMwVkdCNYzuC/dB
RDcC8urNYOdVI+VGdAede3FfDgXw9wscfTX1cyzJ1bzWnnPBXVI4sigxDWCdMsVf0Q5SsA3nQ8kT
gQZ0mVBzHSnBdbClr0wOk/WwIpHTZqrDcwK07VkwOHao4/UK6K8S9croxe8auptTf0RpolIFN4lt
dUOoXKsXGCeL2ppst4VrTq6mnz5uWyA/yBdXB3bjl/TT5+U45Zo8dBQCURRD3i/F6GO2k6RsvddH
yIDve4BUuxnGie9yCgbX0zMon+e+cMACCzJqXuAXt/0p8qBmzd5QSCskDZzP0kdQuK4gHzJrN3yn
pkvaRclz8qIy9dClFIVpasddExIs2UoswQeo8NOAvVPTZNSHY8RfZphlCqMRvh1qcuOKet4371AD
FApfQTN1YO3ORCQbBKmKbHiXaKy3Ixkooq5CUSKbwdkJ/7Lsfm/7oSPvHwcI3ooZp1LNIsFfiUq/
t4ao86a68cznkKTamMd0AYo14AIR/Nvd3+tSjyN8Wb/6o4aQKDxsqPAjEzqytenit6KgSKlq2oDK
TUk+UxjxMZmN4sSzNkWT1VZd3U4Cb0F7uIaVB36DsN/uCkCBi1YV54eVLPRqsDbsAtWNlVC2VdrX
5ZRDU7JjJyAa0mVbgHsvNVLYyfmRbGniNUV6dYRhEHV3OFfcpLGNz0e2E3tvUuPpcNt+Q8kmIIKE
MZyH9Wl0gVrVjIwkQgl1ZrbZSdK5FzC/eKtBTdj3Pv/14nHo94xm4QCaGbiJZRpqnU5xxHI8ORYJ
g1YT6clphemL75yophoiHeGg0gLw6gjKPm97v5ILsJjKowOmWTzAJJDcnPAjpzdXwfYoQvqrxsz5
XcxnEQyRDK73x7Yiu9sYdOXZmcCa3TXcaqSYl5OzcGSdqPycG4nJWEiH2YUv/cDILKya779C4M6P
xGmFxrQeI/z5zAEZNDfatddA8+o5d/7MNdHLY6+K+DeMbsN19PqTSlaijBzLWMrR6R5X8UsXAXZ6
wKzZsMTQyVvCrsGMT9iT+o55A7rwdLgCDt1a0thM+NJnmw7x4xEKguilHW3QDLrKGPORfKYHRY9q
zGdYmleCPt04LalYs0PdOvrTFa009W7UuSmbH05WoGzx8uZpdHhSsFKfPDZytL3qyQPtQUT7koz4
jL4nxBKTQuaLbnPAVbaqZfbXZk2fjLukTvcHMDnksw2oaZiPSbNFPmCPLPKSLjKfeyg7FmrZ1//L
B8vQIQ9bXVPEjt4ll2IdUGx9KX1xYUdqDs3F46FCfgG9wZHpGzE59LJt0HOPqi2AjxjD4yFztlrE
9vox+Dy+Tlv9cLXT0BUS2jIY9jqwvbloMsARz50z6HIXycpDVGSOT30iM65pcqNbSJ/Gma7leATg
Z3eY/9yPqC4++gWBRy6AXKtdtaimsAHyljewJg6CspyLna457eoAeex1Y5VARE9Hch+0kNQVtPmI
7j/xGKPD6XKXibzO5qmyFpLYWZzET1bx0TNf2552hbZDC1hamAsR0hqL7H5DPlgAXewH9aBsEasz
GQvPu/5gqEtIRXvEQ7rvZ+VppchzMdNZcvO/OouSIxJTyJJVTQySEo+9AcgaViJGwVpP17Vu8IF0
NMtQQMcp8IBfwknks9GfOd437L+yyqYGJQtboWtiyUA+gh07Wdwxyc55XkpYN7+DWcmK+tFPQR8s
ZTFUGH1MaKbtdoWQeQvwm+nxIgXJ9/Na9pXEf30TlsZPj4rVrmkfD5zQwfofqXLKzd2JQe+dxLl3
6dokY0pHj1cP0vKswfT6LzWO20kL52R2HshkoTFbEjkkud6+K1+jxmCRFjOttbMnEn3sFJ5mTX2b
9in5g47EeWmMYGRuYXDHWGc4QCc57Z9hEKJ/FvKkkaGC8rf5DDh45BF1Goih0XXQOjx/3GH/u21F
muzKqZ7fSV+z8XLNkK4BIfW7xO8l+2GUFMFUJcYwpoYAs4+bSla6UJAttbVg++XVCwiI/JtR5/PP
df12ohNCbyKxzb2CkstZSGIyOOGZutpAW0jMey4EVK7ZQ+mCjzu5fl1liMTEijghGYXNZceDGGkn
I4vc83Qv/u7/s4NOaoU1d1gp7zwkMSqUvY9Pr+du/VbGaSY8B0NxpjKEGmkqrHbgYETNZPOzRNy6
sVjz3TDZpjxewBahoqc8j6yF2Sux3F68Yn79NpNZNGen2uO+tNpAFoX/77FnLYPk8dlG5O6uqc98
A3QLVo/lmuYJ5kO0n3ezEhPEPsglolwlWQuh67yf510nR99XWsW+ei4xO1dqTKBgWcao2bW5TqtK
dmeehJMbDc0Oy1N+kSAiiEnV2bwKmasBwnQQfHkPDPRJID89a5fwA/KXD2OC0gBZ/EnKWccwJOqP
BCrfj5obvSbDxXA1klQxEcA0C9R/ub/ao/rZXgATo5iwX6BNBtsGZPTYNQX3bnJ11vPHNGP1jS6x
Wgmugx3tPqqSJ6w3WjaylxMemBZ2f6lqAmAbqWsbNimnIRABni50WE4/kCyqm7hSNxbn9T4BIUd8
4627NkFZudJ82O0/lGnGpmz4xLFzgCpFjIuIxzlvy5xUL1u4D1hM1xLDL6Eh8YaY7k9TULEzShzz
DxRlN8CgnuF67GaLjr/AWP0+ZSva0y5NN3SQAuwz7sbPySPYKFYUpT0pkCDufq0/C36aVpyJRyZx
g+sTK97Y1DfmoE0J36LDD+fxpbxe5H4eiS3t/ChuUmSNX5lp/R4ZZHypbEmI1Knbi/N/mnOwMRjc
qGmVK3NrhBdi3o16rSS0XBuVJt8XugdsppwgvjcDAeG2exssgOyRR8Ch2NukZVaVY0cMk5S50sN9
pk4At2XKbVD+Nerbdc7ZxTfUynrd5Q6bcoU4urlmnrjDnowgNfQ6Hdxro7H8m7C0T70iftdnDXw7
UddOqh5UBPM5LBbSiSfoaXhmvv+H3t0SihJBR2Ti6NgXN9VyRN+rO6O3hHVIbumYl4T7wR7CEeVh
O4QFu8/x3Qe9F9hVRCDfL4UascdJpVH12y/QY6pW0yx+z7NYD5gt4xr1ZdI85+am4sEwLS7Mo7YU
N0NWo2W5lhgtcMSjLLcC4CHGtoZRtJLdMcsnoP4GfR33824rLcsjaFJ7Ap6YIBJOxJ9+31M6oeDU
QYCRDY2BlPTK7+l+xz6JPMjXlPTQJ+t5I8NVj0aaT62dG4ztXS9OumThlkSbSs99pwq9iCktIQqY
HfnImrTJaDNlHo/JsvVo//GETkSvqjdKc69aZrQL+iuJbRnx8bwrUfUXICFm/u8Tck2lx5ngEakj
slEZvNiBe+l/qCleoeZz1mQrVPSKq8KD5P5gioYZACwYloyerpqkXC9+IO9Zy5U7xh8YbMe9UPzm
uDEn+oJs8f62cLnkDQJQgzGjYqYt7wlPGQOLCDsPJECtQYqu/zawRDfi8QWQfS8F4fc0pOt/JkO5
HfqcWw2QBqnSuhuWkfm6tBAlQF4EFxvBkNoXpfLpgiFH9wqb7Pyj0ZAXulrMYO+hDHtlrAcPz3t9
7lxfWV3UL/+ZrfrWFJ4rnjUrDvzbFvGXZ+jWbECJi2rFFxHap4FU/Vhcsg8NSf2EtFhVepBI6F4R
ImUDa6wcEDH8A9+nJezmtlLufl7xzAnOogOlj6hlBW2J9577Y4xoAmD9GiMa7aUx+SJxxmRYhcT+
6X4BIDx1B4Juq9Qu3HhrfNxM1kc8cj7TERl9DWBmqZmzeVqMnYhACtWP9qORQEi28KalKXbAAAym
Az+tscXK4WQagb9UF85ymzGP/6H386GOyIlcdlzzyea/t+DF8D3mFunsfp7gqwOZLmNdBV3kDbcq
XTiXIhT8gQPzLSj7kX38kLtrr8Y1ievXvADRlNp0xsOSKDaEfbwtsEpyhKyDxqEprTOUDftoMBFc
ImY+fpd1wH4QaC01Hds2bKktfduVeyLe9ph1QBEn28DQhDdCQQqr1OMy7Bpwxq+mzCIvuU6oUxRA
5N1SE+oMXthTJNchZeEz9sHNXzPtL3YSJ7NyGzZ9bX3TQa88p+8FvFY+jJN9no9BddIwGK8e199Z
7C5LV9BtCbCnsu60uUkZpJTMBXpVocmFOzfQoP/clzwElLPNx2fFqh0eNVhsl24btEvudgFNbkwt
FD3fqJXVh54tEV0t03Me2nJWN/k3wsHn7+jDHLdrb7zptF1vi79hPOjatqzL/HyE9/QRfdMBgATX
ts62lMjv0Z3TDO1xjfhpJ90+apARsq8z/ZRRjHEyzrqCjlYrwGahYbJZJk4gjXYxoH43UKUFPSvO
fjuBSsKTFlVwzw+9HECp7M/oBIA8rUdULpB6xaDL+5fS2E1TInUEtqMk3Gn1Vnkxb8waIc/BABYn
a9IYWTNZH22Orxyqj4aL/y87o71SfiX2J17+Ag/CVVQKXVnBgtXW9IxL/9pLwQHJP8PHDZ521ZC9
+mCoxzEqmvl8wofapDFUhs9hfsS9STFFyDWJpSeNd4S23ix2zc0A4gL9kJ1cKLvvvZqkCEUzwtW8
Utvd7pblnfDXnisJ1ntnUsG2eTfVlpzKsyt5DYtu/Q5wkrB+ypcThHOXzYWnaSlL0NjOd35Q+Unq
dKmS3yYemqwmASTR1UWca4qTcZCmeQ2YRIKA0xz2VHWv3PKAU8tfZsEklAPYhl0M1PbUACWdKAm3
4jvdSqGJ5beUcmKZVHRG0c2vhBrwEkcIqzlBKiCCmkpmdapVQdcjgc8e2+8YjCe2K15VImG2qsM+
T2YUzP94PNZaXaPZ4eFGY7Elfu6eTImXI4+WKHVSuiTwzsn0WorKohfOTOoQ81DY3gBK53jaOpdU
8sSZLHnOhl79voZuxF58s1gs0UYa9V5r5shiOdRLPmkUjh3Hqazfs0MC25G2QUEGXEIVo/PQWT0m
+XN9qiACjmVBuuk35ihpS9JSyoby3lOqy8HzU9mClL1heC47YA5980GV3mCL3FxLYbrtUvUi3Veh
2G/kSgDEt2B6dzmS5uuzn1KPuJ0fIdcz1W1PvSd6V6f3zorEt9/BAioQlTntdwaair2/Yjk4/ypG
IKHMqd1htQzVPLH/Pib1slPGarQ0GSc0WcsSSFG2JwyxAyDWCAshiRVOnXU7wc5Jfk3cOLanUTgm
mTJzCi7c0N3Oa75yNr10985dSnCKAozvgSk+zBZd2V7h0LqGofY3vmbxfNF+etWPInMRZNPPTmDE
zPQXWJnT4kiNOrV+CCQikshHX9jswnGASAX+ufs4jzjSh5Sh4MA5s6UWGHfLjUvU6JAAecmnUpTU
/dwWKcdys5ZIn+bZdM1w8YX/KMgzCbLt2ihDbh/CT/SGaVcfpijlP/twj1pyIDazMWsI7GDBFpIJ
/xkFREzkFejDadqA179DiDAiP+lQ1Ryr8C/bRiT6JcN7sFiWESibt4iYe2ounT655eJbPmAbA8So
2G3ZBRsGreExTLxKWvd3RBQMF3wbDCRGE2pgzvcFrd1diY7deDDE9bXvOkHRh1vlHdPD+F1pJycc
tUkAJ28OzuD9/4wIF9yaYU9j4u9w0luygpssZlOSP7tm511rxjILWBmuuWiCctWEs3j9qu+i5GsS
h1nWgP2w6RhbI0SgyN7tbwzb7slFhmzsm8X+CeJAm7/faaUjDJSTzJdyW6Q01hYzeqeXPS/B+4lj
I2C/Moapzo7RUrLKXEM1rzEI/zy/AhV6Dh9nOk2uoNqLt/TtMV9IVnW6J1f0FYfetrltPOyShLPi
652831UA81Q+yQHLn5TI/ZCSJONOvYnURFtYp1VeqiZE13jEBIByLnQPIYbYhaeAC+6kMt7OXW5P
WniCiFQ9ad9b4mt3Mea4LpQDzRtquPs5opLrl9kGXE0ko8oTdmLZun/u8I5RR/Nsj/KQUbVEWd7y
U9D2WpmcO+wLp9wr/Td/+GBzuY63Iw+r2eqmW0X2OSfRf1bSZ0HtLFl9KOozcDOVVFjtISQa1hy2
yBC5ygaJ1hblC9zHaAnNONVr5M4iIzJNOoxj3EHtlmM60Vj3PasAr2M2PPw0fK9uZG/Obq+O30gv
p7D/Mq/hIA+uUuNRlODmYAWeNYLr20p68Rz6q+Znn1wKqscvKj91MhHmafMNGA+sDA3fl36g0eDu
MpaedUJIduBi3bO4pdBfD/niCIdjtQnp1ar4Y6TG65QsAlG9oxx0qdaJLukxiN68EkcrQC/ZbQ9N
PuWtmBMnhMxrGURWXEQPrJEaYzMFgsMMmNXbkgoxCpcnqsfpQsOHtQgieu7FRB3mu1ROKMqRJ4Mo
uJcwEY54ZX1StMwbCZOMVkPpTfqK1q/vIpd3quj/CrDOWIxnZaLvpbH0alo/Bey3CevqicTzuKpD
5Oc9KFHZGdV3wiAKI6vOTrb7/V5BxVbIWBt7UarZGLRQTHB7BXSPTOq64p9FdabyAUTq1vdefKwb
QbdT4gJxCIvCiRJYeegC4qwMIibi3nGd2RODmW9jpzSA3gvG2twdpJV8tnJOE0MJSeCilGX8SAbD
BRaF9zC5NoC+PK7CT9qS2xZ0+35iBqWqg4OQIeeVbeJRhwUGB+bXlLhAY7X8XHCAs+Szejvp1g0F
TIA4awIH6ZxhRTxJtD5N1NAOP0vnAOsYRKsOXsKfNTEUbcIC8UKycedUzjc6eKIKpxdaUmUVtV5t
PnTGMvvUItSy4xWZW+3xxuYT2oGBrMecP23g9xIEVfL+8KDlsRCRHetBWTAVq7klGgkfZ9W4xYEw
OmWcW/WuO6JOzrhCUlu9v6KaP0CrC+aF6SGi0loljpmZDhnrwifc7aeAHTeLmQcftozt2smNbxuC
zVDc4Zqzw6G1OshchFq3jsARDP8eAW96OavAZynEIWgxoYiYzIL02XdOl7XfD/Zoi3hCKPyGMS5Y
XvnSkQOvS5MGpcd6OeebgTBKl+adEVdhuKPALmdn7EdpxymObpV0du3DXh66kxM1wmTgz53lHMwq
s+NuwbS20AmwFAxxBGSyTA5PkVH9BT5rcb/Ot1qg30uqNuYDOJ3UB8tw1vo1EPGcD1QjyiU7tIn0
FJtpg37SgbyaZaDpv4GjdKXrylAQgO82kzquPHUgHoZCg06dCqOg3N8Jghn9azDb521IilHvno1K
j1ozems6IuAzeQUmmkKrXMAPcgU84bVJ0ZnDKeDW79sLeMTRJuiG9dvxF3el4CbtLWNb6JHBvIOx
2NoGEM2GEyz5sHpoNKslmyAYTbbrsdSDKTmdCL56svf3GbJm2lCDFw/2jlWI4Z8pFFiJz6IBnw0q
FlyLlWxk4FWacmWG7l4Nosb8qs2IeVkxaenwlHaDXJ5vmbgOBbK+ZKJ+TmHyczIkDG8MIbrQoDUy
8f2YJebATnp80e7rpdjjBGCTSQ+Xh9dIj+exVPFfIxjEBiUC+C8+O5TMwlYRSEHTRrwD8OL4Ju/E
jXXQzvOxn0x4ij1NV8Z6fkTUZVIJqRxSqi4hv4e+2lBcBvRzWPSLtqe9UelrcCGzYqisVYPrJ5k+
2HP2dksQchSFUIqtdp5hBjxEukmTZhQDlWCiEJv6742oceFXEZAXz+yqLc1ouiQ7l8oX5k+rwVys
iK1ouU5J6v5ajyHPpV79Mf9W1rHQoDn37fTH29CZ3cHHvbqoTm7WrCIA2s5+MFKH7neK7b0y3Dwr
XxgEpJGb/OD6j4TaFhNsvhc4qYGgzoZJoHbGr5Ph42AyGGBP/OGFIOT8YIa4uvG7AO+f1oZxBR7V
VtrL05VV1CFIxc5AgaZMWA+k0TJFTUQw4QfIhfkHWBaNUT20j40uDMjZQVj7pVEgPCdB4A41wmyO
ewRa3gHD38JKUfdfw8KDni8qxWXRqqIZCq+BQkHxXMU0uZM7uE2t78VNRV/JPJk9boxK1lMxbtU9
LlA4hC7R2FJaDPqWl8q2LC7Uq8BLHFQSYMirzbxtFWUeYvlqJCwbseXOZCMqVj6yrP1U2d1QuL5I
h7tgmI8vjQ5thoAX9sGjIR0Z035oAtsw7QFs3tVbKWIzpMPpZeCYjhPua8tgiK4xabPM4H+PLZOY
fRKfdSqoJ6IUfEKPGGcdhF64Scqkz2K/QmAXIhcgOZMuHqFo0n6p0esW2A6ugHpcxBD4nlSq7UMM
jsMOChMmbPxzssdIR+6ml1bepNxFpyKbfKR0n8kqxjM+g36SqHT2R28cKEhQqEIGrWcum1O08cGE
xGAHxyoFYETSBraZ2+NXm8YI4mXBbN//Wq3EVopKGHSismUhQXSBszN+1gjvlLP1uINTNSDgcvUI
yuH3IkGluFZKk0SiCOK9K9d6WHoey4Gtglkzkf3UWaaGDhSatyx7QD39GeJvV6Kjlj3Jm5z0Vt1g
V7giWowhx+wFNiWeFkJ6rnLjYfX+LRKgNmXL+RPLOJDy6SHwqWLvIeLJr5aCnSpu1Jtshq2RkioQ
FRnHjPFbrF9WAnKHum9udAhldj9j02CisGZNiRgEzTwn/5vxty7R3VGCi+qH7xNFkPZ3bGFZE2q7
2ul8CrhsGAQDGPPPd76Mniu7C04WBTyGVFf1kQlkzQ01RfRJB8kygbsoVs2QV9lquf0Gm+ehzhgZ
5i2SkYtDEZo+thyS0L+C9W5+udnVKv0wePv0pYsxGIGs3JbEZUS6/yYDXhArZ+dTOd9oTiwbgWOF
FlA9JbMBiRBie3ZZORlTKmTXvFl4czeTA4Vs3n1kKTgwDHxRRItE4SuzJ5R2U9cyMagmUQmygMcw
/iL9rd/jkhhCddwMCs2szC6eohkNf7h5daFkGAq9N33EfFBlj82riydkgtgFmLO1jMOTzEL+pW/4
ts1sn42UFOYZgjaAWxzdZtmGnL018B+sJHoImetkSvHd3kVow5QCg1/4EGQRbSS8zozAWjr4Pzd7
nVLHdkh82LUSxhkzveQTe3vig+zKleMOcFflg18z2HEg0AGcF0bOKLS1XDGqj99NNI/OfpWX0kc2
6vAKsl51LWL3wrYs8PLgv//uyKMpaOvbUok0/KNgyk8RTDGJgGvHDyVriXhV9LA0W369pco7bcJq
xh8l3Tt0r62bywkki77ZcKJNMIPoII1MSROF+fEIH/Y6iv2siZDhypycZqRFq/8BhbVulk+XjK5D
hen7hqg1+oWd8rw7lwHL1o0GZF3AI6qBLAy1qI4hl34HqZWBFZKCpneAA4bIIIFu3uI1SJ8MRdTQ
PBKWaWV78VDEzXMABuHC2QBo2E4WehlFo97rPyv0oe9yX8lUDUozH5sXqY6otuBNIZoQ99KxowrT
aKtPjOL+aibJOyk1GolO8qZ89Obs92VqzSoLODP8Zb49/hQEI8o7l+FiIZQrnIwvzfWGzwH/qOmm
FpfUPDtK0efrhX81SQZBHbAN1dEEUVpkg3OI2UghHRbsdwJEFqJ3NYQXtQevTzBf+fSMCpk7uzXx
0yRB5OEczQEG+etpJWSfvSgUKlrLAEBRNrj0eKfR0DKp0LF8A13WxranbfrAeduDMANKywKyC4eN
ADGY3UUlb8sSPt8GjWE6ufkmr+wiMkUQfY/kWQypQuxmPsHvivzwfs+OhPgrxLAFIbKiRv63fE55
rQ+B9PcBdh/0y9zjvfYyL+fNDJ0Q7SAuXnBWzlLkIvBCV4E0kpGbrKz0ZEpG4GojQvbKBmPqVGQ1
Jg+j7sw8bfQyDSWnCiYk/vw9LFXs/rgSm27B5vKHobFh+z5oBUcSTxEu89DpmeRQf1NCoOFbVJ/B
dPGnol66TONFhwd0KWGy9FVS2iKV8Cwt3qgM353Xe/eEcZHAA7f6oOgIu6CNGIjlbOeQJDFAl0m3
E+cYqGTTMbUs7oX8iJMrUTXAHOGb77J2xnlMYvQYZ76LukXdiwe9CePzdi9DVfE+Fai6xfWo4mMM
w0aaXgy5hsx0zIgtafO6rTGagzU+9+RwnWMhUgqpJpmqraVG2pqF1Kmxd9IECpjn2OYD6haVlmdB
ZF/7HGCRTWYJvFipRuhJYK9sOSKC9xEHmxcu3NHx0e7BO1H/73d9pWWgPWZKCk+bCfKGoiM6lEoU
Cef9pa41xIccWc19YWRWrPtd0RsZL6Kja1nVkS5OmGpO+Gy81JOPD4yBULB1gW8wBLoWYjra27eA
CXG5IuoBaNlu7Fc4U8NMxseVxU6qdvs/iPXDXpdax1L1EEojL6VHplPr3TFEhlD+MFoSUWKT/9vJ
CHW1wlPdziNesFSn3T+MbrosTiZAkkUEwtXbrIVC/SJExR3yrHJ210QmdeSAqTcwVI3+w4RCn0AB
KYz6ZPP/S1U/AXKzrV7Bj3SNZdR07PVF1RQ+w3yTh0Bfh4jjDv7CpNJJx4/g6k5IH+iBUNbTMOQZ
JBuiYHaW6fK7gBAvFDnBS+8kchx1HArpE2F4s5Q/ZclVYWj72XaYhWBRuL05i8PGIDlAgNIrz7s0
p4lAQJrCy7Dg6mP2JSKStU33m+ghIAo9OiPpmfs35I18dp8boGcr8fAD95kCWFqUdZt5XjBO/m7o
/BcwN9/nXSKbUaqACATSQ75EOyo2q9eBerkg5IqpL4KN5zDPqmTqCIHOgrlJtI0eF04VexwXrZOA
v3SfN8Kv6dfBfNrtrsRoHv+Dz8F6XMynMjUmYaCFnT1peE0IYRetXA1OfLgkO/oLqDcmRATZbfBo
nAzZz9rfqhl3jvfrK1mMaU9Xtp6MguP6haQyAVD3DET0soWw/X1mpoBCU+dm9v5g36VwAWXhTszo
9nMG/Z8KdEvZEFagqEgIIiEAUl94NyAAoLIjyIx55iyDqzcp9FXAiCpWasb0jVpV+8wNX5dkDlpA
ct9rdo4NyE+9GAH8SDO52jFQgl/dMwCSy9ZnByB+mP72qf0IgfP00x2BDVQsLIbkzwQYqf5bAO/Z
G4BZMrt9gH/MqJpxZu0Q6NE4AqM/1S9bIus/m0Q/RHVZDwIPNJwVFZ4ILzvSMdwNKlfcLOGCHJLH
mCS+n57IoswrkkIWAeXA6Iiou2xYeeO0nyqkKzRBNpd/NV/Y/Bl4Ma80BXuV4KiGcevFaIGlxXak
XRNavAVZ/L0gGJKv8lhICdrqsX9voYDBPERWGCRcWaOswH/3Hf6BUsnEP6lWNKuBmwCR99rpiZrF
L6wJjpEEAAv3tFkW4DSzW7NbNQHMedKA3TwJtJ5dIoCU+chQvTMeXQiHhHojMbkdno/KyDXE08Cf
JB33PJYTjwBIyjtRO3Opq+xljXmah7npNQp7/GjSU6/bf6E80s6J21m+juQ0XPV/4PbhemjmNYfm
Ng8gJsIaYY+yIZa6tWh1ysgbDtjNowY1Bh/iGCD1Mm+ro9EdjU5ZD0a4MAiyEBd+rszW3FMJe+UB
sct7NtHavIJ97Sn6Q1B4GkvecFLIS0AUxclgmqFkl+uGi6jotwRYPY20aPKFEOno+xviTbGs3UVD
ajgTdvVgLL2ht7Lp3UjK2aHE0vMHV5JQKF3o/ezd97+/Y9mdTB7tOYEAHC6ZD6Rwh/3tLBmd6p82
i1XiPmD13WmaTAw0w7J4/9k4J1lJfigDnTt7ImNJxez5mR41Ch3WjcjwSL2+ipfbR/byae9tDCJ+
F+11q/zVEeMKrq+jmEjtg5DgRA+wOHkocSt+xOArXVL4/edzuumUPq1aSBqJv2QrZHooi3ZJmRdP
9L/+SYvz5oOxqOV7gcdhKT2zf4xYmB467DpZ7meeCa9Shx643QcDseNpcIpkAYOWFiz0/PQKVwRu
qVb7k6XqojEcXUrPc8h8zwcce08AiXomAgNOyNpY88isJ3vShgsp+0sL8EMosMEg6R5eezZKYoab
xMiObb/U1c7QPBMecFd1MllGokWc2ELqp96LkoZOMLHXepxPu8V5R9YnHilPZZ7hDGJbImxfv9DT
csG7XX2SLyQptj10gvAxmliJrV4ti6B/s21MmahdLNLvReYz+LarHLeY3NHIdeV3U4GKxBZ/koWv
w4+JQIMtYh9E5YyBh08Wy9pHZmctfrEQYk6iLAr5kgM4IMfMnA9OL0DnRE0BNsDX5yii3YhxL9aO
1w7BEUkU6RRNodjHHflcp5WovnLi5Wkm5cfibveR2KXAmaQeDaKJ2w2yfsu/gwMsj0shN16jDNCr
6ip0sTAT48JKjINKUkrK67ICjeLIORTCqtY5rvUyjv4/Ieq3vhyyGYzRm+YPb/zudCR5mD7EKnKi
qYzkgr8viXWeSNAMFi+ipvvsMXtMcJ6ywYv5DBdB62LIlNm0qUnBs1VH8JRPkzSYcHb+2v0zlxHy
2A+AP4lghf7H203g6/r3XK3JL6TqfaEB+sDuALdGOquDscb+nElOLC2QtDJ37DVH8JvtWubvmU3y
FETCl4nvqjtbanrvRguhrzizcwuli+Ipz6+Nh17Ar9epgsjitopkFR0ecdR0fi5eRH6arC2n3CpF
YcPoOZK5aPgT3azy5xovnc9F+kCEg8Wb597vridA/wmHUG0mE1laDpWu4nyWVKdqk6a5hdbxFfnt
K6Lns1wLGktniB2MsbeDJ10pG3RvuN2dMu/QLpbxjznPFZ/zYISHnNbLvM/3rptffabtPgA5siJ3
xA8uN6oe1C4H5HU1OUA5elhqLcr5uAGCLWXMCvxGKysyspcSk9C56QKj0UhwD8wtMxxLnWSGr913
9jeaTEhsM67c6+Iweck00PM269hwXEBlkK3ajsGAS/y0wFoUlz9cU1VlQTEYu8F7SM9q70bxDQdi
2LxA9BSTheccwOC2V9UhUooVEF+WwaVUQU+dBpXhLZKKUkaJLO3rQk2AOf72V2fo5YkM8opI/Vl5
+BPcOIh9trTOQRGPzcyP+p83lKX6uApAoSvrobUdWMlI9hqId023jmqVdYPQgnntQOs4nIapfjSn
GRMay3l4JJGWSwDImt2TW6UFDL+XaeHq9zWguoQhSxxHti8ATnWVxnqXkgbuHjrtKw6QDEvBo3E5
/wYUe24nNgiGbg+tlPS40bXwNJwVRpKFnrXrtUJhwlkW58xMlZHJS1Ra4RHX8Ms0f9zDn9tWBlv5
cBbjHFia7BEZXfqU40Gakhah3AiFz12xAFeKC98Q4IRoaErgJTzaP13OVYU1fjpah8CaW+lNCcX0
037vGty8TBcqb5NSZMwolA0W5auHPwhO85VUnQclaeQApGNWP+h8lxJpsEwElwyaReW3VuPkyMwD
7YmykK7sv9pE8NUKkg8mLJqIX4VQ5vdfUzDIfGrnJuNrv6eHxY7rdFCgOR4luwLEzOA2gcMkGCNS
jLX2Qun3rdoC1Rb6a/0XHrPAtPSp0nQ9Jr0lyN7HrldMhnKntyVLGq0p6qCbeKPbpP8y2LME6yL4
OBjfA3ap7oW4H3sESl1xmKmoFL3EzUGPJrZbfhQehtlUggqzCw+yhF5Wo7e2EuJdNQ0nJNgsScpO
r4Z+/+Wx3nChlblyZd4HZD6thK8JbQN0mbKmIGYjYup5ElJTjiSQQ5hNycgvTu27NHHpmJTt0Gid
zu8NuUyRc2PJxAknet7JnMwqHyXoo7mwXsAqu+Sh48T2FxsuYxCm/NIB1CrOkrEZGoEkDjz2Pukf
vl6S2nKJEckM5Y5786SjMVk/GGQy8TXbf/EPjlJgJxJU2l4xnrpZoq/AnjlGWnk0XyH5nV6LZrRN
gMrmvHYD/H2o5xHanAn93odBc4CFSX+a7ADAVrTwOd5UhIqVgbdNnV2fnuuokI7Dhxa4oM1SOIMd
tZIOioJrcEnj597fAAaEDvWN7B8OfF0UPXXOy01RZJiPBEboBVdhLzdEVpuasgcbXTImZtEFjhHv
/DUOWp1TlJjaUgyGi38IBRl8Qx2ug9OzbLZsralhnPNeqjPPcB+AIN7EqIeQgcbxtTShRpUmMsj4
LREnAKJjSJ2s+txat9PHwMSWBLocSOEGFQ0+RIYI7MgMMcC80iTFx/I6ECGpYpbjdRxcrQDVh7dN
DldSAupkIus5z8iobs68aldFgrFsynPRkleD9EWlJQqFNTawYq/lrEgQ9jqOgNe3Q91KJebCd8sj
ePfYC4ZESM9D7e7eXUQVzi9TBjNXRJ856h4R35nEHJVMOs/Qu6EO0uqkaTIAa5mQf4Ri5e7Sqpp7
I5RCh6WnzhwjRdmHUAflU5npjRJ9NW/1B7K3qmvGNHhtgYJNILwXLg7aD1+4MqslZsqfpUNrry7I
028SHDD2qCWNBABy7Z1HHuGyiFpMeRL3354W3L1A5P8AJcyrxBxlQIIXy+ODAOEtXZ36vKvfeDhK
dWq0cmP3NvhGUPNwb6QWlAt6xc37UfACTRqe0aUC3j8tUGVfJpo4gj+jUevs263v3B+trj8EbmDF
cNLRmn06hr4MQhn06s9iqC8mCOQ/eXqUF53/UpBFFe8zQqLLgaZkBIUfcmGqmap3ldI6vlnM9UOv
LtNr6y0rmmZYJl0U5TR3NWYfEhrmBoQCVgo8QuL4ufvtRzQ2vSnIwaguk5Edri7cbGgGWOKto1VM
K0w8KQJQ8DEYbhGi8WVhiLN0urV7CsqUC9tG+lac0o1PJJgiQLlOVpRYKwH5qwvm9MTcDLU+Devj
fK+SM2o/qZ6D/HCTCNBV5/QtPcCZ4Dc56rKBjWNPmU+Uf4S7+V40Y6lbXSSf530i8FHMHnOo9WcO
gKjrRVTBn0j63s57rGyyJulgwnN+BE/qPayavnwsgLYMxjKg6LyHJ2p0eqAtQOo+GhnxxaX78Z2v
JbhqLv6J/yY4m9ski5guu7A3G2vQh5r4PH2j7ptdJLRlD0J7Ahcfs/PpcUsFRwneY3OhWEKwZPuT
M8oxq1/5xV7HQn+WeyDfYSV0Q2op3ggR2//RN5hqekjz2lSE0jKqcuwhpwZsJcI22lB+7J+t2JBu
IbGDdxPXEJxbbMpfhWH79WBUZ8wwhW0TDHCuktqIrBqUQVuVOU08NUAAVZZR4jbx0DCI/9Vl9buv
vBlDksluB9NVrOh9jQnSZjbmYHR9W2r3dEM9VXew9K8X9RtHLx0QBR4njnhcAfNE+wFY/kk2jjem
jVOxja/5eUVCQzt+x4hJqxnQMuDLb9JQXwrh8GUqdlSbvXWM4pmNciepzItI3tAXPqgLOjEZ8pHS
rNJkCOiz08Pzj7pviYX0TGbhkr0nbVEVRahbjPmJ/+joQOueLRrr0qQqybI1N9BL3gGYnBkV+Aa8
OdMwNefHebUl2zMg44DG6JGAICq+9CvLoRsKuMcoo/fk2CAyyEQ4EWZ68EfJ41n7/T42X/XVw2/R
WqL3iR1v+9YFofxH3dN0kV88HICRwQxzuNJBmXFLcMuHkiBCe3tPAw3XROnB1hVUywsJTUPAj++c
cdKDbn1S5ytH11U1ghrkslKa5z3ln/DIUxncZYPE6WguM4KUlcsQBQrRbVF95XeYo/YAz+KLQM3Q
4a0UmD4WqpGQzsAgZaQg28ISfuVRLs/bfvteakiYrIXOwB1tjFE2M76tLlo5CF1bMMTTrpTyNgw4
jNL4ddnj5YHgootsi3EXUcKi7ZQYtdSl4qH/WzGOfrWAlKq7+EIj4fMqgH5xbfUVz63ezS8Rd7R6
RHqffRliP6Wmq7aFwV0wqiT04bHjU5B9lkjRtgQ4JzdVLwH2EZaCynf+wMixT//2Z6Tl3P1QE8OX
Cr/P3SUhwCMszYQuZxt6x6MX+FY1Nn2Z5naZBmTi0Ys+pZAQ7CC13sED6JpJn1M4i96tjiNAw3SC
JIiP7vnrHUY5Znx5MIxuz5vHABNq2UC8LTRYDcIdtqX0Gg/BpwPiJlWlRbtHgyJXe+2vpdYyelru
6/ITqbBxo1Nk4Ezt6FxTTbrEKXZOuQXW0fJPRScy18cPr6PkPZIOpB/h4eUl0LYSewgOUf7pszNb
Hu0xsI/HOdf4cEIlnrLnnt+v8obAKnV8h6xYVQud0eLqVcE6/sZjSS61fZTVgHRJmY38Ib5l+FMp
kegl5I8ZH7aRXGac8vuyaScof/CDFi2z0tAuEcr6tSrWX+32Tao533kvSAH7hCIXXcEeBrrwaaPm
e8TnWbd0bOeAHV4lJUN6CtD+AhTqOe6biYMpoBo0/PQaFDl4NSsy00DR3OwGkdv+J5vlFVJzmQcc
OVgypc2AylDDgNgT2O/lMOeDn50029gO4xzXO+5sGM2kCmxb8+JiNzHx3o30ar6wlzD5Tbqe9OM4
y6zeWusD4F3phGbgP88JnOHSeBv68IfZ5AK2O8bUoDoyfz0l3tMEC82lWnqJhpJ6aC+m6DS97WjW
/5JQ+ulHC+cb69Vr/SE2miy12IsCSdXYRhR9r8Q31lyhL3HioTBZDcQgZe7a+C2WYOGTmiZUf9xQ
e30C+MtV+GRnw5wjbmFFYGzzJhSLSxi5RbzUU7WkQTcgfUu2d3UC2dqF7Vy5xaS+sEGkW9JEqeHZ
kXO3SSFM71Pdj7GglG86ylZvEv4kFFQvxWVsYeM8bpxs1CpZRIsHMXv5FSAdedYSwtK9fZkCNcmS
Gc9boNFe80+6loiA7LGb1/aJKnqxJoGVOJlhs//hsWu2skZcf+wS+BjQyaTfIbo10AMh64yb9PVF
e/3Dm4bm2pGXrB1zxycF4KQxs+ohB0QYj7b+Vz4tI5A6x5q79BvZqT4R5p81x0ip4mNfLSSWFnkE
LqcNQmtVCXrrhgqqzH11FHjTeA1+d8cHJejWDrf9QC+ZhYnWNCOK8KiLgMicvPbCsTiL73nI3c5P
YipPVRz2TzTWKpixxWl5zQez5/1JsIbXqcDC7iyk7XFXkFHhYhMZh+abrAeRPfYIMWBySU0OH/HF
o8a40GqpSMvSuF13YXp+KExsYTaiQHV23u+krZU5faL/ZSaAzVGcRJPvHD0zod3PUtk4MQDEMNwI
Ct8nqsp+sBugvz6YIn9yYFraoypODyAI15wQvP0J3txAvTIguamrhX52t3hIACG3q6ESyaN5zxaE
SZtucZG+zcIwtuaCDkpi+qJ5MijvpP+X4YxJSGuymUr0rrMKOmoM6xYHhfzabRAYCjaV3LyLJ0Ag
R/ogf/PJ8eUnyYPfHivsNr5e0/NApyCWhbAhnz55g+cl9kNwQ4Hmv0hywglXOAdgXBXYa4e3eE7y
FZ2J8oA1MZcJ0eYpBSihQ6p1auGef8NrfWzp/zzJMTDV91sRvODWeTjd4GuZC4U6FT6MfVnLes8b
8d1kPW6d6GJh+40M8dH5BufrCUt9u2LhITzefOOmLWSjKhyeczCk8+wxRG0Zf7TUWjK7U/aFKHWA
sxsGPAV5N020L/X6vmV1hCWlEhmukGUPuuqti+nK4l89BuU7sT7MGkNZtjGUcyd12pS42Iu7DYlC
RMfwG9exroyXQQiixp2Bx1fGhsXUWOumhr/euK+8R6ZhFTyrw49fjYCM+pI1KaPJCFQnRnL8iy8d
T4DIzum0xWyyrld0rjppGm7OlHXG/hkYirlgDtRSX1257SR06yqbfb1tokAi7JSP6zOPWY3I4K+V
XtyL13lwLYzBSlIAntu6/LIRYWtwA0hZn/ZwRgCj3WFSJ0ESfMf66O0b83yzN2ip15xhpZmWS4Uq
xq7btS73kcO8W66x+QTzPng7zRNyhVynznq8+MrmlGvdkZdB6E2eoL1wUfc1lAf2QiuAZfrCOeE8
ByovncmSVrPYm9wjf+JKgCo+sugQ5iq242CdHLgUYbA8OTd8cmPnNku/5Mqa03vJSAfUAI7yf8R1
ZhPqSWHPww0KjIFCJ4QoZ+q7CDc4vthVvY01KfGfTvGHyAr4H+wDbEDq7wf6AtXKPz+eJzdoGPyQ
5P4cVsBWsX0nivsGXN3NDKsGk0Z/t9MA0zSECb2+R0LkT1+6+mS+1VRplTn0MLjqml/4EO7Ytx1Q
rhdBrgrIR26RfTJKTbAYOmvXD5DtsX0kaJ2zG8nFgUu0AcOk7FvDl/pkF7550CrwxMDJTCtNDTNf
Et1MF00vu+hb/v9Q5BhZYtc9j1grqpNJzF/kfHc57Afmz3qJh8enV5J1gZGKHY/kKaJXDCjvzIoZ
7hop3lUrpTrDbD1FEutMe5JhixQx3L6vfTxSu5yaJhCxGzknGNNhduzAUEhjFcsRBIMWKStascHQ
i6GgRf3eImg0IckiTeuouP6nXbvsrEPclWLZ1jh2vbY2IctowFkuXlKZdLgo7BAhUNRGVWizZqFD
4p0i8JhU4Y+s0/qu3Xk6stRmKDBpFAaUIPie3AGokMxj0uzRljPMQ/zp6pvQwVHML65oXEInRNNf
DKVXffp3JLNL/Dwj6LI8IiFSGFwkfINuvAH+dxIu2iqAXyzkL4rLnja56saii93x2eKM0oIqf8cl
iZR1/bSZvRcjh3au6oLpr9DrAS7Gx12A67o6Qf4tHAwl5I2fatBYdZ0oHtyc3C8eVZYpejfHn++z
81BXAZ9kA/t8ua/fne38jDZ+Ow9ympYaoM4CU+iK8Lrac/G7b5qb8qJmvWKo63nlQUqEj6ytSiq/
VHqP/1bcF5ziMPzElyxd8LnL6n+LOgT3p8nP1Me9EDjQnZi4Kdh1lLytwPQ7DFCjxQVmLmixKGt5
euyTECUNQd6xAMHv7l6+wu4ghxbe1wFe3/C67IVwGPk8nqrTRXxlCB5BXYabWjz1Qaxfxv2naJES
fAaTxAmPAgV9xYW5zJs0GdCUmZHqHBvHNc75J/Sj5n1ioYcYI0CC1OngPphzcKk1lGxPjlP2y3FG
oWoAmX8wvstaRgDRthNHAJ8GmFtruYQOgy9F7JM6jEtu40dOfP2hu8UTfhouZ+C2NraLBs4cScbe
3C8GLfNfqNxOAMg6zOzfGSeTtP6dG/h+an9kkVcBD1BZuCqxLQfRA+I0K1aF8w7Ehv2a7nI/8l+E
nZCOJmvrmgLH0OTOHXlYUZGVptbXk9yBu0XbJdg1XcHSGBqOPDkpmYdaZp5Qt0tLNhUxTCKSYPlX
Z7qArjC2EathzrYMI/CHuBD4CnmqDovMeQutvPNbEGwlWtOqACVdMGrm9RjdOIPU/potyaBMXLl3
8l2g36AmZeDGZ5mrZDPPtyPr2lc0OsRnKOHrIpKLW1wJG3oIEnr9J/1rhkIaRP2kmaBH+87OfD2p
XfLWzuCYSJnxmDJhTvivyagTN+jsbM3ZqWYdi6aFYw0gDiFeetZVF5jzWs4FxHrsghJyoLvhtE+o
UafSOMRx2CA4gGr7dDaHdECPn7vzmEmM/W9e5iYqSq2L2vwtaKpexFu/023twzEoOlnkxAn0yBD6
QzluFk8mXva+8feB+VJ3zpbqH8ZUZzaEP0LbqEVUVDFisvzaHs68Kcczqy2k7kIbvNxXawzEMGPZ
Q8AzEjlZLM20P6m+o1dA+YxFarxJGTvRsfr+uP+Gqa7NRh95h5URD8vxbZWTxDNO7Lhh8pdWMb49
ENsc6jnvBqa4m9X82Z3SuuRkwcfkFIhZeXJxdxpq+4iA17Xmx1dMJ8BjrGkQZv9oUMHGLGbRg0tT
vrq13isFJWWEOH//nSp78mzbCxY1+hzGzPrj3IGiCLc8yL9VC4wUWl1owWtPYqzhMuriNQLmfdkq
5/GskXox2fDO1WnvGR0El6EDeht3J6B1xcqxl7JXqNRtGGvJ0VBvDWRVqkuBvA6rb0NqoVdWNb5i
v9XKq8A91CeyhRA8vaQgsNXCaiE9slQFFzcvh8M7i4UF6qQsK2lcGh+/lN6EwM/ZnkN0T47usd2O
cLvZePcxs685l5IrvHiRWc5GoIBa0xdp7CkB7tuu+E9mylhucngSOOtQp4amJCewmFE3Ud2dglc2
WlriBKUtlag+d9FUiwmV64a5LqY/X0Dc/3HyR3JnQpny23q7YFxZN5qTLAzkc7KuFvOTgH8SSLDR
zA7A9h+Z2T+16AUkAifSKVXhAfzowz+UpGv0TnlmDxpmXAFZ+nj1KTu9Ypdf2vgA/QoBRfjOrctK
UUK0O1S9HhWp5vz1orHM6AOEytAbackxf7c4y/MfqdB46LIDeohn67VpKP8IQE8RWrgy+1WcIkVW
2Za6zF+31XXgng1lUAgYxrIhx2M3yE10KzyT5kNUrkzTtSdCf4X20MGzrWRjQZxJ+olTh8PQkwbN
TJqan9xeziLz3is0FKVoyunYoyL60hFOlZKfjebVtAIfHp4SCZzHOYxYl9k5W6yZOIaxuVtyxw8k
efk4Bo1HVtcIP2zNf/jlIqFC5rl3FtY00M5Wci57eFbrZaAXUpLk+OJ4ke15aZbDZJnFmkGGoKbG
nOzv5zgrOmIwLr82JGTGf9tFPg2wSaR1a8MKfsSJ9kU9kcGgAB7fwImZh0mvXJoCruou9dDS5+yk
pw0R0iGyyu/SnC0rYTzw01S23sSeOLl7A0DiiflCt8hsmy7KdsRvplVjaOOnpCuMn1105ouK/XhT
7KR0G6PohN6YtoAI3sLV/Dz5iD5ldbW3CodETTP5/ELRMYspf7o1ZnoHOBs4pBLeB69RNpSUZ2du
IJZGB3/1MDT3fwKPeRYueulu8E4NZgjbnaatJVjwTbVLgXOz/mmi5dl96tzofhynWYK5kDUKl2q6
+XSQlg9cOsC5BvLxLL/BCXlyn6aqsDkAuA1sUegl/w8sWjJAO/n+5IP8MjrlppDbNzjc1iquHX5D
nNxfgy4I58ylP4fHp0prQEyORppGObViAIQw7w34rcTBU6DFSJfSCV09UWqfaGKtu3JLm4Ny9CTg
DWcLr18J8l705GcrtWGkyAFW39R1uRI8a7KaO9tLBaQ1D1Wk2sNJ1FvTwVRU0ApmztggNIMdStz/
oPs7WeBZq6416nCRCvS/rBC8QAqUkE9NhNafcKoABWL7TviKlWXpRRpwSqd0AV13EwKapzh91GJG
mgzs3Mi1H2CY/kn++eXlJ05QRI6V93w8SsGctqxa00k3QaM8EFIoKM501E/hsUhQLq1eEd+TcWOz
ScHkLB3wrhVkmYGhoTVCsHH4gGOeTfIWbYzQD3K10nz8LVnmY1CxTpFV9Or9R8rdaLoI1clBs5eA
7UK9LEc1nD0f/7zqeK7860fXBLmE32AOHDXeCA/srfIwfU3eOJoSF62z5fVPwx1HtQ0w8QK0DcdB
hsvIpTH/IcFJp44FPtQz8YRT2x0vw0Nz/ymqqIfoHjtzmfOipdC35EZ3GJF1B4/BnePD5i/qiDsm
vWdVStAcjGNifBKtAOuoQ8rthbNI8XzRyhQFCfXNNLzsP9yAj3/THiuazc5SVssD3M6ApCf//4WG
o8Wf3yGVkZr9A34GOlCAeltRneclC09br2xaeP94VQnEfwRAu9zGBBOz8WF/Zs2HZxQT8nWjeESA
04F5i5tfWNS0iQx4D8IHxG+FG0asLJhAgRRug6SXopbv9YSeZIt+ceUMI2Zc+EsvivPBFG1Oya2l
cqF7rBj6R/4dDSGXRUvaZjNRmfw1DjM4UjFtJYaB7iA1BR41clRcYy0uNd8XEPkXgzTGbQ1qvfGW
XKhQ92EtYC1ewd5y38GjciMgkSCSwxoDB9KnkiIpecorNAP65xSVuDC/iLJGaaB4Ms+N4jiZQ+dC
GPruPGCgRShPJrx4chYM4gjspE1emqRujqlscX3Vk84w3oePpe2/JsG9Z4GGj8dgVDIu47W7A3k3
8/xor+fA29ukDdtWCkzfbZkSzDCIF8jlXiDm/DiLysU9XRro1sIbyf50qm/UgR+4w6bRAxEXNsAq
HWmVMVTziM6vS4p1Ikcl52NQLhgAiB2UP1reAbTD+y3xQEHML0OeIxLnLkoRaOCIbv6jpbauCDOL
erJCFOsk69S8lElpWDRFgWG4R40nhuKQUMciZApBKB/9FUn2yQF8/PpsznlTkXRGi3pVKMJemKRH
SlYBS8BuvSiPMp9V9CnbYqg3EPk7RMk97h2X2/Ng9m0iLpR1q9iQpFGY7w/GevTEK5aQuehFcN7T
1HOnqJuqqG43o3Lb9k3gUTcz8ezjqpKkbUPVzhe0wiFq6gii9XDsURu0dFu/GHRB8s2uqseaPfb1
OuE0CWPoDhLg4fCXlw6/4GVxMnyhOItELf4/qj6x4SMIjN7rM1Hbt8Zf7zcdZMJZai8k9qXrkjEC
sWfU4NGp+3uWf0MCIeZEY/sINvNq/lo2YKvbT9x9LyxLh2XXBdaM1maUr8cF8kqBqS3mNK6HPArX
Gc4EqzxwELxOd+CiYTh2+Yh8w1V3l73lbsfpkQRN86wHxkOt4m0dl+7dDfvLpIM4SIo+AiVV5kNc
S9Bxht+0FM+uCwmYnXX0sfRu8bDmO9qd90qbKd13MkkzU6we8NDLDW4OIEryWESeYFf3f8R6XNYd
Rn4nkPwD9CMfyQuMJrhg0VwwOxO4pxbLdlW1hrwX+QOgzFSVD4DU4sNtt+QszmLMK/r0KuKLY/Am
UG8jpZVroHSWBkqwbUFoyiYFiYHnZs/ElA5BAtUgrZ+fCqhSsuDnpBCHIJbpawcASI3YkY04reMl
ja1CIncpZrBZpZTOcvtjBPeX1fovznNU+HoucfIE/5ugyXEMhUUytAyPk2eF3kypqcyIu3folSHa
jJq1pCMJvBGkbYubzEPyQ7ej6GIVqAm9JUFLrXiY+nCWedZWTT51ERU11fbTIVdWZdrhSC0WzvCH
yJw9KkTTP1i4pM2O/aMgKgAcSBoUUi3HjsG/+5gsGw7XyP+kCRNasLCIVofA6Dyj+FEahFsoXrC9
gRIA6RyDwiHIaqEJN1SqtNHTdyLLGoAXKnf38gT1HT4XmmQHuh+E0g/XtX+ybPkh0IQnPRB9eNQs
/0E47dVoKKiDtecGTaR4nrG8wAWS2wUsPxZENGiw6v+2/LrVaQNw1YtQrite8RrSWGWGuabpUACk
APIjRovpK2DHnzhXXqLHA9GaBkp2j+ETZXwRDaM6/8kAyVwWjQvTIK9ght+lNprdmAGIPp7ZApEX
lqK11bpbjdxbLgLVjg8Xc1VAbahp+hg+NgnDmMwj5Z+L7SYo/D8R3DOd1PjGcX5MNdedVccpgwCE
NSc2nnnDEmLkcZI5h01RAejDVsrQe6xQUXBv2W3mjJEkIQefXKcbIKP+nzqnPsL11XAc7l9LO+VF
nJvWnaattchN9T/nW7NAwg93JKx8Whm/FgvdfFX/Pc9iQmuRZWBtohZzF6TLm0i94XuGDycOwzrn
SsXPX6Nn34gO8e/it6xrieQnhr7MIb2meKKx7YjWtlp1JOReRRzLJPIFrXP60Xkf2iEKuMfjBQzo
7mVzzlyebiU6RS1PcA1PgVPpjXQvwEWwslM5q31bgtAGMBmv1SVYcs9YaOgUlNznORbEJewHvyWL
qRCsS2Yoj6ygYGUJT07u0stj4t4ctl7c1BagETP2/MBzSRM6AB1jSn2XAqZyXmvp/qtDVwbY1baM
AIT6C6iQ7pJNN2zVEXD9qbvAFdIqd6RC853hTnmQl/00s53oM+fjsJceNwLQs+C0j00+SZPhzSZA
wfajqbXTukmMwbvj6sFHQ2xRr/2Q+8cnItaD7HbzaRJE8XgJcKUI99p0DxF/pkJ0xP1RMQc8oJ1a
7xkq2Ji3UdVwpFhtb5p0TrHSjpq2sD3oYbq7kV9NCzAuIBJLjXwvxJYVuUFzUNg9gXcbq9zRq7XG
0lOpJEqxFB/SlE1nWSMIaC1DyZU/wVKtmUdREDPKRMsRNmsbZWJkmydW4Ho1oLMCrIveyHx12ir4
ir0tTvMitYjLLokwVw1a7C4yIgoNX3lvSnZyNOwahIT3Z+brSrTRC0tUpJnKHX3y57iZhaPntPOi
ykg1m/OY/9C3KFNuKc3S0olux04vjZ/OPh12Oj9bfms6kKx+VHrNJjJdAFArYtfnwCBSP9vPY1b7
5X1VX73bTEZWRZNWbqU1qoWodIY0gGkma34jQ5ouGMCtV7XS9M2J9caNz4CDfjCDH2cAI4cN6sec
cV74HWRTwJiyTCB/6dcVdroLqwIhWrYRmpOZsivH/MQxf8QCXzDYNg0xdpAIBd6aKrnraBK4egpT
nfoLIi/NOrpWWK27Qx/tqPIrGDfzp2pin2X72I+mOhimfDjcWL5leNeqyna/cM5FdyHDvPWkV2//
eU7RX1UhLXIPp+fieaGWWBPy7GoSbf59CkHQ2f/fIofwlLktkDGOXMOzShJa3JBy9SVbi8APoYAG
dW0Q2q5tLa9R6fqNv75UiTFWignewkGYdCc19RMC73TlOyQLLGPHAede9bixDogGfh6+CPXqFGxc
WAelmVF/BE/9S1c9X2nC2p1b9pRQSLBAQMWe8VDcMDa4x2fW8oqPw9QKq7hhshrQeaqluX0o2mJx
jMl4aPJbyaLDqgjL+hDIuQwM8nx9n6OGjeqmYVger7BKa3dpnlE7ZjGjAimrLGzsHZcEBO47FMd3
AlctTbguvYd1YczYdm654+zHML3aGD1QJ3CKlj6C6cxpobwQHJmhVzc2sDabZK0UMs55p4YZlL3J
5iC7X+FwWzYSTwaHH2nmGcIjJptpd0jvVvch9kina3fwdbqhbdqsgFTLKFzbNxGnxaMFsS8lfsP9
IFaVhYgTL9vvyKIsc5kb7Azc5TWmfmgU/X2n2FLdbKE4yi2wQhImKK4HWdF0wiJwAVSeVKFarR6d
i7Lq+77eM/D5cr0f5WSFmmof5j3p+GhWF0LUhwHLRoSlHRJQmLFc2xo8crhIFNhpeLLTZXj0BqJK
ewRJaV2M/qZ9HFrM4I3M2rwJLdo182/TI+x4oQC+UsFD0Gkoo2Wa/90Od+JslEpjp6f+GXAEFSLp
YVU5Wv6ZCqI+MxpMZjTI/quBGp2rgsdwjDxgf2v10p3KOHw+q6MASyyJYECwiwmHY9wqQXQ0xESr
2hiUoZHNLmj50cOy/ZHLI9iHjVSuUfjN3JeLopKt85UM5GbvL97b4UxgZ6bCYNA0y+gBVtMlFcCX
xXKTEiSTsP6z8bOGkJX+5/ThO176TR7yxuvb7ZRooc9Rf2IVxipLAxXP5cYMLQJtthNic+gm6vvd
WxICXxqy2dOMdjL1mcLX1Jc2Smvsr5+56kAB+DC/nrNuHwthjv77ALriv8o/drz+rpaDZtobGO1p
7glcyPb7YGEJnb3wF7r+sFtxFFwi/CMx0ECG6GPwv1MTWI3+fw8jwEeuUXEDfkMPV+YhL3rksDhd
kVkUYJ09RJT+Pq94aBu0WZCwx/NWg0sO1IcirbdPeTfHA1tcHyGzWD8PQKZkjR2WP3IjCABF89jD
21owHTw59k3PKpNrkMunOLTPTPVrL31BnJFIZVEtKBMyi4yaaf1ajzo+Yunc8e0EC+kniLAMlEjD
bEZA/Bi3lLS59vouNfBevfCh4sYCmDrDh7LiqPjHzxmFnS56QF/uJkKuWB0qqMZvOeqE4IzDUDnj
zPe+o6eDKkIsGVjpL5IzoD5ZxT3RWnv4pTCDMF2ms/FXcd0TbIHZaUtzBFnyxSHQpsbsVQxrRK4y
+oJHVVIFyovNrmLyflbUuYPZmR+/b+bmQKDYnqGA/zFgL2492s9xwPQYnxTUBvKdv6uB6eARAQ7u
OfaPpTX6KcpTrMImBcISxOQn4FPoLdUY3U7+noi97a22mylqNFdwSM6/HUYoBM+S+9gcZy7uFs9b
kciccxZJLznFPM4TikG7GjgOxFkyVExJ3J0TWdtCwlcxKVZ8WGRAImJNOLiAAv9JYmK9S6L2x/We
64ng8ePfr8DcPFmPCDWF2PRn++iI3kg10FiRtonJsq/K0IDUtHnjxItY1cuUN6EdHNQn4+EHdtTN
nFwykUTV6vaEhBsfzy2MvHgpXBdVgH5J6W3EjKlPi9BI8r8C9PM/NLPJvERT3a/g4vcKXN3/o7+A
8RnW77jpQr8IQ/uU0ZhA7ghX6+U1wtaf+xgyjapONZLDvnhQY0cMIb1aiT39FM48Ath2KLdbVYmo
AYLgNvTAwuMnlY8niFEUXQrq027zI3UxmIGKDlKL6gfbAXVAxtIe/AaqqLIzVtBPHunaSZNjzht4
dHN0W5vrnedWg38KoYY1+ExpX9kVYi/smphnqhpNxE5+dl/gkm5VNjRl7iY7KN606VofTLFqMVCO
GwTBYafB0j0reiXwIOza4bpW/YPxLk/6FUfuPicJpYfhMXx/RSo/vLp8J5KULmIctnD3ZTxCuiew
kug06XGaixoZOSsWyzOlN2Lr98COd+kuonF1pzMdPoktJmpuhQgLQxTtfbDh2jXrP7Pg0QkAxlWH
x9jcgHl3L9qVewDHiiluW3L4bM5lbhpimD7XbZPJ38pv+eB0BixB/Pvez8jaDpSeaeiQ51XzYt7h
BK7yZCVZKs6hpwuPOQX3lDioYj+//eyIc9TTNhLHqZFji7GUiJw74dfEnscZhmn44WUiwTTPAyFh
sCuZt6sefiocn+HDDnYs4IE1QT0QZ2e6Ptb0wLLzHSpmpX9ew39SNp4W535BEaAeSR0YDDmlJV1Y
R/2tfxDi/dXMwfoE6LwLOSlHuUtuZwaOBAsY8NhWviwFcoIpU5jeelG/dn4Fv+DZjmCQAoTEGkvj
vcD8QU3N08eyECoLeqe9I42NOiMdMNV3EjJGdtdvncr69zdMtwEL2eRYz4A7vHRjaoxS9cv8zfBS
IGXFzFxK9rG+IWVK4nZGtYOmWN8W4mFwOh7l/V92ed4CQaucSoAZyTVDmNWH5+re3vvczi0B1mdX
o2L46yY9n6zHTs0erd/1EIHfKzNqD62SCPPF79/Znopy191EdyEp7n8QD3r0Lf6ogr4cR4/DbDlC
EAmPWS4mNAIQ1qPD/JjLxLdsH90TMJg4xIfTCdGKw0cFh7GUJBLJrmya99HurdggxsNJH7fRu+wp
9NrLoI9sFV3dkJpTfJXs5c0xM974I4vcuNdT7OtJoxoz9XK2DUWgotqBdM/mPZqV/8/mgG3C5KSl
0yC+sI9NTLYppLwDCdDRWo3MpwWhW7cashTnOqklUtdDZdkWIH62ocLdUgAuu2oRcUuzxnludF8C
jUVjtQGt8yzDtbw6UnXNxlYui9cjGCQ68BI4CytapnFsL/aD5kfLmWJMLvXsWEi5i1WbbUD4BFnO
EDdjBQuCtEM1NhWbIj/sTjYrg+sRX2JlcO3GESdawD7wZX2hgrZR477oMBjQUue5jvebroeO87mT
6e1S6ZFy57e9O7BvJS0SZ/NaXytiOe0GHhBZUkc14rHLFQD+APmvcP00Qvm9wtNiHOJQ2Y7BKa/t
mwsYtgZxcUBWv6/Pn+Sl3pGnUXA0NaqqpUw2cfxya7x8o0gQvSiRpH+8BZ/z8BaOSlmhJ+Wq4b0I
haUhDyHb2UsNv4z8PiTA2loPnyiwSY3QrdoMQFmbW1lzXtKDbi6a5oBAUgkMbOH6Ijca1oR2DnzF
xaYfk+xLeMGO833B3fWQP8vQO6boFOg3Mn9XqZRRJlLLbxynnmcEzvu9iHWRbsR8XurIJn/srZVy
zfqZJJ4jjvx5C9Tv+ik/Xl63W+u44v5kwXsWCv5DbyzgsLgNE4h6CkDRAVSWkLiA6Kcejkm9f/QS
vy25BxdGjZDfAlBATb4UK14lMt41i6946IrP12Qt89doWGjAzpKmd5fss0XK27yJNXZVowR9yoLe
I8xwzNxyCUWcMadMcbPUvNdrZfj9LBAyPo7yiN7eKFoqkak1GnklRUSCyeCo0uFaKoo7pHI7J43L
Fkz2yyYlYOxtjitlSUqBSuRppfSbIgopFv+PdayRCgFK3hn8SkBckL7MDg8eXVjXsBZfcsMePhCv
3Je7OY9BjJtrQdEUwrV6ZuR3sBWcqgleBziTB8lwNIfDYKNg3F7c241KFEm1ZmFvxoUw150GP/Ew
UzLWeDHQHXa2UHSey26VuadrNE0qO86gX/iS9X+8XUH/2wbN9UW5f6mXsxe/giMDljCKgVSEVlJP
KuAjdo5Tl/5vDLYTCHFZXwGztUtp66QP5wl1IXQMivlTatuiXHzKRKuemiiZdCirfJfV65ChxQ4q
iuD6o0pWvUGNj+KNZPVpR1O4s3rFOg0KkOB83ct6Sz1x9ZBR6f0/YnOfnfzMHvdxrsS8wia2QfoW
8SMeAk1MUtL0N+STW+fCf3+MQ7r6VXMZecOSPFDwl/KYNNrnqTjCqetqMbl84IqU3fvxoWjfHIxh
F3QLuZMEEjeJzfaZp1yF9+vusHGHp2O3xIf1abrTVUSBKXwtytA4mCIgyuJNBoTwfbfVF9SRSlQg
DBBPDOUDLncJZRJlIHSZ08SDZQJOnjeB7y/19x6W/iYcjKKApeTqaGxWK7HHwM7FBCaBYw4LBCv1
Z/9rjMb0zZMHeF5pn/uCpUuy4oiF944BvsF0oV+gLptkPbifte/DgyPdreZFmD4o5ZIiaxeVteD8
jT4pH3u57Zjxt4dORFwEm1cAcT5DQ5SVQfMu/wiepLkeb28Wp4vvOpjnYT5stEK1uzjNHhGoEa8u
9JEhgVVWIHtWDSCJxH1lw4whXZBCq9yF6kb+N17UQr8LkZ7AF3VlzEaiuTdgMTzADx+utYJ3YH4n
Poj9ej+z9eKkSPSCu7W3/JbzUZEKhAHYlgqsEB1J/Vb2JjoenT26QdGPBHiYUorGpFXjBdfXhS1h
jfOqpJrpRddVLjLcZupJHSi1Mqsmvvz/Pu6znyoMVILWSg0KNKTsh7yz8r7VYmLuXFIKeEvc+fTn
MV7guDqBEBs1wcYad7ZTAAuWCoYmmcffRlOsqnAeHGTw7FN9Hg+HUxp9Q0Ykgb5yLxoBi0Qx4kEk
llq4PXBGAlBK/KAR54kkO79NQrsYJTqjgkqGURDx9Q06ew4hQK9gyX+333ASmU5Kq1uP/9Ceup85
mX4g54adX5x8+TGeMWTvCPPXiqM2EJojYIp93IMY3lcE9AG9Rwi6TS77MPVkdftcgV73OSHYoDrr
fZ9ea3YeZUn0JRDQ0Ymskwd7iqV3rZBJ6CY2H/UKVb0EVI9CMSapH7IRwNOnb830he2w1Rc8gvZL
p/vxLU33TrGwtp94zEQO4pSnnBbVijD6a0LKtRYDRIJQ34GgXodsFz/cmDOY70CQFrKTZeSKoCbz
v5rPTR8obmS8xvWcNsqPlCS5Hyk3S0CaUPsyTFGe1rxT8fwUfm6hdgmTHYExE8HsfMIRXAMuTzuR
xqu4WbQiSe/yuAdcXsNionR0qUTN0MOW38oui6+ehTltmeU6FRIpTm/DBubrAAR+mOQnKxxZZO59
GxtRNWiiqKC0Z8v5cxiNWYstO9BOmDU75U2F6F33vPPpOGqaPjwXvA8BaB2BIAzVcF4QokU8KI/+
+I8IYGs4F1sdlnYiATym0bRnsMWm4t+ZCXWOzfcIl7OTN1epSzhHbTHSRMcilNHr/3+Cyro/WTuC
kuiY3koNTtVLEFxI/FwG47raqRSFuxMw0pS8ez8uTJ0w6sS5KuEhHu/ujs3zbmBlpV+DMe388GzB
52guuNRkptiI2XU94F4kHKVF6fXjIJQe5wDZG5lb4/4bLVMU0/g6dARlAhDTfaak31GLRyBz8DGY
i4R2FeY7tqtgkxq2Yb7pXNmw7gKtgZBMhecy0kr2kKXPZUnNx3IE4oo4HHHqhZ+AvgSeSktDssK1
g0JdGLDjf6meLX4cCg7J4x0WJl+NGPDLeQwMbpVG930Um0sgtVUDfLyG83W4yQ+1g1h7TIQNayhU
A+gPiBiUCIaKS73arZD8u3B2KS+0nCb9OWrdNvSEP6oI31/SAaUOJuJmf+7VrfIYnI3A3lNiAFrx
FkMEZ7knhYpCknP2DK4rlRuxJ66k5k8IBXFUIUuHg7Yqa2YNm16AticIWWcaS5L4cBR2aG1mkyZG
84BHnRT5Wett8gCix1fJOxvO1fL1ACznT0+bFmXfMax8VpUMhCftOrpqeL1s9bKM1/jg3GeR6pdD
VcsDvx1BUHBHiR27KCK5Ypi8jeuzUiEd9dAZq42VBMVQMwadh5n9tvTNAzTyfBowasbM8lYLv6lH
Zhud8qLH/wUMM7RBR0PXIlra9IFqCw8gSNKLdupaIDEy1V11EBOfCe22ByoVzE4YS6DdL6At4Ui4
UzikQEVniE3R3MytK3pw/aQIroujrGjVrmXOkxJSiSVCR4N1zRQnbaPYe7g9rMzCV5zBZrKxoIit
6jMfvvjdn9F70wvuKSR4/IANP6RnN50n93v7Tr7K1qY5xDCdrNkrw854LNSm3AtrviJRsTpEFGyX
outzC+zvaUuL+KADC20t12p3whSZ88biV2xOXUnVHuVnTFQCLbMW5VscZk5umijjabgEnMCO9qJp
g9f2gBYfVBTUu7ycfMSl4v+z8DYbD3hpkY3jQuuPEuj4RAqRe60Zxr3SvBQ4wLsCsHzbSSYR2vNQ
9r1RFyLIB5H0lbTfyRq2Ov85fp24w3XcQyobmvy0IIqd0/iSu8zWv5SRvl6z/di6dqjiO+S6W1Xw
64tfsobQaRFssQU5l1U6yHlSqTclz/wqes/NoIfbBGDjowH7eWue1OuMgAxROKA6PMpMu4NaN1YV
Atq2gQDLmB68NZMC79bYCCsavqkdircXy+1FvSozeiCwPePOt7+d6IRzmScll2diyCkpC/cM2vaX
iuTMrdoGQ56XTQRZYjxGBIJj/wZkc+T8eE3qtgx0xnO+FmbwioSP8HHpuPdUJVaFxqugMv0vv3jm
Pz0nWLJk3knZwYG8aD5FcgMLIEShReYPU4NrxxvvSksYguw+on7AAvd7swI9ZFgHfMwlHymolRs3
nvevj56met4dYKG8TZOc9CzJv/fsrPr1yc991ncik9pMx8DvKDVaImZQEvrVdG3HxE/FE5MoWAWI
oR29haenHO6NCn4pwBsDwnR3xxjbTHmMtsA8z16UzSKTrh0FEzoLVRxRvCw8AbNOOEqy8h5f9LTj
E7Ra96bti2uyg8mmezZUn8PIw0vlDf/QGUnKslJCbhTSvkCCQqOeJEefE+1Ub2s08iJnIAYN9Y/X
FtP3vRRIKzKf+hl19GQhDP5phb3+nKkV4TFTySPzWByWOof4SpKXjwEztfcq7C16tPBmNPLYnQPR
xOjlo9GTDNdlhEA+dfKWw5EX2vYRfpA4Jy1MJZQfLskYL0G/OoD7I+mB/ofrzfBguLzTHm7T3MrG
3z9QowBVuVljryQlw+pvXoivXlZ0/BwqUuNz+g60GzzD709pczZQO8/VKRB4f6ruCEflTwZ11lzj
R1ggCvLRTJcUMMSspMF/Uf9v0i/Kx8u4IA5Rip0YLsH6LzvWfKcd0LdS8ZhcowlJfW2qrc30SPJy
8RA+DosMP9MXCqJAOmpxzm/tXqumOhWMBfJS4cZQ1zj37BypJtDFe0xxaWECp/X7LD0l6XoV2QqU
V0+4zrKH2BaeoHtuijf4zxyP/JxjoTOnFqsH4XwRZE/r1EOhWmmiWF2x4q6PQ3WnJ5yVRl3CEA5g
ddOs1/9W3XFqQSEvFEohtjJNFI92alE+2fzrTjVlEqWfeZYktzv28hgUpnK8aJOCG93y+Fx0b5++
1qDRLmznKx+kk7l1Fdv5Eag56Iu6AyIKZjYRWRZ2M107IprRmdVWo31j4axKJOCBQeP0TyV4lQre
AQXGjGvtWTW5fJEzEO350xaeV3r0wk/boeBkjKmfcOSP2zQTAqqAXxxXY63MqorCYzlEaKXUwgK/
nDU5MOtWCwXd1AvxHYEZTX6jMX29CjD/T9wet20z1Hy+byYbRLqnnP8C6qg5LvxQTfYUamMMKDjt
fCEvvp8tECtiUjASoBZ4N0vVTeBoE0LCqFHv6E2XAVxSXE56TqxR0Jfe24TFKuyB3v0kTPUcdoUH
G69/eXA/vGMx0WfBpBfzALb7pP81qPGkf8ECeV407b88bJMmsiFvQJzrxplBkx/7uu8jkZSlBv1Y
jfzhLraEUIU6aAf+Xqlbk17lsx1w+jBDQzrp8ZoB2AF41ipn8+AN4/9+tzD+0t00ReA3WYuRRbHy
XETH31UIc4dzq0TQagJCTHONSqm93C+3o7VfubmEvRvATLROsxLsnQKZaTB6MyecH4GeOYXsSI22
lxyOEZFBkkf5hD7x1xbNNLhaqt/7iI6U1A6vc5p30SEMnlYYlujnHrjnbU2FnUe+D3ZaEldOUhnf
cNaUip5U6cIGG2iKpsMZbWBitXZtswc08KJwNCCA0fqMFRA8MBYkUQFBrMz9fxDtdY1PbQ3iqNj+
n0T3ppqQoWGwe+adNSB87Yl+WgBqKDHK33ff6s03Mur4HHkOmz7GphFRDjLrVdF6e03s+PuAMZh2
CcaHBD95Q+OZqymIlX8NhNXJrf5FpfmB0XlOn58oHcd/VgR7XUrR1+TryrlnYrBQznOZHbaKMvl2
TESVLgZE6aU/hlaBBXJV4YYKW52hecc38vmukcRX3Zkgg9ienkV3bp4WKTnNGHtJ8YL5yS9j23vG
8v3q6Nb21xDxZ3i5gaCFiVUjgxSQUaNL5CI0Wv9vu/Vxp7AiAS1ewEEj+CBX5buB0Gnl13ubAx8l
V+JJQWFLqZgzeYpX6AsgvIlBlGmuluA8Ry48RWOkPTDKBeOCEFjiVMIFg6jaOUQAenDOLxs4nVVD
F+BFAOK3HJvnVK4ukxk1f7AlfHG9wMeJPEKb/x15haeC4OTLMJTNrBALNSnWYcHQ8puaCOi1MnW8
nXVL+2PXivlKK9cfgKvpoGmV9kGVS3eB4F1g+Ss77JtA2Jp0pFi6qKofFU3N9g1h9zTI5ArPC+jS
0wF26DzS5WnpRwyMxdBPjTEt74fIK1SRg3kvfMryLre+y7+AZM61H5envoN9HYjcoMbnELaKdN3P
+DHGpW1eugSJKZaKg1JXjCxxehwyuzKXonk61AENS7KoLOLwzJfjl22siyJuYuBt80DSo2dvwObf
9DnGiWSaLuIrkJJ6AfvVF7l2wx1k8qlzQN6BzO521baJYVIbWwJ95Bq4UefB9jQWX0brc3RARhYA
0GcJLkvYUKtEqrOkIPBSI6L5aDblI1VxfBGSgoq5qa1miVG6E3sIGnWC+Emw67DfNPkcGPTg8MF2
s7bu1tOXr4R1+0xyi62SDJN2dM8vV/2JRc1u31coPOu9Z7zs99UR468r6cBy1LW4ftWCyA47CJpO
KUGU3k6GMiFpeNFHLsGzniHKueMDMco0tCKV7WRmXNFlyxVYTnoVc5nQB330tus61EA1BdCvvpHE
p3d4+qA8+GF5jlKiZV9kaIxwSC4uObxYYvMlyDsek4RSH78pBUVLL6iaa5CNg6V2N409irDz/Yta
Ogo+R9LZRLc2KwOGR/bAyzxD0mnDEXQ1teJsLtMZalBU0XYF17nm879nHZ7WS9jowyYOxx5UBNza
WZmYFptryfxwsNdCWY+Vpb5rsPFhcFTXKMD6TTebzneO6HClAz/q2RxBfDsjfLKw39ldISq2WEDU
8T21GDucJL1yCTbs6urSWGI3O2UA65k3sWN8Bc+6C17ok9PX2OBXktyPbmFqq0s4VLFrqKZR16mS
RSbJ+Elqw7JJr8GejGFs7kkbBu/eAOIsSD/hBg1p8zIt5zetJ7SWQcHBEE5LyZ5MiMGLZoxDnN2O
mI81mxdaQbGbcTTP3gH21laHS2wq1efhKCP/PgxBO5s+qmMA3vF6RzJp05yOe7CMS86sP5xj+eZh
P/x/vrQJqcDgvcQ/fWSQkPqqQocjKnXhM1Q2xrsZavEmBrXP1vDBwclGTq6saNaxwZX7g7W8/g14
Yhvzz8GHEb2RwPRg4ULeb+3ghW+3pHPiYSFZeEyAMf9WoRt/efKVTzffM5qcgnEYyLNnHc5dqtFc
5+NWShLfEGGt8idxFd+KGmwhSi8OAZdL5M83xu7CR1Goj4ImEbBabCcaacTWO5VRlLt1x2rLAUvq
ClramQRGU/TExGI0Jqlm8Ee1f1S16yLGml3O4lePWBSFeLDHjVqrpVpLtOUVdGjZo4QPTzodqOIW
vZx+gN4WpGDxFPGgZGd++sEEA+UKdlQC02dCFy5Rki5gxr9+6FBbIcnukZ73VdF5fynNP+kopiV/
xHkjvwS2iZOhTh+SLQ8PXNV+4hiuHtgSV5ftw8im/rHC7Dkl/w7OznSIGX2OYIhtdUG+iHXN46A1
IS7F3qAcfPlyuy9yMs4F6wu/+rFzNKgz9yx/rRTYXzS8bTP9rseIa4eeWMr18fbxxo6oMDbWfFeB
GNuDpD6CYrODEOpoHyAavWBZXDiHmqjW8NGf4wyjUTZUFb7W2gnJBnCXkJBzTuNt3a87ohWWT3hC
GRGCx/Q1kjf/b+WNu5XZS5REmeUQQQKK8jMuGL0hpZQI5lO3Gh60iKBju/7J1z92myx9bmHInKKH
uUMaFWPxNftqUCFctHAYxviW9ZuhAMZG1Sai5/FXx0sBmza+mGFf+p3PS95hB7C4wu6JqdEukLLG
wqGOlaN+lSo78aloVsoGE8Q0f3X88+lN+96sXXG27+LM4XT8JJmVGPjDNUWyGk6OyA8koqZzLwQ3
MYjMVgXmxj9+zTJOObyejqeWaF+zh1M2JDO9zc63DuxyRIlzwIujMW8DNORruQy6ELA/a/gDA5GB
hHABZUfC7AD4cik81YiQdujtOhhiy1WHJ7z/1CpM62BCG3R38POVtrZW9d2Dt3scNZpO3YG1TW40
+Uyq5eq5C/65GdCzo/YEtiFZaFXyrCN2aEdWwdUvfzoeh60qdJaVG/bGDmxVGog59wMX0VmOPrk4
1T1estMxEFE0MHsUmfuRdYQwOafuj2+yjzZNnF2K9s6V6V64nP7z8ouYQkTLyh5OONLdJoFx2AV6
LstclbXZitpB0q17RRDNQMdaJ6dOCuQ9bRMRbxaIdmQQjBLV2rMGy+Ypt+PY0hnkv7f3RMKfDBei
22ZUQGTq9BcXSpNukj9fL6f+KG8IH64abK7BjYR7X3N+rsjYlfahz5lGqleRjAt+8PGgmsJ7izdh
QjVXxw3qVTRRoqgPMZBtNh7IYLD/SMbQ+WDLLT4mEsAByYicE7RnnyMWaFbhosbVAgJ/qW1jHJe5
03KfKOzO1wXMIvWR4Vgvfflt5SyNxgYHTlTu/EfKnUG/Bf7KY32+XEbCNgLYQ6msuWckFs+pY5WG
SUlZrUYE3TF57vLNS5ymg+tQSD3B7cWXn90WRXwEjVhiCFyTT3VFqhC7FYyIIGiIXRhNLuV5B9By
LVLA3C2mCX9KqCMQSRYDRFLfgG7Fk3sAaIobB+mAbBOKwm5E8A3YSGBtsP3IEMp/bUAITsodZBhS
Qjwht/wECSCaYP+DNYongx63iuU01XabEdH9ux2iM2oT5RTtjZPPBX3nowEdsDTvqfJ+EX7EvKVO
hazw2tJ4z14l0XU8c5suKzySFjroGjanwKR9kUauBwpjPGtvK40Q0I8VZm0ZgyKoHgHHn3MCjOBB
arVCNcNcZQdnuCTyB9dhBvSp2pyHjZFBCXOopTy3voWB4G6WWN7xiUxu1mryKlHZZkojIlqKeGPg
ep5BCLH98wK084HdMEPMamcVVs9EbQuAfQe5+Ps2cUvigCLT1jXzi2fyo8kkYedobpC3/DjKc3Na
NX3qfYpKk8xkRPkXRpJ2+sU+gO83EAw5GT7Lhm+61u6IIrQ2lci5FNAJAePwSrdm+2fnu3u3n+2h
8F/SAPKFC3KiERzoHs6a14cqgTxYstEKAwxPTDctzuj/yzFJcId5sW5BGR0HGdty5wX6ZbTyUYZf
i902Av9dwAYKzXnFb+GNkBOKwENXfn8UQq8AVppe6ueRjkU/oiGfmocg26bUO/HoNZ7GcdTUigwi
04E7JaiFMQiwdngdvP0X4eP7WWkW9ELKnt8Q0Jlrz854QlYq367sbxJz1aZPkqSIeg+2XebcsY62
CFq9HfyQYtmx/6FVclpbPxxgtQbM7hMTZWX08AlYiToHz4clCZf6g4A5EBr71ii52IbEVnyC9eSf
N+VoQF1r0ncdt994pcIBfhF2t2HNtRrcm9034aRqkGi5DKxZdg5vi8dbEJol+0WgaUjEzZnaQ7Ss
vxcruilQwricTKlkTnMM9EDk9XBWy3G7q2wxYkgdHoxXku7CqWiXTpNlrVged3Qfm1T2PxVHESy8
OI2PoxdRJQxB3D82qAwyF65REMLbyQtUhDXGYpdhr3HvXlakLxY2gsT4mCEPy0+lOBh4nEixlJC3
91cfC8XpgCfz0B89/5Fw6pK4Yg5QRiDP3dXWqIZ0AUUHg/j9vVo9yi9mv6gFoCflhXXViv7HhAhh
U6jAr9kM5v7oLZkWIao+uuodJGbhNb1CcqZEbRG/1dD0g50govOPBqlnyG+iHrsFk+GW0wUWSG5n
nr+cXXFjowxlPfAXOKPyynCSvU/1c9C8LDZo2DJcA2T6XZ/jfD4EzuueL9Lqei9WdDeLHty5XyEA
IU5ct9E5jz1DESEEv70QnHauJMu+43S5U3KA8WU0nrXj5D9GDB+mr8BaWyh22dXBYWYcx0ybcy/y
UckHd/S1NS0r9BABejbLfM2RlS01qOFlXbTSTpEPh/S7O8jBj5HJ2sWOAJrzKgHm69GGTwGgPWWE
tGu4f04ZdbbCrxwBmkbMMv81kbnSafNPW5MGSjZx2x8YENAwsImlBcEgKoGhO9Kt0Af9OnBo535z
uvJK2rh3jlmnKJqmbE3vb1jmlssJoKIrOtUI00cTpjji5yv1tF5jNbq3dRHKuGEzJZ5CRdwdV2b5
nB7u26k/AYjmqXEpUWe27/Fm+ntvGEkUVqBAQimaXvYFXOnxUGUmIntHcSZ4wIYTIRvzEaO4tBxi
fiA+18xL5PLA/AmJhWg6bQ9f5E3jIe01myNgszYp8ATgvJLkiNSxvjKR357O20GSh/IFkJW8h9Hh
3jq/pmtARg7/gLSyzg8nioGyCNRqM9jMGf/TvlCB65tXJ7VIUi5iWA9Psz5lFv6JSXuH2aO/BQfS
U/1fUnEUGZ1nqwFU7ZZR0YwWz0PGpGdjQC2uJ6f9FGSKve5xZQKK+m2jMKJPWF2PW6wMEH/wc/HK
2PcoJC2CqjIP0LkqPpZlejHcU0utyiromr4lpKgDJ8KRId5OXbz6JFmvkHam7MqqBvQdassmCgAu
j8I4EFRrQqq7Tw+/1vOorVcW1JBqlnWZnySTZqhHE+b89fiNbB/F4aV3kdB067hGvCUOf2VSv48A
V9LpFpu+aiJQ+TNy/H2ISRCqexQvsBDwxW0eoUSnJ06GOH2nA7UZwqw3ZKZWdVBnNUUs6KZDs5Xy
xDqdiKp/y436BNotZgEuaKB/Y3IsAkb31ub2nd/SI92QTcjLtNkCrDy4isbY5zc6mh1aIP6od5bH
nD4GclyIcHryKMDp9PKKzC+wJZOy+NMKkoMVCTG82szpK3dR5Exg9OZ3KJ97Dv+hpBZKqecVrYIH
ex+G0NrnhhOQO0T8PzvA23KzordlfDqnNj/mGpeugjtY50w04yf2OMLYaACFYUhv+OCMRpG4BLS9
sBeon2XE7aj9sMMwrrnscYFtvyOa3Cwarz7Xug7z3UjCKVm4Jul/iv5LMv6xCKeCfwcmeXSYC7V6
oCCVkk3ZnaUlaPNpZzrpWg220kv+N1EtVKYV2hQstOgq29fyY/mG4x8yNmVtRnfYqwLLTYe1CPS6
T8OvnFvIvDyUKcepZ6gVvq/aWORrZeAW4ZEObQ9kfdeWc5iv5NHXTjR35jKDq56mfCg7jn7x+Lqx
4fjbiKwvS/gQuo1O3QlqFNxN021iS/6SKimxZqPg7btJsrBakdLigRbmUzU57OO94hPRYWL3q2jG
ZPMuSrsWh37VSwYElq64fIiS67d5r7T3d+ayS6znLlEaHkvkr9/agKf4et3X/2F0xqoJA5GDq2J6
YBJRe+29HM3I11uPqDl01Ueh8YYzGJ3ymYOmUqlWddEMLJ6Slh0RXd7Wc5FyYVHHq+ikIHrI3oPj
BlnUs0n1cJmZWDdEYPDQ3VKcahqY/RxhPa7qnK72gxEFrlHneqw70syJUMS8dQbw1BTZUniARPq7
hCy8mLDh7H8wFmEicShrAgN6vLRbIvtiaK8PZ1qyGD2P86TU52R4l92ppmv8WrH5iZBa7OPgo4VT
Tn+Ge6baNtLHazJHU7qHj64ztvt9suQBdpmRZvVXzC1BYkb84bKYn0IJjTCadhph7+RRQunUOtZH
zjFWylOZawVhtgupgrGLmTNL+yVHpCxstjpbNY9S5Hz/2lMSVlGbEzQupYSeIyvynCOE24fL73XT
XxHf/BeIy4wNmrWKmzTzS//b1agzvsQqXlEXns3uNq8iSJuNzbq8bIZMBzPOF1lqgpFN29gQwW6S
Ry6yXMIySFRqG3FxU3pXpb4SYmL2pAYQXf3+FEieHqa5JJYQZiYZgBB/fmWyE6VvqWLiVoCQlxuZ
H2AWoyHA3lafIekLnk9rqxGzNuzvVBDwf0Ynw0Y0j+T3Dvn/mK5whX8zPEp2NpNfpXT0U4k/8kFg
eAWg/er3NJhEAQ08F9h2W438khizhptkDS0iYMTthk4xV6QXes23iumMYyPzvoyrZxsKZVkqSWxY
kuSezotFNUWMw/iH5bqNjX9GK2GxscaFMO64TSaIwKWjyFnOwOKNqInwhrkAMjDxOAKp8mjdQuC+
byMCi1ZVN7Qr2ywgYfA1lpasee7iL73Nh2greFZA2QSpq2HReJGmqIUToCEpn9MlhKCkgBkqhqFA
3wRQceedxo6+leo9VmiX4DGU5UjHQHgZloyOGNW4WxXz8Dr+QWwv5vS08lPLxFqUIIl6w9/nClSx
u3CR5WMqPO3Xddn1CNjgADx9vV3IKaoHLimlxAFW6fZzGsDchULw80OspDrWp+BysOc2TI+75ykP
aw/wn9oSG8kbiCubwLrtFz9qbOA6PmKSyA6kNCMgNE8HU0ucjpeMNHf5nsyzdQDf5e4Aw/G+Y67S
NWqrqfaSagvw1B7F2+85Ysr2b3QQC6cKgv+eVmt8KNz7C81ijH5DNcWeJi9F/DxoNwPL2mLUWlUv
BGVyvDcs6Kx9kuzenxUen5wm7cjpBg1JSvgl6OyIbJIOJrX+wPEyaL+7/uHUkZuqNL3Cz9Ub/Ya0
yjDSTpv08CrZ3CoH9DnrH1Rht7khfKvr1l/v6SiBfPZDFQEtVRFLJkz1xfA8lpSmx2tknqFXo+NJ
Kg/HdgZqAGCwlVgx/9Vm+o32OVDE2a7FhDuDjyPoBrcrCtWVfanxu3WpGxFNNhppQlzjw6HlEB+0
lLwRoggbFRoZ/7g4f6/8VltJD4qENbFPYJ3mUalwjCdRFdt1Wp1hlQhG7jigqXz6xhlNMfDRjS/D
au9pycqoqK1+cvvjwpImkhc9PYUShToS5FlDB6d/Yw+n+rm2VjGrdgM3XeVIPrZXsHrJmHeliylA
5gOTfY8eQC7mU88cpI4JqIx8LsFyWnZUTlB7XpqQDNilxX3/f8w+5GsyPxXsDOrYgMmz5HGjMjgf
ZCfHLsAvYMuuhrgmySIG+DMAxleiyhkQeTzgxttb1Zx/pLSRueq3GM2C0STm+hQuiI/tU2YgQU20
hUI49QjZrj5fvYO4+iv6QzuqiOPy3E+DjGbwFgZ6NRjBHiKUsQi5mmiID8yJH/tFnkSBHU5iHdJM
cQv71wraz3ct64cse5n1mzUOnAh6ryne8pO1rif5lxFQyxj1/fT32VMQ1se3zgJHiTnFMZTSd2xk
ZVmSgdnBfPX8bEdo+zW6mJ2yBV+giLRrqOf67QKwqDhyhKBXHMf6TGZ3weCHmwdvRqYDfCDB3uW6
jaEf7du9w31Q5pEPXMlDu6RaOfG9UBNq0gk2Nx3BbONorUJJE6cWRiEV/DxGR5dOpS9xZH9gPz/X
qrsyZuYXDp/yl3QV76AndO/xUDgcufCVtKzprT7f3orSTtbmhZBYuh08kxfTbyBmIx4BUgMoLho4
yp3ncF3HiktinVRCQe2yt/yICns5vnoCCDjjlvcsDt88/Fhs1I5tlWSlfxUO06z55vcixZAzbb6G
5Jn+ZOwla2uTvh95o7cq7Dh6xoyvmhhTTllS9AR2IJJGFNlnDCekWWjhRk7zaO10UofCmXmXjPw1
axxwp2pPDUwUrOchlDcT9O5rC2jV61luEZcU4RAs28KrH8Uwg+/w3tyQ9rhgXbqT9gxEzEavIYp+
ZbZobqHEAv5ei61UbhSsTp+sZDpIyBXa9HSFNdCn2orNvs6V0tkTvYVWgIJOElvr3xYtNB4A6wms
EHoW37mEnsvaVs6vnNT88RaNMP1sQHbZeDYR2uVFa9YSc8OGowO5IPsYz2tWVaOVVQhdrGkxDlbl
jPgfbvMwxxBVDJgQW15uhQefOUhMsfQwBDGASFm7/hKIL3/bfF178tTcxBWTHtTnit4mwGDA4Ser
j0PjH3z3mRXQ60mfywuUEPP6HhzAxndFjgAV0isUZNRB9MpgmkYUJaXnzkUtdy7xU8HrV17ZwmDK
TS6qF60VxNNDTihPTqmK5libYvyUpaUyjb0EEAW2H+ZMyVfrpFL53I0EIHPfQMfjx0dc9U2W7WiZ
HiJeVHQ0Kd4ScDQxNy6iEyEpukHAngJUunUFp6/4+gG6RafQfXlZBMgzkOcB8o/jODhge3hAQ+ie
A6iKniUwYs/9Kee+sJqxOe4Xs4+iMQio4IERkCMIEDneuvFIv6Uvn/ogY2/Jr0VDQiC+gSYYc66Z
HdmJIKX76JznV2K4AHlS0zS3bkpvev7rcKk0Y+YEFc/MgS5t1LgnVFzV5v9W33SJ5+9d0a4XM6Kb
zv8t8qr1xPsoHAz09LB2gIsQeb4sMOvcOYZfSW6yoQzjDe8alFK87STWZ+0tCcX3nIFPD4iMP6/Q
ebIuIzHMwfpJqKm/hN1zlsGhz/4JgpBdCjUidDeEEBTECt8U4zrwh978JcmkIbDZYK9v3MVCc8eN
RnXj4vJYU2iYEsYiOUiyq3I1pdJK71Q15xEPWlcb9H+EaqXoWSmkzePK7fpcY97jVR69CApze9ua
ZcwCPKB6seCN+DfEw/R1jYoMlKxDWFm4xb95c5c7XjwdHXwrGWN4pjnjqcRfy+uhriSaSH/9mka8
VNPMObLl1fwMnMX1u5/kV1zhaU6P/WTzYgjYPX1bmNUyOZK9821BjNDe7Y9+4agRf6XxNGyn3Fpe
o/+YnoAS+ZbwFKKoVQp3VJsXxTxoK+Tt2lDBWYzPvnvhzH6Iu2IkMpdckqRSAFGLXKOoe2x/hJ4m
w+rHuPSvCbopU8yikiK7rjptdyW7ZsoW9qkOmVN7/cMi8ObAk4TE87DGmkpV+llnYgmJXVE5Q0v0
ARl1abMW9sMnrm2dKr3UkKHelk2IDaazZzqKrYxdAhDy9IgsKvkcwyurcjTG35Q8+vnXDGT3ZhKP
3Ngr8pjJILw3KRdAY0B/JoB74hJFNgZNlWj+x5KGurXKvixh8pJ98+wXmTm+you6zvK0mi03+lzi
dSyPH8kywrQMW7Xr8f2s8Gn43ZqYWj7m0uKUUUG5TrGDwlzbxnZQslTk5jjsxEaH9F5SD+4bexEu
3fnpuY6vBzqRONEkI2TxRuOm+QJdKlRZ9Uj+j0WW7zz7hGDo2ClrAdbcPHNUhDIqFJ1Mnpn9QtIf
Q+7EO+sNGZnnu6t/AyTeGwsf3VRy6AAkaaoXHzwVnaWqyEnKrwie7h4YuoaEgAy54MPQ8f3KYT8U
wzvIMfft3ntD57abiVq6aPuHXtoCpL9BQIKmLToBe5yP4Y2CEirDk09zC8sMeiLE9ylADKFKUoOT
CRrEffZuwwf/QceCe3wbDgaYoU5bDp77ieMlok5EGmL6Ykyfe7t7KheMT2MCgggyCR7b5/cJd8vR
w5g+biJlrgXRe24EucVauOzcxwn0pIUsEiUqw8KGGxlonBH0U8Qo8SWtjkwwZLn7PCFoyde7QjWq
b/xUC1xUBQJagvrOQ403AJA4M9UGNiW1xiHS1VOvlA0L2tr5K+JLuf5zt45K7fDjAI20tMjk0Ejw
GDtgG6HxdrjevllmlSXJ6NCXobF7Nja1UUzu2r+0Kuyrzq6607eggOP/0wYcQDrJPfhD1LGd6n3Y
ECF2p+5hDZEbWa5xO85XB4QfG1wOrelvxr7GPv8LakHLyNARL+C86XQ8yoPjc7iOD04uTl9hrb/y
gRoEMQKNCGuiMlF7uSJd5aFkNRXn/RaHZ+wvMCi7n8WCTPqmnkR6yysGPNCEDTSj93mlkhGC94IW
odrwfwE9ZJW/O+yhMRjueYBaUPIHo+Zyn5Nz9q/lYU50HvRNgapemsIV7ptd1NrVOMTbZySTU/zb
iFF9OmzZgCTGAnH25I9V8Hs3Hf60B2owU1Nyct6h/7D4IwVn4+U0k6tRdHi0/3PdcnQ6rFXjxxt1
alXWjRWGMQ9nOv7u6aFyuvni5Mg9KrFcqr5IkC0614zZaPLhZtlLUp7oH8mMdKSWnkGTTLySyMwn
zy5nU9LTToBB6HJQeCTJjTTuIPmn+G7yoRJ7CLmzv5nYCkpMSLkfE0pKPe7NPLeiSrmh0GQdJ2QF
lwr6tJXb01Nl7EjYErziNwAO5WUOCtXsOmWcTuAOikeHrX0AazdIb8OMCaNYJh1Pf3b+PCJWIxIR
pu6/wxS9b7lhtwnMdLeoMthjutj9FOx/C8nUYBJABcyL8abpJK/emo1HOZqzDz01i+WVUPbM/6ff
NygS8LEhGb44s/5VtDZ4Kko9mh3ErWyYSyGyr49b9lG7TWKqhGWOIRaHHAavwCnrhddNtclJ9RhJ
sZKySsX+yzezk6/i6KhwukSD7+S872KAhCkPk/lodsLAbv6hbGeLGwZ4d5dG6ErW5WuvPVqWjDxT
jjmyPb7rPEgLsR3H3CbNN4tIEMQNElDpRqWWS0t8hwIOFPVJdQZ6cM8WFCyYfhfgO+cVObX6FJnK
hMq6UqmxlPNA3YRVkjXD7w2RP/yQt5TGmXl0NCHmpmN7HqHgyKAPx1i1ZPwJtcwPAqRaxyHLriVF
AteMmM0SpUiHesC+a0/Q8Y/S9xCdRMzTZIaTII38i4zX6Mk/yqX/uS+NTok+tEmfTmTZislrAOm+
TzV96TSChfSXCdXFYF3sZ65adLoxmJtWcu+le6Qv+XrBH0RX5Jrht8cl8C1odtjR6Jws+dMbaVuV
4RAyhAzFkdDe2gjeR6CqeMK336ASfbe0dzjgpHBroxbcsgbmZtdF1J/Q6+K3Ky7lKHLMZ9mF7QKi
JdsS9MkjJtcOQUlYGPQMwVGI1YdktCwyor2EOga7Ntfoaj3c7Ysi6bP2FvmaAcNk99ZhXrManW1y
IsfbinKvQk7CMIptgEy5CU+AVpc2T/O+6tcNFIwZtlk76X8KURcdBMsTvxn2dGAlQCwj/xuxI+Ds
MIeKZiIM4lbon86qqLs87M1qH+Qtk9vd2EBQQT9oejerqilaatCPTPpZ8SmE9eRPnghLKltW3vK+
kMg4qvRKCIvangHZMLX+/Az32R1RVmQupP7SJnv5OlazMD+vdRd+Hkid+IntQGhiPn8XxUPo/zxX
JweJvOrYhtLr3KIfiVuRN+h8cH1QyKo0LvKztuaJUEEiWRHCtidXMUXcFabKZg8clWp8j7dBLZjY
hLAu0u7GGyc73lGlqPKS49aHhheqx9bJoZ3zETEkM4MT8/eUqHGdAaJKW1XxF2um6vO4zdgIYhBM
tfwIJKtmNREFz2Fca1OtExzQs61B+LCDOh16vQLFFbZcr/VSFBFUnZAjvQGppJdtZou7HHpv6hAY
6Ym6Mqy1Wa5Ypk6N6D/rGQUJF14RDYfplkq9xdJHMi/ZNJAPFEPY8p0perE65qlH9WuixvftZ39r
xOi4NQDeXH7LBkerhxaLIECUxQZa1+/XAPcWS0MjdHdPjkQvtuM38EtOEFcjCNhRoh6dq4iMC2TZ
f1+Oek6cH4yurBp2BTjSj/RZsZXsJa4hpoNO4S+ZvG6dhm8cJ1Q4Pg9vNyrfYO/bkNlbHqEtnUhW
StOiVzsKqCePXThw4MNQZNLX21OEuGE5iRMCHjkMnxczY20wjpAbPusLqERdKwUEnE3JWPODFssf
O8rrbNBuT39SHWxPzHy+F0MQOvpBrtiO/Xu/Btt3oIkNQ9xc7y9ha8uvXpPBBtsciXafit4w8ddq
nE0eV/S8kerJte3MSZP2o8MjWe0InXXKDL8tbhBVYZFQHOZYxpBxhXNZdas4iWqWMvNJAzkyxC1K
S1ZlEpWoOUvjDktd25w4fPj1j6I4VwxrsdjOFRw9nzOzpXh0lSTGHUKGNl1CeoQvYNXV/A9foABh
eYhSgaOH0LfWegxQbkzMe7vfk+ZnrQhPzFdIIjzsGwDIH5rFlOklyUo7DwvlzliDaMKPJIMr64nq
mXOpMKg+cDOkaz5g57W0FSZQL4mvXjTwAe96llW8GRAP9FQgYyNEE+mz7nmntI+xcIfLSWIDW8JU
1FE6NXhJXokp6mV9crQ+6qZ9S0MLmDF//t2fFLP0NTEtWP/3juU6To7SsCbFeQmwc46CAEBBoqHL
QnDOuAj6MfzxharPnZz9PNoA/MQmL3znSIdl3XsqByExA8/k2iU7U3Vu/25tXHa6SeCtS64n4ZlW
1YHkbzeXe3HEpLsq7/Umf7d0fnDZ+EKxQNFm8hxmrWFAhyc+kfRQUj4EmZf1RipmV17c9r5m3jq8
owABxPbSzIZBOpcAUmZGRcJ9HO/zu1Zf5+WYDV7Ssz72Z91sfn+ekjo/NG8Vpl5a+Aa6/nQqGNUR
iObyz5uSpnO8r93JtFC4WGrSWciplxHeA0debw4pAkg8zHXfFYNzUVKBec5iVYfRz980jWA3MvBT
/k82F211eE7V/eXqxXfKY/+eVR7Nj7C45F2B5ZaPQKHKUn53uMaopZLVywLnbQx0WrrORC7aC+7L
cU9UXzzLciQLvt8nNkcrWS7eDhq/ld1IZ2W2l7tFmfnHhFrgDLSZ81BW8a9UX3yWT05EpJ6vRMzp
IXixroW9VR8joI0taONrnxyWu23rsfVZy8GFDsPejfolJbVRH+HdPWC5DfMV1ZsMDKAm1aieQW3D
LIrpz8PMNbXpNfG4gksTHjcJXXi5xqveKdE9G1JnXwOuvecq9xCmfWPRVBg/jXxbms+ELI+afjDR
5ogAOhLGgfYUjCkHAkAQqixd86BV0US+WfGj0gMbLr7dsw1Z+sIjiIZsMYUq5HBV0WljmTEZrVlS
EA4X+Y5GMg0JGz/Vx6Ldn5N+Z7So0jwUB5VGn8UfVWSutVS3hTlRu0yEZ8k8nglsxlTZqm/dvB05
aZ0iKhYxukyNAyK9AcpKltNPPwGC04gL1JRUZGBkWTHGjCGzyZ8pZNif3r7X9+ZjsgYA6vC4cbXq
TqkVureN93doNIW+uwW8jtEU6aBIYySeDFHDA9T5DvTmW0M/w9mNjL81x1lFE+5S6h2vjPr5Gs1N
xZAjNFRMKjq7FkRUq9lAh8JX0dnr3D0e/kz1rAuh7BwszgWV5r7dKMjuatxXJLrisLSR+PRnWRKT
Z9hXtqwhw16/xtryujBxttoY1PdoGj9ZzuIuvNfNPS6BgSACbpQ/M3SCQBplAaXyZcfrSjLb6gXe
LW12tLN4Q1ol9JnYBQ0N+6IjUeZqxFxURmoFs7Sjd/W0IphoLMBWtnVefnxjXlZFSpscmZLmuGOL
zRLxQwA5bGS5cviRFK76PJAXmRHj03bKrf63YE0fRcWFgCZCmZShkoDMD716/eImGr1dzaa+Ufwy
i3uvj4iFr396Sczq3qJtnakPs8HZACAtzEhHHIPGlGd9bZlGcLOHN5jiE3mL2U1NOB6VrxQkuERU
nl2NRZZDVluEbqtU3EV7xKI0oGfCPvDhxHVNmJYg6Fl+QKQaUSy3jU9Mb0yaUKjkfZZTsCWaTax2
mFYbg/nDU2xTtWgjlFZDyonl7pLrD5wpKXA+3EQcNMmITOVjZsjeZwYtq/9594MVmkWlsqReed49
Z+NYvBBOTrCPfuH/TujLuipXR9rsq/P50ezNPjW0ylHhmVb6viDxw/yw8RB+a95m3tAdV7Xm37Uf
rjklIiMC5pUPjjnRb6ETGjT+KKbiw3doZvHnhkSvD6awLnLk183IxgQWeZLr+SbUSKDP+KelX0cP
hZYpGEHqXEOinBwpIEL4dProbOPFZntnVlcNXD9eZRIPzu5SSaCcCIGHrdObNhX4jt3sizyQ9lUS
NmPq41UOmnE7sGlVXleOmmeTCfC6KhRJ7pOUMb7l+VCxEfVzRHbO08aDepzOkbZALZFRlVecUGCJ
04Ib+6tloLcvcb+mt5wL6mSfUOKaS9ygcImADgUiL57SE1blERWqmhdfI6O+oJvF1EmY+Xp+rriC
9oIooMqQn0x2oXstmnD68mHAnSTAz3mbdeZX7e12zvT1EK3cYU7MFvQHQjr8ptDvZVhC/ObAHBLg
ubG1FgT2T2Ef8dPQAZWKNFQNhxYxkhNOeCugzwLaATumwP05Q587w1GIjcqTD0IOaRQ0NBuvUxAr
U7zPbsk7q0sNZtmufFzXceyQ5NIZ2nWOuRMT1IsOwzaykx9O+B/j/x2gFp3SClpmpcvyVmfWmWEF
MNB5e2qoeOMQEfzj6cut4Zr2uO0uhLhVudn5t7LGDRxLeyOdPMNhV7uH6UIqZLr/xJUdMVimPW0+
It+N73nlezjJnu3mr/Du3S5HnyfDvcXUyWLsXwy4UqsCt3xOqw5kdSugpOY0mSpuRX8Cb2sNR/L6
Vj15bd04Vmxh/5mOa5nFezNpPDxQ7SI6v1L0BvlIz3nHTunEM3xzbBFbHHDWVA4VfqnZmnLvbnV4
DSNptSXwuMnMGCoSbUMH01g21j7Fr6YgP3013huHXjrecQLezWI0ymxUt0W18f4zbhPwdgyxGq6n
nh48Y/WORR5RsW3UfHiH7rJFqq/j9AgifDkZUCxbVQA3+klET9uGQfLlnLFSVvldqLhgRb+cXr9H
1eAZkYBn790vXFuVLfuA1jboYDTCz8BXqVjhF91C2DKbDaqwJQeg9Qmuv7XJ6BGdfaKQcf346QAW
X7nkS10buMa+fXq3KjAkCzFjlKOGTZumN/QxHU4JbO9ncdWyy2BRxsS5jgIlaiBphdu69MjjYsI9
zXyo193klFMcWrvqf5BKngX0rPPCNNjrYEM7HR/nPbFZq/h0Z+des7QdYRfHYiyLZ+sW7HTEUa6s
pOYB/5zv9QbQyV6kOESE0KhEampdcf7lxstHUTzO1yYbfQmRpyobfhyEkHxaS92deoQacYPoVkKk
OES4WO3zsLE1KfFvBCawg5Nt6PiDaQG+zRtWPK1WJsmJ5YYI5rKqe7JLW+3xSdLyhUDa4hxklsiy
cgSSgH3m35HrP6uFT4zuNY1/Urw47iJfvn2Kl2Fv9icpFgGrVl74M0lKBWMjwxcxfHNPnKaKeY3p
p64wg9B+9iNrXDY99zSXZW0UJIPI6dDqscXi/idMDGBNbN0Ad4sm9ZQMFbK3ARecgKm4ddq6yYMQ
YY2v/Wt9hE19uw3hQ0D74kh+TLchTP6Y8z/eGhQ76+08ThfqSjerNzZTt6dK7WpsCSuTDETbeDg5
9XwZLnC2uj5HxiYILxM6Uf+LP9F88OGmdyQ7fl4tULaXjngTDfuXKvY4nWL+P1sH3K+BNlZna39o
O09MLuYdKx8RI1ODRnT4Ju+lTv7MD4w7+oK08qEqPedj1y8xK3P0t0+XjZHuMf4xoKiNeCIefuYg
yW9puJgiag/cQhg8OWCPkxD9hoZJzcPe8qWox/XQ/iNEZVU7Sgarfdl241w1DI4rCsNe4Fj6tS6y
h8gzJ2vENOqhEsWnhLmdYQ6L8vnCSUETbNVT7b9oqle41itf8kvZE8ThOJLuVVdZrzb8GYOILlUg
lGJ4qBiSTV7G7AzD+qQR5rfp5LItxwKzmq7UREWBLCgubd5eyBF6dNh14CeV0nWWGbSlUxyxxVLZ
Y03xJM04hVFh/lmXb6IcbosInDuMlGtHXxNbxfWZDYM7QpuUMNODU48vEyEAn/i5YREhBHje0uf3
EKFHsWUSh8rKXB82ZAsaWRkMh+5KRXWOqOCaRABJKpymnOEkiHlJN5AMQiVRpMI1g/HCEB/LKZgX
dO7c8N0g6E82W62E9LHQpj5KEvSb2P8JrhqY78+I3W/L3CP+t16UmV6yPeOKRUpNApQ+07gxzoiy
FPb8Uj5qUI7mInBpFFJ9Q8p+yZI0+y/6OxSxWTEJJgeCtsG/Dott8Ugfk1uggM+uvFOiEXQbbuaZ
Oc9JN31kuCufaGs8I2ZqCzrtTHPAzJuQ/gmZeIA4JHECFLWgDfVWrC8mrJPhD6mOqUIn8dyLl2VK
eWlLvkKbNnm8FS4pPHElSRF+UfH3n4uoOw4MwDslZodQmzH4PtpvQIO+1yOQ8ATHnqtByCKcsxtP
g82DAHfF61Zri+GpRvOfJtEmApAkpgLhE1sLs8uBPelwXgebjPvdPCKNNnQ9HLnCPeRyUSr3i64c
VdyYaJ0V141luLm1r/C1dpj1ij1mG22UNlDZJ6ePXM/RA3tQ+LPb/ZEico7CNhgVi1gHmsgI/8Tk
cPydQpgnrjNxew9s6/rkmO6MS5br7N5d3BSU47GfgUDho5ilNl/5/rXoczR1BbTEmU8xHJeXicje
svFec9rgc29dHKIb/njaadGKgzPNuljz1B4W5EhbUAriHGv8BaKw1n20rMshC2gIROqBSypLWzsg
GmoZzBV4IjJ+8z6I3nUPY4TIWEaXBnoV9SAUlKvOiux3HDlDbGEirtPibKe4HNf7A4xc3XVOZdsW
QNXdLlTnLXjuMJ6+HCWI62swaGZeH6cJcFuAr4Ks9m2oCM8XsdAXtfaZga4+rVFok7W/G036eABi
a/HVySG36keDxa0G5LgmMHlbmj16GTCzdbeT9Vj+UJLYJKaaIFgf+XEvHn5B887s7htrQfcSoffW
bC1F0bkU6xJTwTYSBPfnACd3wj2iCm6p/Vl0kKCi4vv/rK74HBUO8cKgPuCQyECrO6nHVs4qO9+m
MZ2M8f7tRC8rT5PDTYR3noJln80ED/+hVP/1soolddjt5liZ7Q+hYQ1i4SjudOmp2vCvTl+o8nr/
K+lAagjjs36I0XGmY8G/oiQR34VyE30sXqfLRYKimmgLcqfTnNukJ9H507xvXuC3S9AClKOqoSkq
j4tL1SGfJs/4zmK7BSRUWR3Qr3OfknlY66eRQX/sQEUJEOEyZk+rMtqQtd9M4P7cKVVQIGhgPcSG
KPpupQf3Qw5chATR4azI+Pa9+KBkwu6kyDyoUm+M4G8kzl1un2dklt41xqbO0imWfs2Gl40czuzb
tmH6JOAi2KROAck/FsOAeoiHPN49jv+Qjs8Ro39IwFjTgR78XmPVwxylX/Z7tvv4S1d5Gn8Z/0lw
qK2zDYepc5UPInoEOzJdYQ8z5j3vCrCNdk66amg/3GpMir/opaRzEGHgK/ZYu8LNOEG++IPjG6cq
EcaOCg+vx9DUTCgdjq7qQ1OJQ2HjbkW8OUxPt7Y76xD9UIC35q7cufxxoycz2Vm42WMkpfKHJpI9
agwGVnxAo0++AGATiXeRsVGkaLxvyWeghpyvBSAt4JCfHctIdXwKQOAl2/d8B7utXmoNv7WdS0Ie
Ad5vO4wlV7mw0G0PC94k//6m7TdgSW8JY4UEY3OZMOaCSYAwCtrmHHOwuC60locdlBJHOdz4YMww
azEIkbn6M6we/n7RzOfCOZjdj5WYASpBUAxIq5NxIiWHy4M/v6NyrBjbb8B64N5YsV2OIxm+0ZnM
bfzMok4xFARRkXrPvsvVH5HSOvRUSbLHHitdXQyPfQB7wLCV+YOqhK6wEQBOGLdu6jzGDNEH5wyM
0QbELPlrSEzlkhHKmzsMxIHlXdm5+09WKCMR4ZQpUDvkKN0CJGX5IPaw1UXEYJD4t2ZvANf1DoIC
qWM6QtJhaLwSBtdLpf3OLL1bSMBvOaSYNaRBsJlJ4pb0joVlSzaMBdGwDIIe8iVCeLoHf0acS5QD
Krx04RUOzn/vXrfvMTXiwMGQ2oscBtEgd9l7NFuNJC6VfVCs1eFxDO3rB58mL2yRG28+PgwIfjzT
FPFFogbfcZt3fXWTRI3FrVtF0DcCa0N+M4qy25RX+i+rMwI2dXsDwIAS7st5LZBIdGRuKVqk+FVA
n/bd+85QKsr1S5H8jlbHYHRzOsMJNxav8frtdAPEb2eRp+89p/6OcYSbTc1S+NdnrBZ4zrPAT769
s4+K5qBDR/EbuBhi3xlXuv8/Sc14RNqrqoZjXnHgnWwyEjBqFWhzWX8x6hvc+cuP2uRdOlZDWS01
9WyPQilLyJW1H6D3RO23W4ZWU6keNa9FmZbEl4ik+vb9xItasjUF4HWAydaiLctfrfewtFvOwQ6w
aBsVLxl7ISJ+m/cYIZ+qm9DEjHTlkGJfq2/YZ7h+b08tbEF3EzFqg3gqRxiQNZV2id6BtyFRh9e4
EtggkqrKm74TJIH4HGcC8hN2xou5DpNWVbMVxt5li1zwyvjdbsK9c5cCQkmhPW8EX7gkt4fyD/ms
h405dAQa8iXx9R/InzYjn7t9iWIXZMMk9O8O2GwJixdIkuOjGU6FNRrIkFLUFViEs9rF9VnqGxtI
rg2gEgOb13L9LUAAKUU0sz77fzWYO8SnpdqFq+Ej5MR7yWqf8fb7a9hAL5a/Hum+DskcAOChKc8o
eXPQwBJ4IBnMizp4/NwYNUJjZWzR9VexvLXO3iP/gaZh9Cfiq7LJVRQ6/9C/Qqq737HctMWB2RKz
/dyrQEUzhrWHKzCi968D5JUbebcKUbfN9y3m5aTsYP5H6rE0Dx/5bs5dokl8MRJ6kak22LZ0NbMg
D+wNSL8qcvD0I6MY9M0QjkhrVYOm7l2rUaO1U2XWeJU0a0C82VtVNIzNTKtoEDR1TpgDGMrj5oep
roylxd8OEXns8DdFScQ1JVZH811lbu1eYv4G8a5usfCe/Qd8Z4LyX37eUqy0mUT4qDaiHpfFtxIi
gd28Vw2OZtjknhOi8PV/mw3tTb6QpfllVrKD28JiQp6TLbVcNVOckz+w25qbhGu4p46ypcoE41fF
zBihTCudhpnXlqhicPxDxkX0LI+8pV9m2xGCX5qIRgo94RcuiPNvHZB0UUlMyWYm3uwxcVPABijB
HMAaGV2h2ecwKBYYICyEhrhx7rBGTEFQyL271KNm25huw0DdWAXcB78qujNOEI5mkL2xbHULbVZz
C4NJ01oRzMAkAqARZF6jpguvCytjMCYdgrskp+89Pn9VFAnN2O8JYTrtWs3hZ9ZJD/+jQadC9oMV
6V5PrEbfwAU+W75YlmXbx3oODpGYlqOeDWoJ0LrsJrK8p591NRhH3fnBom0PQnWIIxyLTwM7pviE
zBg++hryuiFkb0aloQedSuDQNV6F2q+L9ZnJBkswNCfBhKDpNox/Uqc2GOw7rPjMb7W6nz8U0GFi
nQGU6X7012PAQ7hsjFmtkkVS2fbvFap0vte5fzSH+RPzT53T96vcBtyT0VIj0HjdgRNXB3KAitJ2
f7e30EXVuAO+yLEVnV1Fn9GolwvRkyjJ/atfZDsGt5QmJRA9mdPiA4k2Fy8ZHt0knWL7ac2HIul/
mjqSG4ShbquVWNGBM6vt9JalINGfIWA+nCpeFMMZYMWnOOR1YDNAdHLFbsrKgTlsleVouVDRv6Dk
BuIk3mIb/p6lRdF5EOoVcOMRgmOp2POSPJAb0gJR6i/B6KrVVsB+JnuW1CewQEINoGzLmWt2o0z5
EhiIqnbcJptvOhyEKiXCEWSdjsPORe4C0AK6XYzltgoy+f+GC9nFKYLWpNrAbeUK24xE95AyypYb
3T2fMAnC5lHPchaot8Fpe7vCqhy1uQmKnRUjFPSLCGi4lhI6rWYC/vetq+5ckro5RbxtQf4Oh+g5
N3XTycZ4WabRXXQKGa7u7pWgXVZSMJL0zl3KIYBKbnJ5eh9Si6i5KFLIKeA00fmb8y3QjrRhBizo
PDPXTN10NNYFNVB6IpUBfRrVf0v6P9jB8QqkJDzebjxSE4Rk5sKgji7d5ziLFbg55uHfOZ8fJsLC
W6W3RcN7mcvFDyucG9GfC+4JUduqnkD/O+apubh+0tCJa1wvBkj5djvocb/4QBIEJo9EzGyMRQgu
gJHFzZh0EXq/mnqordYRgeaTCc2TY5aAslEYk36OSrJG/PUlVS8UUW4RWsrQ8K/Q1nAQKtRGyL/S
4D3VsG3LA9nYkIobbo4L0L5uWkOsr8QJPVq0XeLecJAHjrXWA/1XUs28hrEKo4VGhh97Ku49JkEJ
nYFP9fv6XSyfaQIngs5/dkdBHz2qq1OrRHBY+kW3AI2+SURjMxwMqF1FJCNaUdcTpS4Vh/mIlqoq
ofSNCcUn38kHZX0A56ScldJG7NxNP0dKlR2Lwilx6RGhA/0ZdtH0dJWLxtGNFUaMI1rNbh5krKuj
tDa7JP5Qn6WAUFMODBUiihZVeHZczNk6uz+CGxV6Def/isjfdBUBDgsCGbQU6mtFt4fef0fqwtvT
j7hf2gUte9AxM+7/LUGoebJ8DdgDRIIS+Ph1b+xUXMHA4MTq1CIS6YZ4FrEYKVVhEhoLtkhHprQK
lrAOgZJFIc5N8uPrT5XfX46x8qwO13wSFAUyWPUfEcviDsQZ7OE3r78AAgZ5ydAgSzFqvGc3+fIU
Uu5ixpcrxJ4KOR3+SXmLz5TazdRDT9bYgYQPRjgYoLvHbEC3OdSNQ5Rzj+OhlKv6dSOa4IluCv4T
HYA3WVcAjm3bghpI5Ag41v9Cxc94ypH559fdmKPVslkjsRjaq4hLnAhEzulUhamErG6uiEQk4ysH
8gzUzJemMVsM/BZeto1gkIpLJJ4bw0uS2WwT+Om+Op1bpjisroW12pq5fDEJCOx7EVHZ1u3ot/vH
HVTGIQm2GcomNPqzDjEP6IPhuMhNumz1bccde/z40eMT4zB64xC2BCKQLQOfyoYCzXZRokgmOIwL
SAs7Nwxa/TFyJTRmVg9WyiqSKPVqc9FqCjMKV1WpVJ9FhZq049xmKrO5/1bCnbvCnnBm7v/trdX0
1dKiJnhSh1reYGAil5eCI3btK8NYa105zUZ3wTVppKF/hE5ec9bjwdtBTcvj12Fomls0fRfMbUw3
95gj/bWqDLGhY3eUeleSkUKJ6l+kZZGgQaXeq8QF3qCPVrLM53Y2OW2Ug1rAkLTPMoJDeSysai0r
C+9+OTyHjCu1fm6490M7UsCb9h3a2yg66AJA+bunqiurFVSkwB2EuRVOGq6QY/zoQb0MFW6rx95U
iORFi6Hwi4aPD18DqhQT6rcdA0o3pdjLm7JXYquF/zRRmRHVNxw0C1FCjSzEDIf9vxShBtcdMoD6
esEgCQwqn0NOSVDV2OCXfHpa0jlL82pWEhipd0zb1IF5pnVWmCsYilbiZBISPF8W7+rII8xd9VhX
aOnbC470R6PvnulYvr6gVzbxZmEyNPXQqVz3gEh1pj1qIksjhEZNF2ITnrQbvONunFhUprpxWRee
Yn2AxZTmbxQRL27UOgkKPg0R7PCHr3QU1trNf5eloywV7Oi2XVZBBBDbjpRwuTobFQWerckzeDxH
s4KQpAYCK7/KqDqerMe+ZZee/gkXBru+pJtina/BWrWF++4MGinSCg21kL2wufkg8mEBbFW0NJju
Nz3r520DQhw661pgq8frqWL3uVHK74bZYeNmrPXGRSkm9O16jB4RO7lIfw/3T7oFgE16Cv3G2kyw
O0Tfaay76cVFlNJUgUxvNMQ5+WNaxfWZTw1bwtfR1vcURN7U8TNVDjqJ6af1L+2MLbbF9CM1krYN
i1hWLOQGO8/XXqr6x5VgCgYaNbvzdza3bHYqf0rdd+HpCTOuhBdVZlSJxUp/LFOgqxr9egpOitJh
7D7rdSy+u12M3LT7+vEAPuB0rnloaCroqXiP17lz6wdap9mzN4XKFHtt/bOSv5EJ9HIJE7IZjtUv
+Ok8GgwMj9oSJ2407BzPg+uQbnrPHKjw+BFfarBBzUNmz66W/q6UKaAPebrRruc82v4ohU6BGci/
TX52/lakcFKqwwr/rGGB9/agsNkvuXRp5PNdfWy0XhNw5J0Jxi5WNSS24FL8luyJrQpGczNhInsf
Uh5bPLhxty9jwrQ46dvXUto1yYoxuz91PJUwsCYelP1eCYF9fKBWQpXFZkfG6Y5detsmdFT7q0g6
HZZWdOg37FIeevRoxcLpRTd3jqJ+h1JpKwKeiI7UUs1o7gJJlFZAj9cHpTswpXzVKmO/qlWCqgNZ
DyevXS9/Y/aA9W//FyoHt9ejA3aSdv7QqebdXLoyxHFZ6Ta62+FXV+ikDFwPKsBwPoor8j+I45kV
qkRBV4IBjG7kxcDNUK47JjYKPzHn1OL7tLGlFgU6A/vKh7SkOxakEM99m9XSsefdEMdVcuhu/sbd
/KyvuhZGNGs7/j3JR9OAwM17EkSByOgg+4oWpTuUmF+I8Lp9hyZy1ml2vFywcfvzSiCVhGVX6np9
6WFC4D+irMMXDxRCd8nG4bSuTns5dOujI4qDZU0ohcFdLVPAnnxxW3KkRallFc38Cb7Zo2h0/fyf
6Cpc1NV/i/GoezSprzFawjAEKMdDk+XOFTI1/I2T2WhjBQWHj5wkkHeDpfZy7fYY9GRJ6iBVPL0L
lKbAlpws6qXkkH4Tn2QIl4iN0Hb64X0ZzHwVyptmopU740dQcCsiyaG/JdrRaaV22mdreUJh2kGh
lqpYAbPLrt42F8oCrAg5AL7+f7ZW0iMceFKm4jtnbJEaMTvCC83DvcuOlJGBp5xUdX1n22Fwm4RJ
OQDo5Q8qlOMnCbvqkjT7ZyIJZO4t0mKa/PGrdaD9ZmtdZIsbGrsVHM4/wk36K8K7QTnFFZYU4Fwl
mfWsWq1aaBJRgkLFmhDo1vKLGQJ3KZh6sj8OV4F+rJRE/zjC09KGwqvD1sq03Yn+uxx0hGQzC73u
EfiWsWB5SxpWPzqLeIU+yjpzUyVUMuyvmG+FHrY58xpvK1lH7FuZMtTPXE+vqJEpU5UNDdYp7fx8
IuScK/eXDOjLefKmKNs9LW1/adBfeA8CAHYXV6TlX+MgzMxQe7xYY0MjNw4mmk4t1ppwuUzSZ68n
t+5wn35fZiqJu9KPFTLa7kVWFBU9C4ALKF5PT9olUx01ZxBgoMf2w7YJWJXGuq9vspzQ2VrSQgbm
QqtAYfnldTB/EOUQXDHa3CQws2b2L9gbfaR8A+dFnaeLe+l8OMuGCYSmI4/HCupK+WpTVM/99ZFn
fwX42NbLcYKrLHNgXTQZ11U7uU0tXiPKRciLTAMr40950e7rW5UJ04+HFL+IdhONLMRZEX21X8Cn
G+Qh8dZv84QV4+7AynYrc987jSA5kqLHmw3yyNroHil9VdssbDbbXFgYQUDDQDFOqoDc80tdt1nm
pSX6y2x3b9ebkzRBlSHx1mU2F56EJwe2kczH5eWtgMWzboD3nnNQbGgAdOcs0//xAgyvx4pFS0RL
k6ZYtTJ3fiS1u6Qvkul70PdxPtoZWOmJXGf+kaJ1gpmsizHhDAYQN1LGhwoTsbphJ8iSzm4Qm9Bc
aoPPbA5Hf5bNqFdxP25XIklUBJtoZ5E6OYBU/m8geZwxRZe3jqSDIz0WNu9gmzlp9r0QxcFYH8wU
yChVtltGahg+SWhku8rpJOq++aBsNEIdu6ehrLjpB0IrzFyn4oaBw1OZbVWczjydOQ7nmrviPDfR
HVR2cieAJhz5Im2qkDjB1ykl5t0sSOb7Hze9BnGy9EHRp8HrQOrZRHLrXPB5fO8bdFZ4DaqUILRJ
tWifEtAGzfyNanJjCzaU/g47psFnVD8NtfsQskewoFkpKK8OhYYGfGomJYLgbfyy38Z1COBcPlSJ
KOdLjbx6QmgYZUJegFOh756WD5jzmkZd0w04T4g2GXRlZ5Btt6JF11zF5afYtALsTbWMxfcTeb9J
Q9pFCcqKqfRwyNJznxI4OR262tf7ypoRgae6P4tvuHIFJPgmJkCmn9MIi9rJ1rwEj3LNUbeU9Ecc
VnCTY+PjLfzlNJOJsP9VWF/YjPuoKJv/JEvHWBfvM3Wy0mD/4EVrkzOYQIe3JxbLfwFbR8kDAYJL
xkgRJX0OeEfcKps2FDGpfuxDHz/yyBV64/tTk7WzyjNMbIufvj58sbPvS8uwwEMBslDNCI/utHIM
BIt8vto3LiFA66oKdpG31rEpsjD2/hOmZlMkl7xrvavTQffmBaAvvEfu7d5KrJb0HiXNsd3o0oKX
ZCkIFln8wr6zZIlwxDOuJcaVNkvV+PXCb8LGKljcZ3CU7t+qAPaBKIxZlolLBMurt0vcER2ZSaTj
VnojwSi6YWDkT5xtaVLtliIYWtns1rHFsktqBu7RB9vOW7/b7IYT5GSxZawjRBL+q8B8lTU4a8+q
+Ad7FUfYgNTR5vyjUmcSFphCO4Tb2CfOLQN0a50btCTLBboC6lWdUQ9tB5Cpo/POQR61jguSXs7f
4MRD3NSXIj2Gp0tifpTdQQ/tl4A2fi1FnoXqWsi9d5f2HbSzPIxPZzs/EccXxYMZvs5F6Fl7iI1C
UGOpbhMS5b3MU5cKkN8v766aHvcYrt6xqZhYnxKRtkApDh1po/zGkvMHlXGgC907vnA4UQHTHGkN
xGiTuKsmpEdjvXzD9JIViUR8kb7RrhrQKxvjku9WWyROaLXqV88aB9Blm8mVAyia6RRi+q4hXzL3
K2IXB56j2o5TwMqZL5m1jitNRuTKCEMzKSAc9WpE3mYTsNJqwVyiYFjpUwDo/bsHJMiO1Qe6umy7
PdxwWkmRP/sk14SHLO4ryFtIHfmPeoulaHLJKQPW52lfOCkJdsQZXX1CovefeEvFvXHqYHwP9o6u
oxiH1eJXJQ6toepnH3VWcY08lcznv30ZokOmRNlyDdndzowdA4Ndw4OYe3UDON0c5cgzoc3is9gG
LIoaxWRCumWp+jc4ZB0lBquWzDlvIxygUl1j7qfHiwKFPYd4MKNwWvC27A/jvUzcHE4FAuSheycN
UNRgs3R3kFgw/3S7BFLc1AZGOpnijVnXIaldgKL8iXiatOMrMLY9GGi18Fh2D6AauDikDDAaBviA
rWyDRJXmnV8bjyxCFIipa4lb7+pU/7rOtXPs5fNn4xcjMrcQBtQgMHWL7a08L9jSNNCeGyT8IL+6
gNEOEkH4KHCOdAZKqOKldYlPE/Yh9WwD6F6jxfYMSoEsBQbTIGa79exXjvP4VA5FnD6IMl1WYCUL
lmFWNFRlMhX9vL8GaP/tLAxzFhfRBMgxqv0avA658jjr4YE95pxvNUtIPSwLUoPOZdaxJlnBh/8T
0eaWKfTYlIMb5XOgvTi5lcyL7dAoIMhqRskLbYsDoELygi/VoGa01bwdFEmq5qx0dMvZNZBwnLPX
mttVYhWc1ZAHQ/25NrOW/gBqzc4AkerFMFFXWeDQOQd/JXECOVXgez1qCt//zAwt3fOB7FfVYc3c
LiRjKdrqhkHD8AptMqJQbE2fp0XMg8UVHadkBb1WzZ3ypReW2trFL3Et1VdfALUECbqGm1nYtlTH
AacvYtXKO0FAQKTpmx4+rgE1DEhr6oKHjDm4fhwZfcmo2nqFRxwwtw35IxYArtop3wVzZ9MelFMb
iSEnBoSZfvDSTYlJnvkX5sQifT6yqLTpqYFhsVXHgiqQz/LTy2+AQnEY2Xpv9bIvetWGHpBDHr3Y
VAGeAX8CqYAhgK1J88aJ/kyhZaZauJmzxaag7oxqDqi4twrswCshS5sUw+H1/GhY3kC8a5R/aiTs
ktcmVZeWuYCj10HCuj0W7g+mmfprmEFh746KlI8nZHqZBBAMsku1JSCSo84hY5gSf03T5Nekb0b1
aFv72lHAXDVh7SROnfVp/HerD4V55Ww6i6Y7b2LSmTNoehvNJ+SLQvDDtbGHuWyVjtICUCbyDFCx
SCXos3xdZl3j5KogkUBdEZxKjFfR3zyk9/rCkW7ilUserdVq9/jB6ximd6n3ebhY3X29i/Pshqqg
rbijwDw+bYX9+aC5YFAr0joSbBLXBdRE8eKJf54T3ym0s67nIi0CgidaGQp3N7bIYIkx6IhzDTGY
Vkr4esDpoWMRPkEsxVyKNuZjhO4+aWFKNX1zCRsRFln0Q9NJtgVeHwGNQaFb8w11OGxIEoYmgYIs
yT0kDLNmmPLhXXqWRVV2ysEp+Afappwi9xWIiltOclAoj4g74hgxAglb/yLLnRRZJ4JMF/CqB8Nl
WnBSwaAAEXuerRB1kAgFPSrdG7gA93w6/x5UCqgrLgewPojZhz1QS+FOtru/a7Ga37iLtPfz1ALt
kOSjXyY4G4KqITW02YJDsNL7f2R3P8lc9M9/29R2E7whBoqE5+xq/vvYcTMv1x2/uqohG4TYDVGe
bBIlcScmyRCioasLwnyIBUSBIs/iQ+BeaLJ/AdhSB05PKOYS7wqs8gOdyTVkojvGVE7+pJB7sRXr
LTXSCnfO15HVFWDE7pLPK1CTeOPKFeJxVYf8370H49a+qDuQ70cf4ddOJ7O+IjoKimyU9tRQjCq2
k+IOsHAwA3xbR7A6tzgV/tsYgcqYr2M2fdL1SQSl9IOmY5U5p3Y1v3iABGw+8Cl1aHzjaghgf4L2
ZGdM9MIeD+S9xqmnaq7Q4Qb1rhSss6RJJvxaLq3cFw0vOlmbIRKk5rlM1dPR8WmjJd68mg+WaStL
EIkJXSDGH/4ojo1MYNYA1+jzPaZhMCLHM+PxTL8mrD5cMB6AhFYbUbkH1YlUnLWgJ5jzVTsGRrfq
nCzsjBDt0HQpHQoQoomZQPj9JA3taIB4SR1UvZh+55/aNWF18nD27aTueTdniM/b7qkwnPdiTw7N
zcAA1F4zUCFKV9XrBVLelHboUsjOkR5/b7zLxZ3iukQuvcwCfB7eIvHthDSxMgeWlzDSpB6DpnP4
jAihuG+4OoWbf8ElfYNQJvysYBiuF6BIFMYyt/N7l5MhsLZ1peGu79xbigJzceg+bPhYBSJvZjSV
lKCf37alGkDsQXzQlC3z+8xHkf7bFsX7x92QV8C24NzfhKk/KiYDLGsl0t25ZnFFPED+VDF8uoKj
igB6lFDugqArtHGTmZ2OVQZ2Gf4S65TjZtWVFogIntCyYQKONJgo0VDSLuIu5IQZr4nOPJr/oi7W
fTmzpudr/lo3W0+pO6kREYkFl9cx6oZXhp1puBMl7rciqhdJPEPRnLoCLMUeis0Pq9WZnyX+xn4T
pDZmYGMCBTrqmcRHVBStkb5YqFWetv5J5fhqH6P0zUaip1humxSNA3R+yYq8A7wOxJ6qSZcP1E17
Ed4RCd5CJmJY3zzBj1sFD32g4EjjXlihaBJ00EonR5sCMMWGRLUH2QrsoJJK9xktcSmT4eo3oMD0
3zJ89kF+PDd627eRxLjKILzmM2BI6odAuBfmAY66gtWKd6u/fflHrrE7Y5U5XuH2rCcRrXvu6Z8V
AWoB9F0SmzblgaPiazYt7zO7f0aaFx9OwVBI8geVQYlJV58ZIQHhZugGyoqAQ3SaY59FFRHr2iHV
0iZaErw+ow1R87swom79i3LtV40V7pWFak+mB4S38smKUZzn8nI/C6u4NWIiTgk9AtASft/XFAob
/jEjR9DyBHZXL4xoGJFVHZdy5griEPLH4xuAhZAVH0S8K96qEzbhStPyGhoIZPg8/+70FDtk8akP
3tWReQE1Zs00KDhVy7Q0bTLu1EikIMtM/44MeIaMnuSsLI8r5Tg9TgMWAztexOvHjTqiy9Ts0IxY
CVWHUeLchbMkRSv8dpw0mGxfL/oF036pe7ZAEKU/n9RY1GxKRuE0pEnX3stUon2wEX51JhMqLULy
8Gckij6VtEW66OuTawD7+wGEgmUy79EqGmHUKn9IpoSDRKoMEdQ1vItPX9SWH+6J0c46CMDynGQP
xDGdCDYrZOyGYfEIku78WDVYPYQNg5Yvt/kaagVy4+G6TL10jLRt8vNV/0Snf3L8D26Oc5CReaNm
/JNGh0vuSA/6pkQSbk7RdEkxN0peqZY3ySnw22CU5VZl7MGZzAMdaq6DUbFH/ke/WVKpIM74/4SQ
kk0bf1SbHzCmGIQNzhK5EwBqhaWAg/Doj9RByUYAfkamN5UOK3VG8R3/p61a3yFVeIDq1BkxAEgY
lESQaEHBUAX/syBZCmDijbCE8ZczICFiluhWc/xkYpBZgaRIQm9X02niGU2l0I7vKedMGzo/FDF3
l0Sl+lEPpLOftTypvM1VdwJrD+ONPaKJKDj94GKPGCEP/vN7wTvyk2EWe4Q2JHG3WoLoJ4p2019T
ubOVumiUlJLSHQIC4pJphTdp8uOgaMkfMkILSkpanQFNkUd20LZBFM7O7AhnDw42tMieZdbhy+iS
ay6ohU66i0WAfcpKzCux6ES1lXAIjaicNzsTRMEET+aispPIsuNlN2kYqgSMYVZaPCVRzlChoetr
oekARgPMyxfpy7/Mx04jJt6BgPfsLVEhsv+0xsf7X60wO9+OLayYEZjsMj+4chC0WZCAX24JXXve
FnYDTKRDueETLxDIBXrfknkTqQlJv/9infG16nW9cZP/qkZ5uece/7CxguEvxibE5t1d67HXoJHD
gPKLknuRte90PqRHzFV8M6GFkWNAuT4sUg5GjdcMIXZuhwF1wXV4SpYRgyMRtI3f4QJRUiT6rc1F
0SlX6GdWnHM9IubTgJziLs8d14FvgdgmZ2xdGRt0zSSnzazI5/I8ppopkdep8CuL2WwxSL8PeSOL
k5YkaeqjNc9ZEKBQVNuYlMLp8veNFDyquj7ouVwwbHSzQn0xmdAhKrgyaMGMtNJjskZkREvemdd8
B2ZTPhzgLYvqUkJ/EO10YQiO5jkdecPLSfEUhbRu0wAYl0k3SKUlXESLDGfgknU7VBI5NeqDu+0y
2syFSIUGbOpMEnLydXqBg1nQvxha3oMCguOuL69anCQ/fNk+tgzV8ZURSOaCaYxp3ZNok7kQ+TM2
4YLKO0lhqBKKW8411YeNulqNZ+1P/GtlnRtUhBe7zqv2AKB4BPU+V9qSnyv6jkIekqvcSFyIuamc
vNp6zzxr29PunNT5jMJmfkFK87ivx43+RpEPSl3aMdjjkeiN5FhgF9z2LHCupGVyRGyrnEBM6gqV
6WlEu6oYcrMonfBNFRx+xC26yKZat7n0Oef651oLesGClCTDNNTdCsbJd+q6VqwnmKHkunosfqLm
9QO4mO0ioI8tV1mABfS+0OOUI9G1s9NoYrsnNDAZyl9Txhxw7OwmgpIpkNhI/03Zs6YfNxvhB7Rd
apo0u9sfk/nHStMPAA7QrKMUepHigPVNExJy3COMat8gRZN50k8nlk29Z/bBiLqeAZHZetRJx1qk
wZY2asAdFbUUhKUh8sS9EjnmU84Jk7l53IJAOP5/QIcRo/cy02b2btgI+TYkRSD3AI6ASOcJxdvu
6+RCoDcnoRqwtz4rqv5IFUisSIJgm83l/CBQ/L1pONhDVdA8IE6h1UaU+tCDY7XA3iCcDFmCOiGe
khU2WBCJKDxI+wsKZNeUBDEFfeJzTIk9UEAyBVMXsGaoAXIS4ThaW5okrcJk6e9EYWHmu52xqL8n
+l/vSRxdrI0aLz2GknoXIYwzPYqUnzX97is95ZaqBM0L5r0123NnCq+nPEBTr6uZprco52f7Ekwo
IpJ5w0eRH3e5uGYcNslTDgWLWeYXQbKOyRfGhBIMTsILMpWR3LhY7X4H6HE8lw5OAk+tsdBuZJNg
Hqul8VtC6lIQXvmgxnZjJFb3SA6PRcXdiib/XJdsEDN6UUgxWtTury9h6xUlZl8eKCjRzmHzJYfo
F+QlwwKaddF7/Dayd26TeMfDBOciNvEbzWBiMLcc6I+z8pFGVG7rkuZewUVQkXeTISjZz5sg3su+
kGKMVl94s/QR1QMOHJ2eY6Tqk6VdLckyQxeyd83Kr/riIFwZErrpFpM8qJAi1HdSzlIlF01MV//D
RdiwCys5MO/rxU0eTalEnjQoaY3wiOh0DRCHs7PTjiHaiGHoeP3A/PXNFPrsyhcqC5UrUXue4/0j
icXZqzUVTsPlk/D5RUWdiPOckEZh7uRdqDVv79TawMy8AunMYA88MnkxQgJ12REPFtswcaiyYTt6
n9AeVAYAcs5IaDU5uO02Dv9Yt/Z0UNiV5qQAI+jGb3oNFsGBVEy/+l63Gkvk7oJKhAt7hfZscULy
c/wrDLc6PS3rJFTTHQuq/tjCP6UTaBNRUrwEsLYH/ErpXwZW2vgm+rCtegxgf0eW6Ckhl1tcey7e
/56gGioRE6TcyRyeNyfaF48C9okJwnk7xC6Q8IY6ycr/Aw+QI6tzUxPPGy9Q3QcEwfg0MF8xEdZq
7/nsVA+V+jEhwbKFcBhfW/HuiqNQwbOn/l/45ZZwF6TQtIpZWUg0UNsynHlCwFXWWunQANO3W+Qp
TuI2rAbiAhyMNvUl+Epp0+7r00xW0eMMpmPbkCEI8S6V+QnTdcu2TpgaxxTrLdmpTCbXG+1rFEqG
XRxM+ksZKtTFSLk35+mi4OtLYxMBAUCQFnajHtMajb36ANJENQI1S9Pc2H+zjx3w+3UbbBF7wz0A
yc7fIAKqUGFwGp2nbWu+DhUby/Yt78YNRm78/VZxYcn2wVLyUXCdgz5H9J8MzPPkSttUFAm2yoqm
iHlYrhlIBfGavgGppWgyBByVkEsg8QlknSiSzimS6jP2rnmbSuBu4cYGATMejPAHCY3ctH3OFlj2
YqIg7jt+dO+8elEAuv9kLmpIiIoPELIdCWKbY16fBpnkY2XJKyzzT7Qvo0k+Hagyem8UjN3HVMoL
dz22vYZZABTUqOuaQYGlmHm7Z3jwcxovHvOyTfaQjIiUCdxVcGlnuxnGUmJN51O0cSBG0w3u73XA
kRzCvNXdYcdUf6ACqZWHsz1V3ZVZj+JaLOrLZQAMLXfpUjfHtxJ7lCq+gE0MEWv6/ivo+TdQ47V8
ZiMmFSU8cQ+wzrW+lOIvH12ZEAZPP2KnFR5P8niBHbGOWTCkzQBaqNskCE55J8SZ7HiaCaxC3lIc
fcsvvNQdlU5DXzJnknMozxBGkREv2MFlf2Rle+MgCf4VPNRh0URT7MDSKFtOVQHzKDVqU7ei8cL8
ygNTN9a4+03fC+WXht9emqHoyPcDwBCcPqJMLks5ZTje7Ztr3aHfC1ECHCucufHE0B66f0ntjkxE
ECYhe3efSl2gZp1GGy0qoF+jKthnp4Um+KEyDJf+xdpslqMTngR8jD9VXVSolXsbtI2EW12yPavo
t9tQ+JY9+jGs1Hfeqfvl/qS0C9OAOnxBuD54i4geAWxLKTa895mM5x7LmY1bJzy+wOgRwrFnQInx
QZD6tWcdTnsuuw1/GIPauY0wXtlHoyakilCjn5+Jmdqm0Uhk76zxtx6xa/8Ki6NvhEnwDLl3nfJF
KVFiZG+lLIsPHUyvRZUl3oGd83TXr/IQJMCpTafVL6SW67OwcimYKwStbozX05vuQpn2Hs+U9arR
W/mQsPTthKD75/0TonarCLGPwfcD5+9OS+Eta9kY391so7Ppq/3KaqeUrtUWmuwonAsnOOseFwiL
RpDFp1QtBnqRWnRb3RQhCowTvkKrwU0UV+CufIFOTjyjSBjirZXsiGIffQvLv10mWuKtCLppIiZi
hWzHWoJ7IO/7+W7GBwXUdNJz8vhudp+Ki8BV+WDjFowHs5GStiE8W/evxMr6elIw9Y97g+/mDW8o
3WfYPYTJS8Q0uYe5lzyhc8telYfRgr3bohTAeewGCFcQNfcGx1XpnVNs5khzVkqQl59aUbZYnMw5
JzsW/if4LGsSLx8JJc3QmQYo/yRol4yKuADN040qajgplfKfgzC/bBLcsNRiJu65t/bohrcXLrlo
dNGF8R/tcxZO1pM21WA4ykzl6W4gRX27560huolwB2BYsNIY9D+WpK5Kg8FG6gNUtlVhglHqkqze
ieObC+6+k/I8SxgciBXvtyau3qxmIn1asbZPGPSBVXk/N5eVLh2efGORJ+OwZt0mzsK81LxIBMSs
GdeL3phclQOq4lDkMlOITyb/bLOV5bVm44WxUPNTS5MkzTl2k9fktXSNGu2nBPdMIqBcLPX8uVBx
kB2lTccE3hCxA5GfboE16MF0d8p9ULaoj3vjTA3E5umY41Im1R3lQweuVPB8QJIJSwGJel/6dBti
f2wFuRAxUVbU4NlWhnLLsu8w9FEi3F3bNVTkW3c29N7pKJwyuvzHibJfMZVoV962wZ+ucoKEL/Er
fn99W8DtCAGM6lL2SsWJp5V+wa5aYouiJGBumLVr8fgHwqdcC2TxFE7qGAiw9bp8O5S18nylgcSZ
9dOh4X+uH7X7eZo8HWxaywbNy+KLZuHXIcJMACNcYe+Zf6btVu80DwLgZjeOMF8Q/QpG1LFDDjpM
PCjvlAK7DaAVXC5tqXaA6CdAr/5DF4yZUk8xF7aAF3hBaL+6f7iFG8oeDR1Odj1ZB0C3zsJU4Xn0
9/NsFt0PLZPTG6ZM8louzH72iuNowEnvNN4iRcKd+8kI+rBZBcglYZbJZnug5KZ6RQoHYO4r4GiF
5YtTfIf7xfFnRNywt6g+BCSa9zl1SeTk2z9eBjaHkUbLrA5hBPisuMqh7mH2y7p518ehNh7g93Nf
BSORj5UHruOoxlb5s+RJmdCpcIw5aEIevGmHz2UCTjSwK98nGEA+OuLds3PImoSccLFujqtXnGG8
NuxcwxxAEDfsQsf7NeVEYH+h2+hiaEcLR+mGbtzdYGI0WLV3fGaS0d8pjE8X5VkkcQxcEBhti0Rk
VEh9Q0SK3NHFQyiaA8y9vF1Z1JvdHIAHsSizbZz6p2HMLfnqQ0DzYw46ySBQzZY0qpSoqYuJ8Vjz
NDNfMDePq4cmYueQ7khV78lsggBDz/31QDyPVilmHG9rPCi/11FF0UMjTPyPnTJlIIykcGYG1toy
I+8ZwN6F9TrE3WWnlPV/XmGzxaZ2nwK/ILJdNTxLa9i2YWPb4NtMeiG/oiwpoet7JNvkKgwVMYV6
OMld/7Fu+w212XKGtiDBJnwxFGzlwGXbGJwc6vCWjEjV7iPVRRTC3dftVCqo0t2/d0BMMOab+voT
CA220eGrOPTSAVCVhfYewjcO9v4ekOZ/HcvZuFAFDkBRnqMP/xJFofKRlOGHFOY7wPbY2P/3AaCC
OwyTjga9jNixn2Yq6/NzrKG1h6of32k/2PWW5DsJqqwz+iCFiw6Rfti8LhzM0vzv+vJnMChH6xVq
jvtWvzQcwa/6bvbL10mkpiSR6uVQJq2EuuJj6wUXoGPA1c2JYjP+ujhrzXd1lU3qWjaYQuzI8X0y
6x+cLo9Z+Cvxvm9RnfSys7k/0Gmfb93DWB/Z9phY5310ugU4hG3HBIWXVPmVnPn4gBNzbFANzPBK
Qw8N6VI9rnz6yEtNk7W/aAaGyNLxbHhRpigT/lUMBQIhxYjyyJb8vYd6Q23ZephIuyi9fF1a84ZE
mMkvK0L+vdJy2ONEoADXkqQERa6RGxUGylxgTKzlf8C/Gof7WohepZnqYOYHBJoosmMk4ZOQdaB1
TlXkop0AucVJCDbPRfrSm07jRijtcCeQQv751bDC+buuMJ9a7YQlqy54qmJBNunMWkvm94r7N98K
uZPWJPCwC5VhuS9up9FyhB0jqvGt/sDn2dWhFSLfwvxTq/m2LFprY8bbR+PDhUyD0sT2KS9Wa4Rj
BWgRS01qU4jmtKG5tG41KXASLCQmMY7fCGvihdRpA86wGj039oIwS1CTSCFiPYISbloZfNWcStsF
9ybuSo/2OTynY6YDuu3/AZ2E/SgCijufnsl/EbVaG65VZ7NNBTvYhBSqAXcTfmpN/Ux0Du9X7q64
nOKW6oUy6nfimKrM5y7Hr6TZoXjItMEf9KW3SmJMSd2nWqtwBwJdCAbmUBroWvkYo9g0sdn/4iEF
PxTrAtAHYhIkk4ob7S8eBoLM5Xt4T2tnEdMBrUoAbA5QfSlzvYJdzBwhDXFt67Hd4bDAIO5kPeC5
oY2xIsIg7Vk4DgqMdt8OTe+CQe2ntN/h62ACEBkmnfhu3gJcXDLKGxegJYAaH33DayJHw63DIAtQ
S6YNv9ouBRngXe3SxR65BwBRES0KkmHU2LNGPIk1v1E3m7OdC0f7rm2ELKPaQv10Wvn483hrxJE4
klcN0z0UTOCDEGBGlPST/1h02bV9qHOnl8szy5Vp3JXIdXIa7H7i1Kp1GC/oogtWoJ93Twq7Dwal
UTOI9NFQDEbdPwvQyjJ4KTQnmnFqdIMJZH7hSqmsGu6RurYHu+Ns2n0ROcmBbAwa9OgPuqRPYPa1
H72/O8DJf8N7Pfj2S13halV9ZgpPkhoKYezE/DZPcXj/NpGbiEiibPi4ObqJx7GYHE1gf+9UB9VX
CXwOqM3TztUu5zD6iRoDfQoCPsBjdUb0P4q1nz3H7Q3/RT59rn9JnqPy3PJmYSJH/JsmMdPDfuya
eeb8ON+OZEzYbFBWdOqobuxNw4qZegI4ezQnJdLM3wBoj7wAd9Qcv7GiFyVTa/kWjwEdhjVEwGhB
C1GjP69qxWTzJevpVjxDA8w3k03lC1zGQ8SsbNESZH9uVNFXSXI5Kjgit/8mjWVs8RIVe9feCnlp
waQNTuZTr2OV6chw2oWxZisIGlGRrutp2h0JEOrl0Owsa1cWj8NsMcZmHitL108efbqE14O948zl
5fGhObimS+q8YxjCkwUcTb0Z28beeyK5NwlSoogt6n0N92G79NuZH3roE17cI36FCbXlR/Jgjs7n
YCIfrZcWb0Pm/s6mzjSyGMX5bwcpABaK6qZcJO9Z06kkTu0zw0olX1WmTvzyYvyKhAfYotj9rnAJ
p0tA8V6pdTlm23HHb7XlovINvJH5icooBlE4+Z+Y0cZZQvBkmz96ON5nYvUyqAAYVRs2sQgBOjpg
4A+MbSU6yJFNjBXLE7GP0dummtl0pDfNiRtt8vBoZdL8Km7MYzL37IxnN01WsftCJGz1iOsSvINy
5dHRrJWsUzwQViiEoC6nZDMny+/M/W8O+cZYGh8wHu0VBReSu06XUDOuNaeXKGXG/CkR5IEZxo9l
82Quw4/gfijciCsgj1pO4hotJS/QiqCUhHxoxoBDti7FNmLGBFHXhmZk5caa0b1+a2qfOdzTyMGv
2DE3TEzW3IcV8haoG2krNm9VSPgl8qtbxXRBi01uf4upvgqEviPcJRZx6Sg/8hrOhywclhJ3ZFw2
qyZerwFutrrCn8V5sC924L/Thv/4FZv8UF/0HN3pC+n0/nRcSSPLYg6SnbUr2WJmcywJsXW3AkNL
S88fOg1hybxY9HYlZiNjr1vnn6i/7TMps6rZEPqWEsHpxP/bJR2iM2R0bb+fEAQLC2sikz9uEKw0
qjtBwgwHfIYX93QbaFBs4DvDZXlnoqqXHXxHgn9z7rNRfkH4acV5SMP259w7C9XP7RU/whgxrgzN
zZDg2stVzNkGz7vy6F87nS4O/FqbvdNP5r4SwcQZAaOCxl4G6xBngAvzAN2DHBbyO4TAAIY4cKbO
cPWS5O6Z0ejAdrZvSy6+jWd+wMgh5jAR3iUdBTGlrK7e2iMpk+m0WOs42kSrL/PdkT3B++xDMGY5
kW8/l2NwQ8764UgfAmN08jOe4kp0sInrK9mv+/+T/PY505OzMvymKS1YQXGyoBgGXlL6zONegSl8
yuCTVSLfk7Opr8ICl3s+SFoeHkRYu7tw04B7pCoRmpPWNRY6uMLhdUn3Xg8h2UsHkdCCZLwbDvsv
moVNbOqNyKxPOtAzOPXfDfUffLCzSfXhjQXukNCQa+XJnkz9runl0T6uKMXVEFzjUcOHC7lb17pm
lfHUbyTmv42Su3EcIOzQYtXaqqumIbRWwqcoo4fOdY6xDJx2i/r3ai0dNm8+B6FlWSG1fyoXvid/
GwZw5d+sw7vVLx1YBf8ZlDFHekdXxg3jBI+gcmChGNI7EHj2xlRWseGRLZn93W3000cwn4eWd68s
BxBjFyPSBd3AouQhinpmrB2/xgLOkzE1VxxcL9W5o4SMVCqjLcUXX8F15gH/SRkEIM+mcHx3dlik
SyXhi+WbhWyw/R5lhrfuTe7mGMBQMJI7KoYRjNkCnlPAlwaYAbSNK+YGPXe3NkgTxx845p4O2JOL
n8qpzSLwzXdJQENb1JDHM8jL2aZLGTexyqHZy5mKd2Tjj8McDx5h8HqlUR45ssGUBb20o0J+tTl7
x7l29bl3CdzlFvfA4NfQT3IRXfunuPcVlRFXFnDCrgfkPeu7zzx3CRt8878KKbfoacj4yYOGON9T
8GEjlT7XJ4quIV0bj6EaB0svboo34RKbc+wec6UGuiqJVWmSNVDc22chIeFK6OP1M6ymYkFmfqHn
NTI66t2cGzlD1LpZmVbj7HfCLxl2QUq8nv1Fo/WgyuYuSylYNM7vLWgUeuZ23alNlKGhI4FhvMOU
SP8SjOmcJogSh5t2l1ED50LPJRdrBZz6vv2ra3WshbyiakRl9b0HTbI+tDo0PbXlcemCM5K8k0I7
c5e8p48yNkqEZnmG5VVVXA1yu+jOyRUdSwGNxZq4021nzEI93xARuXgggJY68w3Bb86e3SpuiGoC
t6mLY8Y8I8SoGTXeYL+c6JDokFWTNcr+OdkBeGvQgmHU55Qg38vB3ParFMc/RI7+pxynrhMGC8Lc
Ww2zs8sl//kRmWvh2iL3ZuftyhOcOsUN31C2Pl2zz56DsCB0lXR1ApzZ/ubGGPMfshWZXj9I3hNU
iUgd26K/BqeiA6JP3mmUWcGeyRU9ydFp1Yq6ivplKzCXqaKBd8G73DK//EYuzrKC+SpuIb6LiSNF
dehCwOr6mXHonkYc1sT2Ay9jfamHdS/9m9E8Z0FT76uVH6qZXO5FHFZJBm1JW3h29YLaO2E4cjGx
4O67HUSGw2Har+ug/aEmrMPrQAAopL7qdQji5J/qd2qTKilhGcFrkn7P8paB5B9ah5XM1CbTgdlZ
33t4M+5ONxLnFbMgNj3dD0jPwBlPMuDo8jJ0L7DhNJVe8LZfdWua7MjGrBJPa9rFX3ItSboTviMw
otDsb4NZqPM8UF5KH37HfwZ3evfhf8IQQKscuqP0CqVXa9ysIwbk6dA4q051WkkySkKkjK/Wbg00
/AqGYTLS/ffbhRXDkCgZy7wxOKXLWkEQ6x9uQAlGLP3S9m7xZ/WEXl3o6XO0lypiB9wi1U3tEW3A
F4xydVhdOt9U9rKloj4cgO+q0bK3LYnZwq9dCIkwzABT886MV/5TBwCJM9oGMw+9B3fPxL/1IqxJ
ejguehjqDNicw8SASjE8yMxKUgSd44vdf/0foi/3BSI45N32eQ9w90M0Bx8PP2fogdp189rTi4A2
+c+6Vg/vIseHvAj9ouINxKrOHh/DDLO6WVfT/FqR8rAUYMy8Yzyjy3Vdw3Pnm2u7771MJJO5r4Sc
SV7ChVcPuHyOaszYN06is5idXaKkEmR4c5abzatv0AYJr5D9ea9e0FQIf2DMnxK7Q7qLGEnQCB09
Eg0y0rs1GeOojmXuJol4dz0pWTmM+HWE/MyGovpUt7SPkFn+d3Ret5Ud08ITDEHds0niS7E4biJg
voi6/KwFocH56vMmR9h/EVDcISUrUF6EB1+S444uw3XERxvM/4eAXsZl+zQUG/KvOt4fLyNijPm3
ezfPeAiPenuygQbT2KFEl+6Z7ddx8aIsh0j8fa09aqKJo7Eqy+pe/b46+aLQFyzlPs3rxeNz9P3V
SzxZ1JG0hBwf0JkAhaKA8RdPTBWVAio/0vW+muWV/88WGVsQEGU6L8DOM/GUPj5O6Bu50rqI+5BM
LmZjSq9Yl5tBGsYKy0/ZDmhByjhP+Np+YSCB0TWmCQ2lw1B0Y3KKoWpyLnzahxPLeB3pnzdlHcao
wEQ4o2M9syx1X+OlXl03t0QOdk426K2nBs/Lr13dvIh+pK3o+10I9u5sGo0mjqD+n34TpUFJHS12
782evjK3o7nuiorpdq8g3ffVUdwNSHgD+mEzo1IKCMc5T4UT9sDHCFeenOrLT4T8MafoRV23D6JO
4/Fbd02DltR0FJ9xeP3DvC/MQqz3Yko09nJWYAeg6KXksGL0nKHR7+CxK+bMSkskR6qyqrZ0T0QJ
R8AYP39GAFK2idDq7hgytAH6MddtnngwFXFQtHPji+LpXfdAlACyj/WdumgT4DDs4DvSLD5f0zFG
cI+WFUZ/e1EV6ySBgTDRfqKLoec6nqpkTCGSB7XVRTY3dnAia4G/47UkoQYfC78fFK71PPTBn0+F
66z304lADJ207uCn/lINI2KAjMSC1D4vBUo1+3t4qx9e3mUutQs/uITfgVpBFMavynJE4m+rEn2c
l/6/lk9tGyvAvlu6hjypmsW1Sr+eNKHx/sJZtO8LAn1+TISpzqHy2RmO1jXaUIWEJOxxGs7/OXs8
a3g93eNaRRa6/Ht6LK3DaP59BtO7qG0rhEzcxUf16/qbRopY3OXGO/xhFUYTxx4h4OK+Ik6+7NEW
cztcpzvYtubmcJhZb+II48MLDavZ0MGnRLRnv7rsscsOU6cxI4ATSLg6SgyuzgNvvQUtaNSdES69
aCMqXU2knqWohbsHmm6TB/+7RyPKPn92Ks+ZinN9cb/ZuLoWBOnvT+iw3x6sNuZuXMtKU8ojMsR/
0b16FZl8o1aRBjpZvaYHdI67w/VXFc8tjA3WKcxd6QuiSQU6u+qFweZH1llh0McC+DPxFLjDLL+G
teVoLw7FfyrBrVAYv2ZgQedDWrNt4afLmgTXXscY6Gac/cT3XGG5rFF910XTu0j+GOyBbsRFhaLL
eABpXg5yOeg21Cjltcicsc2KICjPCMiJeetSS2wMe6EUaI9hB7l+t3BiEckOI0GqpRcWysTawGu6
C8g+YZorIGF2yGFFfOEgxgx92ehyxyEicXpM0O/NRV75/s3pHhyHFKJwbXTzIyhbDFqjfy2aXezq
Z4BYpFrzN0Chjcz5hyL2CN4BRU91JmaroI4OlU8zK34vg/404BEI5UEvc/Vr2nwXZtRWKW3NxnC/
jGEEez2mZWUfqMJA8yJFRr9ctkVIQvkDPgeGBPQXf7zgHWvp7Hh2JX6Ge4Am4YJIJAmkN2F9ppFB
j1x2YSiuRg59fzGBJzzNV9YJE70XyMZav/4c3uIL9JnSo8CGbLhvA4TK/mwgmGFZ+7qgC9PJqkxY
tWg+MeMZndShMn9QNuMXlhmvxPqZrdzpQyBV+jabQfV1/s/Ewgf6RwkZ26wiDEK/khwit8/7psI4
YcXOi4rC4Pj9fQ494IZRzBy52oLDC5BDJ+4+d9kZOkC4s4Rm3j/tOYQvGz+iX92hFmuauag27SHS
bvM3TIwcATTEpQR228p4rnQLXT20uXPBpViX2xD5OEG4OTfKW+u/mqpsLB8FTL6zMOhQgDWG1wTG
phRJnY/mawBpTxyK2O3Wvv+vgnYGvWjfI//zDkH6umZ37pCUcVa5ckSStA7gqzc79KwHBwrxSQQV
bZ57mJMKdXoD4YcYJE+ZfjSNOviwIfdmjRlV/1m5RoYCvJ8jN3cZ3hqCXDR7tm9qel8dtNpaFE/m
ARmcpNdWaf2lOfFJDn2wO0eWGKDLq89IJP+XNCFVI4tr5b32jcrXqB9TF0cBzKXH6bipgFJTLyko
0P4TF7+CWC0OqM9iDBfEZeHtqi/BqojPXWnDDUTbXnUQyrduKJdlDcpj1BQawNc50hI6PtfrtAWh
kkVA4IglWi4OjNfjWSjJa4XajFtxO4yBu7nmQ5mWHRBPhcuugTB4y/eJgESXFZTUerKIq1RL7hKB
tzKgSknFM4WZu1ZRh3OoKnDgAooibdFXEo7ZR8iOo/1YDxN1w8tm8yDpyHU1wRJW+eEWimM+pyar
BRXwvsTEg5aGyK6fR0pIg5xgZRLA3hWvZr8lsVI+qa/fHx8opSNxfluNMnivgH93F79IRj3kkU5X
n8fUQxT7rCWuQn7nDQL7LFleHeo4xjfTNuk0l34uqv6k4SpM+kFWV5dLjA37Q4ltLd0gM9QLmzRu
U8QHrKsbsdBOl6jKz/nK/yJdgZzxmynz08oBy6Hw9GdAk2pWhZ886N+nPIMNb9YGCUZSdh+whFIc
w4j0M+va1wlZag1zrBERxI1RCjNjE0qo3Jqg73z98V/2DTyKQJDfpuMI9EkX3v/wxlBuc2frz79B
0mgyUKU2iLbptk63EOjUHuoAq9MBJeuGuKS8nBA/gSMWoNqcGhVwxqqZ8AKKZD6iliQt9yaOTxvN
FFvLB048lfjrdOwPqIxc5kKYp4Y0cKc1ZuVF6h9J/wcBS5keGY5U2Xf8rMVpyCt5olHsVg/Sm5Ce
/h5ODy1hv05JvjUi0po/vapZhVtMSoGXJSSakggg0x488F12aszxiVKCappEQ+aeln32/0eyySss
2WdGcPD6YFtA8Pjzge7DWK6Yw1REKH/lyIcj8px+mMZzkrMHSoQOkb458oyypU0HJanN4Hp4+dbM
NvTNp3HnD7EHiaigwgQF7vu3Z/nxbR0KWFUSnUTF/kbrBDnhm0lJlia+Wf5M7cXSfOwTnJpaajXl
oqwt9gJNNgZHapsV8wqrUUTm7G2b1U4qgnW5DZ9WbKGJOEbGe56dz3a0d0CPChaxb0njkzTs8TTi
OIgtAGUnGFXuNGk8BJ5RgiR0YCyrtTnjsizSbSNGYs6WRZ4k/116t6iVZTnuB9j4WeQLwaPpY9WV
TKDWMh6zmU9Eq+6oWRAvz7PqmHlwM161TBbN7tVTgBaFzq1idYhi0eWRrcM1sNwyxckyCnQP8uZQ
4VRast+HfOGYyzt/Qiij+G1yuL2H4SQ7PgrfwR8RGCLzRrLAhfwz0O+ljqCgSukfBrZYA9EPq1ZE
B/SW71RPKp7/mgkPZZEcqC8D+dIqAcNvcOn0X+vTTKcLziiumEkdSaD6HyJPBbKcZJsR4KdIvheK
awXnf8FaueuyGWRmAk6NZX/whhMTvcpmkfg8p2UevlZQGfu8Dcw8adQ5M4AJtz89jwV2yqU/Ymfq
89kUABSh0ES5uCNb4VFBKxYAYaiyT8rTV8eWzmNEYoYTpj1BsJBbBBzrBPM5uvu7k6Oj8dIbcDR+
DtdVINKF2MHCJQSV85U+NVOJLTQqP7WGtk+nhxTSBvNfqTIlJVCoQsS990TvFZlJMnMS6+F5Pct/
/Hw45vNXjn+w9Lsesm7JH2kxvHu8q+QXrXCd0aaJvE43FDwrz4SxEjijlmI7ENeM8y5Wq1avC2uT
jnxuNEHOdQ6aPkJ8ejAORmKfBuuLdqIe9lQ7oO+6lfkUWX/DjSl2Dt5jiKNhO6PrsZTw2nXTgyZE
EvCpLvmUmYJM3Vdhp/joM88OD2ydnDU4O0RHOEBK1ek4DssgaVK5Ao7+NVOOi6LnmILyCZdgqn9K
iQZFeGUMjN9ojZBb72IJ+Cmb/soyeaZ2MbWgZ+O3YWGZNugLiuuCP1rI2hAr58PAVVGiVF3r407Q
IZaeKWQuIKVv0+PiVGzprLaS03aAVUAKUZvyhMeOwgbt3PKehq5dhn9LZrKcSWXoqAbsWnnPp7mH
/3ocpRNok5AWQzpUUQjfwSvh+gsgv/SURpxDYp2ZWnEbzKIeiTgKZ0s2mrnDjf2+q452f3ghralr
qnNqbtH4Kq/4jR+VlU0lviyndNg/jZWVIv7TnJh4cpQRqXScJ2juhgtp3U/G+XxpKaTz6tEIXDYi
99fMY/PaIfIvtQTr5+C2tqojM+Z9c+piqlhv9wYL6bQPHp5c1zZLHiMAsFK4dI3NsQTs8in18ooZ
9mUDWV96qPS4XElqvmcjGXcIAtcLL15DBYwpF/kviZO8rqkiG2uJmkvX1uwIgq5qafZl2XGFgKvk
zd1ZD0YSmHLPrjr7hM0/CSCwmUbUwLalsnes88R7G8Y2ZZJRzqStN2oTco/rpVsRWClev6BAgSa1
lDaMsIGxOj9Ns0pO5nf2iEqqX5GLPEyDgpNRPSvjEmtMm2hDUOY93v5/gwjuZZWMJCh2BTed0IUZ
EbjbIw4XBoVgMSYStbeKWBQVIi18v02KId5Ugiaknu5ydCSzNOP37x7QFoqA+HPHx1KDf8e+96y0
UyRoypgWFSCdXPAuKbowjY4sq3vDHCdCAz5jTgsRAKr18VU604jOi/yJz9N3CX0RXU6k2KOfeQ01
Jbgju0udXKXI8nmS/j/jL2wDALHaXAQr/HOROzdkpdycwwMq6i3bfxCiRpDhU1NU+BVFgDQbk3CL
Lo0km78NhJ3X6tzm8KfY388rCcm17EBRXGmnU+l+FJ3gQ6omC7ML+wH2nVzVzexK/aAjFe1oNjLL
VYb8/Kg4kG7Qnzste4yW/N9SMJnzT4NAm2FhrN/Hj99MZNxmasYScAtIqfyZe8Y2ewnagMLLLhcz
diPsbld1D0I7QOP/yq/iwRXi8esbKuwEM9OOVYoec+zQ+T5nm8ZTznD4ABKMzu0eXFCRPrK887CO
tslfAQXyjgB0BlzEzGjkX6POvbyxelphiR//jNNoc979TIh89w5tY2BlQz8amchHJ6h4u2n7sYay
5Z40xasTi8WGDoEUz7WzuYzUUQ7Ei+808aRUbcczo6HDigHjZlb1/0F1MmkajYW2BcFBIfSGTf0l
t0iV6hs42qFy7LZWAyNorWYG9Y1mHUg7u4AxKpm9ZGC++6SPwLnF/UUBj615MH13A1pPkEz/EOAM
aXOzVLceroA7jqWji1C+OhFcB9BmkYHXZvQWXME3SW7Nua9wJ+ZxB8if7EUGclVPpf751AkzqlVW
QrXtH2M3FazVkvm3uruJnN5d5IfmMKV+mUQiZpK0Pg0paCR+o73X4tpY9+JS0m5oqrq0s74rGbEe
7zf8AdJ4lFpmGuacKUBY8I5UU9DlKzwVIblSHyyYUt9h+008toKhO0h6YX1COSIm+TS3Vq5EFjbk
Oj5lPmeWCaAdyxWwN/3RowB2yesSxijxurCyvNQ94kYPR58irU6C+xDwmNusPNBpl5LXWo+LYW2Z
8G0YFoBeQ1jtNHSCRNTo4m09zueyEeVKkk93TAItazdgp7M1/yYhxQnzVqim0pL8972OBSarOzkr
XOhWWXcLutFQqsjkVwPYa9aviRrqFnEqBiNJh28sO12Irmv6lLhjqz3xVuKhxQ90FDheigoTQfSh
wfzNPd4hM4vGvexlPy0CF00hRV6x7EpjIaN682+gUSBBG77NWMCk32sDfxgm1Acmd+UCiE3QYzU+
WBnlmryHTl/m44DCp/Uii6zKwhsht0nhbQih5VyhKL4s0AZTBqui4RmIIJuab+QDtAkOGhg+iKgQ
ic7G2MH/HqJNBNJIX6OjXdTgTufuJ1WCGWomKAkq/EyVnZQyrxEgnuaf8bPK6XnpjfPnJwC8RP3f
zJcu5aFGg1D4OtHqtYmhZsmOjL+lPJMrVNVMJZnmxFzCizqacgN5p1sajHJbtnw6srumSqxYMfdj
u9OYaNwwDqaRIQakVAoMAnGz4/ycAVf3tCa1YtHBT2E3JRkC4ogpgSfLmlWsCldiLhAWNto/f0t/
F5Filg1n60DnbBYDo7/+IYPoYaCyI6UD0TKPvf0b6+xCbc+3UV7ZlwHWAr5Pq7pUfe8uALBiex33
i+C1L1nNgb5RS64iBzujJRzNygUooBwfED7BEsN0+Qq8GkY56Wa4dxNxq/1AIIldHN/M1VxTAxpg
/h7bDQbK5MZzwQc/67xBdIB8rL/WxbvYsTZXWF4D1rdyKjEPiMRjgidJ2Eln5Dgo+FBS/ACrVzpP
obUdz8x/ob3Aw0sxlqJ2XVMI/rf8H0y5FJbut49MC2vd34CzVI6GYcfg0f3rMHQIz9hd9Z1Yv9iL
5j1+7SLRjFq3Ye/51ZtlnfWKbmilChm/+PsLJ9RTEVi/RYrd127fl6+xpJZDI+lckqqq5uCab92o
B6TzRSn2srYFSZFHryHz6NBuWJAveBiaI7N6kMYCjZwLNC11QXA61eaKeyZSslK/hiH/3YLiQAea
a9xJibVOQd3O9zpaZPQL8W3imflPxygTwnOtoVeEsQaohWKW20yjpmCmcFmnrR+msuyVG74R/6uW
aX05u5wainAhnmL+yRZ95aSodaWixLzTiEonbLNTJ7HrnEdZM80eRzGm/1vHTutuQ4Qs/epVCtVa
S+A26r1Q5NysHZDIm3OdBHxSE8rkyIqX/cnbWeD5e6G1YLWZxrDOIJQnVMzml/dzn+U1YJ4aZaXe
4tD6PADY1r18adfpOCIfMrFEYbyDt9oFKXG04uQuOokrIZuZ8Gjoc1fRGn+vOPX2ptg4ikfQhoHn
QToN9LbnNrBo7e84Lyza6wW+ki5IjC7IjBA8USxPHfrPNvNjEsBDmcdNT1IDruQ7xEqmgmjL0lbt
5RRKAp7Qjkbhds1fdA80bX/L0IBXaiZS5qyyAncE9MIQcFdXGm/hvaXg5cdV5LyNgVTBMvlUZEKX
ZEKVND0mwZg4rlkO6xDsve5PPJSFAk2MA4RUpiMu3A2syd/5+4MFf5fOydhbdpjhb4DaCuMtlLo/
fjetR/YqAeUV6OrLv18k60LfOduummgMcEvvQuUnveH9YifMg6l9FJ4/m13dLINi30+/O7N1id92
K6tvSWNnMlnyaJ/o+VTFBRxnIQV4G4PhA5bg/M/r3701xe/UBfHx5RqOUZQjAPRZKangqFD/fNkU
sLrnHWNNfwPuDhYXId+DAniw/kvQFeCvoLEQ28vhpKx0n+JBf+1Ek3IbR5a7OcmuU7lY0h8M6Ccn
m8xqkjBvOlQJP4XGmFMqrVrc6bWjbU2wXdaskWVdkgC+MWQPNaBBfmnD1gmtmfKtMRlaqfzQL2AU
bzmPeBHWztg2iwuaSrVC5wI2FQPan1oc3te8i41pK3m5EijWVqQ6Df0AKgPxIvRpl4skbWUop6KB
0Z9y65MWG9TYvC0b1ejUmeWbGj4VIMdKevDhxNBQmFkwTsVaOAuwE6VmaT5xgD6U36V4khz26uZq
Iwg7qj1tGPHNS9U4m+1d3bVSqsps1Rbq3PC7tebjWA3y2CgmMl/6OVdUDZac3hy6h+AeioR19I/6
817H7ycKLTlTczBRzjI/pnHbB4CxdLKpf+5bmtFmbMaM5URegbvxNrpyELNFh9XRy9AmmiCzPEdk
pWXlPHW/WmSzpjaZPqUz7gTsLw7p0WLkawxV8GI8ikie2U8wZqYuZJxbj3G+TaNMEAgbMWnnRWjF
t3LjUIt9cGnIFsT1WuKilsvbTrQERtTMTHU2hWkNAO5es2MpVLRcsUuHdETwQomb7n8Y5fxfM1GH
IkhQFbOkt4NFvpixhvfTQCIja0nLL2fHuLVcBToqfAeZ7uOdMTHaY+dCLsrHcmY+KraJl8QtQczN
DUQTUQghPObJvD3rizyfc2EHj7DWBAku0tbtXDoZUyn9+haw7YqHXpJAbWydGpwoUVOrKlWm+e8i
K5s+kTqKJK4wRMIrNx8QVMzFLSnUH6yvij+MyIjscuhvKreRQPK2xlPs2HnNwvVJKQqy+FTVcUmv
P9hL22erwdHih6h7eOMTE1eAW4Fmmt77TiX+sSWRkZmM5fPJOjwUwBukpKpt34AFRkGTaUliw3y1
8lJ9ZOShfJBmq3KMAqosKmd0tkRURYLxSX3YP8ccnQ8Dpvf/BuGztBTn7kQirJvxUXgTF21LbQvt
NZNC4IBbop1zf5UddNLhtLiug9xCz/LTxbUgRoR78l26atZ/4ZIwPHI6pUz5rsgUYzFIGeZ5kDa6
MmtMwhleq5IEabFgUCZF4xbrYwdG2mI1Yd+FTmumdYsV5arXlx3b+usF+4ZPM+FqZRsbm4I9GNsA
HHPrsWp0yho3v+ynyvEFHCdniB3WaqpaCs9CXrL/XZrq0o8b0A5FO1qr8a3WkmN/AnUtNhbnYk6b
oWyk0uZQh5LQn0JXf/UicxmNwZG0JPlVu1qW9ZR0DRc/hVWo40Be3swJSKpdeiJwUeg8FfYYlxF0
cKUN+3RudDF0ZM1oGR0yYGK+tGvlHw4vRhm5CJuSVL+aeQPefgaA1VBM0fQS60SXhSq7Y43S4f6q
StHJZiArjloVZXU44KzHtmso+K5MybHqjEhE4LtQFNLQJYdUf3ou0zBSrrN71t7alqT0kPOTKTtw
cO2mJpIZyBY5TEytu/5wEUnXeDm4Z7QKHd8JTYsqxZ//hXwlpaxOvgLC2atemt5+G27FD2PMzZpR
34EY6tJ5HInhUjwV/HPNIovvM1Mrh29JzAwcgYq0plgLxubWbUfr7tvC4dkVT2RiUpVRAVFFrDbc
ZBH5eEKdMRz6Vnao+rM0ra3jlN5c2SE457NLYNA9JwAjP/+6FAbQb1ZxO3Xy8ot6Pxt6hb6Wk8nD
FRDtmXpDdyV1JC9fQn9EwlygZW1Rzso9C0nYk9cPWtU3jhsHYM/t3cw+h2dJZ4ztG/mGFj3ivZOS
YYa/2XZIhgKL/QOz5rIKwZvlCjDQUbLyq9pEAhJ3vz3Fr3IbO+dXWKnW2ZajgGsaLL4am7bJqsou
jmpGOc9LfAVh/M+bHMQHiJok57ula5COkTleWk2OM/TB6eQR939io4zo+aNW4PDy/9gJjUrt3jo5
nQJrz4Mc+Z449J8JPaMr21Y8tC1jkuEuDuFrd973pDvzDa8OjhNEX96FXsQbpOu/J1EoNQ8JJSMY
tko6CA1ygpgihtr22EdUp2/st+w4gU2Q1a1UZ9HYyZ9CBMHEYHsQ3kiv75sWj3NFsI39jmwlhQKr
tLNtO8IEo7Yu7UQc/bKH1F0vJzxfpEtcYeiPMBCaTkSiNdmsjTJ6+Chg8q1rgCTDCzgWramx1m63
jkxiy8bfKfEqRc1RhpCiQ1lGxzbsC33XVKoeLvZP1AGzMO16OLFHvm2QyEMszLsZJc0Tz2QHkEOX
YazF27zi0UwiTOR6A9i/bt/5qE8H9MbxSCQd+vQuJs+GGJB+WEBnxn1ifTP56pl6/Lof4l2V7wf+
+l/FPHN8ybHibq/8vq04Y+2DCoOj5PCbqOEdRjR47xl7S+LpKcVDY5Rk2Rwg3UL9sBCJ6KbCwYjJ
6ImJM7/mgnG7C22l/0DyEq3URzB9LwOUGOPwM4ucMDWYT249DEk8M1dqT5WpzZhOeGuakirW3uVp
kwcsWW6mpYLJ1VZ2Z2OHHCb9/iRx8ntZ4G62Enr2TwKPiY9IEOtQCk0lOY5JmfNNLkkCSoTwC9o2
BBaHzG8nyJFLEERTAkHymIJ0689pyayADiQi7CsX0p/hLRchkduMK9vcyHdXce9+hU2JLvId1euV
IQajbKChClTzhysq+oNVmuv1IBsEhYDP7QZGh/9qHekexD8mBU/uMaScnMqqg9n6icJqovDwsllC
S7ERtkoqBpU4xvFrxy908eb0xk6Axxx7ah3DH9oigzUZDL3/aLtqhvBR0RJAOs/gp5tRk7Oqk2aw
y3hA6V4ZG3YE6ZmcDOtYhFky+DQb7YioFTdrMUEQWwzrd9Zyeq54LZybhLFAMq2WzA0i6TOgRhpP
AB+K3jtN4ku9gcexw9TuNuH9cb2n3RBupIUkHLoV0Sl8yZmLZB3qvVtX+UH9S7OUufc8R57EA/db
e16lMxEqc4YWK2PMV+y3evm2GorYCkpu9qZ19+H/D3dGhRI7GF5YBqJIIggrII6Oj2wAkbT8VT0k
lZcd+LPzYBmSjroUSdGsTSJNCcdY920cyb5UZemcDHPkFDfMH9ocFZdZbsW68gFA/7qshlVyB971
jfhpNB6T0CgIW3ss9J59nc39vW8EcVVyzNINT+5HRJoQDMsuhOWsplzLkn4fMAC86z1s1bQtf8OV
LHrbBqGHQPme2BZwXcPdeJN+GviSKxx3E0wGug64xP+95znCynzIlS8PDQ2WjfyliWjziQQJhiKV
qQN+eDwI2VInA97x0NOPcmWGvmnT7w4ZgB2Nke8QtwfxaScEblx07cP5vFJE/9AEikvc200YLxh4
SPItK3FoMccpy25rpyG1//xs8qv1RcnRbyiGOQMobuuxiKaTXivBxSA4l4pJMcIzuyMsUfkh9dVI
5B+Vv3UGzdEaJuwOvY3ZOVf2bYGS60r+FidPbgl1Nfx+NTDxyYrMYTnel+V5QdccTXwgwjYVAIB2
sYnQH+ruk/XSFWo919o7azvpP6lUy3nLZZeNVPUo+pzfbSzJCxajol6it+IglotwAlArCdOkpTZR
47jJeLIMuyo0Qs7SSEL+OEuFSqxTvStDtUoaEA3avi/nmGvfTz4K0/b4oCPeysR0hdDqoxliL/SA
lrJpg4v+1kjVi+eGo8QRvaP/3jNZlE27ta5hHu6UaTPq2aSVtCUX5eM0qzQz95RcOCi1xX74hvy7
NOul2Rvny1kkD29xcv9oFbPBgX2MYNgWFGwDpQ9ZEf/MGscvVRMu4otsHlO52fTmyUbjQiiBhHPP
ApUTa64P6KGKjG7ahKcxnHugXEq8EJqQAUvKlB7ngiCGukaItMkL4ATqYjAmyIHmR3GTmlq4CRVC
aJoAYuDvvc37kyazoow6uTX1RpoXhFAW9eTuJLDwJ++0tjZ+sGc1JjNqEtdZJcot1+hhejyKyny4
fdzZnq36KIgRDdCHIGBtD1scGkT+3LVzFBUgg8mRQhxCj+hGMcZ/BN6DQEERwHIoCbqyciTlWjtE
pYHWdSmBGh+xzITez0eF6euL3GX4E0SGAEHntmCURuQiPZFNMDuSGhXn41JbI85FDhTP3OyZOPGV
zPN2TYxO1OShrry86HeWVyhMqdEX784epButC+46TTRqg3NWvPZh1nfb17EfZMWbpK3wY32AKW3t
ULcFvEPBvjylgfgIxMmyF1uMM76SmEKI8XdclYO6SAjTIfT8oajbWrkd64CNenLBWhm7QrT+beeF
oUcgmDpgyg3UGq1oYdVizhbl22nyfieb83OorKE3LlmCmc8Gv+36XvytRqhsB5tMGnASHiE4uGvs
mxi5QoDn12HvuY4l8KAX2lnYbuX6LYR7GdUKsTqyFhyEtSqvI0ijbClOu3tOTnNAa2WhiCJfLcGk
tczqTqitCICGimKm8LsyLxII6lbk1Uxbq+ZdDR1vDF8O4CZdbjFDuiwOYNWxH3PNu5VWfPhUy42a
5LGRcw76Qmemny+GQGMwv4AltKZLy7psHxPcapoEB3p3vVXgLFEc52h8w9yoMPL8vaaCOokCuCAx
uerxmlZ8Swchcm+myUkL8Jju+rc52AA3J21e4cLxq8UeZLRHyQY3tP5FNngCtW6EeFBapvKAcyhp
sbrmANl4Xi1CGlbs6mFndHBOgSU0yFWUVaSExp80iRYR8MjKQFf6lr34RG0JSD+nxfYH8h1OI+No
ug6ItbfjjZZmuEKjyqmouC4bxL1siKnnohMa7qdDS/rwoZuoer8O+AbWt5jvkwF/ODneK5rwnHKx
tCu4kooDkljAAiMC81nC5MqLzmX4pwclGH+9TuJoEf/E5KDZlJXVbmqB1fo5yWNXgPuFja172W4X
6Lq/y2sMRwhsV1ejFA1itbSgZsXEjQR8umIkNag8TACcNRXHcq5xqgHA5juGBPgZ3HbxEghBVv/U
AoxM3Z9RrcT3lz0kqvP3Ivydzz0FKJAeqTZbAjbprohJgkChgMn35RrHo8oCroNFHQFuaSMQZ/ak
OMLQ/8IG5QEZ6TaKbXhQwotDS0IfX+ZVE9Szjv9OoHLN36ZYu58Jpu4SvdUnvF+DpzqgnE7lifQu
kGTXcKP6vBm+CyUYe1gaVXeHd4OQkbqCL56O0DqYD1sf2rkhScG3W/sT2TAVmJRMOyl7vc7EiApj
Ra4YuwOJT+3a3RZyM4RZzOEbKgldjgS5gk9KdLLhIZEBDQm/RE6mkZMdZUVvrbFeL+2MYNNGjqZq
6CnoTCGSAoN33pg97K5HbdG8+rd/25H+dUdFbOB3cu0QSqM93Y0WvehCKR536tObl17S8AZ4lyIj
Unq9oKljxm1R/l1qi35yeekw2G0+t4NcQRN7UMTcuL+vLgpLxDgWvG3wDxOhWapvtRKp+b8OnsZA
MminLfI8yms16hquarQIh2BQ4T1nLAC/Q+qYoF+NZ4NRRJ4LM+drEM0kctqjCRfyETfuvi6FB0IC
1W1kzMU5FYInqqkB0jyIqSBKFUbw0yryYO8vqP5Ckyj1p3Qbu3QIp0ci1+PLsfi93f4UZ6jtfXOY
ea8qgix3a3/rbdDD+dOS4ac++fBs62VQvxuzKAUF6Wtf4UZhwzuiJ/rSlLQlryTHY4JDPLvQxzeU
vQcuGa9py+xvpLhobI3YAZ0kpZHcdbZJTrIccslte9/uvieh3CykstI8vn1QugcBSk4+IagwYjZz
fXQEwgSIcWIPJsMiDZE1iRL2LzJmIDb3xYmNhLbSr+foQuFiiIgCUO20ZF1yHyB2zo8yOacjlONW
EcAP++cTj7Phn9Jh7xUuRIvovKXIXHMbcxp4Rm9fY8FH1umGzxPQ2ExMtDYBdXgDx0dNxB8SJQ5M
7yfzYti0y0BJ3YOjwiWe81rHHWjgP5/4QweWk570V8inVIDd19GwJYxeM9vKkMFIPXbgNbob3lON
rV+8k3STYh26QKVuGHujrcCYOQPA2Zz4l3S23F7OOGG/wj36g7h1O0ORfqPbLXTk/frGCj0FGbo4
yTDrMX76MlxfW0malsJWid7GO+I3dmn/krNcUY6hX1Pqhr8E/TvClKRXTCi767eWP59waY5WiuBh
Dhs2c9ND2HuPO2V1duxbCT9IFktpae0EPxcJ7g9dTmLiUCKlatY1mIP3k+HRvV/AjH7ShC/delPd
gQiEHaDIHvqPksHYlkf05TBqitaA10HF2DB+SaEItN8g2CSs6eI9jdLNLMWQ5HeGlE2djiEbQ3Nc
PCDfMhNmcKc8jg48H+Hu41LyM1m7Hfnv3/2rA8ETZJdWU/cNdyghVuS/zbWs9/jXSqHXjo7kMZtM
Jtsrq2UOq2fdsjjZLVbxNAAVLwX7zBaksG4iVZ5JW4eZPGSbjPa3j/fiY9XlMRoOiXmxqWqfMj8w
zZ24Bap7680iv0vVZ+uuf1Mj/TCPWxZ7pPPmkg1Xb5S+HUYls0zktMOrxxmKRNQ1h4tA0sK0zcJE
H0cGBw3uwT2Dc8bPwaILuZFlbOkxi6ABklrGJYPu3HG1/tOsPGpLVUrbq6206EsrLT7QT/Ub7e45
8hMGgffRfXbhEfamT83aEWhyFDlJe8lf98RBataqTGVL4xzzfScfJ49MuzHiOEaq7Km1tw6aVfjo
ZsIFOgoWAzTxI2AMeA6Hx9nWUMuIovuiramcu0rxSwyHpatPI/4gePkEx2fMsir9HSrFV7w3KKmN
0F0P2/IQAizXj8PXG2FH4WGMPwPfUqhLqsDo3lFSbIZvUjuwpKAxUxohOoRCCESBsCgzAEJu6MK5
P1oCTW0oq8XkYXKMwlnH2XB16hzli84fjDC5qk99/BxOm9b388b34btEFCE+f9+PwANace9VI29c
z2XzlfAxuDECF3z3rzNwyiH+4Pk7MTCDxyn5jtqTLXuA5zNMAv7W+nJm/od+acFbgyGobDJZRIuc
2D6kEGopS6cPg9Jd//zxrOb9cPqX0n6r/gQx7C1b3ow47rz49Muk16+5kcQDYXI5Omo3KSFztV7H
qjhrXJJ0WJtZyaLPIVwmZHdT+iENtTTgT4lra5q16HffuudImhJLxu46SRZWjG3tWWtzPCwzUbH0
34dmrunEhde/L5zNfXIZrygnKapEsUaQ/Fm78eC/kIQK+NQ/9bdbTGZVX8CPuUY81JkmfHtOiYa7
akzoxMD5+prnJdNxSr628TzCQj+bn452rqqpAjnFPd+F3vLROFOzREmW4JjTv9Vro0JVypYk9RjT
txyDrqdf0KzemM2eC0pkZlkuUGVejtJ72g34n/8TpJZO3nd1YE+I4F92qkGGHSs1ax+mZIp5GcEv
kiQpEO/ctoDTJtRKutiBK6eJCE7yhXrs0kiVwwDSxiqP+DRkKWGtmRUw6+DJLNCQS9wxKilsMxrB
WMzlogP90cuj2LHyv99XoiBCPS7bUSw8fyh6tPGMCe9K87TuqDjMnC/DaNGNbuR8225p3SD0qp5r
sNzI6JGAkK9uK6NiQXX1E8AxVMjhhfRyV0aanGgXYSQE5h5X68aZ0b35piChvVtkkUDQaC0W9vqu
B5ybIooT2QwTFQ/sgrNMf3o1r3qbNSteznMBLWF4RyfOlNhn+P3sQF/T/w1gDf2AWidyfpdvY90n
crZ8gv351Xt3ePS65Bv8NvrjMihgwPxBOOCy1Q2YhqHjLxmaXZLB7Z3a8J3Eo08CKY4c5HMMKKkc
ygwiiYcABoHur5NupjDq6FALxZiNiHdfiSS9WsEdvr6cuyLf26H/C8noP4L7JMtR+sKdtkg+BqHT
nASQ43bC/9tDSsZ6U/u10FbpJsvdHq56GPZWTrb3WJsSUKmp0PYkx/eKCPFQ9iFbWFfRuf4RAPt6
37ogci8P2Dg4iKWc3FNdqqxrjjh47w0uW7dK2CB1d+MDM38EC7f6qz5lX0GdhyyQUwIvNGWn+LDo
OgonHlUFi5OGaxnaUYyoDlV0T/Ce0fX+lmoFSLIIIJk0gzUzVUG6bdZIqvhn8dXb153sosuLPazJ
j2oJQdhltf4AV9j4S1Yzq09xkmOUa3rMxae6xYuBpJuzZahOGXgdE2xatDUdfAzBlEOdwfqT17d/
AEEkNu0SHfJDuGHPMKT2qq2eWjVEsLMeCsMUA+HQzH+jO8HbbjkBVJ/Xq6GBA0vZyJXmbngSAk0P
FnzR1xSSmpQmjXunQVA6wt0CmJ63QgoR9nwe/NJBpvWOsD4JSrBoYvQZ4HZz7bzPKC/oZR1YqmoF
YYJd5vCHaOyucRJG6Z7w8qc6T+EszN76AemREi/mHAVChcSvfxMzzT3yeLJw746kf+Cx/JvCOXjE
S399CesckA9eIrduq6s2pXZsaRW87cihMqxjSTd8nqNOA8/wlAIWaUzIBRGHwW/JRayiTji8TafD
pJ58VzX7mWGofTY6cLjDwKrhsVaYpN9ZqdOlX+UVSTiRcJr3P8ioAnO+nKEX7UdaGs+crqCW0QKb
A9pDhzgoLKRxmbCBvFiMAhdGvLaiGgsePPVZlKnkRqgsphyHSRK5xfBUMH6pns/41dcQtvxb1ZO4
YekIfrsN7zOI4noOc56NuvJFSt2zYslKDf/4nap4te+pbhrCe9en+qtkrvKDok67+9P4OHBt1zJT
7KaJj1JCXfJ7LGv0H4rX9KVQD4u1B+XOFUsUBe96PnOAWkZUIS50UeWgkQGX01LUbvoVaRBtFaBu
RaY+EibZFzaNcGZ3IrB+1xFcnJDBmvTLQA46tKjQF6uekJFBSftiSn/ebKWmdw+fIj3Wh/nJyVLD
oJ8zEqWPDQua/Q3bKcrYEHH6wpJQZAKaXyLunO0aoaNDJKc9fPCVBdHww31xgKd4a+eOrOTh0e+C
eJHurRAofyPin8V/aQg416cDi47ulq7kFW+9RqNUYMNZbFKCzdPy2u2XqVwViPaIGoFNrAUMVlK7
ER55p30XTTX3VzcmyD5aJpeTbDwrs+g/np7bOGnalx9mpBoM1HsDqmVW9eSeYWCg8Ru4d8SEL5Z7
/V1taKIm8Hf0xPu/XspzgnbSz01q5YXUpoNANRyx6FECynJehfgoynM96mSnopd/UNMKkJ8c1IWX
dz12g6EVmfq42EgcAM6R15spXQjfRLCfozk88YsCfp5OiJsnnOGlkg6ClIP+C3VZZYsPA6l9XBer
e3mT8pwEtVHnYDLVBSi059wLNXbNQ065Qumpa5wTDMBmGVt/DNmOrng7bjXJmsVeOLE5nSpqCz92
1gx6ZX0bEtQGIT7X1+lQNf5tEwBhWzLTikZzCnzlhZazeLEATslrheasv/CpK9EPNsvfSbsog6Mm
CQTaUdO+mR4OsGDf+BoPDlMEQBnkb991zfmtH7/CVXkOlqNOfJTriloPUJD6amcr6PkwestGIXQV
TASZ0pIEvgMjyqMnZ5NnX7XIdE3WOElWJSIA+taJDz8sQAQzjJx9AnDPxsmYx21O07Q3NNoGsFCE
Gd6vI6k7LyR1AcX3kqubKTdNPSIjlmMsp4/Ae3APTCllW7s9F/cHvUVGrfaC/RdnlRt8G/Gg55rH
gT6auOjHAMIGqFKpRsOD38dpn3YG2/z0R374eZJOGcDYWyEr9t7R1tah/TvCuZORjjJhdvuttJDz
fdAiL5L5KHeDaJRFt5/6cSZZRwSMUFmhbqyV1OH1S1eavz4MjfmCDy0l8B9FJk8NMneowtVxhN/H
FPJ+lMuA0B0MDSDoNWwh6Z9mfX1b8cL8xIu5Q7HTR36LbSZPNcJHkzAt/pwCXSJtkra1qnWz3O1t
ctgtVip+hLmfEMK3/8rY0ZtdzeIXDYy1bHetuvTrrjBLwCaeHNiRc++3CM1hwvVHC47R5SGRCYH5
iMa82MZwQWiYvjPInzkSlk2kcJVq7xwuXWNVTPa2knbX4xsAyA199Q+XL7XwB7GfMJlALlY4DWDd
kUEhHbqXf+BT3tLtRiv4xt2LRTWj1PeMYFUmRTjUm38yMt65FK3VK9kNcluDNaWHt39uLV7AjeMH
mYJasQKdpnf7BJGehEyq8uFj+rt5VAgx42+spsjr5FgonbnwA2zqFt/EsXigV8KEIseJJWH4g5S+
dZvxgLfDTTt3diitoNI8YUbypHB/IRLghF2yG+dAo8/OQ7wdHw3bcupyHPQbEBOl3vdxjJ3RI4n1
j1pMb0PRXfSBEQ2ltKRlzDCLdXUcUvP+hnOE5l1gDNWUifVog1nO/9NU41XxYd4Zezl6bl6i63pE
VH+sHkgdH1/8/p41K4qbaE4Ya4d9BxfTByjb7DH82alx+V33dRAtCBKGxQiV/v4SMeQJcC0IBOQB
3ZviQsoHhtBXmLBx6Z4kdtlkMbrKDtCNK9CON7ibxhIAYwM23Jo1n2QEPwyId/UL3YPTRKdLQW/d
GHLOtI/AVYEcDjhcgsmFvqWvbwDEeM9IDgmH6anFPTNwpESGnvK5baWZV4Iw5AfBm6C3oLnTjzok
6QE/uh8nmhzkAXP3hf38fDU25IyEco8nSkaErddZxeeOj/8+trURl0Qf8o0vNg66JpSlDV2TF8+s
TeT7dY9XmVeuCx9Mr8fFO/sda6UbaWtvqXqxs0Y7Y6GeeMr/IKcPDCZUaawi654mkevQFFjKgjEc
YWzu1izJ8KaS/fFOIgVJu/uqt8qJ0WbX7KO/uCBy1E1PGLtacwCJ73ScvQyvyawKedAuwRR0FWbM
E56pghhOnXCSoWcvR1vAahFCEPaectUtzFg2p5OAYAuHemcGQ908WWm25h85p3Tdm7wyknA8GYrD
7TgMnlxF8FcGMLGVoYEPPoprahc0nQpkxdkTLJI0zRZFo6sZuUckBXREr9hiUi8EJOiCeUUehrT9
fKdE0poXiu0gvoWkqVgBdO/1a63oP4qe0GqlR042uDgF/IXMYUvn/5uoV54ZDFzVTCMQHK8ejOa/
BlsLIWvokFCZC0xMW9ySF5JtHkEF4H7EFZUsE3mrtR6vjU7TBJBR1KtvyFeFaDNLknHLsQfhoDmw
nNFHE0IpPXp+Q7ud/doA4wY7gJWwKqE1unQ5t3aj2P8SbxTgs5gcsBIxm6pIXkMuujaK54VSekvW
WegIcEq1w83+9+X1lrf0XPijOR53wL7ldQzLuyqrdzPgFW6iLKfjQL0/ypq4YMUyjDfv0CJDZhqI
e9ZXI5L+pQ1DyKl5tMnl3+oMSIhlr/mUdtWK5TUc373MGKdFM2upVFXGDM9I2zMeHp/kcXnl4H4f
DDAu+Kotmf85g3fze7+AiV+00fiwCyDLyQ3cg0BCgf49eK49vZk5HsZgquGnZk4v7/vrrzmoGa+F
Oxxe+J3tF06gl8NzAAZiMxmE0Mth22oqEt4+u8/faPjQMmU14Qhg2TEMDt+JPHnnA8CvE6he0izd
TpAavLvOxgqfMuywBpQwvh+YP1Z0oFGd6G4xphZvqJAEMlrNAi61VKJ9TLrVjMBSUor3+1MOJMx3
p1XyGjSFCuhGJDwNhZ0WVopjbtEW7oOtEe8JrBrmXnq7yIqF2Tb06h3oCh3pQsTjTJlgNLIYIJCq
vQaehYAllIzx3XW6RQqtJuUlZCBjb5IejPIF3emY/sVTemPtAi4hPP918fSO1YnTagwrHqBPiItj
5E/MIrDsv+OhA//UrvjxHLg5e/C0M35wkDlRjeF6/tm/Gt4RZibxs0ycRTqtu3rPYZL3h2LONs1l
+v7UJurRnDSEKqT+H9mEw9taajiNkgfuQ/6Ue7v0T9jDbAVBxR6XJk3mkadQf2kMbLHEPlzZeCQr
jSeOcqIJnk2Gpf8SbZxfpGpdkLsKjb9tPk8MEF2tgL9moyEuuhqyeLSwHNAQPU5YpeCQI4vCPfn1
JxGdaaEzeodFhKkL9hnOo1SY6GtUJxHpLVUuLn3NHAWJnyrT+jO3WtThVZTxtko8n8iUtJ2+ZRYV
o/JT7HlSX701DSy5GeQd6DgP992rjgQGSb3/4YvEIL32QRPijSO0LTrIIcyKdcGvy79aYi0/pUau
1yvFfmleIxCaqqlVJDw18bKhZ1G2nd9u0DTkw6dItP43NhwyCz9jYKbskAEvJG5wfpxJPrUmWt2k
gwotN/KkLvdNrtieMDZiLIOrtze40lye8lLoBbxCJQQuREJVlyYyOqEBBRPR0/Kvt832aiak+qpm
InFdxCiEeeIVz8xxaJjCd41wkMSyUJK8mQ4SQT/1e0UfcP3GootnDgOM9aYRU8mSqX0qdfSGraHw
Es86DcKv1j/gC3QOWGfrxdHCJCt6E8uiS8N6CSQenYdLjcUAFj/1qn7l6C8IXbzCM9WDEmx0MkKM
a5aZ4jSE6BoWney4gBDqHC0Dnm5vuG3S6HkCTkwtqYDRqAy2jDF/Cb77yTOPwsZMoz0+2sa5c/aL
Wp0Tr9LNFSBEpeua9XrKTpSzmwTnVs4YeIvbKua/d7q3SBTuLp15/Br7gB95dcLUX7vkkLVTiXph
+MAIAVoH/EtSUTuN8fne5wCAsG8L2AneKgGurMkr7xMmZnVa6WYOB6pA4KFAAScxGlbPD3/g3pPf
LftgABVGBG/+D11BkavsEHYvktLHFcRBp4b+gtlCii4rK5E6VjPJjlM4VFJ+UJb4Q/cHbrurZ5lm
Fz+DjXq4oRkTAQlxyOCJQA1FuA4/50DOTXbGY0BeAvzezMupAA7mTRSbyV5Rlw0dQ4mzgIYYBVFe
4zEEBiU+vBCIqQPh2ZwuElQ8t7I9I7jieTE3vWPzk4lrf7veHG+sUvh1l/P4xedX00hZ+4en2WJU
rRADErTuDTArQrCAG1l5NMjbiTCRSEGlQeC8cWk38fqaB/rsool7mMIf9enYWVWxCFbF04zf5q/M
JX2ljYUyKkW6utF2dxFglxp4phDGQblgA8ze83tjEB67EOxvjtBIPAwMTwD7f9bL78t7+c6w7t4m
/OOxPJRzVdJn1hsOfRfHM6u27YmJIbVB+UrBhvSGcErN9bAywVxLyy4sghOqrmREe9meApngjlJU
G3ZZiP6F7zz7BS7WwRuhQvbcTxKTkmcKoTw4F8YERQzmSiLjTsdsSiT7ptrfJ6YxSSBCMZGZUM/Y
RvIMc31wdsC+Ua98NtPqVbVHVIPA/oZ9t2C0riil2fQXzVz/dKzOEdKdLYHNbEORYG9mX0AjPQQ5
0OpmDn49ZRdsI1alVI6xYh1KqfBGakFbrdov5dA0FLayVXNM8n5b4j67PIgEI69QSzEIDbde5F9B
TJRdkhdEO4CcVpJNZKy+8Ncq8ucbLlNTFkePZREaYlMEUXO4bX177I2aJOQbMGTPe8fw8DM4Oo09
4E91q5sfenjEEopBzliMwaPoCKl42bFs0Pmfd4joUwb5XaveWVCfU8RHlPN4gLrDJ7TEkFY6v0p1
fDWheLAYKkEC8W0EuuUmOUf3jApVr2omfjdK9II+6VWvl3GOB9LgLSlxE2JzgnxbgeG5cPMCMpEU
zVjvCTflQzOqdcXwG1E55CDQ9R0FkziZqf+U0q+C564IZbE2q+fU8jSnEtg0Tr3Fz1VhdMr+BTgo
LqsPn7lBu3UBYU8I6W7jWO/odVAWmtFiYMRhOClaciCHhQronlHEwJfarDZSWTDEl6v5F4XcIrm4
yHIfZRI/KA3ArpkCPY0zyl3pSNx63pT+YwzKA3s2ZP+rZtkjXJ4SH/fcjJCAuTC7sclg50eM7DNT
Q+a58K3jBRcJT5xpkc3Lr22YOb/hpgkjADy3qRxruTEvVApVznSI1lpga0iRoLd+mjZv5U/00bLc
GcsxcZedM/jx4Xf4ZSUpqCJKmrcZkqImBRRakKBvnPvIVp9Dlnhs4FiG0WQID1UiLZUcXytUd+L8
XOzpwqSvs01rVaW2BREIb5nYxiO0drxJSaxUO/AsYs3+o07CiVqx/FKKBD2DAUTPI/+oPUS+c0ag
Jw1TZYjta0SnXNN0GAfu9WXp9NaaQB5BXIETmVu6CgVXwPWC3/T9ucXUuBV2Bg+15thNfMG9xe+e
Qt7EngCeYxxjlq1P7b9lRQuW4CliF+xRhQ6NEkP+WfAgkAJ5OoPKiInPDK5m7epxYzU30Jra5vF0
LHN2qOMzSEK0yTBsDz71PrYPV0LCsy4XYTX8FpoTYN7TUnL0ZNlgOcj0szB97SnOF+CQwI3zSmSH
5Y4m1E79+W+QwD6hGjHkrp1rHS1Ac/G8AJHmDUmFf17SJ83evsWGw3xGyJc13MCDQREh3wzgDBnI
YXJRETHX+QQo7V553qLskBmnV3QgfAWO03HGR4L2ocuJj+4UZfk5oHiaxncHEglTiNeI//chaChE
rEJeGOlHLbGtGvqi+7d+DoqA2cRCy3joIyw45zMIUygOgA/0v3wuGiYd9LtdPN1IBFjpvSRxjT8l
Ux8ts+TGYJZhV4nzW/OPjfu/UZ2/pJCOupd0XMJHH/Il3A/xjYPXb1qO2P3CKpvcM/jhLk8+4FnV
GMPJxuS8dN17GBotr048WPScC8RFSogJO4cUOIsCi7PLOMwpYhOJ+s0NwP0RsTgwbBW3qjjiJFAn
B6ZgpMLfAbPCd5l7Bu+HFjtDQo1zNrSe3B2Om7k+xFz8IlIXhMkw+0makp9ZnPUaMtiIMTENQL8T
Fdx47TM+5QdqCtaHXrkX6Il0MpetZCcKr4BHbWX8hYEgudox8eYWChiPkLaWfQ9IHQ/KGl3W8Y/L
j/ng7V3725tHpcd2dvMgpkkjZ7eClb31H9CrcPLbVsIKGiNhTZGLPzYg83iNhPPbCYrbtGn2lqZ5
NdTu/fS52JUsz3PVMHdiqWVwqnwTaf9oXOTA40HW5BiiH/Bn9KB9O1PkFqsJvXuLDd9p/mWNu8Rx
wAFsoFEbTwP40AkSgpMIyMKt8GDdqw32rTCnOSw24tBs9LhvntK9wLvx66hbFPZfoTRAmM8KXvW/
arfkXfEwhqCjoYJRc1u0SJRvqNeF+K1LGCH5Rknk6RuRhzbt2KvuExu1AotfYzCIYJwItuPDHsDP
NfgGWhSdig08Tpv6LZdvIBE0dQECFDjKH0KCD8I4khvw4tB8tAXavgSbI3VlZvEd5GYwcffZftjY
kWAaU/I0ToaYqGzTHL62bNFPgRojTmSWp9StPY7wgbpdEnVaOnGAbToPwWDc31w0JWsMiTCLiq4P
k5c4TKln8J1K1zkdIt3VaGZcQCQUlFJ7u9Rhdfs64JohzoveF3qbFChtSBShGi613bQMDmSCQCZ/
DiujkOjxi+WHQ/QdjbYHEPmt5WI2QhaV+HD/k9Xzq9KW7pqV5hfMs3d1kVyDvrA6txodKZkO03xl
wYxiMdTJwaJ8XNY/d2+EBW4wQB6pKjqwcJSOBRVtw3AuHD7dbBGLOlr8iPHAhLvxxt0Lv6lgyzm8
Hz91ts9c+rTXLJzjbt9vuZClbnFhut3YlvGXdjX1oPP6EbIJjDHKlRFc0llt6jDmDxNJyghDCOfr
80sIZUoaRyp18nGzdNXIRAGXtDQi1WFWJ+vf2yIIBQP6YcfArMvHz3/5t1rjzRVwqGneweGumj1d
GYP86Azs+JGvRtXVfphiQ0hhGr7RYqKaKR8yNssG73Lvh6soBSUgryYhr/Ufee6w6pI9QxuAcr8r
0VT0qKkZoDxxWCU8C3QL8R5Ch7suMqqP5HS60TVmp+jQS5WEm2daj8JW6eEJinjY1G6JYbNT1Hln
4QmhIwoixYbREyeCGoXfk4zf1ueQOZuUMS2CZLvIFivIQ7vIqF70JI56wjEnw6/XS8gVX7XKpjYP
gLWAhDRiq5Q++UyDVt4mk5MN6AGNcYfLzA0QARid26i4s/l6n9Uyu0AzWSHaxoyO9p7RfE9GInxr
S8PMItEKEKDiyQW0DAztI1lMB5Ee8p+TwYj3T25XtKsJw67AC8Bo+355TayV2+I6Kd2EdAbq0AH7
S3uAdDl7WsTOkFxNw9+/V7rm4xilaagVNckKeezEzlmGM3DroJe/rv10mtmMw6cxR/rGGAeT6zkX
OaqUULXqe7n2ci5PGrdyTY7E5c4u38WDz/WJMuwtNjVbX2TRXA/UB6lDlS+sm5KnsmfWCqpUse10
ysVymikQfitkztJbF6gavUbLZ00Lk6FXozZB7ym0Yp/Q9jMnMhOi3uqa/jdvg4HIpPxILMg+gusz
joW77UOYcZ1WsaT/MeqMMzELcGv7tmL5QxBVMLAd3yii6l8WTKcjbK2LiJaEw8Emnr/15v9+f2oD
22vc8/Jmpxy0kH1pGuIaEleaqxds+TKNf8PtFYkt6rXWZWNuYz1V7uD14R68LHZQcizwc2w0vW22
INLwCSprpitEZGryWIqnVtEEzIHybyMQEnoKke0/BrsKjJdj0AFwEWyRfihHhmWqadOYa9yZlzFt
DaG4BjDX2GFxJXdfdDEi3upOsLODO0f03wI91euMO9SZ4zbmRfB+BWF02QvD8bKTOylAW3+LpqdA
EaQyjx/e58k/x3tfA+ecIMlGD7IwrX5DAz9CLLVvtPhU6EEO8i/s88EWezjEmGWiLzZH8vDZFyNE
15lv8l0NKOEpEDTcUgXBlYxAeAEmU/Ri0P38nPR1bn8kVHFUyFIhRy/ODoWuuCP4qS82DvSB7lpB
pRo0LikCnaShBmMkwXVKzOK/yu2YCewuAXsq0lk3wg80zYf4fI4UuQHQLbeQYV8QvY84tds/tyl/
nXcZzL/yfDmLnOfagCDMCQhRurppRPoULFwN8C6UcIY0JhY8F5Km/N1DnxqkS7I5iLezseY86kIq
J5Tgh5pw/KMhsfv63mJZXs76DhrodPcadKIj46vY2FCBLsc5AQB32F28UO32aArDhK2TLZr1spkj
dD3rURku0foUEOgoxf4UTpvZEuARqpROsRcnREyUsTx0zHB33Lmj9fNX1asXTBte+ApxR8Y95Fl1
pTLtNDzXpEVcvnAwoANDWS/JYusyKVEslz3n7+U+c38WWF0jPYhQTdRYOMguZ4Y/jloF9Mpm218l
8SyfubWDhDajUX+cQgyDLkfwcP70J2GSzNNzexH7/inyNGlUoCSyqt9EhGVORI+CC7lPeKnjErFK
6pLOKDcxBp8Nut7kAmKoMoInglvUG5F3DK4khJH95vGuH1NGSp903e3YPZnkrcisnmCeCfjTC/1f
ZoKBIc9TFmkr2XRLFWMujugWDnaTwDwddL+TV0asybpQDtmJhX0+6Ir/2/dXhPkeSysaMXf9qaQs
ZrRYEwgb6/8GydgDOM4mo12m7v0kpUg+ZVnEEenAhcHCOwB4jtwX6KSLsX222oe9b4Xg5hd35cHk
mV3mr2AG0S3Ramw/oZW3tqXcmaGTYY/yIk4CCCyP5cOimbzZ2p5TvLJqRvOp94psnacDrca69aTS
kmJbOES81jrHwjyTm8O8YSBDchrtOXNRmvngDvUqp6pQUUDtGxl2kbxXjQehOtlSB6CiY7/aodx2
JDdh2SDhqkiZpHvTacqkerMSNXBTqhSQI7I3EOAdshSqyv7NiKPGIV9KNqOencqf1DQTsdgzG4VD
1G7Fho6K7+VbuhKrg89bIPDgV3Lzl/pjEsc2dd0ZbgONClZUOVJHIP8CMSKbPm5KxapUcb6gexKX
715M0fpS8JipZfpJU5iuV/EuUJDeyj7kWWr1mojo37425KamsKg6okLcuSCWpIqsWUjBWN8mzC4o
ohyf9y5GCC3OE6UxSJeOf/LYNRjwN3z/YT8Ris3UyRPp5hK57K7aCMENY4rjY16JSZHxlbU3/kBD
7XSAASk1pff6DR+IHvemV16GAiKbXs/enB0sHEnbzuMMTqq3Z5JrbJIMBYF/U5PKGwKfufp7ZdeB
4xSwbCJZp9m/pSuxNhV/Z7k40sjQ0f/Eg9wW4m+xPmqm9kSDBV/aslNCQ36o79ED3mxffpXEsJUu
3aruCMZprMu/yvv0m/et6bRPqiF2OW+ocPnfk6FZQ1eCxBq6qqAe+VHC/fuQmtSv65UnLBOLj8Bv
+XT4SkdnuHGh1CCUE4xlwD0o/u3a7o/WPtfwESv+Hd3LejJK3/IeteDaSECsYyCsPs9K41XUYBJM
9qcDeu10TqQh5xYO5niWMybcQwcHwF3o1aKY7aLUoccQjU2bN3UGfMsJXQW+yeB7h4hfu7Vqh36R
11xGEh1eQuqGu7aVHeeFDnq675C6dbqiFPIUrO9JmgFvaseNV37DbSKh7aGHgtRtFEBIz/erCFtm
cDZ49hBBvw0Gd36GIKAAGdhOhPqkmvQ4q6Zk1ZY1R57lrgaB9zHQMy8gmjBYDqgP+QSGNXcy5Drj
SqQ4fWDNoIBhUarPA0rxhYzAebWKTQ1pwjSv8VGdeKqUbrE0pmvauNmkCtsvfSh9SZxvpdzRBeaB
iP2bybJSGZ5nFQQSuip0xQRWJZkVMVLYybIycYplElUktAoaUa7w2N6EdecMaSHvlzL1DMn7KweF
iVqcx1tS9bfHwuQ61Mr5UZ8vk/m9opUdTxWz8tjOyPQ7pCRr2yz9itzmZaVL6EYcUJtLs4k/i8Sy
6Br0CKVYtWNfPYP9UltlGMLS6c5umqUH80DBwNXAEF0Xs8HAPUWlvg5ultpgJmvPMKY8XXL8GQvE
WF172mXlHwYPD1SLvVFsDPgs+6Sw/vQ6tPCTCNTHYXG8XheYhRZAtMh9BDZZM4+1pf4YMZxF7JEZ
amHuPUBqW3qipv+QRLeZI1UP/1UeY7T5tULl1Y0yQxbkP9nal/UzUj822YQZ7J+m8Ag89RfZZO3B
v/ER0yPIcWQwUKESiEv3on+Oi5zOFW3tna9x8FMi4Ap7b+2i5/WKAs69wr1it5r2WItbo3gJvdTS
XqPua8vgE/DcA8Uy6vMMMCux6hudHpZsZCHGffdRSTc9in17keasaYAGQRzk5OcWtddTRmCyu1Fc
kG1GgovtBtuU6mFV+V452OUymrHzmdtYhNHv6kOqR5O72J4xZEiJlzXNZYHK+q+enDmXZ1ZKX0fE
Vq4YpiQvDaRy8xxmX+U6iHlYiRFCHHkGWZVWWWPzkvZKMFCG/H8JVqO4cB7LA6qRZfJFand5UY4x
ZJPV0FtM95eUvlSycu67kl/n/6R2G/fjPfqpBBYM93MYv5toisPHbXLOnsBCI9b2nrvCoLAB0eS/
fIfOWoZPxKraxK6hHc5BHdRVBbWhtjigs4Nh0zNM6BhFJiuxbxPAfs7A/rOcxqXxSOo8MRNUSPt3
TncF6zb7rb7Rb6TAiJQSc/tySwWzVbK8ICiCYxFSLZkoRyHagkT7bu/LhcwD3aC1OAR6fjh6weKY
db8xe925eW9+Bl2GRYIkM8+4VpZSHy3LY2gGq6PwHXqHWTQytB6kD6lbQY3YOy0cR88QkhVYANEj
tffmC7EDjR6RoUzGI8ffRvYpVvi+AcPTUDDZ88ISw9AgPH117NIfRIRQe/ZbjEQaFBbleDziG6qw
qoBeSB7yG/2LGrJidUjEgBio0qc4X7ZpYiC482PEJz3xw6Ofdu6rl3r46whtSy7haS10X/09Li4e
agdGlqCn4ZJcAUA++g4xoZIDi93L1wwrKBS/Z+/2OJUSNyCdAT51s1aXPjaNNfZ0jUrbvwXu0CtW
paVgySL7G/Q6XsJ2ugdoIpQ85QOzxka3eWcQjDP7dYnxcEmAubEiCfby7CgkhbiaOTxeQxAnMg0R
4WgxU0zxWHWM4w8ViGtwmegMX9AEMBCL4eGkBx+f2hdyJIKGJjxgis2lF9IoFaR0xJgjxr3cj/yq
/VlQG3sJXlQD7Xz+C6ObX0dCq83G/t33tvzIZsFvIzoWmKKHNEZ3aTLvuI8lkPPhhOjoyRDAJwHx
H8WwYcxdhRP9wjloLynRc8DJqj1UAGBV8hEmWLY70QiFdA679oFdCGLvD2c1LJ+PCG53cAiNvhin
GbAgENaaxN9UMoRaCWO9srZD6hIQWUbkVotwhr7CT3MPuflvtipm8oBvW6Ud5lAi4tM3ziwbLLuF
pm//Nn9SDZrmHGMcnW6VIIeQMbzQpPd2X1MJf9u6pW5hbd5OaVs/BiPq/KNjAt4R4fAmcO5kWsgQ
OYp+If0W1sVbIc6VS5Jm4ddPbo/0m7zOMciWWPtbMklXhHQmlKuZKX5OzGgwaoCb/DWo2zrojJrA
GT+en+vW1LMsikNZjZCMxu1rdo9oPfpK4BXR5AFKpzjmZxKdx7Ze1yndlkoOemnbBdLV4tl/dqbr
iW6E/MXgK+3Nwcxs7my0yQePZJA4TOaS9+YzSyE6rZ+6NXO3bvBFaPGPKR3GtlLEtnuU/IFaXNFN
QSMbjURl4pJJ4x3ZjNe7PXWtm3FGTjAnLvWDh4exf88sFo4WAs8cTKhn1mCPQBqFe7mPe3Y0aiKN
6cjdNlB39c90xdPZrXSXMA7yyZds/0i4rnQt0paFgEoPq7Y/MGHv1ZE++B/N2LuzYESv/MhR6Mdo
pzKZ27RaunwxariWoSSfBCiDV6LTpuMXFIsHn+6GXyWP4GA2pel3h2Zzz+2nA7P9JU5v01V+oSZA
zUL4YlVa9eIjhRQuuvDwjT6+N3zJdz13pBm49wsokD3doswufQntHsPrp4G3YUrzI6nrx1lrqi/D
7AbObYKRKNpeRqeUYePWr5KQPvNLHEq8yiNHBLrU33ggqWmQxFSxxB4PS+CkV0n7Jw07x8fSq5Zh
lnLtrds5DZtOQR5rheGz82Y1TdVyqYBqjc59V39G0SiI+tap83aExlsXGSko1qcs8HRFyVUirbmB
/bTJpiJ+XbWEhNL8z+TpkQcK+rbMx+h4Ih42XtcEPEw6+1n2NnryDw45hW6q7ayPwTYWK79Ydz3L
NnCGv0XQI0x46xg8I7rfqwOdB9DsMrHlkbwGLRXSDMfqxiK+f8xgkTxxPa0bcw5asceR4YCABLAx
agEu2NatfAsX2uOMZ7n6OmqvHUDqfjoQs9m57mFWyF0WUCIJTy6eMG+qO3FLN4XclryPoGSZHJ6I
e429StEZc675thKY+UASJA5jOpnEBOGSnr5ko1NvrDagHodJbfLrQ3jLEYFKQTp9nVggiaji1MEs
+o6IKHrgPSzozc7MGWr33363Of+S+euuzCzEfHRNGToANlUyN9VdINkT1yYyiJSzXo4NYQmCrKiy
J9ytB/jxs5aWlFRftOAH9VoNTyDuGRdzAcTo6uJiV7xKXRJ2hpMdKc84HJXc7pY3ZwXi0K9G++Nf
Yzg9D6u0XV0EXkEk7Xhg3z/hOAu+NxADR/R2L8YEo/LoH+ttMsV3+pVNbxg0es9ISPGSHKR4OU2v
8L1uatqG5+ZeU6BervxE53i8eocO0YIT+1t8kocipTl6JWbUgEaCsUi1bOgglwj/AjcydVIxFKDx
c8HDBzKVc75FLjOHr2fwLOOfT2Y9mCl8jygwmkHhIIjKVOxfAV6Mq395kYUmfA0n9W+dFCC+ItJa
TByrfT1sF6ppQCKxa09iZktkumoHsI4ZDm7X+h2yp1K5UG/8BdkCbPWYKuw0NzfXPQuxan3kbyPy
8V1+8vWCAOrPzmC+reZS6QAsdcv+fOyWfo9dtSCrvzMl+DWevfKKiyRQrW+ihOkJaJ5Vd3L7djoM
9CbQwxfXws+r1uLQUXdyAr75OMf3e3Jj7iD1VJX0wwYGkDqNYFnME0dGnFZhez2FdozpV6lyiU/5
4cczimh91uPoSeaoTLu7zMn0Lbp43U1Ocsp0ydd7HQSoqt3jiTeBcwEJljEQUhCt9Qai+DI0oxxV
nne8GEvzrpnt5acqDQOn4DDoPdzhZ/mofxaIV2sdOx9w7UmZ9IITKuMsnnpcY9LWCbij+mCn3n8L
u/3rSI07veZirOHEwZxY97YegQo+9ZDv4ciHIFwbaxwPJrk+XYYuSjktlmStMfIyLaeFA4Vvfy89
CjVAAYc2QNDmlknBYZe/0dKwvGHVUIoxOE1nWbkphEMl6IV+FZyjzCq3rvok9neWq++lS0YiKsHi
R6LsXOjiVSfwg6KVgVw82imz3cr7AWR0WlfZ2mLZi5xNCa+P85HTu7QV8aNL4ekJTUbGxDaygvZE
P8BNVJAN0myZIxSFxzV1/4LpJZXMrd4BpaGuH4qulZhHf03vMtOxA38vBYlhN/huJgAKEDKr4l7X
OrzTcio1nt+cxv2bbO1mi/dAHlsNMyRaS3FyduaofCKw9KM5lMUrCVGfsvDGe5v36IAFVprENGX5
fg/Sd9d6KWYbY6P8tPNuTT0o0k1sTXmRzlriVk3OqEOPQKFKFEN8j85fZ8sWvMEHVOwlARDlULAi
pn6Xb9CQtwhmN27P2TGSbtGS8WuFB1IxXqV6H9AMaizh2etBp9oPUsfQBLsW1d8HvHTGL6bpbm90
WDjIAcyC1XoHz6V5kvWYBxUwwGtX7UF0pnvILL4PL8h8NTiz70ojHyDmQrlixcv0C4Lp0sBhL+6d
5fZyIQmrLFwUWhHea4a9EH/Rd3l2C0fUYHvFsRT8LnkhuvgigPyexXdp04EQtUQJpmX9QPO2P1ka
y0OPWA/EXXhIbZOcF4hg9fJGxMRnvK+MZydlT82lfcF87Ysc4oKmhlk8TB2XzcV2GPwLs4Y0Kbzr
ow+MDVaxP62nV1tYM3SGMvYiLMsQNBY+WavasIKXHb+BNrdLqXwMFlGs8bGgmP7t80TcvZ2Hx+9e
Nm3F2NJ2BkN6uBix680lAM0EmoJ44cGuvVWZod5MKFBjodkTDuXs8KTdy03HMfN8uePH62gqe7LW
WAkmQqzcB9zgSk4zqbCoKDSWhDL9RvxMFsIEmP3nOBH0AGYpmkroVuSpRX9Y/wg19xur51JbrYQO
NeI8VnFFs2KRPMu4EYWQEcFZ3aTTYuBQCjL3+weDrxnjmKYFD1bWq2dZyugd5QNHD/BWK02H/zHK
nun1YZxAwt8X+QvB0vfGXZDc22+PZHiAu3yb/83GaiLnWB7VgcxyLItIjfNlHLS6Uwtoh5iz750b
8aRaDlQ/6gljGWV6ufm6oj8TuXJFTa+U6yJtnkVdaeUsA4XnKzyTo4TpQXAoyNxz65pgeZfMil3C
0LyX2DVzlkG6kKkTh24WKJRBiPYoOIde/FRY8dFWYGWIRFvNYjuEQ98xnzA57j2auAodMScKfUAC
qeG3d3BQz/+uS86WFJVya2zjhVMFUhiOn8xqwk4d/Qf86OA7H0pnQ2PdWjESCAsoAAG44oxw6e+X
FG2YMcXzDZT/bAh9D6RB5GCDYFKpfl1ocITvNVOoYlKUnX7TbyI9sUSQde7F5mqZA4ny4Tafd/O2
K08e3QUs4RzGtrOo8g3P46MekLbinQplUscInSLE3TeVDQghuyETOhgX/nH+oh0Qxqdp5HyFSf/+
8xDk3RaO1ljNReN1Ml4lA8dBrS86stg4sXu2uRD+hBkUglDJU49ZzjQHgAG76k3BaNnLCgQ21A4L
++ekV7l3Uu7ZZny1IPI5LrCCfMZxwkVt2jmjGFLYdm2JpD1T8m6Tsw9NbtxnH91HC/QM5aGmEdmC
lLnjrdygI6OW9mKmpx2LQ+N3lTMe1dPK0+o7K/QDHy6yQtKaJmkdk/BnGxN1nm28+GGASCVCFAFl
xwHdmvBFH0rwgF9fYiy6JORRmAoIq5lmxFVw9p1siOvuB63i6m/fA7+NAk1sS69NlxKcBx5++1pt
ntF/49Y6c5XyMc9Df1WktpDBujigsFMF+8YwYXE+zUjqPiqWukyZ2aalN/4ZQ60vpZfCKeKivhMP
ViatLBB1mSu5TmQFT+nsBhXubv/BCDZOTSBll9Wvz7/P1n2lZ645GAbTUGxKzdmNKXTl1daUSe12
zRrgD7ViqZfBVdTs+SBBaksr7pYzZfeV1wxzS1+f9zLAbHWDRK2ZMLlFToSKdV/IcJcrkbx7LoGp
D9vaB1fl4MFJVjUu+h0MNuEZqHzGEBackuc8LuCEtu778yo77wI/OJXKS8cWwxpR7WbQJuQ4Mcyc
foldN34/wfszfFR4zQ02VbyCHdz9Em855/0K+HF/o7isuIQCTA1xRDLTgPxnandhg0+b8rPBSNOi
GMzELGp4Irg5vbrgZueTQvBsYSzKQBqdTSPMYB8I7tyo6/HjR6Z0OK/F9vaHZhWhKDWMzhUhvy0B
5AWdCPzpM7uCBgx7JZlpRTtJdYSvvkrXnMGxqOf/G7lFaHoMY8nIuyEpM2ajvpTJiWOcyNtHqSBL
Kbn9EJIMjREJCXdzmxzLfcrGUGCGKNZoPk0X0+L1J9EwJc2wUSrVlyHD6j43LiztkoGJwS7G4UCV
CnbIupBnW/cdcOlKcobNh6NQB1a0gCoeqYs5rJtDqGvjyJHjgf1BzbpK9yzmwU8tnfSfxU/I6l9h
+zU5G1dY6I2RA91CmFKaimkwJznRRAcyPatWtDJUUwR2faaolroUwb1Bf7nkRUbKse4rkRChdq4p
6FOb0Dod4z9WNpmNG06IaNBfmFxdayP2nJtKm93v4KEr083MGmsqwnNNU7bbdTLEjVIhnnruembz
J++wvv+jXh0otNn+L70wXKnPWCF+lQTT8CqMtCdFa+EbYugkHiCiDpvEXfj4J3x43Ch/qUGhs+E2
B5AjRGJ+R/r8SRivofY6Yj5Ge+rYzZ1eY93Zfh6wXxaFmHA25Gb6FHpFXY+9rOEzrvOJFVg4wR/J
ASLV76t93cof2FeCKkWtfKDbJYuvfpBW5mndtWiaO5nWSCOPUd/l2c3rk2NS/MTjIvzHD+hzTo8V
nA8L85tAg0T5G5U5XXm6VCRaKact2VHHjguAewDfs2qd9Y5aQBEqRH0b5X4+e8tNPXyQ5ScxF3FO
x3wStv4WKFsk3b5a+Xl6lkvQGOxaTsfTHpOtw9bS7l5b1IM8kTNRLcXXIUU1K8/HWcwCrd4hmh58
jL2WPglYSAdlfRPVLe+Mn9H4PgEI+aq3qEzPi2x77XhnJ46YIUwoXoGX3ArkKd5bBoWYIWan3k/2
rxyRlb1CF2wHJj3y00XL4dVW67crZQAg7hE66ft9wQXD2sANDY181UmdEMWOqRvihSp/y+zk5G3r
IWg6anJA92gAQ96pxv8wUlgEoqQv3kmFKCpzDbf0iYhO65t6nbs+t0y7Co/gxUOge2V4xqO8LhGr
vhO+RTPpDlvL4OBOK2lo95IX006oXXZNCStoshu6SIhsrcFCSrrcntZh3QYvYtsv9+qcG9aGNG+7
jtXKZV7Km/Y5yYyXLERer4uYipdKyaKdgF1YH6rQLXN4EOvZHuCyqfy+hVZPFIvUJU/KIWBBQBfV
5ndJG1Mcw/HVw/RKgfQPuck8F0eFFAptSdmOZs5+0YMIW1At/qLSnsp/uO8Ja3P9mqSYuOIhlyN5
BR7gAd+CnmQ3jTSsNI5/6AVMVIEB/gtI109zzpaqMVt5ttCGaR17hk4RTeIc7oQLCi6XJyKV6U+T
oJy+nY5cPPxa6K7SjpZ19swCaTVmSVFPQTSbOgb5hN310fMErQWNDwrZTsH73jbEAWar63XMPnf7
rMFCdtc+N/b61DvBQGqqvD5wG+zpCV/aJwlJR848jEr4snc9c6O+g9JxxhmBuw5z0gkaRPaOC42N
hXajwY402SN041XqJP6mMmPem0N97NGAojUoTXxENrbaVhbvCi2ePnShlgoUHp45JEjZcbYP9ASE
7bAmEVBXF49oaMPYvhsAx5tNfCB2elrxhu1HZDuqbDAGhimSp5amNxzStiKcqakEMZe9xIVEG1P9
v4qKTK+l1qq/NxBHbM0NR99SaIKAlGF5ch7x7hjFDzg4iFC7PMAtbKa85uAUvBuje+C0Alv8kd/g
moxGD6Z7LQqPr+fDBQZmmi2VbL6NCMq8NHk5htV9A5ea+vx2bzS7yE8L+Q5VJKob1q+/QEMFUc+s
2vMljWFEOmR/B9/UREC79y55JEx7xuiaPakxJs7nH4DqEyA6Qj38MDsLi8uyV+6hkdN91hqpWtXz
oSgQDLLNJfYE1afd1QRODmUXjiAh/xRZR4QbuSNdtmjDeZbGdj49vkcUOZpp+6qoAxTG2rPO1eWK
JrevJ0ScsiZb2HbLzBWXXXp6V2r+hjW7M082hVqw7FwoRq9X1+/b++mtOxT31EqUqOKfbJv2GnDi
y/PBeOpTRGTJTWa9dFxWwcIBSUufW2DcEd3hHMoQs/k0GixV5REMCePGCw9c8a+EYsoE9obwOFZo
EnbFahh/WBAPPpU8Mbb/Q9C9ofWSXDzBjXeDIrY1YTNP+V6HiDJjQbTngw+nndzgtmACX7nwtJMG
voC0YOjsMGt48GNcxfXXqNHvjLhGilAk1g3DLLg+wNxVOIfzy6Yy8nfMHNU/AeNctnJxAfCgHsRQ
Khm2bkucCiw8ZHo5iT5l0hsizqpGdGM1iBt+mi8Mr86MIFrDKYJgSnX2aOLAY8EaaAqVOiejZ87I
RlWT6XvqOYtF+VpePk+mwXshWnXUfyQ4tCvsZ+KoYPeLZWq0m5KNJW2bDkQhpjwQMZjYOjIDm4Xd
/sa77RrPGEqvqlhW1VNzx1R/aPDTa/OYxS90JsZb+rLNEWTYTqM67B/93B50NWhO1mf+SE59a+GX
CpYe6s0ebGJw35InSE33E9xoHu0HN4aUWno2iP/iQ731RckkZZZ/S+lZPQzUFHcXB6D4YUJeR8mY
h8JOfUhpAgSyjqr5yqftFd7HHtiLroIV7KB/PLwxifFk1saRytkAMamzKyNnsCBsIITAaiQAMEK0
7o0gNQhA2h9od2FgO/X/IdoDLLPP3aVv/OjnCtd3txXFx03VlyR52BJuWr6ZxaX68IZALU7ds1fO
dPRIOHNDRo7vUDRM/cKsVsYP2PbqXe1eGVU+KPvmmjud1QQNTrQCnYLKmBDsyyzJAwFZag1ZSH4m
25uyBRvcKg8yvUtdLO+JnrxW6HUrfLA+LGVfB/j+8vNIoZIePyOCdM0sjhR/WBwVmM4ZGdf6IAcT
j3XKHuUTwVexH9YrDs6YpUcDPiUl4qjBtfvNnWXHrqf0B0845IWyNYxumbzaA02QgCWedn1X7Sn/
Ayblptx779gFbJbB/dHcAWyGFdzrICmTUbHqMyu1VdjfLi23Fp7Vs1JCpsGh7eaLsjWjACd8d9RX
AdHcxa/GOKX8ncPs4WMkSp5CoE9WkAcw35DWiALOgwM2J91zLQ+PXG7Zk4RrzCrYoWGyJoBM4r9S
iKw8NPKd2Km9tW0rXcKVwOMImaqzIAStc+REsrwbkK1xzszodOhg38XVpP2Od2jK7kyhMEPP+vjP
hKifT+6+qDnW/atsDPB2/yPQeTVqA4viNnY+KaZl5ZWqvSA1FVq0hmeislp+kRUCd9qirUyQpoTd
FxxNI01yN+dy61w5+Rf7PvDE2/j/V/xaqyvR23l6KrsaLZq+LVzUlUJnckbLAcxXkIEYQYn3FG4R
e41P4oEfvcvNmKY4EWraP6D+NGk5pARZ7vjmIz1bStggVoEPqWr7hdOQDYSO5dMWhXjnTcELm5z+
m7SPv9GD75iLsRepsoMA4rASJ4fllVQ8ZbJy/lQeVghOdyX/oN+SKgvu+e67PEYBXaZxZy4KI2tH
enHFqtNPSdD8Wmho9DBvrKcUU/KP0XtDpe8j0JgYhg2rlH15QxnGuECt0Vm+TNuYoND0JcIDEagz
Z3M0J99DiROOwNLSK6ywkyna7VcAClP+wqetMMJQGUd/x01JvfnRwP8HFFzyLjhVDGy/Wlpf3gfU
pyPC4sVI9j8OxzCAVI7ecwpA4SOcB1nfdNtarRuCKBzMlWSha8HJBC9WiUg0J12YbeXPhRoZiP6x
fR/pIBIEd1NgzBGL2p6KMHae95UdanCgAy0f3xVOour6fxXsQmLyJX0mvWKmoL3WQuyVNks0u3+h
ttqhd+F2AVNuQTijDgRbrL4UISWHja9bZCCxpb157JRzzoxdRTInFMbgzvXhrJvM2wKdh4RgXy4E
bAU4tFh8LmFlKHlpA+Hpkpo5qNyTe4YBu8qhSzjlENNTuK51zB0DuqFduDXE6BQ5QlrPVNBSj4+O
C/PKAw6AEC2UyS/TMkwNE45E7a8UcDkxD3SmOtDd+LCGGbepD4BG5mb03udQle2HkJNpsZ8V68Vc
eT6TEUqqLWpuDgicuqsNyMiFfP5tpOTs93N9HYAFs67coMJZNkflX0DJ51DJygtJPvZQHks79jrz
djPXQn7SXuowtx8K3tlLB1yencfiO94BUyInJ3m8oqktqCseNe0lBfrVPFLMH5rERzcavImnDa2k
V9pGHTgGwN9dacggflft4VcDuIMHZmAMKaRY3WeCxwskLqONWSzneg16L2suKWRAD1CwA8WmaC7a
kvSmCHGwk2jH6cCqmSio7NDrJk5gBuaymJbH4ZydkSvXMmnZTJ012x9R/BsqaR7vPAWiyVsuCkiR
7Jy7U4NBhcX3L/qo+yVTT5J6RQcUl64OjgX2JvONzUKUeD5a1i4sUc6qYb1ct+eo2uCpWyE6+EZc
cC2/jqSg8VrhpPU13wZRzhoSJLefjAO2BHS8AmDQnnhNWmdLdB32goijMSDKSc4/L9KXrUYP7N7j
SwKIfAzLgPIgcDQkfoO8Dlw8YA9/3iT0ajFW8wBlJrvNDdgUtDkyKl4up2qC6Cpy+amYr3DF7L36
5/zbqd94NOlxcZNXX+xsIFeJ5cfm7Jlq+CGpQdi8mw+k/rhdzr72FM11q3RmIqRSfWj5lgFeeqf6
D/JVybXE0pwdnLbxQcgGsnfiqCPeJb/mIRK2y4fEFfcklPH+Pfj14/spTHUzy7ioSyZUHw6o5jTm
GzMO2Y9O7SNomN612u0KjFhb5Be69SQXKzTe3crWi4vRG+lt2219Wyu2xeNDby06QCrRNaSkmU3K
+h02A8UML4RTac8sH3LavcQzsKZbck8Ad7rsKNLfTDh+YWDi8Fg0Ga5Ey3gafd2wHwJ5kd7syieB
l6bNGuVIgHJvjz2jzOjWq5sX6ndHPT9yNEUuX73X8kfQ5hmzYxmmbEjp6acP7f2JUIWyVt9P77Vi
+FD/hedWyAomBs29jXLuBTnIQNNgL0phY6HDE08VWDSOnoz50PbKt0w/JcB5ZXCGEgUqWRvCMEaY
Nw72blaa5fbLWrr7UJ03sFjZ5gd3Xa2G+inQDnCyyylHkIuT1hbcsW/uq1spC+WRHNHaMe7DAyWg
li3zMaNAhGESjbYfrzChCroZGV3l6uJD8BdUBAz65alradAhcS3G5+16gog7aGK1xR7KoYPAMG/e
FgN8GWn5zFvw97zyRtO9qZK+xICYSnkkwAVkIown/rBPBYPAfa8huhnEj1mlPOh+I7dTUEeaOn02
WNP6uGRsd37ATdVEEJiuMeeXFvxuC8N35rz/7aNOMA16iYrl83KNcVz7n88Tl9qS731AKEyjVijn
HQSQw3CXGwWBkMxhHf1RRJu1JJV1gOzJ/L+4CFIRx2i0yuz/HnReq4zQ39HC+P3EXBv6cC1ldBlr
tM1ihhPFoAVGyI8UDlXkGma5rr3v4AApDYUZbQGs52TWYXF7H3KXBpUn0J5Olescmtv7oplxgXye
5bEdOE9NGdEod+itKI8GdYloriyyeVDYmnZETUSnmXxjnKKiNMO93Gm+H3z8EKiuhZvGHp2TJ2hP
91y4Ep9Q80b8uWhb6BDv5/Jb8jI9VxvuVGgLAs6kIBs/ZPTBt8+dB60sN+5Yt2TLb+tiBX4zAAA/
67zZG+OvaPncURhdyqS2T7wtQZJeJhQQuy1SYshEemThSbaHhfyF7kcVvS8LOwtgvUjMTCjG0YH0
h9V9/iq3PrPcswUdcjNoA3ePGneS6E/npREsgjTLPcsA23W+i21KMGTNMd9qymwNrKBi8kolm7sB
S31LrM+JeykQABClZY8mZC5TpvC+EhbmqKg+17l1OLoIlOpnXsukp3H4Oqx0txu0yM98ysB2sjpM
crj42YLxZDrSVKb5eeCT+1NggFK4tBw9kB77WGj138BMiuocvamGUXDvAoK17no10WgQoeqZXgSF
pGwFNI0Yhmmrf5GdEeI6os+pROXBQEwtps7lp5JU3KKHpKLEltpb0IxWM5THzVmWSR4+D1AQbA5i
MOQ33NN9PTjadl/g6gjrb5xq/iTMNgyoBuigLtahOlI6ykFCGR8UHvPhauQn5GJ++7ks11MVduuV
E7GRIBYexQfMxKploV7w8YE3FUxSsxjb5bq+inBz/d2qRSkdrOw1x6A5+57BFbrPEB2tV5Xr0YYJ
v2hBlbNT968Cz2Od2MbEhx6tQvYEYeVvCYuz5Qg6Pr2cAInk1x9fyC+9XpPOZ+cd7dOCWJBm9ptG
in1+/d2GYiTdKrzgPtCF9SIA0JxRqAr6t8MnKMHhHwkBC8xn696c+785tw3vH6v6YlN13HpOf4GU
jqNoRyJTgcIaFGaGLQdODhGDYMTmxxAiiNtIjdkmnJ+k5pLiHez/XGvR9Xr9ntmu36UhRX1S8S0Z
xyI3kCvvn/TW73aSBuruYjSHlPZ1ipHCj0HGCrEIFhoiYcgD1HFtuG7ZLgunn4bmJFci9t0In9V5
uYxb6vXO6FV9NiN97xDnPlxhRE74UCypeEs15OSY6EUckESXt21UG6QZiAXYKoJOETvoZK2jUmgQ
43WnQoqxalp3GA7D+OzobeHWV82NYbEj5IU1VjRqDEOQPgAt3AKN0kJeROEDq/2EPl2ZU+QCRrNr
2e7CRW6QWHiTM7LIZajmmJBvqR0ETPjgvRA341vyoTDXcKNRcgdinOMnIkHtmvj+phECKNmfKc6G
3di2rLsxNcw20yAaBz6C8Pwa8WxQp/yGH0XsKgAVzzMa3Z5D/icOKkvp69Wg2MFLmQ0vukd0cMhr
0dU4iDP1IlcMr33LeBOgoopbgoKgLRRPz2aFJPtwVcG6rPGetuKL628ShnGa+SCh5ziYyCsWGTTN
Ql6PbNUXGDFT0L8dlQQk8ioXJMbb8BOgwwdaU5r18EHZSHn0ABXTnSFL2ZiS9m6sQVONhvX7LZYV
2fqXYIy/FOt0S/Nyj59b0A+jIEev5Od10edV9JANNa2kR6thDZy81pN5l7IjSF6oheoP0udussbQ
U1r/A1HnCOKkLvZBv+a8II5t8aLgRS0c5wqr0bYLnZAnLDEjoxImCLk35+iJzoZXU5zuYVJOdIzM
l5rpGlZpdQpiNEgYcyqJv7OD6d7RBu8kF5DQhWjoT7T6vUXcKalTMs9GtwOghMoZTMmW15A0pVdT
FjslV9MCseS5pIqIoA1jiUHXTsZFalpK/pgIipClg7rz7+d4L01vX95YCvQ2V1kOWGJb3gzNB93q
qPau6zfQTebxYMIChJiA9LFutVpEcKbX0kg4Q4aYcbE53AjXrrjI9VscsUhBX/Vbi91gtMf6rpcU
cszCc47lx/Mm0N7hpIFi0d9ccHAEg/M84Tb1610FfdH6yg/R0AI4TndWF6BwyUUtKFQE/xBUD0af
aV7rgDMp8YHzH8SooCvu8wH4n2KMuU2w1ENTaFvBiIXZPPDqlC3AhLIIQOMa8nM61h7Q8hlvIupX
rO6SQnJZekE78GAGBrXOtGTlbFaCtFgFqTYYnhkjFTGSg8VY4Pt+O0vUyqu4YHQQR3Ayxsg1kRXw
rgmUiAkePMF4wWzcPOo+U07w3PKwg5WBbrNzrTO+IHz6dbAuhdTFw2fnC1nS1KTuURBdVCN8cR7A
r5or0bWrZfDNUnhCqW1STDVelNY9Svc7hjrBgFqdojjbyxJ77PtNg6o1RdseLXHZSMgwMg2HdDgV
5Kto+FNfXfkayqPWqdHKgPJjwx4Ynwa4d6eJYoT/jkuJB6ZlGU+fOWK9OkPFU0/l0VaiO+PMHHIQ
rsCTSh1ZKPoooVgagxh+TT8YgIkK5KTORPJ+lhppO/XplD8Xg+2XPgMT1ywOF0Z043bE/cjQNMgF
sUSi6XwuOLqPewYq0dus/iRbutB/9x0k7dCPA07GM/Wv010FSLd9ItIw7z//1ouS/4tlWVZ+8rFo
2z3I83MW/bAMAine0+NH7ElQyHe1W0nKx5nCOsarqyLNLVOoevlEbJIsM7UVuB5CJIRSTQ2b++Y1
vRiP4X97/T2EawG6sTmhJcgslGPp+ehciMPqhpXsgL50+Xk+yhaZ87Xd6YJkMmupoXiOyk85tMqb
NZRxNcXKux33Esir3aTNRL47tFLjbkK/j/TPIfQzPsLb5cNppCM34RHDhtKmbVwRZbLEnP8Ib8wy
F1XACHszFtkmEmgs2gLzWtzoY4YZrwIiQgFGjFf6xCc1qdOQ3oFo1fhbBbsrFHXo8GgIK3EUKzWE
Ivi2XKtl+8Ie8ENuPmxzmstxS3uK7Iq6q4RHSgvCosA6AuxxEk1lXsiN4m+jL1YAoK4M4xNe0REh
60DIAqZP4wup17rB7jCpgPKVSy33KhsX0Yj8p7/hehNAeWTeyds/U9LBCMObQeYFgkOOmTBWXxjc
/SfsogH1yfCpOeXlL4nivZmL7xhZGp4lJGeQxW3p+3HJ32FhCs/FcExh6I9i0P0yVKZjlRknAXDo
q5X+h+KUOGeKA/HK+/juG/nfvy4Xg4eShWux/CelCp/c40/XszJ6mPDounfiC42nO/+qEmTn/P39
kkpCopi024wihmB41JAaRpZbwATBYHmaHKdwpDtvmEzU+BDyMAtlXpfdQgHUhrSUl0VerOn58HZa
lQ/N8SQWglABFRdYPMyv5vQc97Zur/TeAfVAK8zOzGdFJFdIfjpljehqVmtxM/14ukKZQ8lDuydw
0plM0JMHSv6EokcqqNr76fQeELk+jQ4M7BM8BoBeM+OJjJMAuzf0BOw128R8Pgv0r9sc6Pd4+4Yq
auKpnPHQsJiX6/GSTYy71fMjzZEqoyG4crW2jSJ4LXzHG4dr9jJ1S6UH5roBDDGBIllRwKxMFpSa
Wdypy0/NPj4S8IiGFgb9TJ/Kx5qXmAoyWLAnMpDg6wl1Rss9BcDOKs1y+O4D69cvok+HZe1L/UN/
3L4Y/Mz54SImk7j/R6AQJQXur7Zz/vHI/MhpvFp9r7BeMYi1kgxTSBVP9gLXJBLPrIaS8AynIC2f
XdLslM8cElqnimyh5zfWFtKctxKwduNJwfFrhUlwD6by1CZlrEVB7anKwykgX1qyUcFno/vNVGtv
dN4Av7jhgYRyARS2PLxwnD2ZfssZyMR95bleHqRLT3Kr3mn+3j4zgQuu9nde5gHFfn7LbyQbQ7KK
RIpi0hJ+VHWgfT3AYDDvxpk8sDo2OWfjx5blA3wStYWdrxdHQco9AGYFsRk7mP81RXEkniYlkI9f
96eXOeWzGjGSz50NNySBulR/L3tPiJFX93Vbg55Mnz6tStO9IAgadxDH+ZYT0k4r2h4f2v2DP3LG
coeHKAU8SwlEZL8XTktRy3BjaWfMYgJ2+Pnc0B53oQqp92cJwCkiN0YK3bB2b1nnApzPVJz8rwq5
/QXO9xYes9QIxDZY8Ha7MUN6Qtqrk/8HRM1CfNKOPiurphNyLL0ozXFJUbozaJ5ybZVH1aaFV9Fl
WCQfDyXmRlHJ2vW44HJTxIEB2YA0hPZgaBTOwDyJLvRuUndg0F3fWaejtqJMsQP0FPYZCKocPm3h
G5PXbLcANvb5yc0WerMv4vE5fcG/785BbDV0daC9zWcVW+cpw0vRLZhr8k/FuNdOw+qaNDF1HM95
+OIXob63gJFkQgYeWGXy60e8jfU//RJFICN98Wlo6kf3s237uhrlBqdrBoUCO2HcCk2rpnEtp5qV
a1gWeinV0SpQLAfQ8b56Ozw3HeRbgCoqduTe45PlVCb6V4VHmuF30KG1PiCxMdsQnfhuXz2K3BaC
/AoeSZeNYCgXLbGpMyqUMC8YPCCv/+hdiG68l3HiUMF2K2MYreNuoZ0eV4400TVUcVrMTWvSse9h
KygxeRdcaq4iruRXJqHkGNA3RGXISQf7wnmcwzMrNW/uw9/mA24aQO0seo0Tfb2CJ+VSNL6SIonr
ES+gPt+baLI1zSvUNxAJp1yBWsZAUpDAwQG6nYpNjbk1nMkGfKQvIOo+w9NTNhwo6zsyY93MuoYa
mEZwC2Oe59GOqUpkW1HSiCWE5aCgBKPR1L2EUdUETquRms3h1064OAdVm0eJhZRkI1nb8OJDEql/
mko6XFmAsR18GDm9gwavn52iG8m/J5Y998NTCkN31bHcj/D7FrhZYckTl1o5UyEXIfrG2cAKk7UT
y0ybLiimGSyqbB6I4GbJXj2NRUC/vcsrhPKZC0grPnQbnEy5f7rKO6AFtWhBMMCcm/K7I7XEpuLL
PbsjJCZyl6mIRMOPsvFzQF/QNbZgTDLxF14OncV/iwHxcAO/iIZuc9bCRTV7Cj9Y0FkeqbW7AICY
9/95zCQnzRqmtZ7VRBsjkWUloNDJxTYwFYDOkW9dnVnhHduTxsDhLFf8nqV+BxopqoJoMItv0I0F
inTgQf5sg55nfvwbOfTeKyoCnx/mJHyZf8dADOBc0ht7zrgx4vTDThudVP24Mql1lUJX/PAw9o8w
toFG+jdlJqaz/MpRtzwItndtVxWE3Cs6Gq6XJFa9JscZKcmL6eGlUeyqNJ10LB9qt129Cts/WGLM
QmP/69JqKu3l04De5cQ/1ecV55gKy2DKFpWWCLRLYjfPldt/DyehJOTPugYF4XBHIEBj+4GDrbuf
JzrN48fQZa5JYMc9EajdGPyF3ZsYwHLZwOEbGKpqjdi9DCNlE2GADUiUGjPm2/c8AZYaVdFAr+xh
oMzoRZWoTPDtUIPsM3Qv0ambVDyVISUKpLCH2MLDPTjxzrGyK1K8TwmIRhFGBHA1BgiQP2ZAriZD
tlMUGwFc56Ss01VMhxj2Ks3HU9pBD6chj6sgGmIxVifj2ULekCD7wTnu4jb4KgCBwfzS2EivcIvO
T0jEC7G8D72igJNa3owtr5QmkyxgJAoUXyMzvfm9F8j7z7Aaf4bbOl3yGvkzquD34BxiX5wF/L9a
1aHFeG7NRNoVTNRyuMwPRE5fDCJnQ5HcU7bdUTXItBmCYI1rnUdlAoglPTajZUwZ40yM/gjiVFmo
LNB5dm3C1ZcjfwU+5xzbJQbhQOu3CYvVjTmul+QhDu+oXU8iHpk+Eol19FJhq4ZyktjS/QoRc8kE
8mIL11LKr6Ru6wpbIzjZQkiLaUeDIb/KuxCul692uxnirbxhr9YXONNRdInvnjHjiwkYkovs6x1I
aAmFMbB2PZvpEet3VzpOxBH0vy18LaLDj9pbn/9tuqqknqhopPYAeNgNsP+TzXWVTyJGeWqhoPa8
QgkSaeU25uG0F3fLZQsDwgIp484REZC9Xm95OirCyJT7qU+IMhBSxQN9OpD+wIrRdh2OomnBPVM8
LpUm7FWuTHQJc2+QrnPxsEYN2UkfoChPCzrB3xmRCysQaHAMuXT89qXNJFtmfKkumGQj9SXqNsHC
FaA1dF40Q0VQuia1HwoIudyHFfGHVLCWI++YHLKnARmMNcBtVzzETuu5KIJLbGtKVLcPfyd7rzn1
J6Y4lABtjdlQ5dZqrcQD8u12djo4sVDot22jYZDg0WpN6LstFFA0mN+feu3iT18Qf02PG+hH9KVr
lgoKpKh17gF4o/J0rhtQc9acBvQij2MWotTx1JvN08FA8/uMMrS0XVUjT+oYYaVjxHFk53FWNmeL
2C9uQC8EWteTOW1bL1+7XucyVRxtLfIeKJOXZUnvxokias+mjV3QcUM2T2bft5b7zyYK4RqNqLJN
PWmtwgzcPOg/g/6ORmP+5TL83GKmf654sg6qm5ATfSa5hMBJz0lL1LK/oOS38fpHxicUGE7iaALJ
9BqDorYo9n75I2mOAAZLN1EJxN2uncq/GZv/JaS6hEygEzLoXekXxF4AY+QV49P3++5wjzCyS3bK
CsLEwhYmldEVssxxOsiJFku2PoUg32dQEcDLUeNhUKlYIFcK3yQLo3KtZAwxY53PeE5F4t7QgWqq
31knGASaQDJO+GqSOyT6G+sRZmaYLZ/7q5+b0HRmr2ZwzJDNzYtlwjhkbWj4cdRxtbzpMW9okJad
/RsI7El3oXq+EHIr1VSFeXQNSfFZsOnsvqac23DwwU+hTk+HJtMREbVQqOKLq9cxZsSc+zoriNRq
OjsnUCaOvTt5eifGOMvEN5KA8rtDSE2fB3xAMoMEpfzK/HPTT1IlhuATzaf67ZqFRSLYffTLJ2yg
21sOjYpZeJ3ppAF1iNnRNS3yxoNacmOqaHGUyQiqR6/QTm7wYkUQ7GjwTKnLC/MYGtTQts0VBtkq
ZuFqeOfoQ5IKtHGU7ZMcsQ53CrD1xfvU15sx8+ojBH+Mp6Kivkk3VrL0nId999nXFwXkC3nq5ulx
SOu+b7xRGN9W2sLPydvRTxrt6/7AeqImtie994L5loSzihCTR+fIrjMnrKBKuPai0raKguigJbFb
Hhmt/yOLohZbzP6i/0kmjATgj/N/82FaE75rP22dUQak0RQX5CkB5udnERK3IgjmfaAmEJkBmnAK
mvPppFI9LmLysDuVeAH0obZ92er4IzOEnQMfRFrk/0kAbTi5QgF861IihXM3+79KmpIze65zfj/L
RpGUTLB4fMXnTU8TDClTUBxz/BoSuCDig0bwFU2sXZZXeKBZdGROMq+AHbFfO5rOaR0Xd2iwR/0e
7rsfitqwoYKb6638BW5BflacjyZADYi0FOrxktTPvy7tiPC8joYoUcaX3JuoblUMBZHmZ9IPwY5g
NdT/zblT2uZ+2oLZqDNLvucjm+oDDixg2+CnTiA9Yy2c3ipZyk933YC0OW4sVKkLSFkfPkMtDbtP
89AnXb97MsemP4CRAVwG8zOTLwraAWMp2KPHgs8Degh/jC/t8AOgrUzrs2c4vx18MJDyXWZSUJuf
Xoi6GPytklB5BKWuxwf/1xIQQs7BPomZu/lI7Ki2P1r8xy4NT9tTC+9YCWgZotA8OyJd56cck4nn
B5qPcY445g1KJzZZbiKfkfZM6Fb/kOILxet3DvOu9OxxMfFG59oUt+u7puL2ie+9ChHrF2skrOBz
rxyQOppgFOsGIyqoAPXf//L+wu1IYM8g2JDEQEX2J70NOcUkt0p4q/7yKoD335SaKL2kztaQD6I2
6IMNkP9NnhMUemvK7gjBBg5pUvTlrZAHCZ4y/yzhcSX4v6tSqEZtN3W5lDOqW+ikihjU4OJCareO
bxlyPultpsyNDPq0K4XmXC+HmkIq4P4Wt7lAtaboNkWP5vmb3jNrXnbFcPfQvQ8lWxYzRWDJWbqx
uHX63h3L2ISDL7KoTmmEj/WUqt2YQvM1fCDk0dadjzA0RSXgZ4SrV5llEbz4DaXsQ4pvnd72JzEO
8xAQW+h1gG+g0jqppMqvQ37LGcZLpEjTc8vKd82p0Zl8v7WJZAqlmZFe0Y3ewbK4Eg7icJCRu8F+
aOiMt4Ovmp50gOC8XUcGRX1apNag3/IykIevc0/+eBzN6Q6mepqTKtnSXLwrepxVzEpR9Q+n6Qq9
U5CuRDDl4kom+6Y922wpZ6UA+NvRhtT6E2rl8BdV9dJyZas4y/Wtgyd6B62DFrUf1oEnF9dpxkrD
t9o9DIiuUQuLhLbReb7al85XB4ho2ijKnlF2gRJkxd/MZvk+MgTviDcX7sD4nC+JFmO4Zmr+Yx8e
+40tZlPEeGQNozIHvfbX5m0FAOPn9u4LSq25OkOtbKVBz+x0YRVinY92Yq7ye21VkoUb/i+Jmjhd
TaRL2uabr5GXsx1rLs9B7fc0qjMDcW2djBb7+hzPG/V5lq2CYGuV7vypKq2qE4H21w8UqIL3rY+1
G0TITnonKweX6N6zEu85Q+xpz9+3LifM5f4o9ws4Omgw2kw2ZnQHGkh3lUSYra8Ct9CtIGeJmupZ
EY67sXyXIlmM0ipjKuBW6vyzbpkCBhxH/Jkpe2leAldIWb1wIStxhwas3hYw4f5YqF6HvU4fbzT2
5YrfO7aoUnEORgDd0JljsBipvfgtLYAYreOujmUp9zEuVi2orkwXW1kclPoL2G9g7Zw9dtYNF0qE
SPDiZ0YA65vzgzp4/gx7HVpw/UaZXSZnwmoiws0WocmATyIskfe2GCDAj2ZLRdNIoey/a9uQz757
wIBstzspEns1dWpjG+y3QsMUC84dp+tib2HPSzYpcBOn/nskCmf4XKUj32VYRgbis3tfvm5Y87rE
7Iuaz5xYP9ACBj6y1P5WjSQPkomtjS7V+/8I1yh9J0xDmBf/TJIaYBW1Zjvg68Wj/cvZCY27acWO
RGIg/0UzBzmoB68XnlXHlVb9kyS0L2hIDV9mxlNIFr8JcxPMhz6s6EiUL7KB26zI5VE80ks5rhHH
f8c6pyT8z9aA1TBm2B2/yOeylJZ01vvfW/odfQitx8cjmmbRFvpGsvzdszBQhyNmZt7Y+qjftUGy
DIe1LKtly7aJsttVrKpzVYw/bHYCUgcamtz7zBdfjITS8QOedY6tLVK3E/CuSFgBCyEbrpidIut6
YNNat1z/okCobUVg97ikKuPGYh+MPg9WccXLCU2a8vh4o/+R0HZIE5MUdPH9ekA0OXk8ZdvVC+WM
6ifDtBCTNQs6AOumSqQ2dROGAUTETSrlen2yBmK9hcycNgErzUZZqdMwgLbU5YPCiu+AQyTxEeHj
l57h/wCZ0ICTluyuJR60ycnuhS9ealAVA1bg6S3+f00CnruDx/8cy4piF9Gm5cy9DRnp2cTiwRoO
d0SyS9GqMWXBPO5TpO4raS4YBXcLRHhKhuORC3UMQXlk/fLgqrMndQWZ0ZzeC0y353kv4LxO54Z0
RJIk4r675ez+6WD9DUDe/sozqC7A3DscFA431AXbnA0vnNNDZkoZyYYKF9eoenfg01bzIjY+RUXV
/0KghKFYSD+yl4Vb5cap3iX8cUpEphXndUK4CqYOyzQZ7TV7psOIBKFDk7bpfHYJpGMdtAL9F2NY
zFkp77U7h8TPT6/PrBfPYAPlKweME0K6z6H+RKlvuhn7IY8lRpWXKckrKWgQfCgzIhzrNkao31Dv
Psiw9jcX0ra49kPr0fNdt0C5egKgbCKiLogDBUErfI+cNt8eGvokgfldi5C8PtjGQG3wSgzeIm/T
RfBsCJ5BS95JjliXuQ6kTYcThgGO9ybvPnSTfBSwXGqzQrC2sNWtfPv2l8WVnF94ACyoAB/hD/MS
iKF0saTljJmUkgXXG9g7vjg3aBflKWcxODH4uWONLYTn/7A+M1YbDhewpxWxAHs2KqIoOb4dYlvS
8uhK5eFiDR+5N6m2odPPIOnfU3kpcIrNYHE9x57M+ZzYDOh1nKVsJWF4+wDyn4lw65A5r+6h4wEM
FOeSLjG+JM0zAT3Y6cjf0spDK46Eg5J6QpqWhlqatYJv5r+CXyDKgjZtqssKV6qOjXPiYUY2lJCp
vB+FoKGkHBxjtQTbEZtelYoTA5D0Dltgjb5BWo3P+6ojG32r3spms1Fveb6uXT2K0IdJbAtiwbkD
e+IqV+3dzy9i4HWwL88TXOM1icc/Zu/QVGdC9oyoBaSvW36AyzxvqhNeJmRXN8A62h8iLB4HRYgG
DUv/px5H2a/dMUTjsbR20ec2c+a9paSXZ5E2GCkdnfp0W37kIW7AyHDTUP/4r0+mr+QOot6cMtpC
9FTpdCkepvN/ZH62t9KFr4TVog0XNPfw19B89Dt+9LAQ21vLT8Nrtf066BcVozJvh7e6rN/JojsK
ezYwBgz2EiPaZBHsuh+biuZ/wHMGG+SV+1802lxSf5sABIpd/K58Fe8xf5SUZlFi5XF70lCiMQYn
UGwQ0B2npoFkff77podFlHsVSpkJFSqjQCNzz2njc7lBI8fPjIPp5qiuABu+ZSNrIh2+5ipx2/Yw
TV2zeXT1EfVc3ESDqaidAyAqqAyLYyGvHo4K4covj69aiPDz0lPpWU/qk5xO4EXzqe4JAZna4Hxx
Xql0PWzLNfnHMt3TpmPKpxWz2rhQSzBsePHKP9zCISGnM8Et6uSvjbQ77ZpvGimMNUaDZx7zxVng
jOL4tYHtzESVd4oBYBm9HUuAa+NQF5XJFivaiBHE+cFU8NDXounez9iEJ5jbNlh0lSm+QlxM0K/R
sGyr9kUZgkdBGRUqMv5mnznXNKX/ll97LG6JpHWwKKVktyChfQMoXlSMzFhag/Yda5O4Ogh6JB6F
JAZO27BxgBXWvth2GpYsNHTKnTfpll0SBaVhDSDWfVkPEFWmi0TMBciawjGFcO14M2NkWZAoEa6k
ETCn7X/WSUZlTufL0QSOj97gTUUVAqbdSqSGQyhmWuZsxPxxJXKoOEz4osAP1FQh5zQGGzZCeOQi
dkFgEWzqm+rzS7MGuBV7I7+XyCd9lIYD8FfWxUCjxumJzPjc8geITZ30kYv7asd1Tay1sOa+bT9+
6x0YtqnblMAn6abuDmXVinugQX9+L+TMFCJt7VaeF/pvJrCko7YKHAz8k0jzAsrmHubmMJSBd014
cfgymgOw4n1DmmRtzr0CI481MEXbDeZ6nuc7CST08zCV5O/1TgQAvZg3CmqIcf2mUP6Ue3dUafu7
b1OYN70xXwkriEyG6C3R+I2aXyddsMFRMACTSwBijyDdb8hucfKyALLHZ2RJ2BaRySJrt8330h43
dOlUR3+Iemb454T7brAHdFkuXHI7pp7icBN/1fJEpxk2bRtjC1UvMQuWv5nbLaYi1R3uBnE6YtzE
g6I7DLrNloiWnIRf4w6SJDGvjz8hMQcDLyBts6l/XWnYUce6LwjhEbYyLIuqF5gvGBRWxDyGp5BW
qsdZFqoKqZgUXah5CmisY7UQA+lBoFYwZydicfUWEoxN6sKG1ggS1uAAV1Aw8OQ5uqBe8GPyM5wL
p+T82vCtGj37gp4zO9RKNQC9a+xkxj/T8wUWPurAssQYGUJ20qgSwJ2r5xnI
`pragma protect end_protected
