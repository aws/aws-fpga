`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2024.1"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2023_11", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
teJ8nf0wANkUVEl96P9/FBQxo34UVz0++MjrRHR9DEqCCYKUK/toJKB7YspI7XDkvE1vx1FnmyuC
GTE5C5txpZ/GJAkynDOVlj0BNOp03YSgxXau/U4cGnnsJyCB2HBUfghNdHoUiadIftQHGEjOyksq
tbkZI9Ihcu7yXDybYrDry/qkTfjFxpvSTg7TzVG8cAHicDUV5SWhkBcpBBiVZWD1m3xU2L/oycbp
NtzKj/r1DtwbLXv4AnNCFc/7IEceUsWCmxnM0xnvGHQX7OsyhpyCY6MUdHbY/gYOqXnPXfLvuOYk
7WUnGuhMpappoR9d2Vqv8ZVReYMKXttTxsgfxw==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
UxsEF4BbxRtyZas4Wa58J0rZK1X8sfjfFW5n1lMzPDjwkuUdhISi/OoxHk3AfR7o/Vk0zaUoeVuN
mmmugt+8K/ooN0xR4vrzqC+mIJvOz9Yu+htyQpzC7v3CGIBWPz1gA928Og19q99R8lyl1F7X18MW
+9BDc0GLSa6rDAue1Nk=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
B/QfzPn6Sed03EsjNKBmjMJM8Xe8ESuUkam0K1vSwpXYxn7RlhPl3zzMgIB7Lm7m6Ggn6ioerZaE
pytAxAT6SSqL5ZPJ2D5PK5rGk2VEw3+qPbMZVB9tI0nkxTmphFGTv9Rxo+i2SC4T0O8SqnXu8qEz
RCd8HFgvMrdeDB4Mm4c=

`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
hehOgsnZ3Kff2eFQvGZ9dub2HK9fu/lr6tnm5a8ViX1JzYxaDcQ0QYXxJEDxu8PalIgZnRbiBh2a
zvtzXKr3Pw==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6304)
`pragma protect data_block
7XlkuW8+6yWpyXhKgB7bDHv1EniQdX7LfXfmy6ICO4IwRo8Z8eK7FGj2srkT2EMHbZOFJ/g01r5o
IqCyQyNJwfVTrdxhVy3cL/8OYz0T5SsNLfdOWpBbHEsNHoyqKtJ1bSASr8uSKzxAaLbbLQrCHc5u
TKxEsi1yHKaEDtQ3rvhpbQdFp+5rESAabxh/XGRAgarSRQZUSb/Z2Nub1YcV0G+bsmAMIkuVqcMB
KSLAjGEL2GfWVdNr/QE4vvgYryh/fE/BptGAK0QIrtxZYy88qVxKXQSVQ4rhFgTIGFGKyA/HzfLE
5DvVKTcxUD9JAgNxt53LHYiGH7r23oWxcI7xRLXedlgH/r/v6kWBLF8sBOO8PHp/NvcXtcnVkHLF
wNCytd22/cFY0viOaCVlwVQwiq0zlk6M2xpCtW/rR5kAkAStWECtOhP413o+f0U/3delIhDm1Yqr
Xh+49UtR+Krwr1iUtz0dFJlhpinyr6ZRJ4Hf6y6iWS/8GPWXtnIKRcP1Ip7gt8yzY66RPBgZWdnW
PVlrjRpgNFmK0EWGDkpB7TAVCPo0zHEFBxF7H2kkC+ZJOFg+/pOAqFDG6ooV7dSxXQTTwXOlazoT
OVhJQ9fwrpP3e7ce1ugWbnSFIpbfDO823PCxBwo1e7isATjUdySRDw9WCR9/9rAWuSwkfKAyAiPN
dvWcWm6qPB92jyFpPmzVEspwQV8NyziYFuxt80Y9p+hNRC/y2z9BWKXIxMBiXUkpGxnusFQIQw8w
CZP0ObfeIk9PY4Y7LRAP52RWgk4/NN3H2DH6aG6Z5hAB6gT8NrX7ok7QjnceW/UGU0vbsfFfzVb9
dqGvGcjN+wgImKyEgNI+M31vQ2Y0UwrSkydpbNoO+QJFwN09oo3NtWWjo/I4eY3giXRBa8HYxait
9ULhriM5/+AoSN0QI6HpOwTQ1OreG3lOwAtj+EwkCoz4CbGhqeFcMQigcIqptD0SaR3TBUT7m6Ch
x8HdPLcY0CGN8jLf0ZsphniWPtDwh6iFTsKgQsdaiUUaQz1O1UZeFKgZmGZzgQ4Jvo5ZoA8j3I6l
F309gfx3L1b9q+oCYmPdCNkCtVMz5IUcZ0HGJBg/cPV3h3AN/VV/WpElhab5cg8Q7TiR/TGFzTXB
ENjxkWYHusZXge6uMHkzElHmvz9EPn4do2isVSMgL0GkJpjbE2udPwqTeh/e3PYWBDAe+a0lvQaH
xCmGI0LSh5H0dmdiOkyhlioI+YAczhGXFzlxUsTDkH04pXWqIHQEPh5OWHvr6abnV10m/G6hvLWz
8J4qwePjk4b86n+NXndfA161d6sw9GV8eOgosdeLi9QElT52JRXy2xnzgwQuTjLcvOFe75NGGYpW
DsV5AlGLLN3QRg6b7wT6mg505Gh2cpYq6m6FUUBVtg87FWyazDu0bhoz34Zd4IVaTJywpI2+XGFU
7+FH8WutD1jiycAE+PmYnv4fMziiB5hzIMZBOZ79z9oACUQ662ExvewBsaiw9f7L39byMQBOeKaX
MSKzoT336Ye+hogy0FtvmsOYXgiQhbcDTHm01G2wuUpUptmM9NQerAOf14bakzUbE/QJglrlLv7o
gmGw/A+j2zsfDxyA/u/+VqHcjk3R4a+QZOxX1sOdwjWxXZrO4knA7Wen+hphoFrhV9X0S6GfIfPU
nvhJP3hOWFex/6+7hJcOGKa51U0U/8abddzGCPTuR6puOGHrvRvPHjFLuVqQ5SXK5rljQRu43s0C
vCpruxwg31Fst4yZ4E2E0t+iyP5OXYevwNfF2FkE8+q4Y+pniXbExRNrksxbpkF6eo1ZvhI7titw
Uo2Ba9aHFMfiABpcwZy2Tgkq2ZFI/F96ZU+pDMtanz38L7G0gne3Kxw3RAPn6qZk22jZkR2f71xm
v9+fAWvdIif9FJ9drGAd4goHFprPwXpoMeuaVAhCrhMV0RSNnP0s3C9YLz3ktz+Tfx/8uQ39DLlY
wgfpEqn+El6rNyfaoTpQCUi8wP800f+DS9gnZNx+4IVGD6JpKNTcTHiGeAdcoQp8MJiz10cjWqnM
WJH6Bp8xGAN6QA4mIIjTS7N1EY+cuZTUIj2O9Uru3Zpt/GjPRlmQGj68QRcQYQAlx3zPXffSlryR
+xKPVYMjn47VxxfHx4ZBD2ZGpNJWKSasoU5xYemL08Kxu3oAvOOnDfGlHMxc7osmAM65Xzu/CITY
4CRMU5BTacsApk81R3qY3tL1ArjeIaCEBYbsxg9dfNIBIi/6mGa6XuWHxuYfRjV9nL0sgidoqXoG
qy232oPJTWEhuWCZpV9IANthJV7rkJfzrfmrQxtdkcSAr8XytSOXyRfKBQXFerAywwOyhYvx8Zp2
gcOgmPbzTHipbGwzhTSPSWjJTz6T9c141jChRqqH78x34smGd+0sfmg8UmBQo2uJHyEefokHr2ey
imKzKiTbn8mK07D4smgChjHYQ7vGIA5lEpA7rtNymxuwvrRsjwgavFENqI7E0j9lBWSrTnkXGFlZ
Mc1TzO0IL5XtQNbWsZu8NO9Ym4AoHQz7jbIkaNGq3J0Sts3KFwNCLg/4dBRl/IrZl2gwssLJJhoN
QW7y6mnPRf5e+cXe5+C5mKBA37N2+WhKsyDNav72PjhFxAVKmneXIaMujGyvqEEapZDLLY85vPiS
stTXyKpoqUWh+cWvFbg0IPQYIUd5YDgDgx4rFyiSi9ZlqmJIs6IMo1PNndmnlFIoEwy+eAaQfNOK
gwDmslyR1vv5BlLPZOQ/GKEMOJVdHXnxYXCDTK/4twPeovfYLbQysyQVkCwScBhyjNvZ3OVXjesw
jNBAATMKTCuzP/3bUTJC9WWMpyG+gKTkqzb1w+EXHswcaUNTI2OCVByBaGSfb3oviAbBjWd/pouJ
3YVLHekZgRWDECJNYBX25cicgZXOpWEdWCG2CneFqaWvEC9w0YUH+02N4ihFQfn7Y2nfhrSe4Bru
5J+Tklp/YmBMb+lylLe0iMntvBNoi+Iaq4VRV76AFelUEkA/08Sf3OsOoHOy4eOLKj4aVOIpCdWn
wRbWSQWooK5X3IoLh3SvOmRdX73QQSkHBRT5hyWUR5tqUYb2Gp7FEAPUNXFaFaSYNnPIu3onfflr
4Y4rLfT1hwPooMq1dnSi2aoTeaY6/MX8AQzTxaK5uiTRz6ap59jqtoxHZQhcfe/HbWOBCJ1aEViK
YIhVHQBEbn5BiArfUQBmKik2AD5lF+tw/UlAUmbgw1QmdZ+wTKXcGlYN9jPRaPAaswJnD/gfhl+A
1nyvBfF5Y14N1MAxC5xVi2BVDQ7iVqhYA4rGwInxacDp4n72J0kJ6L6tbTebjN+ZeE2Fl9lFNgcZ
4RT2yfipQbLDa/UQgjlkL79Zws8/8J73n7ZZbckpO0k201SsFa9mdZgWWq2i3Tiom/QTrYfsWdRL
RSAvHdhzwE0j6PJ93ujRdSqJvtSjylauE9nlcvTuqqaVl9Tz4Ten9twHzprG+lRmZWP4TJBiGuiO
amgoBrTkaCwhxoKpez2h7vzPHDsw6y/Bquo727lscqK2XS3eAEs+U1IKRRYQpwR2FNTiyB6S7k72
tKPkzYBn3fVR9xnGKbNWfkQSEBU9vFMoQw14h6iTEyV9NyNGaL5Fl99NE3fLqk68Kgm37cGQJQdD
6kgSKfgVhyBYnmHcOdUzO8PPe1zlg717QvOugzOGxBtiVzCaWf6kh3xnyOHgq3/sZGo94kyb/FGM
FibZYb1KMzOJdV7RAlf+XKqFG+k8ziZqu50YH3zJ+Csz3Nu1fJYM2gFQ9t3iFB3FNwJqHjLSZcIr
kxdF017/az8k7i2aMr6M48cukCWJ/NcXim4SBilUtIkHJOhrhgqzLfrvzQbALW7qdXPsAk5U4GrO
um6p7MXQyLJMSQmewgvUT66BWGJdDnMIT95B3GdDc1vUIlXVrPR9tSaUf+18LS0IiPfyvycoJkV1
v/Fv3SpM+ap/nDMLo2YaJXzBvEprgK6X86sMqSc59zSjO4rtN+KdLJ80vUPOJuTxI2uqW7SyPANy
c/7L0FIzJFuxHN2e3CZXOn354C+/T6FNJiiLUzXNBNYhB4l74oAupddKdm6mTF78oJMTY2dE+7aC
CVL6r+ddQp0pHAQQeyIHirJC987o945OH/juUNavyPTZttOiYTeNA+ci43cZnPl6tzZaapE78lV1
8vLnrP32DW1VA6HuzMyFFBL5YDtVdNKHmURwmv2xjUoPUKLsI3i5IvmQU5fU4zaTRKCv3+SIsEgL
p2EFatwwamjUz/qUFYlo0eT+RASUSjMYmEZGreFKpbxg6OWAUV1ANPjYO+Ac9Krr6Pr9r0pBF4Dc
ROgiktB5VfN0aeeRSrfr1rsc59jmPGji7tB9vIoSGNmqg3DObSwHGZhDydfyUMCVdLzjVT4BU4Er
InzU763nJRKrVO2G7lXmSKFgU3QxECd0BaJYOlGKbDuivenSA8NYfjCjEVgHaPjIcXw9ISIydV6K
QJeKPtYxYLo+sOwnJlOl7877q8ZY2Mq+FqmA6gxIgt0YYx39d9XeE97g673Yz3T/be76/ZTE/OhE
85kG9Niz9GM8MnIhAZGSK3ZUJ546tV1mEpEPTUYcp4c2YzaFGN9eWJvySlNqEBFPZAFusn9ui6kE
d60Fitx0EOVlCG1JBr0G1QdsRvScYFyRzjH38Gi2gMm341MP35NZcj2OHQLroe2JVa17PbGMfewD
jEGitGNuPNF1CsT3mlkj5TlJ58CMMYYjZ3owbrCpi2k8MzAPnsQVyF53Nrtqa/6ng/VyGnTrEbVT
hJjgOr6XHaYdu1Im1rKJIvfGicF4GUgTSKewe/g0BywtIppydpet6OHEUqIf03RBw3fC0Qfba80p
BIPGNzJRVqmvgt6s44Fv4fZyk5m9IOR9DmhMAoFw/bxe1m06+6/nMw8PskivGyzkRP9bkWYZztYM
D39wIUP5fX416QtlH4jJhcu49wUT8qpv97FaOpMs8mCvxR93xclnVHVOm1chs171cEd2/YXWVIhJ
Uge1NoBZ4MGC5+YyoSSFcJGkuGso26Z6xOwQjgq7w1ZwmzQElY27j500UVmPzTIpM4PktpSXrBct
zcKTk9R+/fg6+YBi+B4p4SFnT71oAQZ6tBNVs53ztRqlTlwXRdQaQzE9NR0tb85d3o5MwufqtBw2
SuovMCSMrsp0R2Z/30Sm0tkQcYyonR/2hp7Kd5FGbSXt6HshLp5uTId9Cuquyun0mDJuR7Zaaagz
ECaaBJocNetEE7QNO1RSmzKfrzPi9oTNN5lyIIjxsUGJ8OMDROpnP1TOpLi6R+6BPIjEcgSNLwrs
xxVr2Z9wALUQqtMjjDNbpA4nyPLFqhbOoD/CEf4vP72geFVXUOO7FN6iWmnuaAEAvUjdsHs16yNT
4prZv5uVea7VAiH3b63ntp70oCP+aUA+4FHaXUvmQLVFK2y9d92VsO6TcRUJwpIQnuk753WkaPT1
+ZejiKyaQdvHMFw8SXXEb/eraTM3YSN1Vs/msWlfyStQcm1xxxcyuCtfqKTGP7CR3SPz57s/aG5n
ZkGu453jCB4YTz+8Pl1PsrS56e94K49Xx8W+ROwuCuXoqpXUKjZfpb2djruB3tRxCJP//izOK1wm
2YL4LBYp2Zyw5tC/3vOGlTXrygEMz0GCnWP4/IvQczl24enuTCYg1wIU++j5avkgBR+T0BYno+gs
6ljg/qQslae5zzPYKqTFVBcptqAO7+os/vaLrl7lyk2EpMKaQaJxdgCHddFOHqud3VzsWZUfHcOX
H3gPAtKi4tC8KPSTsgJ9Dnt2bqxfJ5H7ndk8syuUlamArPUt3P3byMIFNHL45QEga70UG7YlsefB
OBiUYCJanuznQ9oFsphfqZRejJoAYUAKu19qAU+GwM5zTCXpV96kH7v0vQCEt+kjd18v27F3sG35
iGn98VBT5A/Y1ynF0ESxMVKFa8KZYqGA4PwqjkPMPFQkKX/x3FrJKnRBimmRaExEvHmgyLQ9i1HB
Cu3nj7+l/GNZzfNqAFfKRzoqrQQ54tko0qw1AgxqjCynkQ0IF9Qe69b8diTuKepVi3/B15DoznRV
gVuM4shOi4Y1x+1/a2HBO37GFGjBsh4aWvhQ3XWxX0Q/Zh452mI6SGbYciEsgrdS/9xPViWmy3YN
qx3kW2zv1f60yYv2+VT098UX6XBbofTV0jyjMarF/BTE01Iowau9v/DbrXW0gNXxMb6WWQ6R/b6m
l+9B9VcfEcUJb7/LhpcgC+7OilhzgOlqMPMRnMQJZuyGswFzZSpi1D8XcQS1HwLHpEZwjVDhJAiN
tgu1vyn/DiFBThm5SBYAebaRAtCA0leDXFOSPyGubPPgRP/q7UaUm9v+Js+bGt0Ui3kG6TogOZI+
+SbKklUn02vYEz3YW6VmAlNDVM44jIhMcXUpa9jl+PX2HxITm072zVDpsg4UzV8eYayAxvn9Xi+e
aUnoUtvNAXJ89TXL5ilpiqFgsTNuG2gdTHmteTpUvrGb1QhBbkqHdIoCRPe9swA9VaznMo0DUYJg
uq9jM9Rea5+BKmOa2ETlskp2daeJeEJhU2wvvOCuYr1XoJO5wYMLJU8sqEzAwiPZU4JrCfAgfkHH
kgXI6r+nM7i+dy8PfFCP8Iwk/JzoEzEEfHeCQ9LvoKlvklsDqjmWVkuB21RuG0VFFVVIDmRGk25N
mt5xm9fmUUaEKnvzuXoK1b+c5kzHDL1gTroiUQaU2VdL5sC1vt6fyoWs9EOYwDjLapg18rMxmKCC
xc6HBfmYq5vjnu3GA72nVnAHOFEBEcVYG1xQjVZfUw5SOYHAcCvWFoJ2brkPd44F1cAust3WCVK3
fzLQqiUSrQYv0VxlwkTP+GkUGgPQsvXjk//nqDDJ56H19uDYpBOZgwqQge+a6WobyB43DgESsXfF
r2NGNrhF7V3AAa+VRc2AYYtyqn8Zr1WhIbiDodh/qgh5NvPdnSmUn7VlS2cL6RHt4p0dqRcKcpDS
HXZ8JdC+HqNa4y6x+WUpSEVNw3dEB6zph8yTW1VBaDKxY7be3WAeBWtKdppfKBhZYnXek+KMfmkV
XjzZ+eZjCbpW0VBGWyVlGYoX9LDsedVewruap+Vbd1BZHxgUafOfeDnOKL1zcenTumEUtJsQyH3q
VSfq3+IaqAmKTLG94wcPTcqs3bON6fKIn+GAJZCdWOde2ahcwADcfmp8WO11ZMMfvLBtAPyUn5+x
Oq84CiJhZjdOlAaF5X+bVfO8c0oYybGm0NxpjfNcyyT2bSFgekMTql1a3k3KXYt846zmOG6EKioZ
geemyGTpj7RugP7VEn0w9USX3liqK6rqdfsZSF66AAahusMb/DZQ0SzWKSv+gBJWYkYC7PKKGF/D
uXfNhqXeRtmuBHjYpIQRXDvGqGXz359cikWo+m5uglVNwXFqG2EtOfmyw0TcirOBbjbfOku55X5I
m52m/a1OzLFJZTGZkcK/ok9plqLAs4KZ+4UOjP5Ux2ymgd+toQvyFXQAxreat7jB4fuMdU3xsrOQ
LQ3K6nhnKFrzWW2hnQAub5fXFIMF7dvECN8yYuZ0OX8CAS1B2Kvc6qvX6TRxOjSnAQHmcQD12WTu
czgNHM4lCKEIOs8wwSSfEkNiz88xqyzvowQVTHZHT2Z4MGvuC05fd4NLS+6129LyHEPKcFGG5qs2
sE4DgKhfcVzJfB8G2SVHogTBCIdLmEfbDgw2Kh19dnDL96KpNZwZ5fZo9y7ecJdZZPdglsdBjKUB
PXdPlDvYm9U+znscpKj1bhBwy5yedaJalwWj8WineCXExBZ+BrIHn+y0aALHyXu9VQqJRShaEMBs
RfT4mvTbbJysq3T3NPMeCpW3ULf9QQnx4dyjZqt2M5MvptyiQxpSTvIU+NzUyI9r3UyvMAax8kEi
dTrJ2yjym+1fTEn/rOcK4p1QN5PiBIzviswwj6mno+H/h2Ca1s8dkoaxQCdh81WDpQvFqh/F8iq6
XGAp6wpUKCZ16mP0tuqJb9yYVKkl8NCID07nkOQCDq1APfnG9MlDbApDZ8HXI2RAoX3sp074/CBb
QFKD1KC10fOqEWfz7/qvEVptY/FEPhN7FlSq19XE7HN0YLoXHXUi+mMkKKKP5Nu5S3hH1kYSfcSO
yj9a2Foa71PLOGIoJOTYJHnZYMiJewm42dSMkL+j7B+ELpczMw8fqK/MwzXQ2gzeLPwgVHe6LDvx
YwuKt45rF389sYU2+VEjQtRn02i2/HZXavc8Fpa9ErS2cCylzn18ZkGzgv9KTx6oBa5JS0MrmWLE
xvxj75HrpRj9YWHj37DON+6OiL5rtKAZdjwf6wPdE5D+llc8Tb1fY/DYPKRqV81SsQM2KC20LXTF
yDggy2T4VjTJHAYisgYoP15aBpj/8rZbN6YozXdXzCryag==
`pragma protect end_protected
