// SHA: 43f4f449b937011c34848123159f70bd11b98098
// =============================================================================
// Copyright 2016 Amazon.com, Inc. or its affiliates.
// All Rights Reserved Worldwide.
// Amazon Confidential information
// Restricted NDA Material
// =============================================================================

module sh_ddr #( parameter DDR_A_PRESENT = 1,
                 parameter DDR_B_PRESENT = 1,
                 parameter DDR_D_PRESENT = 1)
   (

   //---------------------------
   // Main clock/reset
   //---------------------------
   input clk,
   input rst_n,

   input stat_clk,                           //Stats interface clock
   input stat_rst_n,

   //--------------------------
   // DDR Physical Interface
   //--------------------------

// ------------------- DDR4 x72 RDIMM 2100 Interface A ----------------------------------
    input                CLK_300M_DIMM0_DP,
    input                CLK_300M_DIMM0_DN,
    output logic         M_A_ACT_N,
    output logic[16:0]   M_A_MA,
    output logic[1:0]    M_A_BA,
    output logic[1:0]    M_A_BG,
    output logic[0:0]    M_A_CKE,
    output logic[0:0]    M_A_ODT,
    output logic[0:0]    M_A_CS_N,
    output logic[0:0]    M_A_CLK_DN,
    output logic[0:0]    M_A_CLK_DP,
    output logic         M_A_PAR,
    inout  [63:0]        M_A_DQ,
    inout  [7:0]         M_A_ECC,
    inout  [17:0]        M_A_DQS_DP,
    inout  [17:0]        M_A_DQS_DN,
    output logic cl_RST_DIMM_A_N,

// ------------------- DDR4 x72 RDIMM 2100 Interface B ----------------------------------
    input                CLK_300M_DIMM1_DP,
    input                CLK_300M_DIMM1_DN,
    output logic         M_B_ACT_N,
    output logic[16:0]   M_B_MA,
    output logic[1:0]    M_B_BA,
    output logic[1:0]    M_B_BG,
    output logic[0:0]    M_B_CKE,
    output logic[0:0]    M_B_ODT,
    output logic[0:0]    M_B_CS_N,
    output logic[0:0]    M_B_CLK_DN,
    output logic[0:0]    M_B_CLK_DP,
    output logic         M_B_PAR,
    inout  [63:0]        M_B_DQ,
    inout  [7:0]         M_B_ECC,
    inout  [17:0]        M_B_DQS_DP,
    inout  [17:0]        M_B_DQS_DN,
    output logic cl_RST_DIMM_B_N,

// ------------------- DDR4 x72 RDIMM 2100 Interface D ----------------------------------
    input                CLK_300M_DIMM3_DP,
    input                CLK_300M_DIMM3_DN,
    output logic         M_D_ACT_N,
    output logic[16:0]   M_D_MA,
    output logic[1:0]    M_D_BA,
    output logic[1:0]    M_D_BG,
    output logic[0:0]    M_D_CKE,
    output logic[0:0]    M_D_ODT,
    output logic[0:0]    M_D_CS_N,
    output logic[0:0]    M_D_CLK_DN,
    output logic[0:0]    M_D_CLK_DP,
    output logic         M_D_PAR,
    inout  [63:0]        M_D_DQ,
    inout  [7:0]         M_D_ECC,
    inout  [17:0]        M_D_DQS_DP,
    inout  [17:0]        M_D_DQS_DN,
    output logic cl_RST_DIMM_D_N,


   //------------------------------------------------------
   // DDR-4 Interface from CL (AXI-4)
   //------------------------------------------------------
   input[15:0] cl_sh_ddr_awid[2:0],
   input[63:0] cl_sh_ddr_awaddr[2:0],
   input[7:0] cl_sh_ddr_awlen[2:0],
   input[2:0] cl_sh_ddr_awsize[2:0],
   //input[10:0] cl_sh_ddr_awuser[2:0],
   input cl_sh_ddr_awvalid[2:0],
   output logic[2:0] sh_cl_ddr_awready,

   input[15:0] cl_sh_ddr_wid[2:0],
   input[511:0] cl_sh_ddr_wdata[2:0],
   input[63:0] cl_sh_ddr_wstrb[2:0],
   input[2:0] cl_sh_ddr_wlast,
   input[2:0] cl_sh_ddr_wvalid,
   output logic[2:0] sh_cl_ddr_wready,

   output logic[15:0] sh_cl_ddr_bid[2:0],
   output logic[1:0] sh_cl_ddr_bresp[2:0],
   output logic[2:0] sh_cl_ddr_bvalid,
   input[2:0] cl_sh_ddr_bready,

   input[15:0] cl_sh_ddr_arid[2:0],
   input[63:0] cl_sh_ddr_araddr[2:0],
   input[7:0] cl_sh_ddr_arlen[2:0],
   input[2:0] cl_sh_ddr_arsize[2:0],
   //input[10:0] cl_sh_ddr_aruser[2:0],
   input[2:0] cl_sh_ddr_arvalid,
   output logic[2:0] sh_cl_ddr_arready,

   output logic[15:0] sh_cl_ddr_rid[2:0],
   output logic[511:0] sh_cl_ddr_rdata[2:0],
   output logic[1:0] sh_cl_ddr_rresp[2:0],
   output logic[2:0] sh_cl_ddr_rlast,
   output logic[2:0] sh_cl_ddr_rvalid,
   input[2:0] cl_sh_ddr_rready,

   output logic[2:0] sh_cl_ddr_is_ready,

   input[7:0] sh_ddr_stat_addr0,
   input sh_ddr_stat_wr0,
   input sh_ddr_stat_rd0,
   input[31:0] sh_ddr_stat_wdata0,

   output logic ddr_sh_stat_ack0,
   output logic[31:0] ddr_sh_stat_rdata0,
   output logic[7:0] ddr_sh_stat_int0,

   input[7:0] sh_ddr_stat_addr1,
   input sh_ddr_stat_wr1,
   input sh_ddr_stat_rd1,
   input[31:0] sh_ddr_stat_wdata1,

   output logic ddr_sh_stat_ack1,
   output logic[31:0] ddr_sh_stat_rdata1,
   output logic[7:0] ddr_sh_stat_int1,

   input[7:0] sh_ddr_stat_addr2,
   input sh_ddr_stat_wr2,
   input sh_ddr_stat_rd2,
   input[31:0] sh_ddr_stat_wdata2,

   output logic ddr_sh_stat_ack2,
   output logic[31:0] ddr_sh_stat_rdata2,
   output logic[7:0] ddr_sh_stat_int2



   );

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
EoSs5lZV0FKTe/cPbFEV/HqGemZrb0bulUDR1IsUUdIyrTkcwD9t2yClkVZG3Key4DJJEva1l1Xa
bv8honbHn+TNghn7p4Oi7pg++fkZldrlxsGcNUI8BdlqlqP4Fp1njYsCWx71tz+QOrsjNF263Czv
BGUoAi3VYITZzYF5ruI0rUueFnA0WUvsqO57diDZfrQWWVgi9sbUJ/SeVrFaMTQkpkUu3vkX8Mkj
t/f6xVbzByMaIHiGDrezS2pyG0+KIe96ooQxRXPlA7o5LoR8mCeuhyiHF5LHK5dhHJ5oXYK37RIB
jAmC2JkdYynh4VZqy+F296IwMfAZbHjgafeD3w==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
vN9w9XH4NBgr+UFq4IboKfmzoA2u+QcSQWXWWV5mmiajZmzRfrswt/jEfn2N13oIjZSqHIPTDjLU
R8/g+5AlPGViePFjX/64ZclfmY0GH2jpE51lN6OqVJ3laGbExEU7j4uso7n/pbTbcLvTQxKoAeWz
L6zO7AXRxQBjsKLT1+k=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
FrBvzGzPvZYY8DOwD5l5W8IRnwWv1Fb5jE0+g82dcNC/0ekB3AB25iXzCteQrAbJXXy4QXkDcdFS
uQPXKWQPfNHF49RZ2i9Z46v5nH7KE5LCTUQ93ilrnC1ZDiKoOunr3u530f1FdORQfnAdhEgkjBH0
Yy2mzrBxy0NO3Ak2XNI=

`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
nrtYsdYfsbrGoauofF8TnpjfHvtYqlIKPB9W8Fwc2MylYIGghIaM+SGbc/fdpu8CSEPVX/y8wv/M
GDxGU3FSOA==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 71232)
`pragma protect data_block
OcDYBRWtC4pgyOYa9nUZd6vQU2WoWcXxy8tPVm/TDz8bxBM0LjpiYXtWiM626MZKrQcvYMtJf5Vf
5jscTvhyz0odktosQWTBFgaHdE7MqcPao3BEq361Gqg0xtrdJ+ejafkurLd0pPBay1718TlAQ9OD
HDE6lHLdc6zbTr45t5t+BiBDZ3N7ht6KeTN75pB6Me8S5lU3WB4hLfVc6HsCKGohWKHy+SBe8MoV
xhaz2niaT1WiQuYrSiYss30umc/ERKosAPCnRr0j5/hdPkDu1UGLxl0ayKVq0mw3DNu3V33Z6TaV
1WmM2RNBeRk5eEkuiFxGd+ZkjoN8EoU5XDqmip2+HwtuEfyiTzVz4YpXO3J36oplA6Pb0cu3Bw41
dSNI7w6IWqJm0EqaGaFFjNZNdKK2zZJAkW7PVCq2qtTm1Ehv+zuaEDlt/bbxeQDOvz0vKQ3z3lda
O5KhFxM9LHHCy+qInfTIJ32fzrLAFucY00LghEufGi4nh7+3UQhOdw9EOZJC49+cXoyk8Rqpik8g
ASjJEhoROD+Vms2r/QuJqpaYpWTQPIoRDZeh+7LURfORjfdkWxkQFZcjBvrRXW+Tod0cuoE6yJ6v
ajmOQ6o8roLqhlPes1bNuVpHJzVFSUCRDQilJSK9S4sCDFzYZMWmRxxQDTWmyA6vaGB5uBiWcVAV
+EjV+dpHVGxgyyeh3XxETfR9HR6uP/KN47F+//xz4bnI0iJcuedet6lIYDw3f9mRAb+dLwdPw54S
7QYk8mijnva5SbNORFzMR98/uOS4uTLIYT9jOrShVtjSdXB9FhN+TiwegHInfcUslanCFKpImoxP
GgbB50EnE2YeB41tlRjjPrLk2Oncg06nUBBNE2by2wdIHfm6nMab2v42K8B1ialYSejzrK7JPYhQ
UPWsbZUelk4ePMqOjogyzhoj9Tm9gaaA/EF+y6M7Vsm9rnDd4514M9BJ1musi+kGt+wHUBx73G0h
Q78kxjx2GYXmQFlngmpxKnWzgEmE2BeTyNwWjjcmCW+k/7eCO12UTpgpY0rw9yk0/3bgdxvAJhl6
y3K3qh5ItjiE+QmXjuO+BCL9YQeqhunu7NoXk3FE/XiUUwL0oPqAlq5Jdk1oSCVZuZ9Mn2ATkkJZ
sTzj0g3CsrE0ixxEmhvm6U2pRqPJdvy+PuzTGNyOcp1SZEQfMKIrXyLAVDtb2UaAjQ0U70XJ0nPQ
EqYZek7DrF/iO57p8qEm+gNOV1iAVo2VKGHitZ3hnkvbOrL6y1RIzIIMa7zFyZgM1QkxzOxvUqh/
TQcFzIl3wUfCZaf9EsnvtBW37wxqPJnN+imFsKV4DDlmazjEuTzu6yZsHOVIJioKkgzDC9ocO/uy
2DYl6tGP+glRqJUn51dL9cdbp8KZCXzMmJdOMBmmBh9L7MMzU15alDXbYmEkVLOZberJSs82c6VA
oVgKBaNGB1/pFUBiCgoBdjhEsmTzT8EAuz+tyYo/HRoXA1C3fO79Y9YeTvGLq8I1BVmmSpKBMkWF
mnLD95EAsrkyJ4vdpcJiiJ8MaxAZYVpR8wwKdcj6e8T4RFVVIQ5xSIdQeM6s0ZuJIiA+9rmlYNnl
jt5TQxtW5fO1yjx1N/DooHxEpsfwqj+7ku7AATjSVwkSslADa+E67hQH99guXWGPx/VbE8mls+zq
pdt6YuuA4uh1dn9t9A/NkIxfsaEyrd7ENebtfzCwNu0Xzdu5NlFthfr6QgdKNs0/fkEgeYHRXazX
ZtUdctlmQTYYnGQ9enrRBpCQF0aiecdGK9s0Y48ILeI1S7N6SNZ2vvGgGdePJcaGNQXP0ZQuwaei
aiFibgPeFbx3kOBq6A2PhoDikoLIQtKKFtuGq5yi56d2HcRAiTFzC5jPPzGuBjNtxAIlDyUTy1YC
9KKCZWoo2dpHZkb3Nso0xcOUZQqC/4upIR0++c8oXWkXBgQ/IWr+yyIJ6CBfqSkf5ZwogpfQxWcP
YvWxg8WkyainJKYKj2PK2Rh+Y6RAFXFD7jqovlsG7E0DtvEH8PZPb/BJ+2Mmc72RiXzMkDaujnHk
C+JXfIYlwmyoStjij68fmKf1AyUd7NpLpgu9rPiZOZuhXvcdxUKpX3tL9ibw1htecUA8L4yu4U2F
iRvs1oOZACe+A973ECTRpHZDHyma9fYyBLk3YvwZ5Lfs49EKQn1BR4BV9M1utWLlc1SVNP65sGxW
fVcLS4BvpOjgFsidsaQ7QexlY4JPOlPSggrpEIPFKlusDhFoatT06HODyPLezYp9ROVH25JBLaP1
jCNcChF51tjSSfiyeZ9Eabh92/kINdsnnxCT7DBDeXyS32lni59Li6TJxCrTXDsoSQhBT4w04WZz
rP5gCm4PM4ZJq47mz4DiNRySTwSq2MowvAO5qS8BSvt9UU9amcRsrKYya1zu0J4YHwmjkCYUf1D/
yJpG4rXgEpn3ZZCWron/vAacrx9UxvAh9qJF5WV5OfAATBT7Cu/7yDMPjxa4jOGfawy5LTw1HbUv
SR1BvI6yxQuCVFvWQ4w+coKmaN2jsrZItwDehe1wrDQPpytLHGOdqkTaT7XAM2XobWw+COus9PU1
FmkWhJhScBLAMT4Y5chJ1YAjPrcGdDtfCPZEkUWe/o0cvZ29hp2UEZu+SPvl+jNce4WU0nG/N6Qg
ZcQXp2lNGSV04SN2Fe8PE8XA42HalW6lHFb0h3+0VyImL7BIwFBPE7Wgw3CqPQe916zVzhPqOTT3
gUyCnaUt6nBadDf2eLpE2/mWJLnAd7YsBLWHJuY0BL68dv7v8jwh/8Hz0+Fg+rymzop6CJSHws9k
kHF3JEO3DzwpoknYMaCc8iVJLVgkTogpJm0l8/i5/JmA8Bye7wRdmziolAW8Jjjz8p6F3kNvWERb
am0L1oaNccgZF3KTEekQHc0NTVNiMFO7lHzaf2EfAOiha7fBV6JgJiwj/0q0cUgZLCFMNmnpvJmx
SU9efw656HxploZLx2nPMUo/hmr+4zyFrxv4hI6rclofp9VG04ZJSPeGbTrkSIvqPPOrgx1PlM7K
J8ODm8hGZ1r7bV6W1EtnErI+whBiXr07tFpSh+Rw+jxqH0nhN6J/3716+s97VH+TX9+Du7Z5nl7S
AFGJ0x0WeoKzxFQkUDNnjERWfbrV1JSDFG7vNlfguz4Ewb8+xoZj+VwtqUsok34tHf3AwpkfR0CC
a3D9CXsCDbE01++1df7LKiG37QXg8YfbV1KoD8S37MMmShATkGOYWr7xyDzVTb2P9WK6EckCdR85
MWjGPzsBhzPprzlPH2uRIUB3Jz59KVG6Z1QSRRyRk2mvsuY4FqotqCLFfzB8sVTvnt2MwHQOS4u7
g+B2knYwK2A1YINN7s0L+YxL4buKDdEZI3cIn4zM7H207yLV5Xq3AKkT3bcbmE73K9HdXP1iox+e
TtVh9NaktZkPwJOR7cNsC2I5UgliMRrj5JLyhBcXiXvlCpRlLKom9O1cBdDT69pkPa3HIZQ+7nBM
c4/Ir1gjJqA4yFvkL4xiE15xHvn5Cl+QIBsjwrWed0PV3soeSS8UObxGw40B7oxcpbI54IVSzRxM
GP4JUjdbTpowFtURY0fnebZKWG/bhciIDq6sF3mhafFcw/PUo50kZxrKsFuXlfk3UuyrkkkLC8CG
QKSYShpxCdnTPA+XxpdaNfRYeTfenJrNY2sg2AHVG0XBpicGPI3g8rCQhZc7sr9Yq6R3+Q8baz/z
dyWxufvrKavQIgRkDPSPLDn1jhEsfao5OVnG2J1qsEfdgrccwZ7lX/GL5ArAsv8Up80rSYgNZCit
8P3q9bFmcOMEO6uroWHCWjNyiza7dPNsvcjWYy695qw8WCJ1q7cSzBeZzybNGFp0txsd/NHtDDLm
9hWnc5507OLHt7BSEVXAo1XeQgwI9f+/zUQTZwDyrzRhdJK8+ckZVKjdZWWgEQzCs4CrcHRZdiwo
AooPHqI1W1ByZcDPW+BfS65+/sN26hAbFNMVB/xNClwN52ckTRR9i//Athue7OdWm3zfhy24q41r
/Tg8tgQsJRuG34Tx8CvqEb9TDxZCBzG7GdFM/DE3N3AbOFdEIHFWEkpLnVd4r/Ibx0tx6Bbg6phR
5kJfKvIxbOxe8yeIRSuK/ue0HKnyaohvEfYDu1fkli5eHf9yPM/0gRFjkAirmla/DxNMwLy0J7iB
ud1i1CQIUd2NenSUj7S+4WUrMjrmZ8pF3K4K/Z0JMGIT4AuSsGwdFOhTYN2WeCcJfOIIe4vIkkUT
q2farxzblEQ4TMootkaYVfDOPyYFyujfJgpvaED6+hp3WWkvLLpEc7v6gwRRGpyG/Ei7xRE2Hgsd
b0y9y0PQWdOmoRq9slrS23mXGqnlx+jerpgD8cHgWAO+A2neHSXoECemURS2VDOk2lit5dvZg88L
TuVNYIp+OAQQLR2nDfnx2OZEXvS+7j8Sq4dQm0p0prZe9ch4aFpCby72Y+cFdHJhInUte+aBVgwV
1Lzpk6yDOoPWDThVZHjsSM6B31hiUs6j+0mTkNwGoDHHp8GfgLRGY9vEUIYau04l4dqLHCFzu/oN
SzUUwTzK5nFC+H/FjVgibQl1+ieXjowcC5MVJUSzMmLwM/Xb0bGpSsRWea6BpR2bqGiOxad91ibG
Ss9eXhdzPcS69dYnqw91XSYH2vmFJ+jipCrNTBHoj7B8TcK8weXK2PQCuUxGfz6bcP5yj0HSHyhL
lfsWJOG9jD2odc6nmEhELsmNDi8aZFz74H6fVdY8bI4JWxlvbJYrrZOJrs+c7leZz7wYV0zB6hTP
27B+r0reJkY0IhPcgfN8liiOGyhCmImM4OpAX/D9aS4M8PaDy0Dj8rrLpWo169hEXY1l35o8n91s
zVpBDH/3QrsUSvLYmnOyozmp/lQHxxEw1v+dxcX6oUr9gSzTucp8S8KT6u7bz4d8XctIXc8PEFpb
c99VuzM26moNP9Na8UIRmVGAQKwx6sMYyWhFQGeywYlLlhui7StoTZv9f5tk3v8EuA2OMIF/jH1T
xiEWyrY+YAFB0hSbpUypK1BXrIo/CeVZMprbreYW6jjA3XdpVCJK9cubU8nY9PMUNv4NyNgeujG2
7iGE7itIGOy5iPSMlr47hD68hJFRUS87g7UVOMX0wnkS68Fq1yXTh56PR5N7jLNNEiNlZoz76yib
6+ovYrF9lYGkLivWA/rSraJvHFveClyf/8f4WFWD3eBF/8wGSdocUq/vNAoI9Jw/vRfX/A56mpcF
LJBPJS1tfJeFlIZaF0+W/8v03Ysp/zHau/v5j2WjZHK8bBcVo6t0KDiGAkcZ3KFWb2e5o0oEFUbq
+kv9KgiTpl39fSAM/8Vby/NP4gQ5XXi0y+YesfSkx5rUjSI6b6TEiVH1HtalOiFGCab44YKV639Z
spl9zaxZXXqcTWOG5GnDLWehCpiPmhfXpqTd8Eo/4kqljpNpZOlu0AqqwhCHFN6sf40/AK5zT2m/
HEjC5CmfW/48HIgRzPcuFH9TZj2SeUY5hZ59aQexLtQrH0B39v22aoV75/AeKDNGrpHxLeSXX9XN
qStL649+G/xkVW3tAqMebyQn/XVGjHRq1BJNhYCBcCb5oxDrbzf08dex/FLz3uRS6fL/BHHasFnr
v1RdvZGR++qkHBdpk/ghdU/WIG8aw9mWbU12CEIFwpc2IxDaPDhp/hbDyFdBYVPZIXPdFsBGcuY0
VHgEl2QeucwpolJeCi43bV8m6SIHP7eQPE3JlUYUDRf3IYpYKdReFpkhtKACKysffjOg8tnPY3mE
GscWQ5gpuqVqLi5/KZNuA6E8i4V8ivU0/kLtouLGL3xciHssM6+U7V+COz4o1ppB42k7PwQ0wGTD
pC93ehNgEqNJlQsVAGmgmtG07CGP+oHQXT0QHMy571ejyR+34w8T7leUC7Pf5iSR5ppp2yOAhi7k
LAlCWheEhC201A6HD8m3tD6Z7vjbKcjwLptxQ86rPNSuLQHumt1EijFGo5pgUiN4f+wD8n+TnPfs
/6cqVn7i7jU8IgbWwmHEkA0h6ttJvSW4cJczYfA+Cz5azWoMk8cQo+JoX+Efu7HMifDRGImgQtGS
GMoqhUvE0+pvfFq4JEjinvVhxtVslhmxb3aK7mgYci6vGZFmJryeleog6lhutMStZpVltwzrkr2V
i/5JwsM/oIwcjKguyqynSoj0zpEzibZPYTM2ZQD5yIai7MG6XS4Btkf0JoPQW3Z8qB8oRqG8BOU3
76/eQUaCIpY9zfSYGVeO1YwBAbc8WcH7uwmsH+2Q57aTqUeT+cVfQUjsAqnE7PNnIvSqZSfXWEdt
mi7iEFXW9hmwmyjdok6U2u/7g0uLibTeJgoQ678Rm93cyJO8L02MK504eIOllJ2rAd5nxf7/qqqX
ObtZRmRaT2QPzEA0IGry9TUheyHLZfNGzIBYf1JD/wrzYcniippmL2Cbf5vF6wwrtYcRthxUXSBQ
f+vPwBe7kbnBlEGqqm5ucEhnaOMxQjvKJ9cOee5SDRH93egSaG+VoMC4N8FKtRKjFir5hnaom+h7
Ym2OCd5XhoPz+QEwWbdnFlpgUPOU41bJI2JKXvmNRqFxMVzbhdzt72VjbwvZD3QvJBYuP35EzDkQ
iSj8ZzF8FdViXbqVVKhWXg+2sHAAmMp2m8HKjtq0kO9rHQErp33o366hZTl0hXYhlA7ceeCoL7ct
vSjkkh1ZVWA7GzyoHgIZxswDbvHY0Is23bxkXgoByAJuhHRqpIKx0HCkHjVDAuTvd2MtucnVqehY
Na3SOYI8vM4ARNeBk95/6miMtp7oG+Svw2AjpL1dfGPfxKNy4Sgxosc/tIh0i8+kCSZOwEHVZ8t2
9ouX1kRc174sh/q67l0q+8ODFtaIaLoBo6YQj+KB6G+KBC3CALjRcdDG+JphLKizZ67btVQxffXR
RbF69RVioj2E1fTJ5ScPObmOkh0U5C495JidiJIV7LRkUcWH82sRWpIw6iMGykw5YZgZBonvlU7b
zFVQy4M8hLaFbj32UNqUtZuSVA92zZLWjrKL6hL7S5S25SZm2nvA0SaZVYv/pMyo773j/VOhwd6S
ZCDAIw948rwb0baVJJTDVq1NjuY7MwarBpIMDOA+ekFLP60xOm/nLZWgsZ/TqdrFqVXoopr/brYU
GzMkj+SuZu8/uNcfamogIegNSFVDZIQHkTQdaZrqTKCN7Zu7zk+LpCOgsoWOVsvcoKt9zLOoyDO1
nRPGTA2IatlxMXHzZkZuBlmcaUVQTc3mHO4QjzJaJzUqwfPX8ljBBIFS2zy0ko1kW5uxD+t0j+uJ
ASTAkAqdkS3Um/F0JQltC1YaV1GHu5Eol5AEwhds1gWVe8jp4g7JJtqKXjM1XM9ZWf6biLRUoAhP
d/7G/KmaWZz9mHD+kROUt5i6Qy5QsYXxxlaYrh3Ei4oXYI8FDxk2w8pq357s+KbC5qYPuWbzTkjF
oI0YPNNzDnFTYjNpiiK+2jHxMRPGp3qgEfzqxq/9RR+7i3CruQc+zBn8X4pu391BljG9VMEtaQPo
Y2ozj9wk4DiKkQIIkGukuxxIuWDZhxZJpYRWwkkIUSLDIK+lDM55wto5pditmxjzAJ3rzQniXIjW
PbiBzT+6vGIEsnrK3XXNhNMZjHzGJc29WctuJ3adXe5D1BzEgseMyHl+TLAo7nDHxa7t2UI+vQBj
lgWNXcNcze+2bKlPybfk7myMU5h7PX5i3hiv6v41ZpuikeiuNHkD76PnmUlDdmnp318HfhD2tc6F
eIR7Zah0T555j6lwCnzxCFXSLwDHREAbB7Qy7Q5DvANpItFCuA7fJGXDJS2hfiKrAuuHpzC6hFzM
IgtnotWPVbW5j200kEzqXXCxSlvQ7pwDos+G9aTWEn7smoffIp1dMcXHhJTuoUp/HKMhfpgGAtM7
PrvuMg6lv3wmdHQbQdteWGVhepcOQRBbAsY8pSgn3bRizBbc/sIeoVUdjrBkVsPUfw4s2nMTMxAB
lfl+uuHiC0W8jm1e9AZPQp8SSZ1sDZ0jOUl8MkOdH7VmEsr3TkVH7Bfelg17XZsN0LRlHyBk+OUl
fZ1HT9kzz3VX1vvwIqvX5Glgejhxu+7onWEQP6Qohs91n7ipsGTzRy6jrLYqihy/jQrZILPUeXHu
C9xMMvpgxsW9dzsotUC/+GAseikGITf/Xy5ksIahFoi9SM16ZHpz4asGyWT7ISsftHf2SEmdG00H
0HHsmphgbpXF50T7cizH4S/JNn9IlvbsNhtTeKqJ13nQ/LXwjsGR/fQYouAeNPQEj1b7HigTCRoz
YhBmFO1TrW+96VE8urZ2XsAqBqnI94nDgm4/5uX5gjop4S37PFdqJRkcT2cCNej4fuNQz+mSM8TG
g4uk52a7LSq4GjozW3Y0O94dbAQGh1QDA1yxU+ez//8waMH7Z+62h9HvZc5Rl/M4bR2ZRcfoJoxv
3xVMyWwUAgxd+QZSHLjfxpmKMeGT/iPSq1XE8MIm1hXcUTFILKgvknoyKqB+KXupbo2H7DaQxv9P
b5HYvR5DZutZ+ymjYAJyHLYEo2ZARWRTTVEeyFNcH+xQYuxl7TKDWPNlvdGnREOGmY47Ns8MCI7V
jQdIQkMXFSZaAcPVajNW5wZERDFrwFL5ULXudtq2fr8YELu0MinRM+Buh87Jsjq7tPxeV2Nja1Vg
mlmFujrt9u0yneGtwnkRXb1gK0EMeZ3K46s7mS9RUWLzi960qYaa206Xh74o7k2kT51D00WQKXZ9
upqVR8bPZbhZbGmIWGnSkZwJyZ01amrZcvvz4k48QiS0UJql+HD3uZblDlsQL7enSooacx02vdME
afNjdLeJe0LWjPjMr8jVcXY2Gk+J4VJkWHC8iAG3r6nCcC2X1QmWfdV5h9AjgfGG96EF7j+i2yUC
f/F3fSOOq0GjCg76UzyeraVNZ+nrKwm9Dfbhct/bkzIg7ZTR42evLb2rh9tZ8BZNgLvCmVqBHhrR
9Mgi7fbSr+0qLwxBcTs3sfvKrR5Kls0icRP3KRuK708LnyHHXGyg76JrWxBEPQ1+jjWlFHGt9be8
OyLwlPh/Chmoq2VNJbMmcb+bSCyY/RwC8m2Z8RwQmCCxM8CYVMrxuwfAARwo1xnSznnKgtTUPb9f
WbNGVKFQdvj6VvX1p/X3dDfWSZm47RKU0964Btk6eQ3MMN/j8ocaOAGi7YWSeqRNLZJEAMJK5QnC
Ib5tinfjOx0MS+TPvgOpooO1YwYGdMad1yV51+KsMxDXv5ljM1mwJMPSkAaFVRVj+Jy2zH/BK/14
eDXx4JGuBhy/6iUDcZbiNle9ivKiwfJYfGH3irVuxsnP6H43Hlgt+B3BF4CDFCLAIHUCGLu20udv
Tl9G+uxAh97K+rJydH/zRHXZa7KW92NhWFKbJIFtr9RLoI24+SjBi5GjyZUU4HWZPdALt/ZcOAOJ
TAx/u7UX/AaZUzJEF5Z1OX2uWwUWjHUOXTSzJWg8GUwuXRV0ZpkTLVgChZztthzR/JTNZQNyCKAn
pDJf0rf9mwQHbdBSq9QUKth/gXbP0+eaHHLzQNP+L7Yh1ZSCUfM4olB0TMZvRvcPSUDcqRYmCJlm
1V/7KrHtlhrt9zCfxDbfZ6Pss1opoQMbg4dgGN8S8qSWtPbR+vOWOpU1+Xh5OKBlaU/fQvmadx2i
jtS4e1Meyc4FEJz/o25pFyKjgUGsZixO7P6qygZPbJXMHZQnJcvtUPP/mcmQTZ53/SuRXmbpIvb7
G7BRAAJ+yqBI8oENiULIFl3yFGlDuPJq0LTDmHTuk9YvOhfiqqIeJOUxntRA3aQvLG/x8M6mTuDh
HdMgJRRoRSbwRlHDaEozlQ/1c8Q0xfQsfjx+mjOMaPUghUnSMWTndoKKzFk22d/EwLYc9sNv/owR
rFfyygre5ApVICFk+q7W+KbGeZ87FsZkwN9AAn9flGj71Xq70BQsFkIj27yFVd6BnQw3VJxyzdvi
TdDt9oEDLCCvZvGqESmuAG9RAK9PX+oQcg54j+hqrjO7/JIi4hItzHxfyziAQg1IC4GDGFygW/A1
nC2orUulM7GjD63S1YFVlQOUDiQtrWzcRhV4DbvvOkUclXL6P0JkWma4tnH5m17ZmysynCa54/eN
f4+O9BirZ/bS4ULSbqeaatXdBQxqSY02Uobt5jv60YoWPRL0H7gzI+LuZRh3fRbHMGJkteYpTM5Q
CpJJIGN7dG+YVAr2LndNpxOz25WsyRH0ewdPZT6G9GgnuiCkuD4h10GdPIxI7yQQBFFsvGD+WdHR
ehcM1Q2dzr8BeQON2VIn+mWfdCFMk6Nl189OBYhPpHdI+lqyVVMYTx0dBAhiz1+dZTnFtNoHdxHF
N6gONegx1jc5qd11JnRbOJxNt0358oEFFsD5scQs+KvkvI5cOU+TGiYlYnIxmwPwLPiTR7bmZuWQ
7noe2Ujz7KnJjfNcpWHBfbs0I3EUrLLsBZpnXbQzPQxMAR8D1Su/aahB5Cb0qJ8qHlO7i4GqT41j
RpArYJwCICRS28ODxCYH3i+7963KafpnitwhoLPnwsS6AL2XL/Ay19kFHzDBVErXHQ5azI0+Is+i
YO1xfoq1tOsZRoc9J+SeZtGapWzwtVUPLKjWLo4LQ0c8AYr6NbXWbignn/CkdgfKIg1R4U4VMPPJ
XGHqQ28WXBOwW6RaJF8NwgGXc75smHqnZKvW1IALY2dgdo0cB/za96zsrieL0eH51dS4QWt8gSMl
CiNgnk0XaGF92wNn9kFrpboECgCzJVt9XP0O+TskYUvf6fLWDOOAcEyUHdy+WDx/GKFPLqEdBTtz
FxWfEx9L5AZDwD40dl2P8bVlarjVJxFFsEwWUEJ19BLUlRoKsgWpbLjc3fhfSWpqsXLBlo0DSjoy
lZwcDpqHkP2y2tS4og5QWmgbqoAMK2HUborlNW/gn0/C62/O9ZIqgXUEyeHsmu5tjcGUYas+Bh0k
KyxSygeFOPb8P+zRNopOQR55EthrIOA8Gvshf3em+n9Uru0LKN9zErRbsKv9GeaeelYjJR/3XWwF
PY2KpG2TILfGFjNdaGuSzeZzSemGkVrDtoENS8gcmQM+LQlfOdcuampjvlaWzOUmoUXwQEoUcqTD
b3pZViJX9mrPzVBbj3r6jJdmj4VqxuuCakGyE5lV0VysvEa+5GaIYmUkxpkeHlP73uyF6Xa036pU
SOK6nUbP0ewLMIhymqcHEvkrtQAyho5IPG4apxuk464++dhy24M1wuGItRBdYNUUO3HyJKVySvG9
RVtw+aOHMiL6ctV4Js1dCtCWTToETwa3k77ij9glHnFrpH4Vu/MfheAJ4PfqZ6HmoTsEPJw/Ig9Z
9D4jwmlbST6bLYUivG8V2GCQwltC158hsa+uVw/NJETFACk7sJnpP18Z1ZLfWqveypOS8zljP+8u
xrBHVUPtyesam/SplYJirMziFP5ZWhNbUwz4SHcFq6RFvY0oIpz3hlsXaUYSP+WgkO5A55LBkRD1
yIjfqFjFIFeN8CFY5dXrGrGdUAtHzJP6Q+PSZlTyPglni3H2+IQihXlKk0mFnU/WrzzbPcp0ZXsx
GN1BjCyIDXM76LG/eEyi6FZcDTqYeLUIdNe0huxQCx52tdHpMlBaUisScbeyttqTOEEz3bTnn/EF
CfVZMg9a9hf8OU8wB9V8hVuvLnQfwNSvvmJZukl8XQv++zQe+k4ty8BZibvq/6LY7o757/2uSC8m
eRne+SGb3oRo2uNG+wXNSltbmIsEPifu8MIlKH3c4OHn3l9kTIK3YBeYZe5Qw9rjP6qaTrPus7YY
ISYY+pwbhFgcaQOALYmXoJh+qP2Ckr3lyZtXZf69NmAOeULcrjw27qy/brtzIPyk55FVwU0YvIOM
BOBc2NMnMSQIImuih/CZv7D87agkT3yd4swRslyrcWqS2AiNWpAwKO4LJRHcnFCBsxW+fwbYuYA3
ZXz1oP0VnUmJ/hkk9QpXp3o83z9cyIEiMqaP0KwEuWtwkIXNHKLfk2lbRdQqNA19y7Uy7CfaS3Qk
ENahTdp8m7pVBT7KXINelFLRHms+v/nU3wnOR9Y0OEnK2keNtnW1z3lPfAXF2YHg3OPOM/WbOwbV
1HjgksqN5tJHOh4Rr50Cp6aPFSF/m95nS2JJG7UeNJjn4gqDIVAnGV7H0XB/wzUtqnBzDza/K5+q
lCqvJyZ48kJOW3vysaZlzJnU4aOlZFaVaivTkTSfNgl0+9nBlJA1HDYDh8gQpEuUAAngsov+imay
IX/++M8jW0XNQTk/p+5JbBPPgZhVuPneBdQjZtxJggmjRJtfb/6DXeVWpCT5K9RCUSlx4/HYcoiQ
NPPiOS+/UXZ4WVvqyFHHOFCVlezHfAVUC3yEhT5CrHgULKMeqXZpufAShr30fYtsLmGF56xPuFlN
HlBejmfqfwQk+RNq1hv+eTzS8slzmfP7WGmNoLRUqMf8rCuqDvXQZNFW28D1b8nJhkjb/lr+5zpZ
IoD9ii7AjzEuval5bY4XYMRhcvu+EYYfNenQAcBvelnxi0vKJexjFEAkFnecBCS4dlBZ4GiRTK56
yfIWCDjuW+n6xjzK6lc7rLE5c9EjKT7yAgljhnlPfWGKUUqpHDBZe4XK9YPL9DCOhw0NAwhWw9Gt
9SwvqoImbQk6HAXz/LD8CpcRERDSPKnZv9R2hEKe6nSswhchwH4frF2z+zF8apnVYoHNNIRN5RYK
YmOIsloJL6ALvvDnHfbWokdwHZXqZ/ESpYYbCy3bX//XPLBveah9vaj90gBIh9fQrrJHwHoOiwD7
zQUnRtneULSX0j32RBt8zRVIXabAanFc9zoclf7UkjqnU3+xhkBTo6CeMhdsRDRMahSVqcBib8w2
i0EJxwMnAdl9C+Qjss+kAiOSnyxc0veaXGN1EPpDKo4OrVp3Zbu4osPAhJEaxKR9AvhVerAiPZ3f
BZ3fbzTz6Bz/cKFzeT4qyJl79tFp8VZvPuQ7NIFsqgBkdWXG0eU+boUEyTdsRUUIaeJR/h5dgkBf
4VB46TKjMHNKWNpTVyN9S4y+Vj/+iMsMjtMns7lVdydL/bJm3I7NdNBMjoZYFkKjjuewSpQQUUmj
cF5K3sybsU9oG/DBDOajOGbx7NNH1wIREKblFLDJx55TOq0bajGUes75r1qghXhZBhQxUcPnalyx
F8gmQ/S2vpFpbhcfeb44YJNmLlOA7X73fPxoEI/0rXv8w5E/fWaZDxKXpByvKU1eVSLj/2lSvTjV
Pb7FbCk+n7Lt4exjM1ZPfZkzkYnUeaJzIYoBI0ED11xhE+UA2O1Hy8hG5abhHL/X4BKjB9fp8KY7
ITcV6NHR6XcIkowD5SjsZmSLyUTyYU1FpBbJ0CUJpchUK8gCiuwmT8YJtMwwbzyeoUBcrCRgBlvI
juDjQwh3zCIyUbOjJnaP5ahrotfOHLSdOLiDRvGIti2iDzb7Fz/NdQsaqlv6RUVQOcg+7qRbLotA
nC8HL5YFwTY0KfzJOu9nZU53XMfZboEPnrzMBTMlL10EvhYF4Y28aTBKJUTGgvzRzXvMb46bxuLd
mPSXwH40ym4bGA39a0qkZxqJVyYhLPlogQXKKd39eqXWp2vfW9X8rC1GiO45LlxS2eyI9lCY39rS
XAsw8tZWNz8odmV5WxtH8RqtQ7rSqc/1qKA/ieuf8WsxAOoAM6Gguf9x5HSHhWSKd6dQzQclI5pu
5BTPiQsbHV7hElCDSY3ei0RR7W6iNnxSYsdAJKQiOc0qIFULcvG6MNbTJh1SOCOJWuHU/21OM446
1CXur97qUgNHHjdfU7un6/tGgDx/qaLz81QRL1EKAP7+RQ2nVy3P3CbU2HyfV5rucWyQh22C1BP2
vyPThkpvW66Cgu0I/aPUu5PQ77qf/iSjPQSDdjwdrvnVC39gJMTwr5YjvCiueYEtKEyfPx7a4CTJ
LfS5SJvYAP+jrXdKzOjKAsOmmVE4KPAjfCc1sgSmUQ+YYuzq/frBJdUtes59H8/WB+ebIwH8T9Qy
HX6BVls+/cXuQY6a5qwtR+tWFGhUbyDMIQUjR34GSnkkfBCCVJ/8WpIVfELx8hgWPnyQxoSRI9SH
LICpu+cTbxCozt1LFIqFMVQINkAXKdspVL4gF/bdle+DsdbIFK06W6jB+OpXHgKsL3SBglZ9OlAU
Is3CAruOXKRCtjisbUCB1k2jKaTJ6D+P9gMv8vkhC1Q4GBs3UKpEfl3HOtSfu9zRWR/8Q7dqL0XB
LD1RzSMlFSxXUw5TsC4/YTUQqvWBwnyR+lKOhorXSLs2isJoFDSm11d32y2GlMOwn/7MhuoU0WzH
/1FyyBZWsZ5zj0VLTWzaMSiX8ewEdlrQ9KzyWLAbBSnz011IaZq/TP2hjaPhgf8u44m0nWNvnQF4
jKZVjgCE0imEaUP1Sbw76EUlPnBYbG4O7X5uXlZp0p0UY688K34LQN8nfqEWpGuFQ4pWG4tZzp37
OmHf+hs3HNOxnZjSNG5yhcf0eqf4/rsKOxY90QoCv6uM1QRTHTrMmb4/T8J/kRkxrsNA2BF+A4Dz
0FzayPG6k2tgPiaKS7NjYuwPhZuIKuE/R4fSfYCc7QUS8C0CIn2hFlzlnyl18LmtDg4LkzrPQKe6
K+9I6k4ADjaVYmP+9ThoPVaKLOKXDS5nQRwKzkNk9JWfdhRkVlDBnpiGviFyyNqnEBci6lHtR+P7
txnwnKpFk094cX2kcJv17gGKlO784c2wFh3rlL99euLNRVt0tqnCvpzRzuxGTKiYNNRCKbKhzGy8
Gmp9gD9JPYv4TfnoNXAam6haWT95/xSsfPnAFgeY9koIg8OZduiqLkGxVGX+E1hPnxbTD+TV6D8R
3uQ/GvW9fsFTkeuvXxnXMGx/TMzCvQ5i+5oRI2p16lis4zI2KoJyXnLWR5Dd1CW9oeY2PqTnvB+o
gHWczDvI4gIaS+2CGrScQ56ywHosRM4T5L+fg35vzlWDJaOVaVb1NepOOrplOBDj+2bIIa0SIAcA
WwmtWCwRMrq8qx8jnNV03ysu4UQg1yWRY2dmkVFErOYFm3R1dltD77RBU8DtPjJzGIBuBjizcvma
39Au6v5iB9YmKn/+i6SbmeM0zTlbu6E81x8ZEcvt/bXqii6j1ptFOGnb9U7eW13uiTOsCFDFR/IE
VPbmSpQ9vitZ/s7DNfw5biOa0aAlOJkX8ck7sVsdqBsPp0WU8G8ndB5+eFmUAx/4mrZoqAswitJj
lMyCA6rddoNB794wEGPb1xZ2O0XmEtse4lY2md3GFViYrkwjSOHe6edAkwlYAKrK5LsE4uhpusqm
iV99ZAUilMqryy8GnL7B11AnBmop1yPiYhuWgxtVwriSC7md7M0SEtBcVHwGVpoyxQrB5rHGQ30D
ysHK0R3JhF00lvchg+wGKwjUxA9IXNfHZ4KsFDCv95tfC2B/Pvc3VjFAdVTolbx6aDXEGonHdlxu
v+yRSuL6VJQbQpEVo6M0zQPSpZXpHUj0R9OOf6saBEB4YNHGslZOCFsPCKiv6ZmeDHVkJ5WbBnE8
VpKqBGBhwq+F4Mvjtuj02sbrWz4OXPRRnX8TExztcNTniPyqzgEm9t5skC+oGOHYDRQSF+3iFYHW
owZ1kBYyV4eGvwpDkugDulMG5odPvlFHrjpCYTETN9kQ8kWgF+xkxfU8U5CtAHR87eCbBuLnJDXM
0vqE3bY1s7sGqJlWu7vdTtv3xnuM4WjWd2NekTJCdfD049PK8vBONlA+TheoPtNw3H29YllLzQJu
neq9QoEWSzB58w+OZiKTzmXCB6JSPhOExjVdRmXwIyIU1LFWj0lie/ZNPuvAMgjiYfyBpQxIF2or
zPe9vc+rRQxGO+cy1BaDZkZigBvEfL/aS7ojGpFVRKNnB5qL59YfHM3Pzy0ViG+IXtH4a+4kdmz/
tbSUAEL4VOp2hd5jkHyb58xc6xHIMJexfeeyA0/BytvOyh9P4f+uFytFThndwM9ZSYCBWVi4fiTM
7Pqyl/bNXjNY8xmDJFohNPraqf1PSKQFKZRoNCVk67AmpWhCxk3Auy+zRJ51rXACJfrG6MyhTP00
KWzs2/sGfJ6MhAfdEtHMOhtWYw54E9EiSDD5lKiMGXy2jOg8NUJXqZcjJ7t4JTJBKQmbhhtOaN/M
y7znyZdg0d5hr42ZMN1XzRqKz/AphuqgpJSngG5AM4W0e1LG+8p3xRyeobbm1oXj/Z53kEpMsEH2
rrY41eilH63L3+3Mwke3LN9Md9H4vd7BGha0sP5Uiztgca9pLxtZ4by33eFmCuaIq4XynisNRCfl
Y6r3aT86b4UwMvGZH3wg3Ha8+gKP3rpQlR8452+95LC/O/z2aP+d0xnFOqxJZ0WvmjQcCjHYO92a
UPncstn72/Q1vg6ccfQxICrbZx3Fv759mFKEE00ZWa3ND9JZHcoP6HjXAeI7LGFN2e/h2jjBsCZr
vl5EId6sBrvLn9XDKYdIcZRYOS1ebKR5sLGv0bdVwo+SiikAsxqLuXnCnWUTfO0GJiWmBn/mLXS/
l6yuYpwIRpfky0rASfno0rX2nV+yhaOX/nw6pDUoR2XE/k8f2dRjpGUvIR9XXA9ZRRkF1t2AWNy7
4NTJKqDZFhlChFHkuO9hGItr5uFCq4wK+Bh1NMucbvDxm/l71w4D9Nq87KrU4QEMSJSeqvaoyFF+
1EcxAfv2BQulc9byhAQ6jISK17cPze88/MOEAtKhU1ZT6hy0drjhfqWBz1Xzd1Ac5ASVLgbVYp0I
RM1BNMe6aJKIleS9Rpqn/KX5Zh0j4Rd8u2tFOoF7crBM78dr4/vNoEvuEGpno7cvldrB1zzuP3f5
iNhHb7eCvmFixdMQQ7mhfVDlM+k6iyuclbx60cIHQc4D1evdUHklDAZBaYe0WXIje4gO7E0RMwRG
3uIimdeO5OXT9k8k01XynBiFf3jzWbGYgCnQFI1l/iIC7vNDrwmnlw6xjEQH2zwLB3GV+Fgs3o9N
j6UmySIgz/kLaX5yA6FPfDz/r8HLd5Xs9Ek9pMraN592wPTmULENhvfqaY0909PwSWKdttlPXTup
CquRpsabo9ibszCzYr8f+pKtS32cqmGhI2txmOIM75FT6ltFQa0jC1AIfFpLdJgv3GIOEOekjzu9
l4+o9vKkLm336TAmVQ29hSicToRtyAy2uwK+sxGL6KPa90wQM3WZ81NjvLi825bIDyrGt0VtKV1W
gp5i3AnAeIk+VLoilq+xGVtMiMWr4ZXES5jYbzlx82pb+0GWUK9F7j7uEXhtJjt1RWDwKXE7zCB9
wGaUADTcnPazp/E2tEtzYIYk7zwyZw1F7PZe6WW9FDtlrBDVol0LQUMF5DEjiq8CpYUtKWT0xw6d
BMr+Q7JFGOgVSa+4uwaBD8Eb83ZJUeAPyJ/CSh/BGKyajF9DeuvWAI4hSAFmkU2viunldMky5Bvt
s6gBMNRzTxvxlxKeZgFbTVSRoE9+ynYFhCvZVOBLzUrZbAiqXHFq6A5XUYUv/yg2rYhiRN0ObqAH
RSLxiknIzkAB+OQ8/1dBLEtdb9bxd69TEipJo0UNsp8LQHbdU/k1T8S+3B/tlwejM0htCSWhIQBh
3NdKwT0GcjAE9C5rouq3vdknEkKfE7LYADmkUjJj0yKWh089Xg1T/vdRO8hk9eFC7T7yrEKX34pp
MAU5xc1UQJbyFb7WV0X+5FsV4Q/Fgjlh7AlKwTiM+ngTdsiu/tvHUG6geMe1tQqfMaz2+5xeCLfl
RjhW+zE0N+iTQPWoVIy8qoyJlmoULrI5DVu9bYVQSRsaCQZ9U08uspoIyyoMqdlFSnmGsYLZo+Qy
qV1c9BMQMbSSyrluwTx1Cj2fIB7xYRB7FBt3jYb/diO2PLkLtReBhMYBzDsFdkV+4BJuOAHsTxRH
dSI139VB6vTX38ZGjbKpGy9g68WCQtbCMOf5A5TXG+Mjqqkf8hzExidL55LN0L/fcjZdZzlPIXYr
bprW4DLmY6YrbUMvQqHhmoLZgtch1gPYmwg1DBIl7IONcT8umcnFCRUE44Q/Wp8u0ia+hUmDjfgl
WEvdlJyEwCNYs3eTpjOK0fEdgrG6JVlr7SYMTyxfRM6Z2WCo5z3cq3h7f+RTRpm6lXHfVHOPJalv
/H9jZf/wY8OfI98ENW6Vp8U3sg5qIYszCHZ7Y9P2+JBwfypZEh1ylfnlePCsICaG7+YgMlvfeBb3
h4nuFnqmGA8w5kUaATF0eOuUpKcrf3g5sF0tY9uFxBb62cMMeds8Myb9V2QgjEpIMmiOmQu7gj3d
i4f8R8N5RvbiX2lDE68ceuxbs9/9n4dJ6hLF+nii4XQuS/coJFmUEI7FjZRVeo09Ngl1WAk6L/i+
1jzQxnL6COLZ+1/sC/PfU6CBy9wrYTEic96LtD2Cc9SVgqnkUBqLFgTTqoF1fqY357et2NI4DFJA
b6z3rf4lRXR9G757WVyy0bmzjbdtKqMgzKFVuFbByQE9C6cXrCUjCQM2rpp/4mSBLqqOQAN2d6/F
/OI+4AQOM+C+2bb518JqXHA4n6CF5dpQeRNrRMwfXqF3TwoPrRqDsQLn0y7sJp1XWAUOX0dUQuyW
rlTiPLwXute+sPzD92SB8NCX21Cl5IoJIAE+hspoiN4vHrv2wGnZVOvsgyyyJpWrrX8V9cwbZjzn
CmOzqZ0QWD/RkYwvn2XBfKb/13qr49z3hCSHh10EzagQk+uLjSVdJ72D3nvFFidPvR7hIrafbrSi
O/llj+Z/DC6AuHeYmYNoHjpJk056CCoYQdQRGDVaifNxRCLtuHCwAtxw26hI6d5VtHQ9ju/VJjmQ
S6OyuCmH6mNwrOvc+a6+bfxdYw7dxjLe7l3ghcvKxp3PSi5c/ux6n/utC3tPfimTImrbo8/xmOkP
UZnfvQLYwnN/RuLIisjIv3FMYRIp8rFv2vzodaXd4I3E6Q6MoIlhfX+IC9YPwPATWkRuvPsqcQvR
XXJTylW87VXsRIjRR8WiKb74jGD5Lme/fHI7xsJSlnGUZpMMnH4IsVKq6162NzGu+r5n4JiBEMQF
BNkhNmasmhIVT5sWxIBWJCyPovdE5CZTLH2MJMbCrL8WSRXMbMsI7OtRu52Hm0s+n8JxK9PdebwT
2yuo0zUPnIp3n7vJUYGOUxJc9Xf0jR7uf8S7zutBA0xzFfsUxJV3Rt8PqjjmQN3Woy6dXnXSSFfM
+uBCVHGninhYjl4lV+4ZKGPxgbMieLdAFtzfjjtvwlS7ZlL9r5XGkmaSCcwsSkrYtqEe6IbHj+tZ
T9YltUc/A6GpYJolxtbJwNi+OnOkmaqS9lGoh6W3Sgn2UwPca+oxhNjEf+BGvOiw8TeFHxAX7Je0
xXemWFCGSqZw8OgP3m4VvL5KTS5tHDsDN/H2AX2i4XBI8MF6A8MC92yhwiqgsScUrkNG3DQKsu91
6BcsLF8vuTnO10lgd4IsT9MjDLRaT4hPK2pozuhF6RWMerE5esPJvaOR3NAJFjsIAKnUIEEQKgjt
J+hqB6bex+fol6yV5zEf1zEZyJfsXk7E2yCsb3x1sLBC8eJsNNaxAA+rhAti+ixDCRiQN8vEk34T
r+ztG51427234ONZY9zrMXIPgXlGaWh+YDW5k41hi5EQmrgwAmYimJ+vsOchcp3EtKcxiU9woPVr
CRBuNFe12RMfHRWD3weUXH0qNP2iOkveWV2dk+HGUB4vkMSlW3WhK59jjPVxJJj69leDtuNuCvuq
M7IhvVFm24ONOuFlRyuZgd2JP7sfU3MGAvxyrTKIZ72dgPPRv9mv4Y64BOV7oTzAlUiXH2Xnf7q/
CNyKiuvXmJmz0BBWaTmXdvTWJagsegCVZDG6kuDGs+xqi4njPk3Gt83mSB6gnzh/YQMJrjSIRBkY
2QCaZf/p/dZTVHW4m/fzvNJR2DRpm3142o3ySz6ToJfv/RFJDk2zJXmtQVGdsiCIA60ndEplL31g
+Kwr3pHbSp4HaKCa/H5a/tVrcfNk0FyGzD1suwbTBtJt2WBXCc6YHD2eK5MWhTGb4vOsohQ3PeO/
Ptn/DQpalJZkTpGKiqaELyZSNf5gwrPMwW4X5SeQUtfkOIjecx+6chwD669GVzyngUkljjhNdnE5
2t58pb9rY4QosgTxhhHAkDPWkzuNT5LFEyCOl4nywA9xaZJ9kTQnDl9XVZ6EOkFxHt6xF2oCPnUc
d0kwEO0emp3wzi8/Tjvgp83DwYuSfbVRGyE4RH7ztKK087E3gn+B1RQ83xS1x2cLWY1ofYIQt6Kq
iR9ay1Y5SeQu7t8cjxc/M77eGlfOMFtlIN1L4En8uv4jGAKDpZp6Vg59msU4nKyOVbKP6L761cfM
T8nmRQpWE7frz5uSvMtnq9Mwi0BGp267e5TZ39/0e70qEbLD4oIwQc7rZCnONuDngW3bog65wze+
pCq7olh3Wfyg6Nu3BhBmMypbQP7axO9wgonQlxDVfC14pa7Gbbyps12VhNntNX/j4eaGvC2JqaIE
B9wP1MfUKom5WMIAnzsoui81I4+TADKlKJFF6hejQwpJ9Do+CkPMWbH0Rg3V0z9X5XZMWHtOEa2F
sapdYQJdaTEOtCOYv+1/a3NnnC9qSCYU//59udSGB0oAKhO52bv+eJrJrNtWmyE0wIaZQbyIkXH3
8Z+p/oODGALcFBHhMlbHYhxHU6xMtQziPlSYU/Dng1XTJKX1GqiH6YijRMAiC3XQ+MFZPR2eiX8Q
/dvAarMVaP4CR3nbvLW/BpaJO3GMW2h/BNSMorbnRa6mKwmGM7xu3LBIGjy9KVhN1gwUPAdbkcUk
a9m55OeAb4nuAMLe3TStbVh04dgrrsZ7Lnz42qfx8iyE+XkoupAVrbGyaluis6lZ+1K8TGde8SOL
12soGVmHbepj3gVH/QN3f2BQsFw6oKS/RGxD+Q9ZWcyiEiEM7T9VnG8FgnuKB0WIujogQwvYRtH2
+KQiglZAr7MISY2PBf7luHlYrM9KZEslOmhC0eYB9TP2ekWpqQjviA0yyCg7JXt6S2LDhEQKC/m1
KljDFKPq5wf5A204vTOVFMpaErQN8xq3M0L1+xdBZzfek/KWNgYy2uhOL9Uz4kBw9sEjdf/58MG1
3f1zgEJJ8TYNZP5ct33n0hU3DOimAFgHIIs8sURhlox7jtvhnfQckeTtpHZ/rC+rKMo+UU0rtkRO
VTsQSJCaAL8MJZpro7elsn1dB1yv6pb9/fk6ejR+0sjdAhju2vuFoJt4PA+yjECHOiBNkWJURolx
8g7exo8KnHpL8w5qk8JhVE9Lz5boEPpFmktf5n9yiO89W2aCB8188R0vii8flAj0abdOoiHpT0C4
MC9h5jnzbMWjAsXg5+FVn4lzyWR85QN85P2tSB+ICYTrsjkC5iIsQilDh4fmtiKlsV/LaRcsA5lu
GZc/UzTFjE8AgASeQSQogy65sCvsjBRob+jC7o40jGRiFaJndzxIdhepT2+4DtSquhPVVD3FE7mI
sqytp3gPLN35GDlopj++tEWJPrOfb+YqreXH4Es0p40N6u8BzdjDAwi3qBQCiGAx+rioTD3Rml2X
0b12Py3E01Ug6ycpRB3vN8vUEzQx6pgKnpTyNQLQRJcNu1XjY5lm7ByjzE6hLVw8up17Ls9HxhTR
VkPdIE5hubU2p+F89Lg3OTFjK6NrrxlnGifWpQ7UNtr9PdV/M3nL51kq2gohTXsIRZ4T6/aX0l3d
q6XAWg7nBc4JGBIoOPUd+QY4oyHgqhgiHgB2AYSYeItLm6vBjm1+Fg5sMZmEVHibD6VBbvnm68Oo
MD8zdcrjp8EM93VP7/kXKvJepHTbWYBw0lW5MUgTmMJ/7xS45G/4BH5OLxZXCFFOXG68f3AjxMzi
GY+gi1TcZP+8RXJJP/GVqylK63YBxwglfBKKFbvmH8VzhlGf4mUPZQL8gvIC0snp25Cij/vJdq7S
qUsk9ZESxK6Ck4sUeHvIIz5NWrdeLVvNpXgjcMhykGbxg7ltX+yvO2hhi3ea8PnyaPyxX3MR6/vK
nJN1gBFXKENW+O6JzdAVfJktxLguz/sj23uiZ8reaUVffjaSc8zjcCwoFeYZbRrjnp9MiE3ti7GY
dTScAwBS0KtsZ/zApSJOvKGhnDEr8PNN6F5F3S7Mp0iAF7sXQ+xyD+3ipnWg/G9zCoj3HhBQB7c9
LIHjfF5CkZV9IzmebeC4XQFm80bWMx7E4dF5iiCqObp4+RIfaJTE9RxqrWJGwetZ9qttOQSwS4od
m9NcRdsYtHQ/0Gueh1vcTNkznMkCn5eOKCBp+WI6eqBvwFtiLcSvi6jHAYG8yqQKtpigAJ9INiS8
G9MtwhJKZE4nEhRV8fef0xhCaOqyVjPyu2Mc+SBdwzU6d6w/BP1Vh9BlM8dfuiAVN/TPzotocTdC
Xm6PhHWxfE6l8N2dY4i3fK8ZFqXEuEGmjnZ9jVfCXppzRqkRB3JXl84a7/FKI6d8E38tdU4On0ij
Wpzo/kUXY8cDQKfBq894qEfnNh1ibPkZiffDOP9KMet9XiA1dRhXaZROBkds1UbKib5eJIvrLXg1
kEdvc6GNmYYqOuX6qOVHJSVw7W2rzRtJFBjj8eghuqvo485TAfUTCtjwu1nm5WA7zMfsjOgEipoT
zyGOLg0kdGVtL+tgNNU2az1jA444AuzvtrfnDca7rBoaYqTkPkfjb4Nnc7sA0YyXRPu9gmIkzSFP
jv5T7cixAXnyBnavX0ZVaykDB1KCjL8tZrdPXDBLP8TptxjsMFQlQ6cg7jS+W7Y/z3hasSvjWAUE
5C95UjKgGxs3yelgZhxnK5SFGTTwIXmseeYQfeOTbUt6fhhywrAk6YXTZ9w6mEqLqdxFGXDCieEl
QQ4q4pfv0PX+qnHEG8r1dfV9Q7y22hKK9jb7tpseQdrITdunFjTzwgJ0wsst/yBnce7iDWvYl9/K
THwRmQm6ETxumRJgO4nZZuJA97tAzIHQP659loD3y5iaADO0xDKwTCpq9x+qp6kWhbf0xbg1Znso
NSZ2soEnH4a9G+uXjdiKa0+o2wIdMTWcIL9ON6ZJkHum3Mp0ZiYrYkCzHwbBo4/QFkBVsZYK8v1g
+R3s0h+QsdV3eq+fU0H/GjDnQRa/aVBQvMD68VEKZdUXFgzoh1PIiHlb7XHsJgt4FiYZ1iAZKvGk
tZOT7cq8XnDp2ECx8Mx8fJs+Zkz+kDHg+uhoYTwoDQ9pduB7gvw3ktolZZMKI1S6q4NEbgJaoR14
hntYW8ZlfAGFXuNtzohcRTut5xCkWnxph7zlIMkhK1oQM1OgFKZyPsMHUnxTQespbNQ0u4sVcX1x
M+MIGZcNeiHALuUSkfUnWNUTlRx7fPVkK0Dw1nTN3FrGBulWFEjtC2dL4XaNYc+Pq6FuTT+9bmJh
ksdefiItzy/k3z8YgVq53FlNpH+5YzpOCS8g2R5I4G4QR7jsq1sK35x3y6CXdDEDB/A8E/1TJuFo
iKnxKOtqw/ZebzxhhKhhC4+PhBaxKUECstHpAyDzJN6uBg+52kNGZK/esgW8V5WVqPlBIDILkBCQ
CZQgPWBqu6aT1saGgWCZe3mm6XuyUR2UtuBiZ1bNsbTVX4vz1JL1fCjUAlcr87nQrG7wZo/itfZy
OYTCUoB4nOotBFM/qeKi4Xm/Z9QWCCu/yr9cGha4ftshfBrP0d+FytK51HC6VEakdIPEoyvI9vFV
fwSrWy4PZjYd4dh76rK8exHIOfIcACx9NXAJZ8/giCMEYFJ0CEb4eUvuEf7j6wMU6h+6rAXAl2Sz
j0mXMc7xl0yyuzfwYSD6dnvWRuE+bP82BcvoBga3jXmN9YgOpfboIw3r/DbhLcv68IXYIgNHe2mT
HftDHVU2d7mCE7ukA1MjkkkZhMVC/MZPjG9VzdBLgOHkcQx1sLRQlnUyVsCiSgoFHpB/9FHFkH39
J09eBDOcjS02+iBcnmnd/UBN84hRheRsbSosnK2AodkdBC96oFluY/fqQgLaMvkGUpPSnXVo4yhB
wwTC08/bSltDJod/skHwDWH1OIeIvnszQlFCnxDVnLA3nDmwOb2fyyvakfZbUCpNQqj99VlVAIsz
wUW2+o/CmXQLIk4DV2ImuyRZAkuuD0fWoiFuHvXZ/7HAo63GlszMadda7NxGHV39eYHR5fP7N46w
E4ReJ5xBz1lQRqeoutPoIlPORQte1QY4rx7vk/ihh/6J+DAjOoob2A24ThppffaGqXkcIfzw90T6
egZ9vXIZpbsXGZtH3WrUq5tQZCw8JwTrENu9GZC76Znrnnw6tpPwBwfecdhrkwDUNFnR+9WtJygb
FjOwMjll+1TAljN918wUiXLkSB1lWZ/rpvQ1ZFPw/4jiGMTS7PiZUFZPmChEiYCtvFhxOSyqOC6M
wHIYaAmgbyftnaPfsm5RoKLuSf+y4RmzT4TBpHl9ECnrgkU58NFKBonuRfyD6I8nMvQ2nb8Y9JbD
UJRtwXW/+iHIVJtKBt/3UWOPVpil1SRIVdUdXAjJhl+Miyc8N8cQqvcQOJ1r6CZtLV6eQtT57EBI
22tKuUbYTdajtaINmcDwdY3G2D5HxYhTY3wq8A+74ewtF+LGckSEj5r9HFlgTSx2PF73/AuXjXxY
c2seizFacWe7TBQLW/GKm0yc4M9kbd/hgL3zvTrb6PwpsXBN+KXnEHi1N8BFbFsKhOMC9rR7LOAj
zkZI+UmucQikYDAagapXi6lT6Wg9UIFCjI+1EIqupUsUTVN4jPOLfwTTXvQIwXNh11m2zpcNZwtS
J+PY8nV7pFIOwsQHj2aSvJIEPbsHlTWDCgJsBMH760oP6ZdJz1z710AUuteKHWnVeVtSud7Vpj0G
a6VzZqqE253GTHiubZsvovs69QJ6r06dAUgP3G+EaaypnzYI0Ro68XReKN8XTwtYFGNmMXpWXx21
rCVF8nEcIjDBPet0I/49H2er3v8nFnLlOk9+oL9ywiQV1r8WI9/nEFC+TYSUBQYB/D9u/licXxbP
FQmFaeamZRwc53BlsJOKSLRNxC5KrpgRhEkTgeTt4sm97wGZeQMHjYS3vzDEpy7JwRHOYGvGQiAs
s1tHWO5EB5YcHNg1MqBroTXybLz6XF4jst8AJTUIJQJI4EAWEbJhdRMNAYUyXgD/2+GsK46iOUWN
wr6W07Zq/Z688xESSTMvMciKhj5/8iJ1tQWKxZpWz7AFHwkY5h2QNsjMMP+4fKNGwdVE38ipyaHs
DXPBlS+y5P40snJb4fA3YnoWmDDbRQggi/5+/7qHARK2zJ3mwimrnXvTvultJ01YNDEDMCsDjWcX
zTin/yb9eRwGrHR6yKpqEG0XDEEhEYFfQRXr4DUVOpmRmFkQxLjgot1zOGGGdsxgMkeaKyACOH1C
cBgA4J4B4sujyA1mKJQlBUrozqPSvbTYX2lw5zBkv0fiICAFe0z4yiLibyBzeVXRLP9cMWF5G6Hp
ChgDesJJM4WDG6PTMXjxPcklALqOHaJT8ZLYiIpzf1C95sZDmcZdJV6mQgS7rIfWvAv996Vn3cFA
eGPmVursx/AeQbt6hCyRL1aZREe7co+wny0R9QeYW0s90D6i7u9PDaqW+EGwMOBwEqmJ+D1E65hO
YYApCvz8s47qKhYQfM8k46qZ2AYKHQjfMGRFtbUzZNw7w495CPgVwgoANKH8K94xTY8gMVtWs9Id
Z+frW4DEH2RzyywlJ02Vy/GtewcYa1oek9fY1cP/rVf6MAwmvM7XQlQNZ2EBTguyW+w1PRzVFxfE
PNS3dVUctpRn1HPkQpz2OCHxfCnbCCKcnHOpU0KBwQMKRmsALZ/Jd/qa/U/jsuGB+kEYRZKG3o+c
EfHaCoriQ9fmeEOtM4mmzmWgBNZzoaac0xWciBpURIAqS5pMg2E4/nKoqPMqBRTdba2srd40036v
RBR6CZ5IVrjm/ffnDx88IGtsFIvifhL+4oUol1q2wZUuzmAI4MgOxHaOLvfRg1tnDxkci8IeoLsW
kHpV5ib6LvOllwTCasDTMP/n8hwfQ8nL0h5tSJOR8WoY/kixChzO2lbgNethb9AqbPdLqv06Kyus
GzRcofDshE4gExAO6ayeRcMqy/QQp0wE1Q50YDXMjw9y/8H8Jh5BMz39y/qb4VTJzXmYXRl54tle
fIfmkrbHZ5BaDheDMckcEcP0luq5qoHiWy6KlTqcyQNUYgLSildcfzzSqHxDy1BNMjCKZo3t2XIh
Tf6tu1pxXkL3IJfXBpD1rRbVzUSBqvTrXNx5bl0cxW2Y+5bY2ZZd9+5dQmvwv1BNCZtr/CcgUqdk
HtziAQTXVuFKt/KIeXVvRQOE9rk+mMZwZ03J+zwzIoPMBkrP+0gHh/ftvYrdTcZfBtveFp2tDXlR
gMb/m/OGifEOldN3OfycKM38q0c3SFO+g7/St6pF90eLct9lWbkkFanyil3SzkspGpbeDYVUrZsp
55eROeKFnyvojmoRH6FGi+z7ye/egnnP+4pkcBSxQyt9At6LGxSEbwfm1rL1h7YozTI2/06NPhPW
1YqqpAjMpwAtH5Ker9pR12gKV9B4Pr1I84bsxtW+zsulz1Pqml7z8OgkrQv8yshiUfolMrLwV4gf
OFR+R7BJNRdsq+LUf8sItl81oEuKZ4etwravAmoArHu236UBjQ7jwO9YoB1RmHepNEU7hBTu2wIi
3YGJlSgB+LpxeFA3ctBZH1rFIwiyemjygO9NtUqDWsmAAY6txNISxiCQsA4pl1NBAFAFArnvBYEa
dHR/gpmnsUEXkqfMIwtRuFhU9BAISAxr3j/C0NZ2IpNsg+6uCmvIkeFbAwYxVNtrwDrgKt18CMYk
kWps8OJGmojHkfUPbqmiyKRmpsYpwITrldGhb32mDQTM/JuC3fcXqkS96CaxPfJpv5UBRokiHf6L
6Q1KCqKRDixoSQb8q0UMIXce3RMl1yOHhF2lc8ukfslPrO4vhE2uyv86Xh+qyWc3cUlU3ztwFEZ7
YzTw6ZMWE4Jm1WGVsmdrmSoPE/tMap8BivojuvI3ird6RUZbYL4zU7FhyeNkrWxdOzXukKnHb+b5
OJCBjOl2rrg+TWnQ6ugjMLr6+AaL9kE+QV5DuokVdlAweoEs1rjJdK3Rb4z/1Sw6ZcDWzZn3BSgV
5wmQ1/8B1C8TL6kdLIeYZVU+nxQzzk9JtU5Xf3fG9uXXpOkbWLklqDMEnwpVP/nIiyDQXj4RT6L5
SL+K4h229cVD6C0+wiBeFyHPSCQAQPHEwt21uiwIalwPfX0Kx8z0nZzaRM4jx54pukPL7W2ENGRl
zkoAVwdaYZd5GYzHPLv+49+Dbb7NCMWC9YXVB2TgqziiBpdNRehPVX3j1GduzMoDX/kpwkf7t23b
G08eUWUXLLuOuymUTj3P8dfOQlXTWbGTX2Gr0ts4uAz7661ep+d6j+Svzv7eIh6QDnVa7zkkvN3Y
SfpwaopyUojUKjygZ5W/+Xluazt5Qw6SQn6KzW/YVi79rSOpjlXUbOoG0/sav/ZP1QmzvjzGLsXl
hnjLqxkG/OYzb3Gt6LhF/OTwlCLge7Ven7pu4HkLeZEh53OtDRR/LaigDmJo2sfJvCTmUjE65/ZR
cqgr8LjvxtvciWojNXH55hKJtX5RBQfj+VfejF1MtVJtM4WB4zT75S6CnL7Cv5pE1FVYu3n/0VaR
sm+ttg7FDnH9jkWv5ecpF1guSpXu8uPivWzVaiWSF+WW+Owp2IYNQ1WMvMBtTKjzoKbnqYqYmb51
0v5PeuQFwKmk3n2bP6GCDiY9ajM8GPHRV/Iq10WIfwIDfRzOZc8Qd195AGTAimxqCIzm5d3WfPIA
JmNEAtE00tpHDRhOEvRGEpP+C6D6r26jNrMxm//CLDCSP5VbktaG9PcTAcIAKOMnX/TlKtInB68Z
/pBdKM/fZVQnRqtbWtWJSUHrxccxkFpDaF9SMm5S4fbmqzIl4R7DL0fLXFhuteAt9OVBlSve/NUD
ZECqCOnkYJ0Gf63CgaZly3ocut5ROw5ItTpUz6GqkFuFDmEv8lOmpJvMTfRqgI8GHIKELzUW9MqT
ryWZBi8K3NOKakqtEyHSO/ZkUGcP1216aBasEqLCFfAIqmtVUp2gZ0LAArKC93NygmxjVn8t9CIz
s1eyj+ERPmKOrWerq9FV29q2Mh5PBUVIEvhpMMmmAAe1YN2SZYcTwodxtBNSnolm7eV5wSql0BIh
/ebZGxm1Bev0vg9CwTA03jjW3h2Bpz1eTjB1gr8tQtkRB1opiL6K4JjNRi89XsMkvFjL6R3r9pDl
6ZbCy/qdSrb4E8YsJx7ILBI5y0R26KLl7BmwXkhS+lO3DrJPD7l/sQOhHSd+VndEiBHdnC2kTRq2
lWq4mjjDhcCM4sNTeJPhmlnYz4kvOtpH1bMpz5ii1Q1R0E3e6kilNZbCqyO9F5YZM2LWYyebESQT
O6aWs40tg0lCNdq6cvs89MME9WeRauiihpPDqgBvOnwbDgTec7CkPZtzWdCv1d/+SemCibIQ6agh
PNgL/TUp9m8rXLtV+ny3i06ZcrkgDabLwvHTr34u9g7jMyqvHiG7OXqR8+2PkUSrSLR9tkenfGEV
DxWWAtmqKqHqDVxyjUTSiGReeoQ33oB2WqUCNfQR4wgSsg19JVQB6/HPQEtktAdtHDVdhdJHIC2R
/SJtqHQkyHbYUm7sszCA6Ym+oZ8Kdn7pqqm/vGWaSdxiG/vUrRrVufODsUaa/I+Kq/+T1tWwLXTE
pPwP/BKI2jGfAmbr1wE2JJ4L0ZuMDXclypXrh9y/cGVZjBEBJsC8ppmMe6L2c+46Oqdjg8Su03Qh
1lElQWpyXTgq/+DHBwzi/uniG1GYq7X5C2wfAksMKD4eLdDIIFuONG/VpDyI1STCy80qkLsdN3r7
AgGbRFLkhq3B1xGaRNqy7fuQqEukWXYCSH8eUdXVPxbH3JU+3JHFIfGZmGMOEpg+fWjeXLxl+1Mx
zqgD6wbpVpfBw/pQGk1UWYL0CHqrc/niKsGdnadORHbj2uHIo9xGXP+9q8XZXDtlmPX9Nk4aQv87
fos8O1f4gmCf2pr5UFZxnV7h/ohO2pYXk+4okh9BfJ6qqzRRtChhEnCPzztmtFFQ37sCqOxs2Whd
AAoXycWK68v+ERTtDfNgh8iwQpoLZlCfXExspb0QBFg7ki+Gs132wZYF0OPE8Iq7YfnxC1rWbt1z
c/+kWvyhlY9m4eSWtlKJzusNP/utWEZX1+vsMEE50kWuWRVCqWrj1ivcognVUCvWWdTWsTTFRoPH
H7B0tEwiqe6GoOBOVePbPMhTfLaCTpBq+s+nU0f7gwIxTuHkSW19QGmJHjmiEHyhOAjqTo9LP8C1
tNi5T9olQ7p0E+pXssDVpvfWTvoGxnlBl+J+gnTXiZ0OdNB2PSfPLaA6JQho2M6IgbTzxFtQ6cS4
hZZXIa3r3b3wVF/14B/xy41c5pIHVpficduZsFeLPdMHogglU7Upjf3RtUqoYr3G75LkKrNKAFPr
tqW2dJcLCPKcg5XQNkdJEFLJZtnBS2DxlK9muPg8GvxzL9KbXfR/J26oKt6vkzP3IdGHK858+FvQ
HEpt1SJ6eXZqvH71ox+jlSmaN5GOhyqq+zM2aRa0ii4SDGMTdbOy0iTp/BnUgrxuuuntTsX9hz+a
so2tn30aSa8OPUiv8h7XvXFIe0K4VSHy5iuI1sX6Q+zn70OdRgBucu0Ft5qEMGlr2VL15MctJF1U
0iYwT5j32+daz1+fzT2pBXP9BEP5oVXTlqHcu20/ZD2qOUc+rGXrjFLKS26eHSSdM9Mr3nB1Xp/M
V3l1eVJoBuSewUU1y+A1VnR9I0t/foZeEPoY19FmqnAESnj0RKiyK+mAlW0/O555mZFiFVW17HCM
LSWVCcWl/XLxi6UdlSpTcJLgcvyre7wWnjuq6S1BYlMziMIuz6652468bDWGXbt4x6p1Ls42QM+b
cE2CmpU523FfmDV8NY0V4434CoTsUkcAx3qRzm16sVN3NY69zr75gYtCfuW6EfrqifHYo+yxqpkT
zSkkR7Rxc8FcgJeTAwSQl5I6+G7ta9qxyJo7Q34YXZfZPe8o8/loyvxsaEs8hfkDoYtoLMDSa9Aj
R+QX32QozuePwafaJu7mO3fnodmMuqXhyM16lybEkMIzEQKyQwKAqb0zPXD5shVxuykPcGXi6Xk+
HPJDSsxvJ1PcHc6LpNUCaGHsJp375BK46Z32JWZAPl5wQ3dyD2P0TUI/kb0qrLoWlzJyIhbhimff
bmndoaiZWMp7v6Nk75z/0oyaKjOPSQwfZ2E0TlUQJ7hYc0oGbKilmFSKf/EYdldHjFchx+t7JbWl
omNFesq2LJ3vbajhSprDqrt1ChAE/oUrbyJsbyjkQ2g3cDADzTDa0GKAnSKEO4z2c+CUy+xUIb7v
qDwaVvTQX1V3jHrO6IK2Vq7abNDa0vzpok0HS4dB0g1I4xjpLSvWjhlTzQv5VYOJMaSxi18iMYwg
EbidOZE/FVyiA/+X5OgIoNcWmd5c6hcZ3zGKHDW0ml2DGBnvGWBmjJsL6qWPFN6HDiGajDW96ntQ
RhtFttLRFPFMhv/Z+qNp9kzetzf5+4mk9/tzwh1OsQvsKj3OGufJDVfzNiWEdPAto7BV2zcXcRV2
ur5pEh2+9u6R2xZNxvS10uvt3wRCi+8+qZmv+ggZ4o5d1Ddk4+5OV99nKa0qFH7jxjz9u5VkWXXq
zGcdCV3cBsuXBb/4QuSljGZIyPSoO8vrifH2SJTDTwHAVRXvxzhngSdDOwpoLWcl+pGqeMUcxr9B
eNd3D7SSbDtIr38t7aOzwYyBUGs2dGfBqoxDRul9R+MF62gNuJgytOipG7vjRK6QK3J+lwXoMcFU
4zTFZngF/fmrQlbs01XDtDfqfIBdaeMgmmx2jUhaN5TJdIUGBKzPxM8iRklhgmGy8QDWMPoCppNh
C9buQvTDSUUxyphkCj01ULeKnTRz/x7Yh720+W2YMYAVdQx2ADfQNCzaGEEeLfTzZkU7jpsr5qjR
OS2LskRDxB0Op9z2c0rZaVdnNwQ4V+Ee9C1x7GH2ZF/ByFStIy5+2Xmxfz8WjIQorgDQcl9bR6OD
MusInjvYjAqU4ne6JtJSft2JJyaNzLEFNbqtS5pwdUV/v/eaX3dyOL9qmK4Lm+ZYwxVmoj2Q7gbk
c1t39JX8c0YHn63H9/no/lIolFg/B06N53vVFtDKWI0iL6BNeDXo7fgg6zUXenGZl6DvY2KsoNir
CMkB4k3HM3wzNf/zPFsWqugxjlBpkGQINp0RxjP2Nl1MsdPAaFt+6Ddu1bz6bTppj4IKT1ru3P3N
BRvCktTzrtxijJMgzukWxXK62aROxb2eoAr2tZdW7BkdoAYkgfSDnG0clMwCWjy79Za9C+HBnzPd
YyqTcctvP/tQ2Tb6Uao3ddzdl7sdqVrOzP+LWlGHtciOv2f3xEKQ/HnD2UIsL6kUU8ClhST/YtnP
947vRBHn3n8PyhT9G1dtiMK9O9CvkJx6yvVsCWvfDdj8liBpSSc2XLPXKvirhjVFPEk2SpRKT/8v
GncHFHu7RtPDG3qV2z0AAbF02uIC7uiGV+oSV9Em2n1oevzRXJckrEXG7qYB+NzhJTHLsqXsGwjZ
5Df2VQLTiFrhyZ86ofbKZoDnbw/A5yJkM7qQEtkLspyDDSlf1QUv06fYS/N8hu/v4fadtPjdQMfE
xTw38tB5E+mPgabXFePSVb2VaZPgVMVFZdgaZQyzpIBYDeMoqeVM1D6IU9UQrrDMMQwXK7ufs+NR
NtyLjUni/R33c1x64Va5ngF+TNVOxj7/qDp1vqytg66bwYpZJlmQrE8FRP7df9hk4SEGFsxZ3yBn
66+zDpV71YKXiBgUu/aOU9osTtEFD62jdIQp/1x4qmdJRyp7CIeck24VNZTjdzz/R1XMkmjFi743
vqt4UZG/lFKKwT4InD5W0lyXn4fvZRm0ZPICxHJdrDOBCVaXuAgpOC3nAJPhs9VovaP0b/vLiQa2
mjzHcCKaaTiSgDLn7H1RdxTguV2zKWH6cdSUUpPtBO+HBjbaXQI/nRxQFKDRtLU1p5bRKglpVbSp
tB03K0u0lko+Zolm4H01W2LPDoFyLKY6vfkfNl0EzpFOmTTaALHhIv8pXIQZtVMeDjxTRT3TLP55
KFRPG6b4JUMAbQEXZcHOjoFDQH92TDys/OgPwu8m4dTEvgW/Qj3exCFsccR7oSQxGAlgx5wGSJAz
G/gbVNcYviXyEHKAs0AhobZOPj5tTe/nbR2vmwQ6gtI+p/SB/xPb0pL9bJv9VQ6gLNz6tiiocsPO
gi6w21ursLVzpefUNwANysM+pOMYzqqU8bqGp/iOEXuxaIHJ9uKJVI545BB2NBfedZG23/Ef7oG3
kvOyFFhzf9H1yQGldHGC4uECLKWp+y2tgbzgJycDz8OeNR0UDrDzmNJjc1xtU2bpkDVL+skJk5YO
7OjMMjT1TzLejJZAUx36bKONvsQU1khIqKs0SEYzglZdR9k7SBpRYwRYSvdxqul3R9S0ODna9W7L
JT+KC0lcRS19Ir0hvRJPooxh3oXZz10iXWpA6pI1l0DIFBIjOwswMXiWAkDKpCtKEqT1jgcEf2jq
RDyWm+mdu6uVBLC0u75PiRJYkLgqv9qbt+jFTyAfbqobvcccNv13i6sJmrCub/jakSXi/EqReikU
0MLFXA2D8e6nzquZJbHE4pqMIZEbszaMe60Y66PI8pAtq3Tue38FyIbKOgpUxCq/0Pb7ptjFblht
eHKGG0MkilR5DSeK4TdJbg2IAbwl4xi6sJFF3ygaL2qa5Dn3nJDiIXpOiycMvqopKBb8cVulaRgZ
Mifkdt8SiDNpi3si1eEEN8wRMwtUlEwhnmYrc58cVVmiTjBKqCZHpm9F/Vk9YAoOKwFDY7l3EqxZ
qpaHebwlZwgA4m9xU5RuECDahGtXiUQTjV8lMh1qm3iQ1T8DtmRp/FoPrEfZb47jo1Anr1kiSE5Q
KfeXZrZFa9eMxcVcjuCd49iWZWgQc9tNEuKTDYO3VC/HErFHUIRp9Hoq1Wo8Bec9Fn0vfvDMCL8A
06g8660cW8dgSy2+VYFetS8LaoFVB7Szbh2ThFdfoAqTcBwqUzcC/O2alJAcRyA95DaBXKokaW6b
Zbi9PRivIUr8j9u9PBMWDZsOgXSBU4DR0jIQg9rToHTF77PfqEQi+Z5Qf/MT9SM3bKK1WUw+76A9
M3axhdqAP+HCxMa1mEI3dA2PbiJvNHBlNu7pK+Ifm4XnQFx2QAzL0Mw4Ju20B1M7kRhUjM2AWjls
YNDJrRKL2P+DHPVr3tFvdqW2xm7wXE5MCvzS3tzZ35mCwARXkEr/1w4ea2hbAEFWEic84Q9vhz1G
zNW2W+gbKqg1cv+disb6izA3s3MG9LmugWCzAhYYQbtjL9UfxPlExVX+0qfrjOhucf0DjuE3QDpe
FJRxTJpU4o55eRffAI1+odqp3HEF8bQ6pzwWyraIlGu6tR2X8goQ0p2+i10MurErRc0CJYxfJ6aS
lzmtTX77fjkWotZKbcak4yywFkPCnFb0u5d/hHpHo7vlpIXC8xV61gADy1x0+S7N/Ji36yJ2xJuS
fQ7i5IvjxdHO0IFvYJUy6D+xT+rqK5GHTVa+LWOwIDIw0Crcw+a6F+sCUpHYgzawNZcirAZ/t1l1
0C1VqWaRVRXhAUTYBnOfEnpVmqO05wGbRCPjGHWezZslGVMqyZ4SnaRYoDhA9q0wzXVCwipIbs2I
YVokD95F0A3OlMP8OmxfEAbUCapZswtNLojd8FFr7pbSIrRgn+Ikxwee81osy9yEQ3/SNKmOOeQe
LvEGDa8n7tFuiZoBbkznT+xf7L2dqV1aX/zTiEgZT4gMKIJJ4tuvUgFy3wMX0fbl2errwnoogSun
katoKSV66kUbFyjvzN2sCZACni3iAqqQCzHU1Rsxwh5WXedl8m8pqMNtWYBE8baDYotPq1OGcOZM
+AmwlelpgoHYajCPTV2Kx0WsyGOCvThMSKZ5UZiuHXCgzlNMILRrohdSNtPlW9qz7bQCM2O/zo2w
EzG8CWHA0dUrQ57juAB9M5GOJaMU4RoQqgAIvRRntLKEsBuB8oaQK+JFYG4MYRrk0K/2yJGGgV/j
gr8SXcsw3lbvIFWWBUwjMiPDFzsD/+GdCZUnIKo/YEOlCAcavr7PhIkJjTlIEWur/i4UO1gnpY37
G3Ew8pJmjGaU9ensv1IqnwMYH5x3GxDQvbAOn6ZuLe1OJNNhjaYbt8haGmCLHNpPlodftCtF6e4c
taW70dStTpezqxtVl9UM2QY5picsimHlDmDeAK7cXPh6tijgD3mi+/LavXqFvpb04ezFDhkfLkv9
rOFrU2l6pGikic0e0n04DbaCAGj6Zu018oIXSFKuhBWugKq7+GQCVLa38pTMYReUy53PDDgKJxKK
2A+Fn/3e6upu0dYJKuqffBDI4I1ldnzzjgMSw+ygVQNJwmlc3WuVw0+KFJ4CeWOOFtpy6AZEo5R9
bx1mpvtFbHrsy9MauLKsc1okA49uw8CvZP5IST7BOTHxjYZkwEASDcgSSO+Eb+zzwFtGx0ge2E1b
gp85CK7VbSZSYDEmg6RclNOxCAWn9r6Wc/j0bnuD6vbzYdFnC55DqzXfDTojbyZhnlHJT3TFE9Gl
CM1eatbaOGmkxf2dyBEEXOqtyX8pDQdJrPC/mTswxdhcLU5eHOrXTdV3EXpwGPUe95pjYshiCcH2
iYFUrMh9kv2x6FJqbSsULIWKB9ggV0xFMUCvhE4aeDNo5fwe9WroBnlcLzNg+z0Y9Uszmn0QiSlk
USu6cdHV9NmlDXWynOSOriY+nh9HqiirQh8yPvZJYEmRWu0PxNPq/qOXnX2ttU2SKDIBTNKEOquv
fZKgDj7dXJr8vnn7xPmB13wyE0MAUk4awHqkKIY4IZeoFfaUw9hJ6DuwEoC/de6nZKxDBLnLvuqs
el6oGdnWQMKTuerPcJLXqEcnMBxEVE95U24ve66TdzfzcBwTemt4NEAFilMk5SJddhzkzsbeudiw
toDzBuaKfKGbn8bfbXDjFRTgN1u3LkHlTvkpv9/Y7Y8AnZGTFcNg8saWqr0EcvuTcWJpSxY1ZLe2
ZqoliUlg3+mWOvefDE/dbF5ZPTKPGHN4DyB47wrw4T8/M05mrPCMomcXJSt/WHSW8rBOkJDxcHSL
u2CgIysHcmXJT2Opb/gu/JH3ZDP3N8Y4F9et8GmeC+vK6qkyXMfhjgftIfxLsKQ7rXX7tnWfGhN9
VDFY2aKwXkObQEUU5Hr69vxRWQ0UM8XVtVthamQk5y2RWU9NrJCp0L3zJUp9c56/J3LSviTpxECl
PwJIYTikPcgwtIUMwKoJFjmkLn4qIv1jVNIKNo0+Xa5Ker6Pr77VVB/u1yzHCfbWdgzX09Jqreh3
KDZkjMk0SZL9zfMaH/1tutbVe3mfqCKzfqDRceNqHL56egOjQOXsilV1nQOzenJZmEcLadgmmRTH
hPZw1hOTAi6i30D/86mG0R8ABVpcSmEWGqOkaL+5tmHv0b1UvJVn1p3E5aWSdv4aVE2/v7VSN4lL
6MCgA9GRsd48dBb1RGNR4Vpik1X3VJpPK/Px5HFiN0sQZtPfmHp/ye5dx1UU8w0TtzVltHk0DR+9
zY07xRQCeIaWdyVn2fWzHAkp/okGrKAc1UyMBs8mCEJMVGIaAY0uO2uNub3cXZCavfNVmieckxoX
s6FJA2KZluaMd0Cw9jRppfUDjTWp9O+Cdq5ZEYxuzIPy1z+JCD0N+T8DIPlp3N6K6kh99LnRnuox
PixuhgrsU7al49LrGdLMKs3t6wLffkjGCyvZprBIM/nbAEPqnBmp/I2K423yudbnLews7AIYZpGP
MaRFquSQddZhqEQoN4BVZ3jsMSnuPshTy94FFA+qHYKiHfpgC9BbeLzSvDGfq3tvqOzkjxJkhKfb
tR3ZTVG1AZIhVyO59o7nbc3tpGbNkN5L7qo9aL+lWWcwNG31C+PqSQrxiUIUdRgNVUsop79L+hyD
TtjP6CjxZ+s08em4plEn0zK1CCKirayQXMEEv0r4300ajHWEjBgtpagVDXpXkWfoKQiB4JM3xLsu
BdP2V8OrkzgAJ8wa+ghILaC3XMKO/8DBdefhbLyzeyRyYaXSwLtYneVuFtR9oa3pK9SuwgU6f5PB
Nm9LYxbqqMifeA1gboZiZu71tWHt8XB1mq48Bd8ln4Qvjgww236VlBJudKeZYT9FCUy/l2WVqMgB
+7w6VQtvcosH1OZBeZ+dKfp+CLPQpB0pBDiEdDUEpQNFyUkYj7HqtuGy0GqlbQa+PIdy7wYEV6oz
eNuaKtwhBaZdOrPsHFozz6CWIB8tb1wfpgZC+olQ7H5emVkVl1TpBld+PWjtjzyKp3PR3Tjk99sy
baa7Ty6+XKVSQWa3UO3/3ddbbgTUTMi4hQk+rmG4xE2PZwkTOZh+t8wTh0Eiw51A2SCXBgE/R9BX
96UgV+KCbaw8bn+YXFqVL2Euq8TXM9fsiDaZ5htB58a/R4SSJP1bxjj1EIfCks1HTw47n/amU98L
hPPaUDzrwLnk/go7bo44GML/3MhdC+btg2dy+s1n15XW4dqj2f35P8Utyt6ta/ugsFGxbnZEEu4f
Y16z5T/bjsZ93sS/1InDodAUXymcke9p1KIdCa+skSJz+mfKupsR6I/LSsJ5gwRkSO2fT65fpRsc
4luZ0mM7vFbfmGFfpXJGGzIpMUWS/ZVvVHFL0c7xy2ODarqeFpXCwRV/s2fHOOFlIoWR1CzzY8CT
6iPSnJNooxypeWu2+kgFF+iDJn1KBQRkTFllSMA71FsCdIjdKFtumYNYjVCamCrv8d+nqZrJLuTP
QarJ/eaOJntDVhFO1Wk+BKonzl8FXUCmQvFNRZKnkPvZ+IA2QdsSlC/3Ib1+UaXUNe0yYOoXmyXq
OwzPWNXldGPPoMh5uFQZCsUzlMSewGxEEVFsmQSPV6BMCtp1Gvf4xBW8LmKfLqf2tUiAUz+NKV0X
7r6AHZOKsv9abM5uQc5eB10ZpocckZXNjmIgNi/K7AyzT+AcgRn5BFlSKmJ6P4w2XGCB84hZwINq
EsTS5Hd1WvW22QEQHdH+jrDq0JiLkZDqgC6RiwaLzWc6p1gB0pfCNnM4QKQeWssjK3J5iBJT38dC
IU1HdjUu1Vsw+XZnioo85yj7IMRmUTYo/AT/MuDGn1k66yWF9NBAWhI2ono+UfJQ42pXt4qs3Z87
3xtXz5QA242737AVx8tlo2aTP7vY5baUg8t5bP7wK3nFkx1WSe2EVK8/sfoozvDDxJ4cvJv8uw3K
LjXWe/PHSGDDLIpEBLyolhW+eh7LROMsFF0OkxNnKZmbmwVF8MkMZZZyJYwvfaAN+DQmhwlY2hfR
J8HV8Ew2kgzhWYlgtsBf4/or8R7ZKHGwyfoOmqpEtbeCV1TNfwjDr2fBiBdTbKfR7EbgH+qHZR9g
9q2IeMeEjc8axajSFxJd+PNoBG3CLptTOvTbM9cYIBfgtIevwcWFb9iTHwbbDfEuJlFy/TWLf3p3
Im3tecjguZz1aUmJ4POdXWcoqsuct1pk4UvxvmafzODqQfUQ6lpHTm/FLaMy1Z+OWqq5bxLEoyHP
Z92zY4PqRhS/Q3+uZVHjZZg4cGn9Jj2aAGv7eY+XK4w1/jsHhZx16sOf5dMFJ27RHqqxx9hnUj7Y
zDhEKipVFHFO9tJeM4pGHoRobMm5uYIM88fdCfVKyYValaFWMjQPN7Hj7DNixYJlT3W+s5i315I9
MIhpne83qWeo8ChkiEAp50HGlxkxcCPaHayE0STcsgZYHTqhMOUjmn9jhXLrV+qayWY69HWqh/gM
MRAltgXNxGlimRFoTnJAzThYHPbukItdzAaqD7ITYgPLDAuq9nKq+zA6cXoQatHwSjkNP5pMhnzO
IySKPyfQ5vrT3cNOCY+X0FetGtQ85uow/bqnYkT4cmGNCOq+q/rUawWkKJsBDrYwv/xt6p6ORM27
97I5JUhkpU5Iu1QZLbqS+BLHoBK19geMXm7DpEkLtkz+j/ZYQXC9+2olwD9YeJxcwWjildisoWDR
Ry6fiumAVc7EZNhHVUe/2TOhVWAu2tABw/7cejAmXFv65jRzL2Q5+COh0h4nZNRlTogiwiicGOp/
R1Q8DmA3k6zl4bXeh1Z+1LyEs4G87Z6akjdodZht3+ruBES0V2t1nNGjzs7kS/2w+kw95CHI1Qla
TgAY0XFm/KRvgofJiSczHC8aO1InEYeChT89AsEcQtl1KXyUYqWEtUsipZDsrAgHjpwt4AZhITRn
UY7F/MiRezC3W5K5ivlefXcJ9/CxeM623QHfICMV1vKo8r2J/l+j1sE7cr6uRayYZ90xzKIFFMpt
Id+SrS3DqDBrLGIav28V7ocE1KdtMAiBqsne+HmT025GRnphTLElDLrM52Hs46Vx4y4OXhCB9Tyy
9f/ZlecpAuhrdCYSb4J2lJ0K5cOPwPurhRDmLWUA1GaRlSk0uStB8juf5f2zCWLdm+5kjcd0yWp2
oOkImiOsOQUeg7MsafkATVZOz6NkU3yUCxeyucQtPUSD9aojzsvCHY3b/1fEEBxZDpZKN6e5d8jU
E1IaFprE+um71lNAkcxAqza8HGC0l2vtO2NYLvWC381lXaF8RXIRj2Wl/zzJDXX+LUsXHVeS4tnT
wU4YNnelRGJwtUNl0X7L4GXY0CEwecMcIb1oKwpbwHH8fjI1UozN7/A/lAAJz/hRzZ6qZns6pYkL
SRDCR/gMTIqJkWwjBIuRJDi34f3hfuVgg8f7GZaxGNhP4nlC8njL1eR31CmXI1nPSFfhMNDONgIl
EuyebGvhEkcbJIv76inJQ78lHB8KfNUTzhGqqp/oAL+OOFw0bsmD9okWmWZEg0PdXr3ymRiB30Aw
mDBDpEuHh+5kojUI0fRL+pKXCOHsFY8DUrmHvFE2OdI2Bjz1p6einZLDTWlB3H5Z9TYFtvwYxMJy
4pkV4xFWY0VQnPeZ+cL42mlM58tlTQSX23sNwHHLQr6JJlkonHJgcIsHY2nWbwZW0ksx0r/un93+
4Nmn6S78mJ9u6QfapocUZgaJbXyzNTE6KhYloNIaUc+pT8L9ZdBz816j2F9kn+OsTEpraBC/PQPM
QAfr3cbkjpipRmW6AbGzGF/m3BOH/jZN5lyISzXNrh/hXTZq2oWbJgX7qCwTHgjhV5AFDLTrSnVy
tJXfVd26H3UDQQlGWixpNRjIrBjgnZxy5zPlT/Y7kB+2tBTUix+OWDnzM6EBwVGDmviOx8eshZPX
WzVkRQvSzMSvquRIauoT5lEb5kmiy5DmaWCnsN33elOi3OpLB6otVTal+bXR+9MftX1kSPZA9us5
0E3iqOq4/wCJF4SjZOP+S75YJb6hAxCEV79KmC4d4ITRiViFoAXZMgvaNwoWe3X816XObsmhXaPX
uZcfyuyRD5AAcSGQWm5qXm4je71e/Rq0C7jGY0Eo6Ka/6NAa+4J/UoSw/pQHZK8rqswV/mrTiKXm
PxW2oV+RhyAsUPAgl1iNdvhXxJcMIHYLrt3sPkAkaCp1ATinhkCGrEutf/OxLszc3lWy4K6OZdVq
DGIh6EVAsWIAcXT9PCD5JVX5yhdVd/3tNuvNLyCwZbQ2vOBqM/s9sysvinnQolLLleYuBCi4o1oK
WuFryNhxPnWp9peA6oX7rZT21Hz6Xq9sab3HlE/nJ7BEe/gfowLkJWm5ekqLuxG7mbSdXceuFtrm
ZuQAr+ByT7hWvvmNsH3VEtSuvO+8iKC10vlgThW2evua6Uina8GruzEveYL20/i7VW5i4sxwp+ef
UxdvGOGZoRJ90O5zSzh2YeXPVDgbOwRfFNmTC/JMBPiEkC0sbnc1+BBezDxJLp5Jk/9xcGmm0AT7
lYBNd/9htwXHcVM9htQrEz2b7zudNhmou7eO+S3kLsj4FN3XqX9MNRMvAsyFhR+6dwLk9xDR6NJb
h3TfXqPATl/stDAjqDYNoZ/iha5WVjaRV7F3ZqzdhAe2aLPdA+Yd7HxcRf3qRwEVkkU+X2i19ejp
yi9WRZViP7hwXpEvzDXkjm2x7dmJpYyR5LaFyqmcaMhnEMHl8y1gL9hac0mJZgb7ov/wvfZYFZ5z
YxkQiFP+ln48FOoPqsccHkdeVq/zj2r8xrW1cY6WX08t65LMcCMU0Z4E1crc3amwRovqRNGrreEr
gsEIC70N8cJzU3WrnJ+rixyaFDI0l8GpVZo52h9NARWeyoCmCELTDHCu23AqyMcXxSJOjDMTa/z+
Iy3vcpzWlbUxBmLYGUx6mYlxET8IgpVjGCamCl7bbP2H15NDBQpN14JTsVdzRkcu5VolCKbTrh45
dfsCtdmIEu+0c3c3ceUQV5ScwWz/ZH0K59hYH5ULwUdCTBjmHs0JJTQq9KoDfAF6kglMQDJtZJVL
/v6ZdUVLYdJFcHB9G+W34kOT9HQ7pe88W/9V9j8CxmTMFQYk8wQpfzvui8yHpSIJxGvRYeYZK8GR
FFSKhtN/xWASSCgcp4vzzxDdOqL0TXWJvZt/QNQIGUZcfCqVrViN0dCP7v4NFosoC6sq/PHuWZgX
bCY4aiofUC/iGlWL70uxT16YnhLEOpMZrRfI2/i+Y5TamakZquZMd3ZMrtAbD1Zlal5As66Jr3sB
lBcEZp3x8Mcdm19HK57nSXYZXQ3zO07Y6ZBN2Squ9ybDxS8s8ZSYlm6nrc4k/QxQxTeBuOgS37rf
ealzRu7zYGoOGrAzcrR+INUm7J/GUMVhqN6nuDeMT7BAbeb0noOoBo+w5CQHkRAusCdWfSdAHxBs
LCLs40lznkzZk0n1WyE3KgmUw6wwYd7+O+DhYqJqbI1QTySI+Q5jklSiPFg4/u64nzxxy4vE5X1e
s40RfmSzDQZ7oPwQpotlO6ZzSCi5vJzzA0g/L6y3S/JkKJPPuCboGTmWvlOAFeVkFSxpjnUTaYJ0
54Rj9GAgo40ZiDGPiExeOWvgTFqAbR0Rzz2H4k6ciznvxrEHAnkN6w+BGOUl2vBNV0rmPdgO7uUJ
LMB61iG6/4lsMzuw7P/932p1WSc5hKVM0IK286xCh89OXah+rdnHZwh23rsyLIj8e2wgcUHx74ON
Y27wjwYbHoLDZiGcQDtW+Al8jxIsSiBHObh5UrwDZiMTlcmSMpW0YLd/k021Wb/NAjd6UUSC/fFG
FMuYmX6e7OrdevXdVHTHOEE595sSSqS6MZHWyS4LQqaoL2L07FWLW3s2eGQFc+z8WN85kP3wcqPk
qSJUTyTJzfCuw0upLZpN5ZbhKtPdkhHwyr5HrA85z8J162xCAB4oHyOAorf/xyiizSbSsnutodkT
CLB9EqYgmnV80e4gefR7LR6xowCdus1fmGDpF8lWiok2D9NJJSMogoT3zpNYYUJqDUVA9ZclcOZi
wrhzfCTdLc/PNTC6+3F8PDUIv7xebeZNFJug/RNqZIzFMgbqpVNulRfoLvPRy3eG0zrQtbFSJA6w
mJ3FlcBc2mSmwdHAqROrJ2EZsgbjemEnEIMAm73D27Aex0nNpQRxZHaOV885hZgEjeHBj42W4NFZ
SfaLh8jlbivdJXgUMWDB++Q+H29pCkGX3ncs5GKiRAddkbCS1oIxvRxs2XvD0cqyTCgDY+nlwR5q
HkysAqD9CG9IyGHZ8kOa4evZbSBw6zRTSlKBqKGXCm9tkGfWNNV5ST77inteIIRWdGd+cVH6UP3W
VHB6sJsR6FM//yyJs2zF3pA5w9f8QuTer34BzpTiQW75HPPjx16QA+/4kgk6nI0SqNHVzVdnjKQY
BoWZsspsrkFKr9bJ5WyeRc6WyVf6ewlr9DSgRMOchRXUrb01s1OpnVEKmUTYkMhZX+c2PFf3gBVl
e08Pu4KuQ5COVj1Xq2CXEQxlfq9vs4ASm01MYX86Mt+BMqJ20OAkx/LvRintCaowuG9+ibpBA6Yz
sz7wUM7usS0UnqVrwDiQrRarUmDRb6UT4M9yfqvnmq+Y+jAlKtYv8DkY3ZczMFSrYaL3ifaJ6YY3
KdPsfnTRnfw4yrvivpIuyM+Iua0/LUFgS/YQYOz8ZCZqYSvBa4RArtPdkGSc4uyFAjsleEs8Zgod
UlZWKfCnH4cIcnx/J7/lJJFQ4bJKstdVPIrhzk9E0OyE1WA9wZDuki9xuZGhC2364JjfmmovqbVq
WVoKOIJLGnatiY0h/LfLrWV/0w8821CMKns8HDQlJ9hz6gONZ4FzIW6/vcM+XO45AR6/9v4+diUf
sMv/G/ddf0ERbU/zAgLR7HZp///7d6tg+TSuNVeYTpKr7GjHDxKxoIPEWGDKl778r8cPYHNYMVrT
dalSdZUzbu8eOIk0TgCB6UY40aIAsswMtABY4A1eQhkyN003tFXgllxGalvaNLQtsyH7N14n/r5r
qB1d3CNvFvPDu0MeeyIsFpl6ofiINeFgjmG+pN5Qz42aiU3ZBCEeTlzOJJWrtblWa4c/rZnZHWpJ
GrHkkpsVUKS4UP7awIKjWVlS774vLdy5hvy+34hB+ifool02k8bLNyUBEL4HyPmodygwPFbW9Z61
90/a2sxPhazcEwWWWhUInE2loWFtRxYT4Se0iKUnn8eeOyzAEGPg1T6zQkx4j+0awGWZyF84cjuU
uBS0KPEF9wx9NghaeCkW2TV26U1oF/nnYmqf4xq1Z7RlPXyVBgCi5YDUK2K6H+IDLWF3wAROgXxQ
35q5xoLtJCSGB/x32oFH1BcdW85ORSiGVVoJQoXwI4iY2CnWNIG6jLz8cjE4pljPZiUv1E50WN5Q
v1wrW0n31/LZ2wnBSOobUu2DkPKhaQGyBE/xriTUuaL0N/ySYGlsA09Pn5cQcep47Ymikdpwi3xd
QB15AhUDH6mDQlMkZLVkEJQ2moQAHiMKdk4SjA0mybWYnGpnvQe+puoUf6OrnA9YBzlKz11fQtZq
SzmwuLJNQD6dlIgV7hpaQu9XMwuKElqoY/3Ywp+fC04VZYRMTTlbeht3x6U2GAfwxY8NP9z9BsfK
0VFAV+sb6SN6i8DCqp3xo8TU1VGtMx/WHGSm3UJALsp13B3QUByuVut6FG3UquLITaCjHFjCyc33
HSB26SStF6cu7hGnlsFWbL90SYfxwxjAVzF7o+szeNBH3sA7/jE5+WAnlvoWns3b9qHjKp4tmC8B
tizqu7i1gN4fJhKBtYAneVRC/8Y3U/y6mhbe890TgYXfSKXGfUxQK7hekARsd8G0vqp9dYjsx7r4
nH6Dj6zqF8hQZwnqKiF11N/8qYC9iDBhZALZ+mWAnFiQFzCnmA7vF1lEDQOMj8pY0SoGV49jkO5y
Of0hyYcYNBwbIG9RJIvHsVeDvCa9DvhgEYVjqisveHzaLRk23ul+G3xb/o1ukGxp5BqoRkqS1MFW
iXmo95WXnerdZX5Ul0nnHn0/yLdi/olw6lt32qZK9YlI0iW5ynXmdJtBBSZdeU7ir3IXg/EIg4ue
UYAYtHKRboexTbo6oL3SBAaCC3JrBoy1f31iptn1mQ0bomJSxNGtxBHZNnPzz3rAIAdnAs2BAzgn
pvp4uZOjVquwRG65etuir8C7WBXOAPY66CDPpRk/vBkCE1sAfggX2iEyuzdfIFfnagrxmIEM4r7k
2oDp9KM1SNQvDnGZCi3xZ8M3X5RCLrziUUI+ymzk2fgVxoDWAzYiem3/JSoWmiMieEX0Tk1B89s+
8yqS5XedPzB0mj3Zz9wNtzu+mSCKR6zdLABTsOmt/cA9D8uqTKFZVflXpZeLucKW2S5RCH2Jh2Y6
rOh3QxzxYN43M3LEiZFnmcNycZE6XLSwPeOvfg4w7B7qWe1Xpckqg1YR7RQddVjodkVBiwFwT4nt
wO9eC84ba2qlPH6MTDur/PfszN6Sc1fJtjD574Vi8jzzGv6IGUhu29Klzgd/E5ZwyXSWr6I9pD7P
AKQ3zPcBJ9iPgCdAUI9aeWBVQnOM1wKWesNUUAV5W6BR4YQ01ooT3tsO1eg0VMe9EqDnZoOJKRCt
aKNK0IfRRqDv8ZBP9E31Gf9n5blx4KgxyUYsH4mdAhnrUyLtBAAiwcefWVPaBm0F0NSCvAlrjz4n
81NTCVV+eWFeDqh4aQnAjHe3PwVokJ/sssoim06xza0kTuTJ5UM22unTjAfgI+Rz858A6PkJmduU
7OpGEIiP29jFA05C+p4U2XSVmOKfuoJeKd1OQ5xS9EcVFnxHH/z1AR71dfgc5T30nHdCym3U1I5g
nZZ3FmB80zpb1wZtvRYUXYSjMUX0TSdyf0Nl4rnAvqHmcZVNTvHklJLQZvtjv3w53ldMCalA5L/E
qHBf6u87EItue8dF4X4+OfCKXCyASlnquYNWUNVIBtBXQHkB6YYgfexESGVcsDPxXjLbzvF7jR2g
BnrO1GTgVDqRpKicBh+xFV3lVce8/WDkp44Ffcx9PpXbi7PRxEjOwvPvUbgY0HChZMAN9qPBZzls
hGkeJDjU9ZIS6r4a112P7YTrkSPDvZxBq1ficAtZGXXFkdik6YyD4UhwqZZB0805WYYB8hPNqYF7
MhrK95VNxNbz84kKtmuGB3aPg10wtlgwlYh4/tv/OVauKQFYa6FV58nqVBHBTGvkkWzlwcAvagc/
LAyUKPTTloUJ52U6YHZn76sjiR3qBy6O4K2rJ+PaEUCnHk1f1WmEybEWpfw2qHsxQbEBFHhpeXCk
fjMltCA2CX44wIVm02ZbVVmLG0usNaCJwMI2nZXCmL5feZ/c3wV3ouYBFpV7LfPcum3qZ/Hw+2y0
zKF4455JzdjwzEP1wLHvWuTKgFWbo8Wt4TFeDypANuiDI7nff7ElxOl+xgCGiIsYx/5aiy9TOFVo
MTyF3b5TxFRODw3c/guTERh3A8XGAdwrJw7K8dktA5GkMsqZlY79ovce+qH64QId016q7adgqO6v
TOsljOr0uauuy5pm52RWxLS0ooWS42xpqIRUXHuslZ0xchfWXNbg4q8zvbCgA6jOmfgdJE+EgsYk
IKFIlzkGi2xyyoSgwIdb33T1Mrck5cGQkSXhkpBSKrhA5ADaiVb6Abz/4WtLpWqNmxkrqyWs4kDX
yG0pV7/U99z0JK/bQfAQ/WoIjfKf2/aBG7wr7EMGpzZ0VCKJ3LZFfVT76menlxQito+tQOG+fIIS
NJcspCnq0PHRDO52E+qS8O2UBrUlo0fkA8lBMOhQpa8vgkX/sTA1rKTDDmGaIYHiJRmUI7OgwUTp
clKRYW9X+rWzIOWs8hFrJHevOYqujePpq78zWrNZjs4P32MeDVtPL0yam5ML/h8JhFC63nLgu8zm
E/dvYylg1rXxLuXcejtvzklnUBV++PDS+sP/ni+b3FJByr91AsG6+WbX6N2FOxoPm4BHSQA/jJtx
s2YYSyUUpVtwTI4VEgMmwpDlgltn7mYwymAzrZo2DvySM5P9xlrmL7BGEgG1SiO3n5as07vdELaq
aOAT8kkxd1opdxkU49Y5Qm6b+YAAg5KHv6jfKoJcfyuLMJsV/nSlRdqP+jOTEXJfBa0hPGZ3KlNw
Yrqzudqv+tJOa1flS3kiUIqw+1SAvuR2TgtccJ1GCg8YHYDBoMvFeO7YvE8XdFs4yUn0Nd/pyh/V
lb8FZzMyOHN5GztWOKH27moBKNw9m3vRNYUd6TKrt/nUx7R4r+OPfFSk/p1FsBHLEZfL90apYCDk
5URsTMFkKHjhQDC7XVvb8G2J5gCVa9Bvy19INxsfN2ALQF1n2hdC/qP941XdPfsTAeJslMjy2W9T
O0Hvr+eVu4YrUyAjWycOVMat3XCW/38mg17ev2/efCH6Y2VtSm74j4GnsYiaJThP08iPDCybQrNP
3jr+Z6mKYwr79Lzl3XEXeN4SCZwiexgtUQHo1Nmj8guc2LvNnoTaTe8D/FT47YtjgYdP1HTiumo1
jSjN0Gk6Aa6v3N7QxWcFnBxLut15V/wbb30dYrREhGzvhtNcjIn14HLLBEpMLoGHs86Fl6f6hpDt
OR4tyTV1BWqzVb+5Ww0TLAX5gOEXjRlmYzhS8p8UDUl52Pl0YicH9Jd0+D+zJNwyl374XNaoBxu5
NpaKX/ruMGHY6whEiyWFFeuUAeSIM292YFv7wFT/l1lnfD72lo9OedPXx8BOcBE+3KZ0TOWKyJOc
jCocfs0lAX1vDiGU9rO19tRDVR2nzHwNCSgQDzEdKCAtBRyNJsqYuobLGbhJBj7TKas14UUoTUcK
I5rwSyxzSv986IAOsSxvv7k2JSDal8hj3ydaki7BfQN3RLhx1Yuvdlku10P1YTlaI/3NgxSkZpGL
ttEJmOLIJ7X6nOOtgt40q3R3crrZOASw0P8aipryXyijbkK13uSWKPdD2nN6Ejs+SgB1UyPCC2fT
HCRZadBbg1Ykw0vjYp8QQpYef5iie5AJwqpDFUZTPs6+ip12UeRDhZpoWGsnkWnfBxbEPfXqIxhM
lQGJ+QHl16Mu71JLflO2afiCxlGuJvZ6I9RSybupTZB47Q7t/EN818p9+dNLoBtbzcIMJEydSNs6
9TQ7GFDeOLq/oxgomBtLGo4Dl4ZlRaCEN3/prfcZ4PES5nHfry5tfq0PY9VFiOZvgVUQzuaTFXAm
7Fpaxc7gLkHSfStJzNfW0neeNYDPw1C7kDO5PStPeOLwHmvv75bOCBvuJOJv4yFaWri7Lex/Jfqw
sB3w8Or/H6QBV7qnNX7J9kP4P1rupHDA/QRGGpUU4w1JLUv/VNBelh84AkylB3oWiXpMx8peiDqO
nqrcNnDxoG8k4S5c614g2b7X5YpT4ZjIzXXYTNyRm9F0XCuTemN7QiEkMcJMwiwmE6e1NUdDU7Z5
5XT5DH37GGHYzj9u7fmUWSDEfOIGHVcyFZMAZR7Y5JirOyenkBm5Cp7EXTs6fLm0GWvnQD5PsEvL
ahdPsHNESRFI8DBwKsXZqueOf+Flfi2GoqQvwCr1A46nMgnfFR6iQMRhLp36Gzi1Xww0esHQkyHX
k5CHVl5fR+d90xPnybXAvwQjKWRWpGbxg0ElWn2ioMMS/dtiePibYcsM1W1GuTAumwuNJ7ia6BCq
dHXxsgAiaXBbXwo760pUBekQ6h61Tb8SoFKYW4R7YQ/6XPgbCYyQpW64XzjM4CT6+/jQBOS19vy2
9vh2eE/EYnYMvmwp8bYDyIOUOkMOI/OEfq+CGuXxrHGDAJqCmTobX2dkCsiYQFUyBAVspPvInaQv
RPIWwjjXSAnANVmzi77eXy18+iK9pRZyp4tWjcoJkJzmyQAzWZnVTgLkuFk0X65xeFAce85nuJk+
rN0zRNGyKNCcOA+hoCBOZIkZ1uRVyZ4EfziNde/Poy6M55hgSIu7CHj0esr/OXuE/xVpuXKgNpcV
i6KC7+9SHRqloZyX3CGA08gPG+QAVQV3fZxcTGR5BPYOjlgZi7vJ31+AHp7CilLKxMiJ56OjSFcw
IYsy3CGXBdn+mGCTDQa6RUpwXMGkBiryn67XXxWayYqdg3zfnn4lyVuEjPBe/rzTz+XYYkzx5sAp
YzlLg4hWxolPFS3QRfTqrd0u5c1/NxfI7nDQbo+67fZEH5QBTd0MMPA8fI99DbsoFiZfjPUs45+a
dTFSuocgCiFMqqcIE2L7Dap7YcDxcsCKAYjlq8+wTmXx57Y2q2pqV67kfI38f7R3/eyG/ZBs2k5l
wt7hoLDauWbRDLUCCgiqIKD8DVdXTjiKvI2+3zpb+7E6QRoRYnCEXo+rCB34Q5gLemK/8T49qoV+
/X1rNUBFB4ZVZaI+dbha1R7T89sSVFsrQpbc9iRfiggq7vtmvLg+XzOudl6msX6Gsem1uTyd9lpm
VfbGVp5YmtNsa15TVTEtzLKERdOqtFZtl3n8vsAfcEhU7cTXCSBk57H/3j941ufhiZM6Q8ZB0sBj
TzbqrCY4SKCot6oG6gyL714UL632+TVp86Ij9sxQZRcM2WEU+g8FbbrwDNF5MQ99eai3dcJyY3yh
u0oSRpAZ1UTD5IiIW0u3tNSeGTRMQU4OS6tBardYbLNIz29rle3BK1bcC6kbXCeSC5WdildKU28Z
5r8iT4szUVTcjvg3ogNBY9dP++L91TUh40wDmV5jtE3vHPW1yS8rJhW5fpf72P+wBRPRgp+5tijK
m4iz3zbS7zZdQaoukGoTNwSznVlYz/OZaL3sRPFYFBf+ws38Z2DlY1NNZORNhjRX7B77ayxxA8rO
CsJbENilhZoQvSf6SBljQvfRXM2O+b97nw3IcSBfahj+o1HCJQCvbD1zex0dXNN1vUSlXsP9t+rD
nidENwsXVTqiNlPEFgiUynCoO8Xw32uMBXm/9+lChnrPgIpu+xqzci5h931b7MBMjYCzMwSSoIic
qHsCRVkLTEd8HXDZaEqsI/vMebUt9yKX1wL3DUFNxjIMqgFAW0VCWUqRAUsFS7j2XWmVvPCKIieB
/22Bv69Sv3Ai8k1k1BeInDmmWnSwfNiP9BK7DxHSkR3EbnMzDbj+dhmaW73TSZZJ1l5mK+mCy52m
P5kKQa3eO1xVRGfNsv3LNgWxZjr2yjAwN+0N4sV+gwFFQ+NcZZtRconq2k9i1dW8d38UDSm4a/0k
Ff1V9AtWqT4bp35NbBFpCgkOnpChX6lnfwMt+ze6RVJEwi57cvzwj7lOfGhOIAQdh5/jF8cZeYJS
ZAzeoDHILPa4qhP+frep+/gIMg06NrbvhHKbO1HSHiIXcjFDnBPb3gf+WcUVvxpLDyfdoBXcuoCu
9rieFmMA50nyhpC/yj0twlbwjL/wRs/SoJfon++/MEy/N8s1tPXGWj+YfhxZGUSHrNedWSNE2haL
/10k9tWZw4Z/gXIcQslckdONcUcbafmrA+oJJdpYfrcubOPdTgtmwxAqNDJ0PB4OukvrmHxK9pUP
VVEoqqew/+WdQ4XmdoBPyNaGfy2eQeTXzDEUOSnwowaAiOfRO0V2yTCYI1fCTx0rNckkh03kiwFo
Dy0H2zHHOSmBTbff4u3dv3/q92Z2NvElCYuzV2l2dfftCbI87uUNLgkldfmasMfx46uxjjIZLxdg
Fo64xwLDrdex924mHF5WLQmcy31gYrwKvwS/2FAYc4Xi3YpqoV0jkDBu9O7ZTRnL5uWF2PcdlHQk
EVGRcB2Cav5UYhdF+C1Z9Y/5cF4fKuIM087VKn8cYZTSbb6IxAjoY5QVCDu1Ipt4B08TRGRy2zXt
wulO/ce69ENq353l9kwPcd1sBJZJI54I3JaCyXPFEih4FGpBt8FVApjT7oOgPrThSMNV/02ltGnS
H/ayxN4cFQ43jc9Vk4pqhQjbEYJPxbldOe9bb/HsqHxKh5CWZrnKVYuF7qYyaJvYycJf4qyhomt/
QT7C1JRgm4FnN1+9XpnUYvD6RH3liF1oPfabZE4NO3ozMxT4Xkmb6r0U54s7pwBYgY3BV1cmyDWN
TMKdTEb6uXHVflKrOFIVaJGM2zXYf4CAND3M3+zY3kqoQxbcd8U82zXPGJvm6ehgkY1mSO0vBCx9
RGNUPs7SzPDkLKn+4MGoQ8O7DQLzT6s6X3+2wbt7uiSrBiqeeJtawUyAkFbH78DTVZqR4w8b+Okp
kVpSgR9ML7mFQWAqSpOy7/JQUstxATbKz3ynt1suXYWEmF/JX7FySUzqW6IvdCu4PRHj3QmBMpKv
RjPFWhmdOkG2pFGS4dUqvSKLs65P7UzQXKWuLbZbdRqirOxA4zA75h2qXuT3IMuKdbFPa/sdV2K5
A1aQysmg4w2bSn6XVFu+ajHaLlHsIlTW5zECg2cbHJA/GV3gbzk/Tu9ad9KpIHqt+XkCIJL6z7bs
bPZ1RR5mBwtnmNYj02ZxNOt9geGtro4vtiQwV5ExGvzIbM03R0Ef1toa4CqtZ7pV73pqDjczPinr
o18Xn51eMxN8sd8K9iW+iqFTrB+HjCnaTG8i2RsFnr129MlOXT2YVGToBsZiBC0A0lm3sxBVJoW9
ON5mxjrFfQO8QM9o67HbL3i+m6e1nbAgepg0MfNUjzUb01imq2aGOqHgjuoymbc+k9EIXs6mn3gk
TLzvORgCcGguBvmvlXKihSv51bH1fzi7SKaKXYsgEjV2S68N6mLbNChvrsa3O6Tx/JKJf4Y16U4L
xwq493waYvwbNE7bPWeihJgG0QO19/2oNG+Zq86C6TtUlbML23CYTP+6viCtFWr4Gdq9IxrNOMGa
Vi87cf7GLy2bIVu2+gBRSpujL2gEiKfNNBollOWP/8M0ftGi7nO1/Wts2GZl3/mzknmO6AKoAUYM
6AREZoeQ1x3k3TgFfYjt3AiBgl/L2AfsZyDznb/0K1dugd7TbckwWqdJrHj4Bl97oDzucs8wN4p6
Er2mGaZ6BqQAej+jx/No5cgZtwrK0lDPoZDt1r9o/LnZbxQyxMgmFtHBDoQ8PzHCq/vgtEbBXrCk
4PvyZEJSkCfi8YyA4OBNe8qgV5+VZFf3q4eTXOKUNNGfrlr83Te+Z4UErs+c8eHh4cbQCgjg7MbD
iwfUvt75O8Hpj3to6IUpPpVwAOfzYANy5ulS+/yektZSe1ljRS2KMDsSy6camopzmk2jrAp8JMAW
y0BvA1aVLw9oTnwuFUDK5JY3pvyj7Y1rUayiApfzC6a8XgdYNo4BOHug5HqAOXp/8yDvDpkwL7I0
bMw5q3DrI2A9bUBVQJJ/xfLnEr7J77Clnl87FQ0cpNQdRfUwyxnNvg3KmJwblBDsDBVx6ErOrQtT
uPu7j/YT4DmLMtyqO+fLqLEAiZuSGn13l0CU0+pXq/3f2INEshgLbitOe+Zyi0+aZY63CJzGMVPU
SDJF2HDwonpZlAmW2MCrG9ZAZbUrlXHfmENXCYw72DQFnVq5H7cqoY4khSyx6J7SspVT5W4BaYFk
N2qSKLPdPLA3g6/baHzn0DONbfEFesN1zgkJGTLJkDiuIxhexdPPYGsMg3/VayLQAthrRGXwD6Hp
SIXrxYBhq/xrp8KJr9IgQDbRCpyTvKqUhRbN8x2y/InvDOE8voGYJVss/gl1iyhxbdlEJzX+rrx8
a4UWOpTdAnjx8UTrSeHdyCZzaDQ+NqU/AieoW8fd/lRpcwHydznDJAGtwPNtntlj0FM957BJT1q/
hNy80/RJOE4SsP4h0GnMCH6WnkNVOHZQ8YvquosjhDkDGURC7uvfpDDPj6CmEV7IYEspN2vKSz7s
8+KTPRItNivPwc1EBiwUYX9d6CMFWoeKQkO+Cw6aBDi8D/BpUyPQ4nbcJmpdwCrLEIpKV8ypZR0+
f7qCLGX410dBDCXK7F7OvI8PdAZXgbLswMHWrS7vpgbrHjrSIaNjXR4lQOvbLwOik2L7YUt33r2t
VLJnfJfEg5HQ6J1poEiZrh8ZNZRiwqyspmhNGGK0EjMhHNmKeHdu/PEpGMHPafJzXwOhSLJw5eRt
GqLfZarjka4YEgb8a5gGws4y6QrEqEtRI0kLxRBbbDIc+D4fQX7ZZ+Ip6c7ejQ5JpHDnp5Zs8yM9
J0XN8MHYPqmGwKRAbED7rTQIzTdtUBpLeBIwfalvhe8/wpBQ97htn2tEFk/aLwSpx/K1Uw0XbpNl
F8E5J6oWjJSRqajB2bdsJreG6KSlGnGvPqFYii19cy5hVDczPrt6fZc/GuMb3CnYf74xMH0yiml1
I9QSZ7gi7Ax0uPq8h4J4lc59EmldQxveby+PPtGwbkJeLqQlx1ljoCJ9LhGhps1m+jgyvuE5TPzz
zA4OnBQv7LKANfQner+wuqQeBHjCWjcnzgEnfsCUpb1i0UyBOKDIVHY5TbYiFH7QDTJTh1JKVkTD
tYOpQqQWeCg9Cy/VKuKSNNWAoqoTFnE2lU5BdCu1w6LjfLaj3bShW6jxvOcmMj/jDQabMWVlG///
+AIBKyB03WfbbFmQG8+da/+ZLKFn8Ehv6RZqAh2Zgj4fxxTNmlK+3ysAE6L6Sbu1JS+a1bKa//qg
9f6yMO/qfg58eQFfWFdADd33tYquPrUGzCYJRPo9gUm4UYjsI1U5FALhLg/eaDGECZgz7tRtU6h4
IzhjMBoaXUdLSI7iSd8wcWiEmq5hWRUTBp2oYZplqU80MZVCrrcUGLItc3sY1YwEkRVZ+YImNP61
Y3/6fnow5O8Ogtl/XDMwE6zePsAz9KdwGNDYlGMPYOo4xs5AQeH/0qrqnsLg/fBZGhc2IfUHlqPj
JLoWFIT4n4yhW8NHYePRFHHDCHHu03ER87A1dsnnmg0eUcLXwQeJwZ54NDJW1bU9WtIC5kEH7Sng
BLzjnj8zqvrGzmGdjx0SBmUuV6h2GA/hKBf09ZaCGqArfbvXlx4inpJ7Os9FeXtEGEkHNs19BUxt
dq9Ks7N+ogblP7OrrEJ9u//72XedAbUjej3p0JqX7SWzpV/E61hINrUb1y/5AeGB9tkRB1HkM6yv
YEcGQzw0lvCvrEst8xZNg0Vcens9re77QEhDe9622K/Xtq9mABlHaIF5FNJdfvObgW9UZhINpKYe
VJWuiV2NC4mY41Y8317yHkDRm2bYIQJ4rGijAafjhgm5hevBzPMu4o9hFQrh7zxcQfYyzBtOgfbT
F63C0Vy8cFY5JhSGq4sGZ6If82LHjbL6WEc4SAOn8x1eERjtDR0coEE2Pijd3EjDcchoDgAW2gCU
XydT00clnSgxUT3e/W/Uj6gOu+9z6a5OPOjcYDvPyCLokgfwivamiyjjW2fMP/qQKT47YuaxO7J5
V1UmKUdqARzKWYEVU1WXRCV00OF6GSWshg8OqxhOkBM6P02GVaXUdeKOOV4roldSfiNtMJftGYhH
77lKWSCvfvBnIqkLWZXTdTYqj0McymOzVuMdKRmz67aFOx2GuwGMcUApRY+N9DswqMfE5fFeIfKR
Wu2XfihD0wIjvZY2V4v8tcBgg82JvMyon3e5DggBAqhBnQBt+Hr3xpDv4zTVp4KP/MmaDxeBCzRv
sZelMXJnU4DBjgHGPNxqkH8/oJTcvvKkDuQ0s4ShcybXwTIRAliuQ4VzdgIKWbmLHiu5CSQIF9Cl
bI/JGDGGPR5elzsM9bBfhUG4mxHArgihrL4Omd6ElYJunh4+Hh3kz7JrRIE40V9vDkgZ5jmKDS7B
kNOGkGM+MNgo0vnsmG/wYV4xyNMoCd34Ied0sIw+GEUpAhlniwpjHv3YhBOkNDJnZUcFBN8Dfg/Y
0Aj7Ub5kMdqgmH3Pqg6Io+tF5yxawktrH/luQHEkc2RWrqd8YWGNKep4jrXnhZV2a+hWTCQlE07w
dev/TVS2sCwEx0GT1hOr4JuBAWO7UHtkbqf7AWeIkN+F/1YqcjGyGRGZHy499x0zGGAYY2yDUMSM
gUrvR9EKdBhZwUe6Lt1R1ItUzKal/YKFOZ3CqF6pik/U4IKwxVW82tbEIbHgnmYJLGJxE6dkrk19
rIeK3CPByGWIYxYejvsjJyTOnwoMBKOrBRjsU51DiVMWmFT22IH6ZsLT9efyRggYqYWV8gMk4EqL
5XKSFs3JvSS3Bfakavm7mQrJQE1luatLUwM21deN+KD78QhgNMw7V5JwG2CCTcrXdsykYqEulac7
jTqWMsyaP7HmTEH/uKIopThQgbOT/rtILkYh5hVwXxMolXu+16DDYeLFT4Wc8v6h5hOYqBf1TV5d
xcx6XaGpaTErQvnVhYuLghRp7kMhzN5WEbTl3Yr3FmzIAN34RnBBAv/uV+Y1SzWI/vlDQ9c8nFnS
jTpyciuboRdL8bJs5o15igXEJnJWO4WGhsiwuZNlqjQ+re/eHSqAsPqyYuQQg6zNBVX+8ouE5w7t
gNKZ1nNBA+SyLVNcZLKEXlyCYn+9pLdYPNg0Wlbo3umS7n9ildvxM1frxuk0WXzIsXtehksED0uR
yq30E/g+1BPNmBONKsmuGmVb3Sd3SM2zARGf+JNBsDQrJyr0XHkBfyTeUMMwoVOO3YyFcZXWkg3m
zvfvTp04P9MqKofL2XXsZJaC2CAMWWRssQHKf9elOXnxwYRqlYjtHcvMeFSaGvDBILYGq0O5IcIk
LR3eN27R3T6q4CHCoQNb+wpioyk7O4iSBaJBbTlU5pgJC16lfhY6BjXUEa51/Oud5D6qJkm7SUVg
+JmyxJzrIY5lbb6WtFTtZUGdmjiIRGWuxn0OmUs31tVBujnBozzisnAvosV0VjYuLdgWg6cE8N8T
4hOw7w1x2cJCz1H2PbaoJrsMS2j32CpQx0/47MfcKMchc7JDvsHoCuLv1yvjy7SfkfBH344TPYWc
zZU/jNIr0vvcdXyUueDfJsSN/O9mEFCnEld4fgci71cZAibaZIlvc8Zh0CfOlvLV/rFzC3aaVl28
Om8cKyTG9qVO5GV2BmrIV2Ika/XEnJP7F0BtpxDcaLZTKwTGlvUEqBeJgkzpcou4dDyo50zYUPx/
/sN9PMmwgf9xkBORUPQX9kq8loSga4oZdnqxC5TkAKHUBEbJruibRZUnOCyHjiT09ZgozdJm9axR
NvPkPhf7Zb5SaCYH8GSX8k4hV2uNmoWfNn7jj4yZRKRtrDfQoQhGDFNiN5KtQQHSxiqK8gBwjDWM
01osfFUHy9lQchPU/DzB3xJqNZCmIZiRpc5+d0aRZUsS7an30B5viFv6d/xc7aNFjbzE6sd7y3MR
d3b7F7Wi9CG6x/rUrkU0OIOZhCmjrVthleV+SOkih3pVJfWUTbBTdgetr/huc50ENFW1IVIr418v
CNeW04iT65HldNOwtIS/Tx/8hCqhyn5QbTYZcMvuu4mV+aoo8uHdPdatpit4AmmDkYnX8hE2F6tD
CYUMqOQAq5mP4VWq+krvzoEpp4k4wcYM6woj9jqm/YV0rdE8R2hs3hY2AEYkn2PZ+/0in4upud9X
ChN6yrHUINl3IphNy+y1c0bkRH/zvTtadzQMzXN+TSv180eNsN/ujuSOBNU8r+8OXo6J+D5XIRGy
uF2X7Z5ExvGeW0PruILA/705Mip4a3wSV37SL0V6iA/82Gs8yXEIALXSQhBangVLVhq4JyGgJkdf
zF2SfDtIIgt0HJhAulx1qkHLsK1tARQrdRpgu9+voMnAyiBfJbyF8CffbMevUMDDpsFKAwfOojqE
/qIesnyfsfJoyiVToNxosvW1i1ftHwTavmmByAsPnMIrU6beNT6v3Si2aVFf6GZVZo98m7aMvdOf
DooMYaU4y3opA+ZtvdnML4b1apBvlGT5OfFwjGwXdV55e83ovCNAi2PPs6qzoPJK0UMdvB4HdQxj
wC8p4Fpl1h511cO+x9KRf/S+Jcipr0VCdhhEXa0VBwkAi2CCXzEILaTV9eGdWOVJw8IsO+47ob51
JMWdeonfTmP0uwDUBJe3qolhtKRyC1xWQKEKGqVli4Iud9TamJa3PtpoOWBaNeZCC0wjYIBDPr9D
6kyDXSBQ4WDJ+caFRR/U1zW+5uEsV2cpZFNJDTKudJ+qIyQcIfFk9TShgpEsNftKIx4k1dMaf3jZ
BbO/h8v6iA1nKMCgIdI4gfbH3p7d6yZYU57msMJH11qZ0b307NYNWov3wujtJIfTTcPzppujseWq
WLkWX2EJHH8WsNDNDQKZsO2kTs+GO6opN7zJwYxVPVawTYDXe0oh995aD9O3J3k+hTBtHSJukpzq
CwyZupi2xyhuZreEXNMrem7LrltC2Ka+5yMp/AKgP0IS1bfcyQylto7yPT4q4gAuwn2Be+8dBs/N
51Po/+cYIZxlL41ssm2kOcQy94rFApXRGFIa/yk7EBtC2F1xnidBdEBOYg2IlMLPymmsIAolb7zI
T8qGhjqo3gItnf1IJoy0BtskjPG9RTjQYItTfxa2xCUWIWpaivygKFBdi5XaJkAno5Je0ooQeaSe
W+D3+ZLdpETpbR5ukXCVSW4N5T2W4EfTDji1pfhO+7+BTkgYsg9JXmWAkT+Yc0YFT51m+8MxocNJ
MnSvMK22GdelIAwHhHEBszqXa1rQfjciVKwq1gALFz5KCGARge5ORJO4rZfkwT4geZH5KKdeIDmq
E1Z0VkHucNCpYuf4NBmhylqwuCtHd6hlHQpQ4Qd9p2+zr9qqIlibaugq4Avb4Uz8YoKiyoCRLmY4
nCg4e1QNYE0C4qfqmjP6EO38SSS3AVeX5KyvDf7CMbTbJQ1jTi0tz9vDl7wWcpXZsrssh54RJLFr
5sKPjSlm2QcBQTokgy9EcgOJozfJSRe6VXv78EvP6uQG6XuYLGXtBO3Y3VmgbeZbLHG9Mve9LSzt
YO5J8tIpeFhYb3rnQNIE0+eHgyib68vkSkxGnnQqsq0E/xNc3QVlL6Liurn6jXCtJOtjireOe8ps
jZ9VaSz8HevRkZI8hDgPFAoqx8jSamd210oDIdXbyuo/lYpiPG0lgPVzviibdmPocrvUYqLnhyQw
S8cdSYXpVA8ml35QZZkF2fcEmWCAggJ3xikIik07AINPQcXBlbHtKzV6L2l2q5bBWzpZaYdqJZxD
dpW9U4K+if6DcQ7VW93ocqylPG7RmB/UZPsU47vHw75GyM0Ba13dc8xEQkvTu3P9d8ac3FtyRH2T
FEApjVBPLUglZ/4bfv+vk508uXm59vFAWaprtr5yrAYQQA2ZVIax9QGUSOSgFFwc6Bha5Srt2Aby
rTzd/lHj5pIsj//URi9RRf1gve38GA3q3EEd2viccuiVg5zNNFSksgbaEbUtfswfvFVAP5iE7IDx
UtzE7CdMDt83dVaUivWbgJMHY7eqsaC9qmqBMmYqfN9h3g65v0fwjHBc2BN3NymceQ2F0UmxMks5
kKewDJ5fLCWsbVhedy1JozxU8PVepFJziN+MGqdu2/UEol8lT4imvlIMzObsTUEhovL6aFIbjE49
4z4atIPtq4nmNm+FJIrH1LleZE2Y9cl0sRhwUhnluFDWvbFogIUlStcdj7v0uHlOmOBx6Wt6VJ5I
swFATjcXgOjO321TKwQ7cxSpjz4xrCq0RrzdJ5bAhchQm9DEnMwpdkLEPTHVC/z+vajx8BClaNGA
m597MhPknuf32oT+a6gcJUOr0RE3nqEEptBMB9Ei3Dsbn49EZGthSw7mCs2LoRVyxtiiPdoIQHtg
JSN0DSYS6UZAYSh4++gHlZytS3GLKEm+j22jMMwPMKoA//LCOYGoyKpFGOXMVjSwGbFRntyhYnf2
eOl2TwHWDfdLrH2TbQRi7ancWOcrWwkl5qI4UoqT+kVZXSCCoMk7UA1uQeNldGdbouQv2k64ji51
o88ZyDU8gJFD2cPi6OkBDwLzYF8f+iE7lYTDnW8/BY8b66R+CtaNecBHZoODvw7Opoizcss8vtCl
df7fBgxf9WuH4E8IQ20wQRl6BRqECpJX8xZqUBVWffFDesPiUITRkkZluSVpGVhxWvfqu7/gTdcc
Ne3Kf7D05+8VzInTbr2TZzLEyiICXXCpjVEAUZIwouTQ/3vFUqAvUZkutjaGhYUERlhx7KndLgX3
MYzHq7LiysLl0BN1GqyMYJ1Tu4dsCfs4tcB1LtEV/BPWmvoUU1PaDaywSZnPS8jzMFZpLbscXHWa
ssh6fdZNhSrLKXrE16E7cDkb/96bUK14fwjWnJ/nab7F9YTcVpsQEQHSx80+gX/VNQp0K7IrLkZP
oJgCWU0bKFPIKKkxMzkY0hjiyzOtW+cRdYba2r4qaC18r57nWZdnUeJvTQS64dZfqDhqmbczwVaE
1xz3FlHH9DdR+COkM6NnpTZ+DhWnP7eyadEi3vGpNorZ1bROJDxN7dz0S7dbqwuJCWg0oj9xs/mb
7lUCw/SHF1osrfeZWQ323szCmIgcoT8LMCGX7arf2sovc2+Vxfd6v70VwOXSDMZZ+/zb42ru72xK
uXkFKPMJ79DcmT4GCnR/tTxJzqDjOHVqrqu5R8BEfdQGPE3dFeO/rRixwciN++MYJV/WFXjcPfrL
dQA3OJk5JHNX9MqnbjJfAvIjUmKIPcbtc+H5NHZSpU8aAluLPRnCBWA74wA4nMnMhvR9XfeWlCaz
IWiKJDGnjflb4ytGNtwrDhEXl+Wg95RWSdqPk/stWNQIaGM5Vc/Mqym1sT7zpzFPcnwk+WfbzTft
EpOFa7HlBij/W/AtQRMSlIte5PtjjyXOm+lOR99fouIhMTwA5Qff5C3Uyj3qLfb2f1Xg6rtUz+Ix
1B1lbpmx+zJwzBjmZdi0it3NUVqI/nTowWyzD7v8Un8SU7Mv34kiSw9483VtlJ8c+A9e8zPGiVn8
NuHB1g95kC85+sQJQu/wx5CnPgnFzsQmXzH8bAOTIiPHPqqQGESBdkeUZCJDnxBBX2Se4bxNHvLD
U20yklwbTRK+U3DRB0Mo38qJ/0vi8GsfLf1o8rztAdArbfMnndYqj+/GfWltokUaUQvI7puKpmEB
0MSSKiJLuVQKAwBIEDAQsYlPNWbTDWRIDiwLej0Irmo6yGRTHARf8tzLEVPDkuFzVam8byKwpOsR
OBW+Iu+qNX0hEV+F0TknjkffgltGmMIsGdhBg9ARGjiT7RZrAuas7ie9LPhjZobhzG4orLo4SMLk
00iXa0TTOKeZFRHxXnRdhEybRAvarUx3nBrMIXl9ABQwEio5UJM5lLwBJim6qmqJ38yxBQm2sAEi
u1UbUqEodIpTr2CfTNRo4/Y9IEXY95/Wm/J11v52acLw7ddWEj9pFkMr65GIy5edWj9tPEI12k/k
XHGFzEGVZnWbvxebaLqpzuoDTFn038hz6a4pnXx0U0bhvoogyAeO7OUpyJNkm3AQCmq9RRq6BJbZ
y2SI8KlCyIB0uL9o+3AeD0H2NpLk4PyAFLe5h4el8sYk9TbgSQe2H+J2Z7a7Glbr7z48CepaXR85
8As8k2wN0dfUwGnxgAR3zscPGYCGQKMh578LQTCuhIBjvSpS8N/RLuz7iB03K5y54SXsZHKXxEXX
oi9gT+DWfWVEwkNonW+tuVtWbxYnMS2E1N1/plu0fqduY4TZWv7qr6Zwx1q+Gjd9Bs8xR23azEJo
GZj0TZyqum0QUKaA2LTPUtkiiRODfbWyhiVsUTIFxi/jwvO5oeamFF7ABk9eOv3GlAUNwnZ3pyi2
D1Dbz9Crtle3cv5iLgeNModedNDJkpWgMypdsw0OTHs0bNImTYS463xuYGJOVyr1TpK6cxIcB/fq
ztsLKzhWep48CFLgOYGsl+419fy1VJnIWeJ1MPuZdMNNs76aaai1+YwwfJqDbrB1LfUsJZrvpmdC
Daeaa6qtKUZv7hBQc69H2vKKhrjeN9AusrPUAlQ2I3zhrD4hIadhH3TLaHskaFVLt4Oz9YTq0SVz
Nz08qdt7krbYqW6wKOLVszTdd2kJRS9Fq8W6ZxFsDWLppptF9VZL2hc3Psyhex1RuE/Zh/0en20K
SSJUNvAx9THGZoE/iExN89mycZ9U63lZZXshvzm0XFH1yHGiOlLeuu2dgOkkzT1mVhAl3McwnpWT
tC3GXCicz9hX29IruBjBXnnscecJWK2P2ytcyTjDHhGXWYKR4iVaESO/ftAQP4wGkCgki9iXRYb5
nXK6r/uFwW69CjSLf/hhuzO+P4j4esGKLuTecxmocgEF3h4GMzhNgb+aGgkswwcOWANIHGsR6aiQ
TDBdSBZwEOwUyUQ2qxz6Y3tbvqknhDSGCoNf9HVQ6U4+xTXrQ1u+l/KlfcjwCx3pY1blNYp+PkMH
A+JFG0/EwcFKxiJQPywldyIvFW8oKuwdDRj5hssa/BisC6V75tkAO7YcHfMUjKiWNyv6R+pqu285
Z1iANk3/kLvZFxKiMPeMmkqCRqSTIeeaB2w7q03ARhHfsmg4DXCgXFntXKl8RCGle2LEuUfnYBm1
H/I8MwOfyvmJ01ufGMNo9KIj1wtB1H6qXMyu3MEDV0jujzGo7LqvMCuNNfNEfGg2d4YQcGj9W+cw
N+CBsDH6O4qedGXCWS7Kwkoj52oFU2p7sPpF2ivHK1auRNe6+27AexesaG0m1ArIB0HnTFHWbC8O
CyIrnglFYsf8lkh+NLYgXcepi+BZBfKhKW906KN8vFS/8HiskgnB2bUNe5/+XEcVpnMB9HfpvJbz
deEh0ZLH3mlJglwTOfLYwhNRtFbHLsytdxQhWtrnrp5GFpnt9o6RqiYDGsr0R6ZFG8EA5UCHmSKA
9YqGqCBAFVBtB5gOEnBTXx6ueNxs9zyF4P9NBq4sPelK8VrNup1fe+2S8kT1oTmiG8/V93QjQvm/
3eUp3lCiQ1ztNnkncCg+jraSMkCMoq762YA6w/WkPs9mfWZqPtDwdgJhjdeoigRxcC+5iuyGIKG9
/6j4k4EknDRBkfgPhMuYTTkW80f6jKpLgReaTsf7/jX/cRkkeROaa3wQeEtGkflqY/k5p6qZe5OV
wm56tzvz5YBxq36q4jLWgP/yIBdlxa2BBWm4aAiClP7t3HJZkvMcuPzRZNOhxebx4V2ZSzqwReVd
Q6tX4HX36BJVjub/TuH0TthJkyho8zox7nA+1IY+xon/djby8reP3xmsZYIeHdessPzDm8vIxVMa
B0k2iXgAyEdlN5PfMK7mAu6L4yAIQl8R13ckTU6AeedzRe3lIiv9HqcjTH7gWfV7SJLWTt1/ZcRP
ZW4+Sllcdq+b6BzJHyKdrRYugztCeTJSKMLHzZ4n+MdMTGnSE7rFj2RxK/lRLKnH21mCqz8GyKsC
GlmdEfqy5/8yVFrl5RXOT/GFPpsXcheSbNmuINldbo1VH/+05LA/T6cP1C9VySr4ASg4trCXeft4
pbX7KTH35TwhS0s8YP/7hoUmWHzvWRqtUZwE6dx6svMMWT8KxqFVZLnfyFVIrBvmajQyLW4DLmGS
8RWkBDvcBOZWXEMch2gNvCR6ZBjgYwxZ+B/aFwfv+3cxSLMMzJuupZSL2NAzHT32KQ8ujpM9LO1Y
s/PgJcQNKw8sVNix+OaEboayM7X2Bh3AFuOZJmlQLv7t4/bWcYLL73HjIQvVX/QthpPXFZz7P420
K1ctaqC6rkugSIy4+D98dcImLnld24rcoaLInm41kitJkbKErBVIFssoFjGSD7IYbFv9o3oa8cLx
l3ufNX4iNlAGFHJyMbMEOEPq3/FWHxvJ8sdoXi6u2SG79xQoGa3vES75q7sUZaX+hMIBOvi545Bu
tjbvSiqhjBS5lgIOxN5udoAfgVo2hmydsJljY7lodAilLOu4y4bKVarHBoulJerrvSqfUZ+tGy43
Ad8SyOs+e+lupRbYpuaAmBB+t2P7RNr/PCrDzUt9f4FCJ5s5ZT4nJpfVUbtHNeb3KxX31D75gSjl
Hq48CmnhDQXlCXWhvnOzE9p6IE/xlgOyZ+CCwA0xa8Su4RjFg04jOhfDTiplgsX3forvcUcMRtxG
duLdXIc8qaHNPKnAFlyUdZ3GMRHzBnlVpp9vDmniQl9GnpmOtyZi64bQRfLIeOHz5sUqovt4V7aT
uM2D3eLPGl4/Ca3KpfdIvSxNgOVrzY2bWxmMlw65xjH1SnlJrXdsL7s4kZly3u768XfOjF+3E68V
DioGHtJMJH1oRi8g11BmqZEQqEXCVYDnIHVorPBnclgs53a/+cRTxMe2g18+p0r99hurGoyKvNyX
WJZALZ0EAkSIl9V9P1gYHulVHfo6duEwCwLOQM1YXdtsSWkx2PcrKcqw46r03vn+0TeuA+aqOMOq
B+KS+umMI2P736AS77oqzhzbr0nMBTmfUoS9y1ZDAZ+hE6IVQmqYSfKreeledExoBSpApLdmDfiT
UFjZkSCSo6NjmSyXOEgugMUBFuWkOSUIFmyiWycXz0EGGYmaUk3UyCYAUKLSe+U6qW2/e0wj5EBs
PqBFMZM2lIJbmP3gMPYscamXhJ7pozE6uXrXlR+5JBhtHw6mPRSRV9aGA/ik3PhzFQ2gOm29G5dX
q/OPJnynn0mgsBKWH3be1m8a7THlQOXhMsNLm259xlKUgHMml2li9DPPXX54wMmMBzYcvquMy+QO
O6izygRe1cNd+a5FxWaUogc0Go1EZ+zMI1ipAOUCPgJg9QnJdjAwHrw7waU4t3uLL8+VmLVJ9kT3
Ac96a8D1xkhD7vbe19X8fYjfj5SqDpu1mlTvu4Pfv//qYFU7XOweMWryVaAjK4q1Bh4YAUdpJ6yc
PaKRMAX5VYFviqoiWqyYiV6vl9cgCgbmwxO6xkLnlzEVoeJiuRxKiRub3Z/EpJpftahQE3VaiwzG
k9wOe8TMzzLC+nC9ToJIkFPMvZo5/S2GQ67ohvhdLylUMsHYlhIoJB60e27yWa/9lRqccMUX/7O7
NjyT5JOflQl2+n39QHCSv4IHnM7fx+VjbvkobO59DXsRXjVWjeMD7PH8SWsqd352DjC1EmfhkeuV
daVHZ0J9iQNmJvosk+FYANaxy8HvxG9IjAJTCyqzIKki9b+BFMr8lrEak4VNzC/OtGuCsv4wKzyk
9PPh8oXpcDWMDmNuEvypsS87TXvs73GHCv4GFtr7F4nQQTCgLTY0OZjLvEdXkXNSPORGqioaxMvV
3/7i7qE4LHX9Jpbz/6stLVGy+5NenphfvAckFUqLwtYYfwUyxvyv9pHdykCf5aNQS6hEkI5qWq1c
3a/bL7DBeZYgSJMGyUFNBVbkMJ0S7SyTdBxD8/RkRkEj+56u2kq8ar6mU7p6YU0hlCRMDoNOI7od
L493Mn/xxrz4BkxPfEvNDQvl+VgADWmlg6sXsUrWjDPwv9Gw6RjdiE/BRUkXHs0F4Vv6IGyTCLVu
tHECWkz8lt1LKWOoV+A8yxb2fzGvx5asSfQSWinSFTI5lRFxL4MLYxeeyiGQ8D3cqbQ2NNkhL7HT
cwTirRWmk+EY06W0fWYkOjsIketsohK3Fgu9MUpc6ZUs01Fv8ICHBsKleiNHwKCFzqUPSQkxy3GS
xvhYPkrmu/+SvzLuNvxqzlf2QK1lA/c4eEaLkcYzpdkwniKXfXdmEDcYMWDK7PXt0uiQUlDutR2o
EyfMYSkhgwiakI4PFqGt7pETBmI9PzHFafGP5K3P9k4idq2wLa21bstBPDK57PS1/j/z4InddBgP
nCkOrQXHto40JEAFbLJ0m04Zjrs0D9Wq1mMaVE1ICcixRm7nfm5eT8D/KPtT73xB7EBiAmuwQ7Ga
Gmwb/EGeUiTN/sY7RGBGEln5TblPaECbpgEYfIdbGL6vxdwzJhXESZdYaXFdsCCReUkY21ipIb8C
d6XeniwPQsG0nUY0aXF4fRBcDzCzIkiG24dfbJQ+8sptXIAanXf2pZo9R0ItYOLh2oVBQF4wq0UR
8jVRF4Bhghlk6QzS7+2mRG0iPMnBqDVbUnFOQERkXl+syHzhfmfbi/PrbhrhPa/wqqLMKYAnqkYW
4a6bwc1ow3WpmmtM+b9WnGX4Gl89l5oW5z7RSbLgTef+0/kT+uaK3s8lasNyaz+5CseQgz3oKihE
lvd5Wvt9nZUmD5aX0gSMeOCGTVpC2y2RhH7r6f3CHdu5NKCfOcpa/dGZxGgxji7vRBJY80CRvkbF
3m7CXyIRojbLiTAZImsdqgL9wmJPfe/bWRUaRmNPf1vuusBDBD+FrIs5fd54D9ZYqom/KhAlWySE
uNtsrHCPZoUBCpdPB/FfxMjKL/bZBXG+If5KS60f31fRqVnU+IQ0Url93EIXBGHbSYPXsBrsi8s+
sALHGUDkijlhP4Kcr1ULQ8i9CQ/aIZugeBne6zWDjc4uERyN5yIU0RIwQQpFB5EKbqYUrPXuY4vZ
Es3ktjd+h/54zBY3EXuTIcaOZizMu/zA5+tgpw2Hk35Somq6Ou5i1QryLo+ncIKxL0QM9uINabz6
ZNB2g5hwFp+Izuq/cxTWBn/35gJEsd6JQYIvXUTTa2AepYJYuLi15bSTLXp5pTKWVl/Zuo4VSitG
z5S+IJcv1DIfBcBOil2bvUeqI2bGLZV6+5jwdTbrdmhLigz30htKLoyEPrSGRCena+uEIkCf65eZ
wcNcvbU38JTrQ7KvEaoN5gdGthnSZlM5vG2VeGUZyGHLtj4pXTJeavHBuD+bqFEMgNhIyrpoDCjR
iGfZUHTBAMG0xU/7eFkYSJUGxsBxtfy9VMnLJbjG2mXIcZGzkeeOllNki56obZDi4tL45uDMSu5I
kqvHE1LuNaO+Cx7ZOyEdEYSnw0afHyqTWUgwTFhiKoo9Qd+pfWgFZg02osflIJFqNRJ4qmGZS3yG
rx69l1QX1TIwEtBuZoSXtSSTIAJfkRP4k57g1dUulguGTIHFL7edBhI6jq9C+Z7tTSkSk/7OU/am
4ddvowoZzuFD1DcXZhfSbEuMsB/XDG7rQDyBHkZZN8PJVvPo8q7W4kt7r34VGb5Bu+Iqat08Bga+
UCT+PD79cLI+7GFgeCGmThVN8rawA5cVoOxpN6p4xxedJjzJxpHVC9MgikdKknuSZ5RygAAEKoRm
MXDVRePBgWHEZLl1bwVrfwDnlYFJaXVvhf6aYqscKrCV8BRiW8yaHMQ1dRmP/ZkTyL9yLxpbdY31
r5BwVGo3K/nZdoLVw1IelzVYzBdOtwV7xFlwQmaxaDHvAOm9hC/u1tMwmeQrCSUygGlb0/Apj3pX
WmF25nRGqrE+BhadX9gobKCzwDVFiIM3ArCguPfV0e+teDeC7xniOJdr2Sdy3/S6wDkvgbeln0GK
kD0XYDWWscLqV5P0ARCSI4XVjx6MFbJEy4jJVwYCXXrtmGpS5LNSuixTGkFVf9Myn4H+quj65WPK
kKQQkEMmfgNbZKGIriAjvfAVDoBMz+0gqI027bWG7hUXdhLdjkz7U0Zgi4n+1LwUnNodMEVsyCKF
ifb0S9e/NgkSfgrDhtHUqRF+NOqbW20QZFP6C3QyDQcA9I9eHUzETmA/HXHR9op/fxTQtAeZ6gpd
Vij55rwhl5nhUP+ZuCC4PQm1XQUUfmU9C0Ma/C+I5fObNUAKIJu248E7Ed0sQyD1RuSg3wICrUth
enl3B+3mcVP5sAYTg3XxM8LQpz4KKzfp8P24qHPncipCSicGGvaU5jR71Zf7gInhLcN1mylwK1fL
TfIh2YY7TbIdskC7rDMNs+hGwgbyj6fFnx+w7W0YtijLBXUlYZjmTW23eo+/lYJ15hYKe7ydL/P2
+rWo8ZCsgU23I881VbcZR6jKvsYhyOC6i4hk1M+mpz3k0N4m7QPGsH7YuTLIZObIspnSy9y2dutT
nPQir/fU0/jhoptjfBFTB+3wvnOIIcDxn7HrwArBSulw1K2kV02YFvx+lhoNvapc/wVr7NkO60Ps
LslsR3sI57iCzm2F+0bjXlEBgVyyIenCqdD2NSMkNltfLeqeelYV+vy1N5dGAoe8Fkc/s8A/eWnO
VWzg2IXqSsDA8JoO3p/oYCM3EU9b1RHXJt9WYbBUbie7qKGR4ocoXBdWh2IvBCRfUvjLdJqBiTWv
ADHiN+3FqZsbMMaPZLifcbgyzFm9GQdum8fgU+rFFCUrAFFeDnjqwmwdhEcUhnEm5kCci6ta2udr
kBWPy/qZG6sh8eiFXCMv9o0YA6z7dU9nQl8puGNgwb6h1vSFlrERLwLsrq0uIgGOnFMTZbKZ3TyU
CPZwp9N/Mm/uYKAB/EEXw42e23ZT1rR3nV/ELwkxg9+WaRrqoq/OdpoSFhMHOLFm34FRsnRZZ7yl
5107uI6LMpMD7WnorSGl/lTyhqenN+u8IJcEqLuapB55IX7I7oeggjQo5exGfM5VEQ9IjUOq7rqq
yx0KcT0ISltenECBetCZnECuGx6R5i5v68UAFdmOnHr6idvWKHw/U7vmgkLXPPTzYagi5CeqkNMW
yrmCbqsnoJ7yjqQffySixIFrhUyknge48OS3ZFfDr4LfNCXpBckpY7G07Vcrz9Db8yQDU4tR7y3R
sFpnKDQb/X6USFaXE9toYmddLjFsKKXyrviQZNC90vzcZNcOx0n8DkCsX5ypqC2xWn9mhE0Mz/ER
Yj3z+vluPotW+/5KOnKLNustWbPtAuvv8q4UhRVseTsXYvmsA0Va5vEj1+ajTXnzp1noaWui4Whp
JT/mhmH2eHNibx0AIJInmxL4LEr19xjuR19xLyvCy+9bpp/tn5sfLP4LUYqbOHfo23c46MawSR3y
Dxn3+0O/xebY1a7/6tJZBtE676OfB+A34Ihom4JV2xnSOM1d2BIfNdan/M/CDwRBBGPh9sKUwXqm
8X6BY91wDSrxAIEIB1ts/MhZYqf5+t2tqEzNT/xZUrmDIBJuCftdsRpjwzGXpYco8id11ouR/Qlh
L93ASb/fiaBjuOUCbotrUzH0SxN+MZlkXsHltneoWZywJYkNTAJ2Z1RFELNlokZbBRGezYpFePG2
RGAtyMV1GyKv4/wP2SwKuMZdVs+BX0Ge1IeunfFRkLZctPMWa77JX4VtE5jaGr+rnBJsqxpWBSiY
FPs7kBDcLPvAI33xjZ2OGjo3m071hgDgXpSPzUp56h0ROd45jDhKrI1Q+cIt5fyi0DyLVEqB9gbe
DqtWKaFHcFaCOW00W74tl+ZCUA1zwKc3QLL5q45ONnCsOAu9Z0Nfg2cv/O2/Hm72+C+h1jbFHToU
MQiI1cxTcZnx09zkuj9iTmXSCb5JNS+misYtXfb8Hvj/0RWT00kQjZDoogM2xy49nqpq1nrgb4jg
hHI2WHn2NtdILGsL/lHS/EZgkF4UEUG5eeIkrakIjiAaWIKFv7robd03apbfNE4pmBXy06AFLdvJ
7NPKbYmXLH3aZDkn2PyClEDCgm6B/VH//bELmIMHNAr8mkM/cnggYHbnwaYcWuzgEb4s6gPiNQAt
eCWDqjGGB2kPXhwdziVh7elJ/8JdkfEAq3kwzzEbmx7f6yV14mdKuAPWTQZDKfhNA0aNakR6xgE6
K6aczT+a0vfRN9bObTaUHEtVs9vxV4Y/G0mT3AceYenUpIIZguFtkngHwB83UI7/avUc63Qc3xSQ
Fj3TKPg5YrUUT3Hk4y7dXh06LzOBbRsmxg10lmR232DlZIj8stYWSlksWaL4Lr28hZhYIYc6eNss
hmB/pRP+xVEHnRcgw4eW9GMMpxPwx8Kx6jXMjDIH4qPksZvAxEM1+2ysWv/4me1dwnhWkRuJH1iT
wWDe0GsOGIsEDUpQYeM63jwFSmmcFxexAPmbDVls/lS6OpqjdqhEt+EJnWfse7O0A/4z8ZvPablw
ItL2iWSf/oNpns6RrCgjQGe3Cc4TExIdPrQWCUSPTywi58DIa2JFBaHcp2KSKnt0nsz3gm2G1WKf
uojrHEOdRQKDMWESLx7pRBUS5H6XhaO9SOCATH26qkMLmyO51o/7ShsRqp+tD/6QU1oIq2g0HpiE
GOlAOuoFHqzosa4x7k9ag1ZCgrHMQBGrLgl5cqAmKARlu0b6NlQ4EN9vQ7AzKn42VrRGvMPkDeSC
LG6zTiK9qz6K6BI989rNEzLvG1lZo0zZTHQ9yFpuCx7CaxmzvLzo+bM9rrpwkgS7cVsWDJr1ezfH
kdV35UK0S39qLI7BKgZKGQ4i4bAFVjlZ8uPlNmOOoiZchNMzmRA9OORgCyMQ8iMFW46CIyz2XbHV
NGqqBUPN1XjQd8qMKbKx38dCDDCJixFjPd7BwqlmzR4iIGG9AQywabE15+ABG1qwtmCJNa9km4O3
fAZFzu+XfMyV9lqJp4/yK4Gp9rJPAdwl7qgZvmskOH+3mtaXN3asrodKuTO8UTw3qDBk1qgWun6U
NpHHNed4awjz0ddquffvchKW8hjRvnWCIufm3L07njg67uvTQb0I8vIzjsG7tBABvBtmz5oaj4XG
hfi6o5u2PJgDx9Psj/258cxbVuvZuHNr3ulRmeVKA83PNn6fluSqrywZFjIwSGIxv7E7jrQxYbe6
h+lWm1xfQI+7THJn7SeLbKTPbz7vwU3ArMYYZB8qR2lDm3ySGSjUy51b7KclnvgPiE/NKsNzmsCQ
K2vvotYKyToaYyAwoCaUqtcWrtHNoEkCydKo+xTLOtrkvY0OobbJ7TuQfSQCyBpROcyTcy7o4U5n
5vQ4sfizhoAEEqssRkGKLKIHtALJZs9zp1E4M2g0sUixcQpj+xcpit4Ca3pvVoGrK1S5xj+cwNTf
jnbOvpinxZqEW9mk6mf7mMVNS0R6vA0LjLp7IJlN/1/tQR6uUbq5FPhw96hIEy65nMlUNvwsinli
ZEO6t8TNAxm8YUA4lbAgtGkGmy4ZeqRzUMH882CC4vhQY3XIhFctYQii6uXqqquUouWoWoqC6UL9
bkncce45XODZIY9HICql2QBdC2a+ytYr/vabgBrlRD9QGfBibFDrVaJWXV30g/lGnqLoJue5B4DI
RCDG1x/lQDIG55qAJfJY789/DeuiUcyE04BLTPRGl0N7cD+gorf/4yy4jntJhILm4GY+owNwaIQ6
8yGT4rbiTbnnkuT6Y/rJPdGjydZRVgZA1yVlHEE8IAbIctr9sCf4Dft7yeE35Vk8FoELnhnPPoH/
l7T0KIo/rBE1b0kBnIYlPukoO0j7o2ZjQtHHoCltycJhUgId6vCRfysUA9PYfqYGnQzL3hfki0Lh
OnjKIjr/cHCcgmhVQA58IYYOjoQdx3NSSm8GwQ/TPVszerDC3/npaOF+wsfQXZ6uxOB0xk9bBpKL
kp9K/3OpOItEDEBiOG+3cy5D6Y/dYviBp6GsNYZNLdVSFnMgR+2JJFn2Epe37ScD6SgrIN2vW+Iu
ju9QzjxnZVefqjCiqXkXDaaZ0dPU3xAfL3iVJ/l54XXdISIHcLNsRazxzAweVv12CiTDAguJ0iTM
ijMMy6SW1WnVeZtEHkwRdzBZkX0plEzm2kuPuoB+B5Lj45psBkAmqZ63tRdqUyOWR2lX9Y2Yw24I
9U+QEnuJuQCDdkDkN7jhnxZXozrUhlqtD+h1IqY44GJcXWTBAowS32fc5hQcSnfWEk/tb31ZKwaO
lGUk2pEAGN1k0lDGsTp3MX0R/vwjwK71vVSGuTv2SVK/xsk8HHNfXPfZQlPIVB3oKudPFne4+cIC
rrYUH5lMCmi80vT6NQVpTPZzDdht8KsvT2XjaAwRY60uaqWC6lccsUXimh37c5ShKKcm3YUuoNxe
eVXWM2AfYKNTO6CVX3j8nZNZD9VQxHthJo1dQiHaxXlK2tf3FY41ow9+z3HQ56N2nWt5wC/sKNoq
ipx5GKFYQZrhuISRXI44etb8hSWokH8/ubqGxvN5v8oZWvIO5qzsoCT364QDM4XFFazOV/XHMm3I
Kn7iIhGTdqx4OAWVmhH4Nj++dN7UZDw1IdGLeLuvgV7H6SG4fzjoUy7jK+Vnn9oBnMdgKz4XHM8U
Lotx3egKfDDQgCsGlSiO6Xtvp97HiIUddnUvr96grJcOuQ5NyNI63Mx8ad4BiTK/dWLr/HYWD2Y2
8OXBCKmNRJWb1/YcDq99jy4hs4W9oDWEGrAquk5AmABJ11+Ku4EleD+S1CEZi4arzEfXpdiMANrH
tWOcXNYaRxIE/bUmxITzJbfUb/vLcRhViDFZwBplZCCaIxt5LrP9X7JugASvmTH4VMTIZ3lGjT3h
tAJ6rwqL+vPmvN4aR0Zui9UW4P2OaOp+1gf/i/PLiwvblln74kBohdiV23iT1K0X1Rnik1aQo804
hgVK4yBVZcq3C0s5cm87TpqBRmVz5m4AJqz44t8mksoDpaNtrKSsYDwyEdypZ/+CARhhmlKP5c0u
ACdUcU90LpL6rHov7iPrMSraQUnYt2BpTzizsdPIYtNX/d2drzE51qbo6yK2mOe8uzbFbnvTeXRs
cPthpgFnvSuisoY6QadY4TlN8ei+0uA4To2pj6JKiGLEJ50f/qc3SDPYV9oZoXoKpMFdoKOXkUI0
KXohpuGtn9xhe8SSCIdfU42pZWvJNIv+gp2i149KwRdGtSSjKt5sT9kR3z58imCpqXlGJ30ekgTP
qsEywzldsz7FNO5i0hDIkjBzY414DRwWmlWBrEZKpQPGnnjhhSFjMS8PxCUdMx5/HjxY2LvOVtx1
2Zeva1e4HuqcE02eJbZuOsz9+yXfKkF0hPkXYSkCMEAy+EwryeaSmosZhotjmsb9i0PRaQ+nAF7K
VENX099iCI1vEgv6VpdoW69XHiwqMbjsmD/35/DHyhmHMibpFVxtzojiCkBxFOgy5I1xrmP+ZR/g
edobtKJekPpV/K8XxqYJ/HnY0OmlvaLiOQM2Y10ZoF7QCVplCoXbOuii2/zAz7y74VLTcFh6nCZn
/JLKNUIKPN4QmWq8rQB6Jg6uianK/1WNaOusm0gbgCCDum4i/d6WTIZ8ddGkPeP+Tine6oD4tpEB
CsE4wCKXK3gOlPF2L4UkKCNGApeRKl9ORg1e5k5Y20GKjDKq0DNV27DRwsfZMNYlMGpoxZelviGy
uMjFqKgMrIW+uvcexRUT4Nn8MxmUoSh7jAy4yBDnAHAe11of6bi8edLaBR9LGgul+hR1EEs+JPfp
+rUrREqWk88TR/BPTex0xgrVVlOrWL+mR9XG4OoZL93QypX7HeibRUlDejD4gg3So874zWMf4TiA
yNS/wBnLrZ+83VxiIug5Zuv+6tBszrRJBlrnV2q8MknVtx8QpTEKhH1ZXy/M+9rBAA7xWVYmWQlL
ipe6PhMWq5f/D6miQb+adTh7m0tkQqt91BqgGY1duihwzShcLhq2GHNXrj2Grm4ElUzc/yzIlhko
dEkvEdPdw1A1V+AlqnVW3a8U7avUIjYNY5OYtQ31ctkJwfDAvPpIo2ZCPtT36srVEaBt/hW9VNu1
c7O8Iey0NcuVWUZcxY/i3RuV0rJqDyoe4gjqLWCHY1BoGcU8+MZdgMlbtbQWsYGgsmzehT3e250D
dGMAfU2eKxQ3c97ePZwBRsP2zVvwQzJ/37s2lFmRB8pI8FYnODgh3AP/WWD1ZB1ewIMEXtwL3BY2
DIOb4AO43LuVnEeAiuljL2mJFHW9w1GoE7Mdsch0hdH86Z4y8Q4Qag/c8z2AuClW0mi1wCd89SyC
Ij53NfqceaqPA/7nXGwJe2lmOIeQusxJe4gaOmf+zGzyw+93YDHtfkZnc+icpTuwoCch8r669K3h
j8vshYdPFEQjuL/oYs9P8yRPhoi5v1HP2X7kxk/r4nBjgwQ8e4IPMfYsnX0VH9oN76dFlHipQvCY
qkQHY7ZVrkC59KrcRhr1sMnmMpGpH38DWt7/Du6qPvQXQw0hED/R9ByA+HWmQnIiB3OXoB69eRls
pNNF8BdhRD8usSqGY6h51egS54H9N2DECaVHNC6wEDr8OYSE2XF0mERkNouKv8eISvlvNkRuk2k9
skqlFSspL1Cm6aR330skbqECYU8P3W2uc2Q7ydn+J0UnhH9BTcGNSkh8KZ8Z+IFdIWrcc/PcYx1L
5WHH3eu3UAiLjQnIvZxHJnWR5MivDffDALM3z0Fz45HDSXdekMzJCr2M5kqaVU+uXGr6agxQtgXg
efGZPYl9uASZYMTi8wL/H1H92Z8cQBPrsrHtoXoacMH4Csk63Q+JQJz5Zh5/rNVONL0ATYmzdfB0
rJp+orsanK5OVuew637Z42/TrypHp7iLqSkw+ZwUcgf2bbvaCJbA1jq8Dz1xYSP2FI8fRvRVk+cX
arRham4197VHeRCRaxXYjuXvbt9VWfxR47tOqY/NLDuq+Ig9zK2XBjfTfY42F8YPUv2fTDfakZMj
GYk8H0ku/H+qF1z2EaAI8l4DxjsZOfrNUHarCkGlgLFgDpNnkjdbLbCb+nUlCfNJ7weVMcIpEDdB
nDeX/hGsbU9Re3FbTd3cR38PeuWpWChqmrfr9lP+qgb1EgS1V/hkkohTRbkSV+0H63dvuTGK93zg
BFhZhLZMcwpjwOUUDb+YTyUOgOsMPG/Ha1hEIm/Mi3dnOPSEUnabPoBVzTiC83QzRnpyRkurxv41
CNUZoJ8m0IbDsyN54W3Z2BGz8Y7zVhyBxFfjWm59T87uPJVgJjZOw9kTI2R9NkjkhqhQewFxG8lT
Yn5SDRvmASsttEoty+oQdOKFiw4MH0r+bd9/zLbcSxX/7Zlre8s8ccjFzsLLWINO1VV7p2zFWUZ+
NOnZBxD/fOJekSVLMp+yfrXhvqfCdFQQsgdapiisTD35WVL5eGXy4yWg4oFlUJrqzGBTJqRi1vdD
u5LroJzRMmEUDAViV+14b4MlznEftZwqEowfYG01Ni0ZNjiHwMD9DxWUheDVHFBlAU1+cJnfddAk
O7WnHqg3Ji76qhHLZCPUbUlW60az9i24a4lppbDyGDCovIkD0cVJsOgah0eD0JzpSulkgv7F/cL1
e22VKYtnZ/8RmF4sxaMS+Glz1xQvhBCgS5EWNJTEqjXZoQvxIHlfcJs8iRULP/lk2CT+iEY8AKgu
i51l6GoYHjKWPzG9TJc/WZKIbfFKvvbOqFX50BGt7/KePhxhCi8E+7MgO3iFa+vj571wMeIMQLIF
FRXaQ0ott1fpgAvihYB4RwuJ2wyDGBYL1wJV/JFc5gPs7HvycSV9skn4tRCNvkE5+zEfJHMXWNON
itXXx+Ei1/EpsNBfmmgnPjbQl5QPAMcuXT7JzeZUdIzqdMGRxfds2qjEKyB7s/LS5jiuB1epP3as
FQOSHbwrSk1mgEkgMGVHnd+DKm0Q0jbPTAKv9XgYhE2M3uHwHz/xCA96I4Ft+TEJky5nKlbX3rc5
Uhf9UOAp/UUApnQYaB7WKkCr5qjs0AKcEF/kRyrfN+prZjZQIu/Rw+DXL+PRRVL+xRRxu2IxgHXw
/PELF998Gk8ZMEiSv5LFSh0iXaFypyCI/yYoBzBMzyhdOoidemwJZyOOZSIX3jFCP9OCcvyo1Cf6
Lx+ouV81UyrPuZHuRZueB2cZTIQbfgM51ZdFGcyp6KGuJ9Y2kiZ9cNtpzhOfGYkIBulgfoMtW9yK
FywBCWX7inmFTj8YZNLzgeVwNDvpngV9pNwiBQd2XNfyjs2+wAvm9VrHjb67eAUCyQ/UKX+JTgVY
rdkWo1S90i28LFMpGUn/zUN7XzNApxU5YwZrPkBs0Vy+nV78V6hKVt4YSrnX0/vplkuM3hJlxt/M
ZeJTru+RdRIPAWIce8bQw3J9O8+hp5RDsWTsJh/XhR4IQY++7uBGsh+qmEDrNix2twNSsVlHkcLh
zyvsghV+H1a2XJcBKW8Art9VBuYjAJIsTKvUUF4LdVKZtQkqU6jNZ2Hz01MvuVMX4VyOjoAHZvGO
XE7pNx/m6kxPbQ5wQLKBiVcpaO3V0iHE1IwSUgaLDdvNp7Ecw/OY9EzO6nhp+f3seQ9hXJHpoqfh
GYe2klkfySu63lAqy3eyC/tSCSwDRQ5GiI1ZHh9Y3ZKjB34Yp6Tn5WvttICQPx0kU8aaa6zfwy0K
0AQ+rU6EdjGhK3vgLt3bP0ObkJfdx4NYfjD6WSQkqcT5mzSZDX9pXWGEsG5esxxItN/8XbCP/a8d
E2+JVE+8t26IkKHENCG9uy1AkGuqgbR1hj5bpHNM5sd/UZ5irSoytod7wPIrP3UUHdkCxJdLbxoQ
G5/yp8T7LH+Xu2kvIiWf4YqkL00jmtFZOd5vb87ox5JGt8FkRiQjtDWREWoSG2ezhncYxRdDQvfG
xWB7qkOPOwHqXNW4PbcMPqFd7gmVLsIFWc4hZG9g64MwM2Br5FeAt5u0PrnPP9W8OD05PGg0K7eY
m446zkX4B39UTopYSajt1tWFQakQ7IIG6IrYqcsbbNY/NrmsB6rIoEWIinM3BtD0zO2UVJnbgSbu
crTgb1kIfb3TYRR5nFWcZpp9Li8M6IGCiqvwSl4sfeno1gleLcM/INQEwBoQbUfRchgNJIeoP4wP
4KYJLcka4mCM+pPszXHWzaBi/MwAjvMDCVNQK/UrhQcQGz6GSRYw7tyQas8c3LpciTS6Uxt5Vq2q
5SZq/jB/jn1VZ0ct3lze+vKXTFSpdINDX2Qi7V0K9OLc4gJiRIFS4xa9/NfyfAp/dJQB7IOCsgio
jZ3curIz8dwjveVbPO2ZQKrEo3dk9PAFvqiHq3Bh+Z5Sf8zT6rXu9j1qg7MmmBWye07d0HjIVj3/
yoNBOVy7Xy8PHuyS2uHvKxC7YAdEud3ZiUZv40xAyRC8vPiz49E/tPqy01PG+wiG/qTwH3Do8qEP
bMtqIcSzyQJbG0zoVUCCNcdZK6g1PCjSViyk7txncSlY+LhTzRuls/KI5NWBDLtJnO0rNG9cr/rx
UsEHSk+YqvGGv5rL6QWg199r9wiy+eqo+gxeHpSWG+FaZCvnvfKNm3EF7MA1b4Cc9/BwP5JI7P5t
DT/5jjYnQwoJ3U6oYI+MzPZZMXl5Uv/al6WbgGasn5aZG/N9NXg8fTKS43MVGRmTFvX3WvtTqgkx
QSEbIrA4PCEWxvSdFDdxZ3NTyUkTd1f/OZRwONe+azWW8WBKrRpchDq4vr3r0nKW95vwjh5S0DBk
kDw2bvjENY1a30IVZmoqpQEW80Xga2OfZ/5NAxgswsCUFz4PKnTZAsPRoyCgTX/wRkb8JtoOCNfB
6nVupMbXsoN7Z482xHLIt1NP1NCVoaZECAKdguUB9KUSrFhUS5PCrAShkP7xaaAaU7UaN6aoQXeF
7dqdJx6YlBXCVTc05d08OULUkI/AMF7WDXZrFrA8GWwijzg0394dGtIfoErdizD/hALwYt5H4Wpx
JGLHEpjN8TPa9YImdcoyMv9IRUeo/3VHUxc2fo0bUK0qkxaqGg1LKW3gqcG3QFK0UkSgQtW3IImv
MntRjUfNbyZmsA5tQnFuDSgBhS59SLN1QBqI9n7N8HX26YS+6Dq6K4w+vR5VIVUXxNqThighopCe
P7zdgOc4ELcXoMCg10XOowrS04k+Alubg5k1mpgHMd7k78zOT73TYsNA6nsmGd6Vo584NaJmoC0q
znYPuwSWpNhs+Em2GfCT3j+Um22LwESCqoXC7WA7kkXz29a1Sng4ofo4k4cU/+Wqa16gQQ9m47wU
fMzDXw4kv1R5j+TPzyBg2el0ksp8X0GLVbmjWSTOZRe8EP6G05e7cJ5Jdg8gfrQYJ81kyEQiW5Zc
LiuDjzbOxrsqCzwO0dbalSAX+TJlLnpQPxMVLbrwkWNmJPanFds63qQ762KxiO8OX6X0Uj5mIWRf
jw3p2Ag1PLCnsqTq3Iy6JW0qs7u7OiAEYyh46X4oabRd+huETGna7KoUuE2pL7S/r9hX4VCeypCL
Vl9+0QG3/dU4zwK2XXdmHnxgoKMvXt/whhsJezwMKB6rxf/acIbKfPHazAP89I1IA1rmlKEq3fMO
UuEq9OQHX6fP5wwSWuxtGuELOsJdiBXZEjZpUzs/UXF7XwuPGL+HB6sPOn+ixKvvPJTYmuZ62nii
R4YICYyb2V6LwAArMVBqQz8wu/pv3VD4eZmB2UxXdVKjWfyru3/lw/2tp6fAthUd99S6icl5CR78
dxrdyFoB7qC+9Z4ATA2ZFauA9B1SHgLbthMreiNDkM00Wi7H93x3GZDVbGwJm3Y98aqT+zCz6Urq
sYs9q3Au06Ehp1OXXa7YOggoUBuZxkIEDuGz1eBFxi/FXZkwq0ZwZ6+AaRyqT0cnSRPjrScZn/42
Kz4+TvWHPy+hU4/D5GgLJI6vX84KUJ7AMosTDwBB2ewwHCyQg3vRTCr+UGqzjMmiBTqnxbZnp8ti
1ZNtlKgLMvV8XFxbnYdIo53P+JASLAeIxzNr1Su3zvBkHvZLDDIl8AwFmyPsP8KZku/OxrGmS7tf
DzlPzmxmcG1T7Ao+vGfkZ8Yay01anfwiYxbvQZ9LgGRt6Adfx7wbmRnAQg9TJ+k9nNpPs+dN3Hec
YMl4PWieP4ok8x9Y1sFlULJFPeZrwmwFRjqzl9v456nPV3FWGsNovKhso5FoENfANAGgPutZvtZk
GqYSs24cTd6418uQakQ+9PQzhGlOleXq8tabd73ht475ZX7dw3Bd0euBhaFlBCvU11dpUzODotQk
WhgEUA7P+RWKXi08u9wahS4ZCM+ia7JSwL9Qf88xFq7aDvFtBH9YVwP1lroT8Thh6jHUtkZiwboe
kCl7rtaMNll9i3DsU9mhR+IXc47Z39BdksW5T9H7kDwECtV71AE+EJlTFod/67R29s5JyvX07viB
1KyZsMQGk1A/cWaJiS6V4yHbiMd0CjGI0vTvVeWi2WzGG2gQ7oQDEaAiPSMNiewd37FM2cgzaNSn
hKovF0mp+zWhLEe+IuOP/KwpZDPk/7YjGm0NbsaNGLEOepy2QVPfXNyDlC+rzU0buVc7viqpKtYF
Xa18ZcTnE5nBDQzStKrrTedJVPQcjJc0B1/B30Yt7pw1FHsQdXQdgv9k62X13NqMK3t3hhrP8WJu
L8USOIW688ROHozbkFJfAdoIqWsPeVYqWBUbEFtaLYO5+uQXE9EH+maqM8bxels4Y7j0/FsgasLI
QfStC5riWy2a5EPIQUrtjxveYxRp0dCJ6VyO8Uj45ispJrTnzDtvcp2+bNKnSP7FpOTFAvXtj1Mx
V+DCght925coPTIgny0EWRs0G1AT4xHyyvojmKMREc4jcCzQXYWykJKfvPBlyUUkLUWfAQaeza/0
qxy6ZLlcERYHKl5FP96dgJdFxDQ7ymLiBsG6NsYclTwRF8O6x8Yx4Ju9w7KihbY8/u12AA5cVHds
QbQ35SJYO2CBAODtlJQoJPfo2a9iaxBbU6OJrOrFosNuK00oJIgnTyWgUAhVcRopiNoqiqwFIK0z
06vchth9UvwebtaNDc/zTxvIV/vvAGRzbOYuYvR8LWTMywalMKmdtGGgbxNDlU0x9OMJTxLmGDbk
ZsaWgNSkVnPEZAdoaXJ0NNnppNwOe7Di11C0YWUWQ8JhO43TyKOW+vPslBXk8uQGI3KGH40mALN9
A5tkgpoIzG4+esUOOZk5jWWu/ADwSD1uYBfm0hIp9Cax2CraEk1V/3v1Y+q1DRxkQepIoCkmweJs
682A2xHJBIe6cI4yWCr155HIsnP/HhXWAmDZ6mVEIXeyJioYmZqroNThqVpoOplA1O+XbzkYye3I
2lQUrbq8drjzBKAyq/iC7uq2SylrptDa+5U3DQxmSXz/lMG8yf65gcIJTqhi047yebSD5R2AFimM
cDcLTrOtyEdV4mtMzQPWKVsdoMVWOpCdZO8Y+nCAFJQkHhZ/PiPdO6Adk/kUbWpOcm12OH75gYBS
ZQo9MUn4tjaZ/OvnHY8bjRLmU934NoX9S+seGweoJC7/xaULJmf8J6yIBT50CoDR48SCFOmDioA+
SFfaQxgix7YpL3EmAC3tOD7A4OdsFioqz/COQnSxqAgvZj5ZBXDEXNeiBQqeCQjp6+s/r7qNmp6D
Mh0nBADZ/yHPfGj6DsGVsX1+/UlSkq/cyGTVKN0nWaNB0nW+2eJ9ww5BU0wSWAaPv+hR/MRqK/aI
mfzdDV0m/Vrty94sgwhHPFZZJSOBXlHGVfhX0crlenSdQ+lImRQLvnR9EHBAUWCQFtZLJHkh5Tb3
V651yV/YOsWhreI+i52tSQ30Mlz/+frXHhVwdZGUOFwEGZTIE9smyeCIudKUp6KsqxhVDQYi6agb
KQvfkC5TLFTbSqnAs7UPSvZPJek6Ulo7TwgDiKwPQt8i7vF+OwPho8jwZonmKmjCt0xrvLAbV/ty
T/LBHq1aVofwg8n0PnyjTdabJhg9FPK+eEelBZkCaUtn84cUvaVN3tk0Jn/XxnHEunYV5BIiwNEe
pQfoElAZJuTWmWCfuH8sgcGGjdcVemTtrTGmDWp6cnOoftetWgG4d/As0QUMsqoUrU/lc5BAFdKN
G/XVk+5ChQ3NxNuVehD14ezOb+I8cu1gUgsOhsxqn/Sc1JEZDWeSWPmM2bCYZKGpcbUIb00DkVn9
z1zc80h7GdbpWOoZqOHumL+VwW5xIIMRYpMgSUr7guIPX7RWqtkE++7SGkT2yylWkrvKgoFTioHc
AymUbaYHkLxaS85aO39uXoHT/UArPA4/cckQqufQGu2jeigk9Pkg+yFqQkHFQ4i9AvTLo828Bwyc
awsKgaLVaX5wdk767ImRzRtfJhJ4Yve/VwKrLN9azSdyNhon4mKR3vJ3y0F+mrq62etSYYkWXtjk
4j8lEMsZPLkAkTBVVifRghaukOqRBaADkfuq00OLzl/TtBVW0JE7rAfvj23UclxmLkdPv3xZcx36
EgTIdKYQS1oyne76Awpogjv9n6nff9YbawfS1zC/H0ltqPEafdML3MX8xtQSmiLLbxgJgbGGg5wf
6SGwWJfjw34O3qhf2ru9ZBAKBZE13xlrUyBnW8Uin7Wq2zuvrX202mQR0Skql6bm9kHOYqPgm+4I
+t/gebTQtCygS2CD1I7T8yMdB7rIGz+HrEkrwU6A1nD+Vdbo6eGsqE1b3Yglk4LOxyyHU1UTCFU8
1eSG29ZPfO+SM1Ia7v9DEO1jSsHcAJ/OgPfxshho9ND97X62+LyCPzS6QH7X38lIGfDVS7/PL5yJ
TS61S87ez3ilkuoqcwSuktX4QTVFctD2O9YKNjR+6NQoKCP9fmYl+jMRUYcnn7Olve4qXNwe6zKd
4fsO3dthRV2OGu6UYZNJxMXq3HD+yzV78YC8S043Gkb4vENi6KuWCBcPRAdexCzpcU/1/oBrPdhw
KOCONL2SzVUTvS3v/zJrxMDtg2Tu1mByTEcUIp2XKPKfyRFsMajb0CFVSzbDneFp174eaVP3+c3U
vWCS5cSpBte5SdqqegPTIYmzJ5WaCnj21ca7fV9MyL6XjeO1x6CkKIdrHGaSzpYB4Lbugwv9m9/a
1E6MWkLCtengyl7mrnc3k0ux9+KT5Y3NNktibYR2ZajVAC9Y/ZAPWorXp0pgHshF5ay8TvJdeWR0
egVBYTYKpje6Auf8yLClx+v1rx0tYpExEsUuMDeKWx2m39csgmMyt+FUJicIgIZnU2vuIqA44nc4
GQRcT2xX979oZ2FeWLtY2+qXQdDFd9hYCVxnvPC2dOHq9D7OvTA48SHt/TEjA2PHw2uI4e68rT8u
2pGDG23xBwy3a8QhSH8OYFWiI+ND4hu20Ep3PuaUUEJzgoTQ6I1ZCvodMc6MXSerb05FM+ZpZeZU
h6sP8QoYcbzTEQvp3WHnx+gBtFbqdv/AVVmVpPI+qFlKCix4GC/zNptKG868hV97FK9unwOiJxLF
CA3OBWauvUOWO+OZGR5Smn6Z210fvLTCwAaPIhzhAWu8wlzr5UB3/+xRi3oAb36l0wVmuUuKnjAs
5wcnrLU0yNerq20ZvmdC+WNwI5n4kthlJP+Z2I7Lmjr5reu4xkBBsYr5M73y1Wo/J5L1UPg4K4Rb
D9pTbMX4qzZSJAjBsxAOJcOzGJLHdm12n4RnU6HC8Nd8NwEtHp8QSgiLuYYicXNffns8jDPOSklY
dg18+b0gqGmWslpf8P+taGpgOeIkXVLxcqHfAUtPavMSFPGOUnImilVeeWFW26+es8kVfW14Uznq
eq2wT1o2/9a8+SXS5V/gfAyvxPtNAsqRG/bESenU+2K0sklkkXbNH4bn2G6PRoGd6Pa1hCVpLe2d
EnPIKIqiC2h7sMy+P3ddV7LSes391sRPN0OnQaHPfSL35xHWjXwptNJorwO+lUnueHywVbmcA1xo
PHQqwXfeJwuUHtEawND4CImC2NfNQwBsSlySRYhdZEGufNk5urYPMZPBthqVsUwvUvd7SrY/d8NQ
B/qkVkgFce12IZL3JuavEfIxbQ7VY0Y4fQMsjHADO/qY2ZfnpVj913MkSxoUkJyQFwiMjLbYJyPo
5Jy5F0kiIjm8joOaBdxLUWNjJx3D4i7AbLC6mzllU+oXxzNXp5IBbf4aJ4YLi7TyKKd6oXyY87af
mK8oq1US0E4Z9Se2Yh/q4ncB7yfEG8q+nLPHcaR4qYpfKZBS5by7XvuFaJzmvqBZmot1t3VCRIXT
WO2yAVfMGP8GfDGdmfKtpIulJlp0UmzttHYpqfX6mU0vLKR8xALCgHiA/bXsGcRQNyi4CNBRXXRX
mHHGdb8FFIKW7Z4IZ0bJai+fc+72r7k1+jNU8hTQCW67t0LtAh+SXs43opzHikUbSTf8UJBQ4F1G
Dhf90aDT5WuFLnpBdY1Bs7Um1MJogh+BG9zVOQV2rPVOW4s/x85LeJToZoE4UEAMWDl7CY8VdZ/e
frzSH+MPMB0rjdE4Nju1JG/gWG9i/PxnPGYbtzAN+3sedLvazF3/Sm+ypVAXhzXazh9PnY8e2tdh
3G+QP/StpeUMMU9vsuWVEqx1xACGMFLHIpV/DXGzLZkSIPp8ZfhS5bdc/KLrZkVPmCCdHU8Q9lvY
+Q8+1juXOESSPbktOEc4tJvroPGakSYMRjz+0436ymk8ROliDZXhHlSGrU/Hu5RqdqwFNPdVcUCO
FhDLSYBMfKcTZSI1a8XkMflBvcnW2QbSiXFmAzYI4eashlxaHnB8iwIrRJCQhqYeOSqlIRECivfE
0tZ7C59jiFAlmrBOiPaUOzUfTadUBzqGdIzJaQV8ruMFl22rW/vN9AAcTsOjiBFQoghuQuyiSatD
yIvKlGCCVhKOz/G6XN2HnImv7hy2TszkXvEdxlrEuIPD/duwRfaV50TCOhhJohNY65E83LtrKaIL
l4Eo1prOV8UUtiUUedG83f6CU2JFZ4W4ga/AzVARDUEbFENc3m7+f/Ntk/oL+GfuX+0BxK+GtFY3
wT0G+EnCIrqYsQdeOY/W7bc2ZgBQbLygRdgqkKDj3p9R7/X8wq3Fn5KFzQRZrF71q22iY3cqA8xs
Pot/YT2Rgaj7t1IErwf/UCDr90FAJZ3b786ZHLAkeznSeYs5DiJ9v/D1EgpX3LqFpq92cWqR22ms
kYdS1gtOt+AmhUHycvAql9UZ/EuOfigL1ZzA3OYGKBXKA3AdUfTIldUO5z4Mn6yZYVykqw85stHh
24ZFInIQ6exspUgy0Xqt/tzj+zDee9UR5UjRuErpr5GY9c2ItjhIxeZ2I4EF9fJxJidsalKje7z2
cCY2on+Bdu5c8yh/5GR/RWlnn675Cjc5ckUbQiZshpwygN1U5cQiE5cPRLg8KOQJ1JrtRUPigK7u
z6FcE90F9Spo2kYyJpjsryjZmUvTnQMGRjAn5qKgzJdjqCEWM7jCbFGXguZ8zwhU5lFYWDJioCOX
RGff7V7smEl+WSjn1u3LtGk0vqNcc/s19Z4qhDDzJAkAKX6wNlbs0aYByLVgr5zXc7tcDvjtvRm2
SZx8PZkGYlYWXlhMJk1ape2btr6kpa2rIEqAYaINfLUiW2yHTwfCyz4xsiedAMg0jgepvje5/cGF
TpM2Owo+aAD0ouZP/pCRnGQJ+bOhfcnrdjjB9DZheb9U0YCMmB5fJTN86f6itMEeXJn0QRO6aLEw
ZRdx5mge4kZTnJnlzJuHBH8pJUSvvx3jVCG+RWAB/WCc1N1epXIUozH1YB4HAaxyjIFKKtr/UhI8
EBaJFXJ3HEyoLRzO8BjRDUczNP1/KLzsNBOhudWzkNj8a8uDq8mBI8SEP6vR4CYCvL7c3Hv0hN4Y
ahQS1LAD9FmF9LJmJCNEYvVgE5OX2oxb4vD3To0macnkzYJw877kGC6oO40p11xQnIi8/fxJHocG
u4QlG265inIURA/MBxDdvm5vSnQ5LdUklT2XPfMKBwQEm+n7iMxYMS/zFcBtgcA/+JRzDA3l4/4W
yUvKyNK7H9asFJFJAX+yM7vtFXFb4bDyEByJ5tgfci2POWG27wUO7DsVMW1MUZ+28YN+vuS6I1N6
LGqc9BG7hQdHepoYkLHMyaBIicbQUz48Cw7xmLBUw8l4vI9QReNFJPsiC4m7IvArEQJCJTeXLxh7
F4O26FhCias6MQ+X/8avZrJgNzMC/B5IU76YA/K2f+T7Qwe8DP4hxLtZUR7BRBmUrvKWoKbGgdCL
viz2Aal5jYtk8xt7+6y4x90sqpmWmeR1cY2/ra/oOK/T+DBMxnOLKIfpcmzlxESD8DRhA4mr5gLh
WkDcNgSa9orF9bajeFFBWl2Z6Ubys1f6Nok3wAGTivmUqD5X+g98MK04SrYaBvbFxN8sleXBoBWh
vy+6kdku+Sjpb/BMel+ws1meimZxJsiFZLydsy2SJoHt8BohVej7qhhGKvIsuLZlqW9mmxRk8PSS
dHZsHs3jOioUQ3/2DBH6TGVosAFfWMQomz6c1g8fogsFIHc4V3alsHbKl82t5G5MTOoJr+8WHGxB
TYsNJmoeV3TCjzOr27vAlrGEEsBcxnZQYIq4DsYWORLdiM+rTIb0pkHpIsh0CeCQV/fskCEyZfFF
4P7bLWt0kQIRKLDoYdMOUuuyMEvS31j4b5KWIoOURq9NHZrzhXY8EujjeziOxXc20Xc65S54jUNv
LvvDQUTSHhUFrCRsLJuRMDU4zum/VG35i69H/Fsl4ksmBa9ghLXdizHyRBCT7zZDuZHLwtci64ht
US7TyJcKryKO9nc74d699tDDff19afYC5BBkspQ0BPDgmjG6z49zuR4ha4xtAWUMiF4ZzF7+z46h
zMWZTPn4Ctz0jk1cBDiopinw3QnLJul47eiqbE8d+RUe8jYn9ItAReVXR5jA8TzxMdN8mSii7/5D
BUZepFrdWojHPN4mAPvTHwF3FZdT4BqQs4tCVnjM9niCBrVMMTXdnS8Vy+xZ3UapRtPzeGTS1nFN
FEgzV5BmtxSUGfarU5tItNwJ+PPqKV8hqyX9zrXvokN/KTjGEc/1opli7lmyurfvNK5rPEgKYWSd
EVTn9Oa8JduIwQ7wYmZPtHnZ0GTjsVxChYkXbQqu6QGAmNdb8N80ZVuwg9meRBmtbV5RBLLLPpLH
4YS1kB04UO1kKS7iJp574OtaNSP1GtXEH7ooxOGMtmTvWd2SmoxzZWGiwyq/z3qQX8IpFTf44AGl
4ILXx9dg2aMFZqtuasT6AJ6fuJ4tsfOzAnQVLpLxUdF7oq20+BsEYlG71j3sO+N1AUL/xoOpDZPt
etyKslfsXWsQRL1aNSAS+bwhBiUcajsaOzIprdx7JG+db49MSDK1vStEfG1u6h9n0QnUmgxCmhpI
TOkpn7HfkNxFnviX1ycGO7gYIi4Wqyvk7aLctJnidyOTYX3ZTyPKkqENvp4Mkm816or9dixXtVvz
9E/kpcYrlzDqklzPSd8WfoI5RcD4fRXUiZMjYrvWpTqs6WyFGNDFq850/ncAwq7TYbDcBr7aetdV
rM1XhihgDWR0kpIZ3GyE0iTkngyl8SVBXLLZfXjy3h6kcbxdGOx1zn/kfjbakyPPdOkvom2/t8Wx
pdtYOy52ZRW2vzoa8C5CqYjS9BrUqYdmGjxwOraxi5gjleog9xiLT/DhqciVwAnvuWPdaDQnetyC
iuvJvpET9cvv6HGuW0LMlxJ3sV5YvtJfwAwHf4TEtZw3bebPttL34oh1xu0ZAXxqukTbZpcQfekl
wObqnj+YykJ99OlHE0GK0OlubO9xxRwA/RF4/bpN59Tk+Pe5BGdRxuv/FvI9l1Zknu90ksalkKUW
wtEETwLlrFKMvFSbtusrB5xc/7rcTSm2ZIBtt3I/bUacT/fE4XoSLZ0BsHKMHM63s8cHhIC75ILf
Cbw0agW9yTnR5zjpGKwLtlrWlPOPa72WxAtQA4EMV4Q/oOfcNp8gxetjtpnWzvLeL9h4jUjAQh6z
leY+1dGmI+wZ7eR797KQXWunWwPLxCNDX8/lUC1PFwci3ORJqZ2sLZKySkKqFzlDmLg35JawnLQX
tBl3hEjloIMUkAwvNf3IC7vZT3tAR96lRfA4k+IQADc4BsK1W8aHcSArKRWf9ais3DTG0hDGgBP7
wWTaS+2nijIgUzJ+HMY919dp2HttxdUS+dxSDU0lOAV+FbccK9jAWVt5ciu+i0Xx+SRsNRb5N2TP
tCAhjlgJB5O/6zgkg5tsyvvy4c7ZWLkamgG1Y15/EioS8SwLgwmCFPN6XeGFd0kudBQmGOtu8y2I
dwuGQN8FhzmwrwbyAN3T1Qd07PT9fZtgKQO2MQ3mpKuEcWxVBSgShpzdxnrBRY5674QMBFD4VNb8
WbzsolT5v2AfRn2H6kNxK8TkbcuqB6OZzjp9OcnfUrcGeFhzORIO2IU22XJ9rDzhPhfG+fMt+m4T
/Tp5U9s9WVwBSLs4Es5LRvWsMOMPwbwADbVW3XI7NE6tzjcncAczvGCOPA30Ti+iEv7LJICLmaWb
Zpe8n8c6u97jtl2GOW3pNjLn4p6CbM3AAbbiwNWM0dIDJm07I8qZ7Nmcjhyzm8dN7Yu1SfzDscD9
H6HHlDq9eERNW33A/DtTHxzAj07Un7ILCQUOodFKWzG4hkOm4KlatqUF5WdYXWEizaHEGZIZRIri
U1d7x5eb/dXkMdioXTYuXKz/zaPCWrfEqoqBVWr29N+/rfiG3b2Iojb1K56oVTMjejZ5DeBWV6s+
enW/TmWcI/leUuw1xaJJj9nzIF7WZ+hnzLXYNAI1S/EUYaPAjjPztpoj/9Z46vE9wsL1sHXunAAu
chYO8D/1/XjFTx2B0UqYm+HkUNUasMREmFRv9RdhPADBX3t07MTapSyRVG76E8/MHEATKkw2CMUa
lotJ4UzkKBg1I4+2B3hK91BDw0rwqI++ca3zx/COh4hhcN6HMnEi0rHLXB4ED5e2ChUcHrsqQIG7
NNIjT5blI8P4K7EHsG5npgZEfKdiV0RDVYqSBavLwhMOk3kFC+O5+pVHsX+t73mvns5n+lUMighh
h9X0nA552be66GjIKVIddlCmynDrfvoag7VExVNCtFor8flAn7hvTJOSA2dd0fBbLicySIvcGkw+
ivmHo/PRxjcZGQlhlvc7GDAzg5bos185HNkCFzQ4GYRSJYO5WC4OTth0GTlcklKUQhOgnE4igHXq
n78HbOtCjr0ff6W6w3G/3+RqLnBbVjPigb6LbCJGo+BTcd8zp6TZLU5jBKmEDciNMusGgaPB/ELY
OIBIedmYikNIy+bRPr4jFR1HKHqwIsYiqZrvLDkdr3xD3mFRHd3DJxYrZUJkR6wBSKwLj0DZYS8I
Xoo+g8yRfcD8DXR0QH7vJBKEvG2V7pCJOpeEsdrFhBqwKo01hEgQcA1i2HMmwqaXg5elZUsV1OEy
Z6IR0Q0nXamgfI1KTVkBfY5Fe+V6TTBS7PYf7U6vHU9eaDT4qnaz8DCt9bCVJ257TpwX23kXCIPf
ryq33MxT6p31HRsjDhj7/CdkAR6kIvedwh6L3qLcS4vAit3/DpjJ3/sSQB0zGxadjyp0U6NAdGEt
Au/DylBBvU49KeNKsLlpYbMUeO/HbyidovaCR/6D+Xex4Qxv0O3zWWO4ZBGaZLB2krL/EmM5ZHPR
2hrgoiy/V3LWaMKheWavrVy/Eq9nwflnITqeTFmNEujTCjQwXsrgca0jmPKY7WJA3MfRWp3JWlXy
dzyoRXLk5c9AUTwHbeJw6WRPZj2z7zfebNPlYomTyk8vZjp7k9BnbcDD+W0A0m3yK9YZ8FQ0Ze4h
XntKSWY/RBSIjRFOhc4RmDYL/o5fv0SmJ/QJ/9GfJfQAaIwN77UMWLowoWR8LRdvQgmHZ/yviUyR
ANgIeo0QbVfzDH/r9T1qnczCIE2gIwXcEQRJ0Ax/uaT1iWxMI72rv0Q7AZW9YoA4c0rERBNLUVoE
CT8ac3kPlgS37c6ZUBmuRzqNTELV3kljr/z6srv0vM7PVYnAxH1whMCoB6Ev1oJ6+fs0OTbL8G5v
wTh2DZjygC3if9LV25a6nnG+dXrdZvdO5kPNBXtXqMzgSkkCMd9DPiseRY+Nz7vrzb5taGAjrqdy
uD7Vr1/Lrst25oY8OrO2FIQezQYncjYeSmfbcWyxgplNnOE56xlD3X+FHtlCqifMQ7SoWXDIUOh4
syWS0GR+THuvcxJjzrqPHCIflc4Mq34WPRGrSk+xExMN6tobTKiPuT6aZDtxN5kW4xvO4OUQ74Hu
XFFJGTf4luUSoQFp+N8aI65yybD5VWtWYtjzSmRvcpJJIYBTsHCwwo6HKsEHNqBFElK0TZMv8E8h
a2ohrb3c9ZDExMVvqci4qQfwOxKa813B79TRWYTMvZiYIb3H6gw4t/flY9O6pH36p/SuSbZhONi9
+tA8D6ulHDfxAkcynXUK4YOugcAoZYZCllUhQxdT8Q8ytfZWwpAPCwNOy0rrJFagqroNGT9U6S7x
X2WKKo+NMENrCS+FoYP8ZHZ3F4kt/4mMLou1oYlTF/Bw6DFdv/30Mn/7WEVm8PYGRRqejslzdC3S
7UGNjox7PNt+tyG3gjBokvXzUzQDmUh85G3Pbfc67PJ1f8aapRIqP94NCvRrxYmLAXy7AK26iBhL
HzWxZmtTt+QwgdbJxxEr9anC1GLVlJUkQeDQkCWFKhVy/hzffrOq57XEcvJ8uoVQ0ZL207/eNwJH
gxceHJjEWXgkCGapqq210+iyFH59wG4L25zNr8vThXyANSuxmlKoG1FGPnAtjSkAtf+vWw97GUcP
lFYDt0wXoSSSP5m9kNrbzGwqtGJdi8036AWTulpwADp3nlcTvT5Y5h9JjmKmHLksXtjbqWAbPPIc
ve8cN3VoMWtuwvAqJSswmemNQ5lmFxtPNw2ZbCKFjNEIQJYhHzSm+Sg8yO0/UA0A6T2KHEZh0HBq
cbkL9YUmp9/puFiDolsblsai7eJSVT7JshDWwpJeoWyw+4QErCysSOFPA58BkgewKUi3/PniBHpJ
upAmmESU8y7kXOt2oJBEAGfhfz+9WSur3Jl1tdtARiqwm5+wIsxPnEnPA73BRVekJ2MSwA/HTR/g
gt35c44RcNu5rE9KcvzGLKWNF0ttp+3dF8CKeg2hWG5PBH7uPIhI1aMTF7O2Sdl/cE6Ha2d7eIjY
F/hXpZYJ9V0118tRT4ahL/rdidyQvlOQJPCy262ydbKJedRHgAgNjAfUEpLkPfosGuDD9UbjFYfl
LTDnm0Go42cwehZfbnlTEStm9iURY9AcfqRnI6s5D4LN/ee2z37iLNDT8T4/XmxKBAxlYcMJxD8w
84b6t2SknuRrp/9KnZpxVv68EWXWTcEwZScil5vNSQ1oT+SMSDNLPsgIcE04VE0nkmEu2J7iO8rK
jH99Sy9tnK2OwTpoCawvF4Acx1A+RNvDOP9DsSgRMrt0XvKlicF/9glvoYOgBV0grM7P9nBUFHSM
pZo5/AN/+ZM4g0W5WT3PlJ2odk17sloxyxiH3XdLCwYghE+xeJ3hNcVFE5cMlAF/Qzki6VSE/1m9
XcwuWv1Bz99KqXMtReTtrnbQkeab8oOAyWu0U+5dryKiOG440zlEmdkomQKJ0mTeRqw2U3OOGfip
1tw/+maERehD+7iJeQ4gA9gwwHRwVqN5snCHNz/6dzBpSHKPkpwBN+owWpi2P2QtCxt2pbsId5RB
TYtFyhFLCrfTzDpctC55g2+8M4U3osW4kCf+Sjz86mwpgsfyVgeGgl88qW0JIBehcKLEJpIoLzBq
JCHBVkBvuysAzAggA5dCdw1Zw8ykzESdzzsgPSuq2AMa2KhCZ0sA5Dgbx1M6MWwHYyYKsgl+xjMq
PhDLEJTKma3vibcnvGQr2qS/v0XO7SUvXxTO+EfQQejFC5UbwaY8QSGIAZkqKPFm6JoPO4zjnuFf
M461t/C5a331UOJERZR1Yh5h9CoSeTFpHY1Q4t8z/kYDgj6WmI3py84xKihPIoUIxFh5kJq8K6dn
0BROYd1OOmVD13uXbBwXy0IfofWmMgBe35pIJFNDgE7bpiYAlr1+drlAUjH5iAJ9hmncO8trnsYb
ruDxZsDbadMCNUeAaJPbI9G2z+Acj7dQitnMjcZJjuOYEPP8KxM63PDoPQvEKyUCpZK38swi/eYS
wqRY0nAD1n56nVrqN6CpWEze+5pFFdJfp8VU7wb6Pv+Oy0jtbc+VIq3ocBo4Ylx1VggPtR2le+uc
P/lwxdW9w+WIZF3z/3b+QwMbsuxnjN+UTOzpJ2s8Yh7VeIsjqWf9I9oZaCKgG0To+6LOXPoLvR1k
IZnTjRtSjKKv9i7oRM/K24T45RNY0h2aQHVJJ8IDypPQJvjyVMuQfKUWI4tRjeW1mRuevJmimlkg
yorFOdk7GSXtGSTxEdDOKGZsiNyz+o4eHMf8k4V3tVVYqzKhsz8/eLNu7iKAEA5o9n3uAwyYkqQN
GZEDO+9xmbqBReLZAoY+eBHOEBCobhsX5SCQAimwlqPNpl9qJc6jH0PQ3UnOvKWzzC8KV4B3z9Wk
7k2V64M349hJIGHedRdc30iQXmIqSOwHnhCdHOL5riFngh+wiBLzPXtKeqeQroam+n/n7iObtQEE
1B0EaPeP3jZhdWdaktkwVsWpz15FUz7InssdF9mhUoWwOXiGefw6hNUoJxYxjf5In51Z27brqvKw
v7i2xyWGySbX3gBHeiAkFsbaoIynZWLCSKCcy7mS/dYW/vUGmUZBsIdhMYz/q6olqMczdiXUqInx
KoubTicjGs6YBD79euyu4Jq2NS6E56IAiEgS7CH3Sbk077XlHZDYv7lWJ6MX1WXcRMdlCO0lZHIB
SKHHRB3/OKEx1VS86jyzTAnPA4cviIu7TpbyYUvpoNIQZfnBX0Mr2w1xt24pjX2KDRl008QZnegf
Qskd4i4j3VgchbQ6IxFjfX6F616r11+Y7gqxs/IMq3Gt70xl1ug4c8KIIunv4LuFS3up0HMDcp6k
bh80FHFrKGIOZmqpIciDhKcuAKFL0tFMjsMD0Nj+LA4UqYKwg5rcNdH3cexeH0y5wmHBLjc97CSh
QL0aPBNMtiXFvi+XRkVhHtip9fSiWQjiGfNnJMS8izsK38zgtTQV1i4sDadZFI1mVDppdsPCWwf/
Df6iD3MEpB5PCGh4e0et2g92hoNwMzVGcPv0qb5oJ9harsTQANRSvInrNHL2+vEnh9CYBjSQFmwM
CzzuitaH3R2h9REn7hTkxu+CwjCPXaBvPc+1KpDrtBenW76ypP7iywGi0wB5dnq2BOoC92X8cfCG
X9bMTAWv1anIUtahz7nwyHNUA0nvpZK+MGyJMqwfOcUQcoQ0zR8MRnxLF0v8iRbGpdn5Igp7zZ4S
wvGF8+28vL6Os1bfPhn0T/OSbde3Xl/+YOJvdCDhEr37M53lgcV63fVPEbvIrlMltAvKiEtECmfX
pI1eeo9tJtGGZIvSTyhTjxNeH2j7AkUl/5axJLH+Bm9wH/ITqJxObWxUCbibwhb9c55uFsKqPdqf
wMWQlEPeHbJOnu5sEFTXOBXUuvL7EmrBEjZZ8VpA5JpMTBK2HxK+WViCnPSG47oKD5YlCDIikPGo
NuukOvYN37OBsutoqXaR4ZLNZLTIjl0dEAsqOJWAYPki5KSm/s15l5SiTOArVKnNaBG23xTxAEHR
Ez0nI9Sw9F+gWvBZer60HTpUP4LwdislaS+AszsDATERhmVBvhCkW2SodP//B8HFHbbOz1F2X+Ua
g6lk3NN5BuWxs2i1rUbzIaGuNkkDRRsxkdHcMceMEO0r36/5OnVG9GrD4HazCC1vz2nZm4CRF/TU
ddkwQVzzcQHYRi2X3rsR5+Xuc8Kn9qa5EJgvwsaL1Tjh1IN+c+oRJqIhytmPcpsJDaAXoxoThpU/
pEzlAMQ8iODrNR/XuJ2Z7zT8E43X5fQGeWVg6uOiVOVAGZgkJJo3ew4aJC/iSICDYLfz4EDvxFxR
CZSDj7l3I8KIZSRzmoKtVbOLlqH6mkFoqAmmZutCx0ZrKGKLjgW0+zLRQywVp/bVNkWDvmrT/4fZ
HHyVgzHsv0QELHFniyp8CAftyLtw3e2EhSicRWHPEcsUxFP76581r/EEx21Q6RMKXu+7m6fnVD0T
HJpIQQN13Cz193zmKQ627VKkamUmBq38favfeTX8zsI6pK93o91px/9I+HqnQDxLlPR+ZecwuQct
0HFrjTiULeMzTEcUlGaDUrq6/yAmvgOXPTk1sOEGaWhXQ4vcWY+CsV+AYscYQR+Ljnk+AWGYdj+R
RTLFBGsRivy3iyEfpqns2gxgbS8TzvwQ4CrBIZfdMDJZZvmscxCpW7mSSg76ZhoJ/ClBn+Q/mI7V
lucpnq5tyTu2oGbtUiTQZeZH4Tf1zV+YnJO8BlISAWebb7vUSC3cFuTyPe1ID5QXLyHtC401KGs2
nb/4q7cqSMPG2f9xvzNFztdskPiFoQ1Ie2gcD0mg+x1qxp7SDtHXuEgvNkIadzUBHIDIhlwLXx1n
gOr6AlFJw4cfoVW05w7T7u+Zm13OjS4rlQhHmDnJjVKXoc52y0BjYVdx6Tv6cpv10IvsVi6Rm6fk
oHFvdA4Lz21++gWCQjW/IyX6l1hLDp+7U3tfeRT4fK2PpxhIRAjZp9f8hP6Lr5v00HD01jm5PD4t
zDGF2MZqGeRCCBr+wjNnq1z7Ko3Tg2qvuRI5eM25gX2Lfw9pSWTKhMyBDQpdM7HyggMXnOfZx3sw
09teU1oaWuaAefeGjuHNaRXLj3obObVvZ4EpuZwtpxTL0NVzqsOkj5bv7QNn6EBfvu3AC5yZTgB9
Fd/HH2jHoNVlcthHLidCOXQAJtlPiwTdTTKQLVEuPAgShbaMt8ZITxm3wJOx2/lJsG6ffNAlmYA7
48VJDtYDD/ePdp/l5UGeR2ewK4nt2Zx68NXphv/ZXH5h7oWtaMV23reWTfoQRn/eG4cb6zQTH6Vf
l4Jkm/PVdDXnhhptJUk2qbGn4EIV/oj9pFbYmQ9g3r7D+KqthfSrcsuvq/bs+f/ZmufOFK+ccRYa
cibiP+eiW2E5Z9oR1B+AZQHAq9MVXRk/8hZciqU9LtabwvYqRuZE7ZkB0FJ/m2CS6a1m4LD0XoM/
44gFlINSw06lPrtjwfXHrnnUA3lkbu19jALNjHt3pX/FL8h3qqKDLxj2JwtoBl+NJZIkfR9l/455
EMTcTnInSw+tXwsVF+kreQLGtulgI2iOns/8VDS+HxClCBN2wCpGibfU7FAeXu5kCQQTM87/mrWU
g2axmCZ2UOk38T0eosAWd6WvMMF7zkAVywbdAujWf2Mo8iFOwdi1f9zF3caW3TrveIwtbSVse+T2
fXrFsRpc97lLYbsHh7+K2VU1HwgoSWK6MB3x8qNMXleXfNDx/zjtFZubSylf/0RbkCftZWMVDES+
tOkmb2SqqbR+hweOO0ZGfc/y4frYKN6RI7GndecxVEUVl+eXd4fCogTEFAtVuMkMhy/BSpt+an6x
ZtYQeQknKV8xvO1wtzzxdWBYqs3o5as8F9CmADP/LSehKOxwWdAFihp6TTApazPiWuyjfK4lwlwE
BACYPO65MyjDjvyiDGSqlXnGRMkkhvlZHJYxZCWPLXeHIzdOGlTUQF0IWCJEu414aaQhO2bae/DN
YGqcqy5QbyHtr0QhhIRpx35qJ8FGBr/HuuTE+MMp+V/IJzJpbGy/yKQYRmms/1/DrWIhTsS3+zcP
ZsBSYLjDko5x6/JiRqQTI9lX4R979/3yvqOnT4WsRTpCJn2/v1X7Z+p9nzO0cb8k2mL3lJpVAoqi
KNbvh02gj2uO0EktePeaHNWp98UZotJePdl9Hq6mQ52Z/U/jRImD0LVruXHCw+U/m2cEzDyXMzMY
O6tzwo9CoOmdK/FcymZOekLRV3g0TVIJq0Had4lciyrc/r0MelbkpQWwbEMeqUQDR/xB8WYLBuEs
GgEBuwR1OHZx2CXyebIm7NCGN+J8oas2alT2SLrVlbhhMgY5l6Z9HMPUxqLhn0K6s6ekcxErovAF
LfKJx1d9a4I46VJe2P+ySnWfysGyaBuaVKqJppPWbGX75c0LDnXADWhIBA+acSLx5yyUoaNRheul
KBwth/Zc7xHRt95H1LeC+IGSvLZAd208CGroqqPkr0b4dVxgRVyt4zKU907eS8vf1Ef0DFAig4gS
HyCXgtMEpnzy7yBnhpWdn7Aax9JujpcDM5Lak0rnbNNKLJ7o2KNIxLbH64QPNx9uAAtBihKKSgut
44oyI5cPqDxs9LieLL2LInjimRWxVCs68PXOqDlhxHr+rw4Q4LJ46CFMCw3xchy77E2+0sts8ylq
3WMgLNLxiGkKfw7DPhaueqYQg8dK62pq45bFa3BdPWEKUFbXsVWoBeoQAYCyewwuUyKH9T7N8kTs
qsfKcNLCZSf1/Umb5/ix5aGFzqlK1G+DQtQrE9GhcNYzTdjFiqWelF9jw4dOywU5WlrkKrub33+I
mUAfP0fSIwLm9Lpv1RYe/aeAHNf0B4lfWIImun9JsIdslb2ND4e0KvjRSBIavdVykSK+keTRmVbW
pld6NJXCKcdNjq0HL3rFjcQGIQS5Xb94sV2DWt8TYFzmFhBD9KSnD7f/5tZLS69X3LMLrnpfLDkb
358IAqLtL8S6HPNNgY8rc8aFFynysCUyoSPf+uHDZIOaNvcY907EdEBNwYMxrWqA6/cIR5aiJRgA
PBEXOQoeVbcMSz4eWEHVQ1ibAIK2pUkFPNgzdVdimE1eulq6Y442+tTNU8A1z61mnZ2xF1O1/Tax
aqD7wvuqVhwLy9KFuNkGbP10cHr85vyJjnTGq2WVfZ1s1C1Y3ik5+q82ECb7ivAneak2WxkNONim
t10OwbgC9iNGU73PK8a4RP6pkf1ln6SXyRiRKmNCoHpJAU6LWXv6nq6T6t8ph23DiP+rOJ2ER85U
ONMaU7REOgfQ4w9ASsmJyq668EZ8o1zmkhxNv5mpSpVo5AanFv2jCyYjEfeN5ClWMuLRIw3PW9bs
+A46vX+y9x9bvO3FSpmcWawM7Elu27qY2FDIY+uzeQU9pAXNNXpdfQ+dPOHbI3+WhhatgTAi2hta
nn9zlFwIO2ULZG3IN0naTw8Lm1QLVWufcNWfg9bMuZix9Jq0wWIDzBDuT9UV+WvvmuVgGpftV5A3
ZsKUDxnJe2vG6EsvxnmMIUrHETSGCQt9gZbmXsj29MBForc7BUkYl0AZwY8jqFP/lflJULy2qTCq
+Ffh9+WPkG1dsKPAbvJQezVGU+ketwvWRUkr6l9Z3rWNB35vt7jZas8CQKGb6MVelAXD1offWsk3
H4f9oIKL+VlkdFppN9nyQ2lx4jlS0N72kbCYOCbtS5/rO6GuIPbrhJTdVYtzefDeSuc3JADd6eZY
72Jp5PNQ90DD3fviMVe7lt4N/sEIC9iFPxyrzo9dZrSkswy/+PM4nL9bUvS8HRe1+1YTV8nn041S
mz6pmKTKsmepfVkxSP5lTMUA5GXPm9VY1YPLgxyBn3e0jhU9sErAhHDK6hrHi5EulAJZDFdzH3A4
0OnAvEvkxssGY6ZJuDzs/QGM17YdLHmAkfW/2X4LREOFMBvuu8e3tNgNV3umQbb8HNvPDgP8xs7/
0wIxtOFedR1c4MEchrnl8YQBSxujIeq22MGUFgZQQLaB2NdQ61MYgDer6XLJBZjdK/YkvhCn1LPq
CcI1TH3fJ4og5B0Kv93gsp3mNVel4XmJVDAILXesrJxVJMm7oP1AeXUj7D1PhkGljtpD3WXsfuKR
QGF4eukqMB6sNTaz5uh//CNddNtXrhbpD3kQVtiKCeU2+pmCSformWeM+v8cUoCg95N74MFLfn5n
xUQ6jNfjl4wtKB+ZFNO0muAYhSq9HIFj9aXIcRtETehOjAPlXH8mWGUuHAQ12I3d5/FimD6MOwRP
8vxiFuwWlF0ZlH8VzfTnHtcgCc3EFGG/E8Qs0xkoi2kF2m0s42s4C94y9RbceHVb5v2kmnFRyaGC
5fw0Lgy51HdJYTDt2z9v6xHme7qVXrf2diGW9ZT05U3I5Eu7ASDmFpzpnjrvqopuGNUJegx8TSAT
x1Ue3KPRycyDNJYY5oV9xtBNpVH4GDMd62xLG0TASo8xfJWquTu/GA9eFbzrIdRywvmuYzQ6CKfl
4rArjzXlWT+gr2rO+4x9oR9lW6Ley+ida4fkR0/BDQNPLld3Uhj6ktjn12lVh4RlOdA66/cRqi6s
edR8JYFT3NdBEU2OI6GgRX87R5W4liIG8jkowT/I0ZS9nebtiqPfReh9vTssUceXxMLaCOAlgCoP
08rFKRTPaCkNoUKhe8DSEdMq3x/yjbzVK4RDBcuLjRTJ9dQJZWaM0JLIW9AVyDQOtkCeC70iJxKU
BeRVbaaFseTqDzaDVpabs30FAbOlgO/MsuaTZFlq7RGg2iI1hZSJyiPbtTS/e1OP9FmJ5SStUGi1
k41f/TPWAlBsuqI/rHXXyAINhctjLAHy5qPllw7MfqsnJJXi6Bgmr9c0ffskdRyfE4Hgo0dG58v7
2zBTeqYV3fWK1o/EYbwkxiQQJalnUpz3nilz5LHMRHxXWQZT8tOyQU3s+VJLa+TatUDwmlynIlOE
StUDOZJamKiH0z90z8CzNR6QrwxqkBcILAeMj8Bq4LD3NOIny5Tsg6VUkANZ1l6mwzdPkPW8LVdj
mS6viMi9lyHDKWZyub23FyhwSVbUzz1YFp1EN4dr7REZlTvPzrgK5U4CIh6eODgjvdsgZokKxBh4
nEYExi/vcljbGGj9dGzOETquFggNH1KYeBeQ5ru2aZ7BHjPUd0/DbnNaUfaJnjiF5J1NllJkGN0b
OoX6CwFATUtGsaPY5dtyLtXAruQmX2LHhkvemOG2JXD0y6CDmBvm5awYkb2LdlyCFiylkLyfga3L
eOnJsyXCHkKUO4EjuKy5Tj9HoYBBzVKc5abc+5PMKwGWpceuOWP5o809HK4toERf7cAktcMLxNgY
/NRG0D+zceOEXKnuXdln0/0lJvzzip0SYACSl49E6P+BUV2uKcsq4TrryxL0SLqviylYnrv5cx38
bkY7v+5KxATHVi6LQOKJdGTLJBoBWuBlOjLzp6LMTVL+RWqQ4zNNNlD3jAYqbuJDCkTrw0LpeQEj
fEuwFAUSmOwUw3gPihAmXfdh9ieSD0CGkQXHbwQ2GeGSHQHbFTU6z5gzyTFmJVqKTTA31znXrpOt
h/LMpUiBr+j+pRTIxcllG2T/+ZF3aMWXtQXTCMGJ1rJsYbXkLooV/PpfMUPh//rpCryBXAoad14t
9Popvi5T4vN8g3egEvK/jPwivZls/c/nqc1pDEk8bo3xgu5G14GAwbTwDzoUhKNXZwmiCP5C3zwc
XDWEc5RyuFONlEc1MtJchmn6m6R8Jl3hTaxqyT/AXLYQ+zzW4QcyO/V634QXVS7XHOIIciy5zIJd
Z30PY1boFVYEWV6jLXjXCTctp5iiYRzgw2jTeQsvVkBIG19hlctQRUwJJq03L2VeuLlJ7Tc/g+4N
PFPpJLqVaXB4zGxcLKNE8J2K4XZm+Ng8nz2HjIsGTkGz37r/b1Q8
`pragma protect end_protected


endmodule
