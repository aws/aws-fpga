`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
C+IHN5J8uh92tq1VwoEDU3GVjJqV30J1f+6y+lBjBC4m0ayCEY6d+mmoO4mWXZtt4Tz80lMMVYVw
CEnkrn8KEkCWN16mze3V0z7P2k+HwHlVw5Vs0b7ZGvROtb2AuiZUoHYQs7O6bTe9Uo8nHtyvDPP4
CPk5H9UGIHB3TJxDpmIZxA7YcGt0SMxsQ22b+Pk0fS1TXdleCFY2tNSlcBke4z9ddxV1ZPHJKYsm
cxmZBjO/ezwllX8ISOkvuckKNiWvyPr9qa3sCoeV0JM1UBt/YY/wvL/IecbPUETRTYIubH7JTHOG
RzpAt1hPScPWZVUsEqWjrPiKCU1B77g3Ls5XpA==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
d/yBEOcadhrzi9mmx2yDHWxc1ngm6sfQbwY17OmJ9dbKdyP2gNI1vRcCYrUhBPQrCaUQYNBmO3n6
wN2ic8P8igW7WnRgkv9mY+MEibFE3hGTI1dC2XIpHQ8u4hOyhgPRGVGq+T4cQBx0C1BpVq4Qt7DI
paq+dL10WlRikpw1VVU=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
F2gbL6CYm5LHx7Ms6usjnEfkv3ZfWBNO8em1WAHtZBw27Gc1ttSYCF9DZj3L6Nv9aOW8FT5bW9Uz
Yf5T1EW5QGNOdsdKtoJa6UbFPjp+Gy2FfjndIg5Sz+LPmWM4jLqN5MiMNeRCjhuMRfvO2YH+nEXu
t1OYI7QG273/30e02U8=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 11184)
`pragma protect data_block
t68oR+rXqcpiW6eTUV6VAXyEHvJLNFzlyBzgZZW79TineL/Z9Y/Vf/vGli/LK1M0bvb2RmTj+nkw
EnMEsLI00a5PZOe7FvOGLQn8XCqJK9yrO9qc0mDsS0efMBiYBRlSehRHTAaXPz4hgLURIOcXmMCa
vOWScS1RA8cw6xeAV9ZifKVxJGb7ePs+D0c1GOUOOLK6nKedlv8HXGddp1ttuz5dIWrwp8uSQuYT
Sh7nwa5GZg0RMhsjibnKHm6UX/aBX4/t9LU8/u5roDshnEal98qAJPjxxDFBYuMdCHaBDzI5daxN
JGr7yU8nPWr1dBL+nGTcUV5YRHUXLdF1b5ZWBDYvGXdKYk4M/7VoMaKnOB+YwlwVdRiPyQDqiLKW
bnIhPsrJ/Kp3icjcwdl4ViuRKoaoMpSYZWrscXdFLNDpEF0J848PRgWanww06VqYGa7q6OArh+tz
GWgfYJFNLDESN+5z1rSSw/S15/uxK0rU2hafjB4PzaOH8peeOiNWfU1DwbGYgvjSpt/ICLpXPTGc
S3QnbPHelpQ2mFvrF2fWNpQRHqgo5fY2ShrGtRbTAkDfBPIJnjtyWF/yCWl9KsxSZiSU4y8sKv/j
fMnlhhKg3f+UCNVo7/RndNNHjbwGRn+P/nVrHWyFXZE9OHPchePPx6j1sxwKljzdd5rSaz4XPifP
O2k3H4xkJP1PcawZ0qSFT/YpaYyZpMLQRsHWqzHoFzLo7atWtU67YNfl8I5t54z5NKF+QMw8Q02h
566bvsXGCEjSN9ty2ZO+dvNHX/AHn41iAOmARfe4pPd1279KYbj1aXP96J9l3ucQaup0EGN1XEtX
UYwVN8f8kM0fFRuLAF99F5jCzNbmfBBxkZvVdRQRvDB3VqdVgBQDHjmVxosyjc6BWDIwt1RCfLja
mJf0ng1xDWdA5jSn7Ck5Q90AsWFYEKbLgzG0dEyf0m+bmEwUR+e+rTstxlrZxSpTKEUaHF7Gturx
ro1MsXuiNFTb2DnspXS5MKfVVAzbnZiW1TXi/8qXjn3RRZZN36GYuNwKtuADUESKsX/IOMd+0c7E
Z0EzNjmFW2McJjIIbr1Koo0IhmFExjS+PYRMxY83JbdHyNB6LwoBw2ha3hkN0XHzcpA+1nt/GuSw
6yWGiLyFHfF8/Sf6GNWF4dV4vj5wXoSgIDkbBI9XfoMsJFQvR1EWT/kYptG3T41/kNMGwY8cFnAo
IrU3P2vZUIgwA1B8yvvDrpmqSfvLNfcQ3PWLDbRsgBp4ob50TWEmqGTRb1di4Bv2wlnZhmSCpMgK
pzDuU342+WsJ/TqI9OtYieOlSQFhSLy2SPsupR26ktN05ykJtS9+IikR39gww7kGVEPpjbFHPOna
dTiTdlWJm6xL7yJU0UX9pjg8XgZV5DDHWWjAebKvhRi0GOutqSwHG5GID4ZThFuHF+2HuwkG6p4u
NfZ+15DjHCWahCL8/qLwpP5sTsUN+EQ+JZh7Zafg0mw5QICqAKPSTvwP5puEbXOck/M4E1TJtehL
rJs3biN7LreyrrM+FUWXImjyAH5DGLwrwF+v56kuwaU3DQ0W/GDHanP11K6bZsAYqRvgx65HaFki
3hZ9jqxSUvLdCzJ/QJzu3MNLSd2Z5ORJZ1HNO4HVX1wYLsTiYT5u1lBEuVeQAV25rAJ7rWYY5fFH
MgUrUaWUj7BQZ5ca9QlOzLr8YmTT0ug2CSsBU5EX9t9y9xaToCYrKnPlrKFGqys4klQGer69BDjH
yowXRSLlSp8Rj9TKzqFRyK8ajGsi7PnhjQ4ZDpiLDFZrvBZE8+wI0odbxyHp6qgo34yEqnlR3nfe
z2XI2OAPGjs9cK5IuhXvXNRIlPdC69eHZeNktK9PWNrA0ybNheaBIpwcezWUTeHUqx3BsWtc0Boe
sScZ/D8l1Wt42kRODcGq598boohRF8XlAKiUVxdrVu2qdX67Dpesmfhi7A4DlhukLgWzNXLm1UZc
M1+qBkrfVZc2aa1Df9fImCNoiXr7UeVqhOSSYrlAvG67T9vIGYd16PIlCzXDz/d+DCLFdaGEJzbO
uZs3rCKvJv5SO21flDVDOeCXkdose8IB4nL9/ubCj1l6L1I+Pmz6TxLJU92yRG7//xRut0c6TsLR
AnFswHtz1s0fhehWKYCsebWqGoEg4PE+K+Kg+CCP9/xcp8oyB8FFAoqoOO6yB265u9WFiZv6kpyD
hENZWHiwVGvSjMHTR4yrmsaHzazXTFCXvg2yXem5GZIAHaaAsqbQVvlgJJoP9Xt9FRfpc7NTwsqz
bDx8EwsRLuF/bQJZRQ48xE2KcbnGIEhv4m5T5fC08mc5hiapUkRlWtLssmeTNZuAj5trRjgXBKff
0wt7YEo2nYtmrWwtOWWR7AnNjQS8tUfHyb2TWeauHc8IEovn4KOjwbFVYWhUayMpXP5amHLSenfQ
Zgf7Ma9L2RdB6P/iVqESfblYJ4i4VEJvFqDvi+Uz9/K7NKV4e3WYPAFMCkSCstl/z+BEJ1CQXl5n
pzgYV7GqROgWAQkA9fk3z7AZ1Zx5fEGbXdLBVF1zluXm5vLSwZgR1dy3NMmCoPbjt7NQASNWYtTt
9goKh2yeICf/83FqXL065tEFaVMiCNe2vQWeiqfYaKZahSeqZ1NVpBhwpApsy807ihFtz4JQsAlu
BPrHzpIsi3R7p9OdWl8t8ZJZF+lBHoAS42DI58cMbSgH6AbZDnkroUNPxcPuqQO6xNrsXZ9e0FF5
svtjsw2a+Yr+52ymh6vVi4nhP3fN03wn8g9HDZmPboVOEpR4fhjVYvTUFFwHCGL6GtvXqyv2vkeR
IIzeGgKk3wcNhTFWO15sr3H0VthOnSWsr81Qn7nILWreUCz6t3+3nNOpaJ4XR/OBWe2d0CPgKudy
qKT7ywpfKQ0S3RjfeBMHgJJQqixOvfS0dcbqFBoFKfLyBxz8QqWYwn1MpFinSfXyA4gikveRnIdD
UAf7m3ICvPTkLWu35FgJBSdCQPn1ro2Ep5aSZbWHmZsqv24urY3ZqLXMr00/93UItKikYf3Ha5M6
sx+Q48RAIjOy0WtkSxz2vQHlGHFZ+tSDQEqaQYm3wujLvjr6j7JkmR5ZCuNolhV3XHYXcLVTxg+8
ZTVxLhY8wQQ0+jAQladWRrN/K+Ywx136TxHzOkTprzfTHXAThTy4G83YORW8bgU7BL90fIAP/3ce
+0qvuBH8nAS+EOMoqOmjMPmu9zbtk05OUkurRVbRg8bVzrLeHCeCBea90NVlt+R8J5i9z2haD/F0
IgFWMQVRxM1ObmbmQxvVL50EoLJcX6Aq9AcQdL7tQ2n4qySDdpxEL0Eg+fHfd/vQIGRfUHBlOqfx
JSxyzQWNr2eARQoHazbgu4vd3QDmVYmmY1w5sJl816qvQrtgFvNnnOtK9a0SHWYsaJEkUB72QJU8
QmGnnZ3Eb/yt3k+Szh9XrqgtJHC33moGw5aOp0+KwXpvQQ6TfT9uraUUS2NtBh4+4Qx+xjew4vqi
pFrZgcarkhGissY3PyIu+H9H2AOpttRYTod17rWeMhxGFmXB/X75SEZ4u6Mtl05kTD7q2rRZUDmZ
bi4lEM6R77UMaUP2H0nCYWxTHX79x/ipBB3UIrUDajX/b2m5ZU4ta3fhL3G33qSYxBPl7LRKuQA5
mEoVrPC8pPuzteyWwie++0q+ih9ZSJ38fVjx6Zu6eOE0AWuFzM6INbF6VX6DuyaSd5pSNjKPJ3BQ
588tmooLuqf6vC3bXpZFFJr8TTsWpcFmm4Vd6C7cFSFhEwqO0WlBWJK+LsDk2qOkWsPvqAlKbSK+
gm22GtsLjRvphyY5YRejcN9qaPUuweGTQSBg1NXglBnp5Bk8YDVDtRlf9/iqTGHmWiyeT2UASlP8
CcGipvwVkW3dhkKrAXkvIdz1qnLFMzV5Eu+U7598fEK8O4jeZX/kf/98/zDIwZNgksUt2ZP9VM4N
ywgf5WnJGG/uXju3L25rcSGeLHc8R+utI51bzE8bgQc+4+y2Xk/CorWH6SlylIv6UP6cYSPLsg8l
JZZHplE/kJzCKKkc++pgjeUU9oBp6pZERYbsf4AR6ECFh7qOb9QlzJYF6hrSLucZriBMRXr1KI57
KvrEf1pC6CB3thzla0L4GyCczZ3iwjNF1TAQWlQGenDFpH9E3M5Y3C+I71taFeqIaGC5tOvzgegG
q5j2IWouWW9GdPdvzyl3oEjK5InizteOD8w8DWptIKtRYnmEVVK70ObgbgfnWIcZKgyNQlDD8zVw
ZMzSKdCCVe88FHflfwkTwNpVnpHZ+VmQyGt6FHK4xfaMZcmYMmDMK3ORpU5kJA1pt/fZ1QZ22Uec
Z0MDwcMLrEl16PpthgMz/u+mkftviuGKy47LY/1WuikPqOVtCs3IwKdagh0YjGz7MLj/VriWL0gn
zK924aE+s1sv+MdqIVVjVbieZ8k7v2ruC71gEzH4EVG6gOKmHI9NROTqyONaGGSNZYLWJIrzf2c7
CLdK6e59rxsvatCMgBErWo0s1I6V1ajnXu9/q8mUuw9X7pnNBgCdDTQBq9KgMD+O3OVmY0vH4DBi
5R7bf+73SCY2lgpkXnOVFGIQNSmLsFhZWLpi1xRcxwtF39AeQpp2VwAYu0WLGoU1998WIzRQMKya
urygue4G0vI/b3mtKwl1ON5nh1uBfrVV5P/5vbPOqLGBiXOYuFhlKDeM2ixAjV4u4ekfRZOu22mL
7b2c9/dJaopflUsCQXX1xP7jPRh1aKVaYIsoZNvcnK62qBxYrciMGNFY3UCjt0zQy9baZByTLAo/
Ai0ZmdpFIiEcRDAvCctuU/S9kBnXgMaa8nxwYuVBdZOwfIv/lFDduC0a3dxVzKTdKY+JTwb6US/+
gPJeQ2kKS/xBP3WFEvsp5FmKg8hy0wGC4Xbqw6MZ5wU++axA6pCsn4Ti3QOg5WD2ThXsRh6/Vu7q
5chUs0Y4NY54N3xaEFx08rp57O3ZRMVOzU1IW45iR/xVBuuj/QMLx6XJw8InMofwidogYftugvr+
eI7FxAkqhhxA/DCPjgt7kJbQZ2ysqhyPusFM+akncqvrNOE33Li+dqOgfjtV60snFKCFpEWWawnn
1/lkixVbd0JtT9Dy5t1Fr8ylbqtTYWyu4rkyIVNg+nYzpH8CwKFvzne3BiRPfa9wymMy9lfUVU9q
GnQzFn1hPimNurLsi9r9gps3cb0WIWmwVHoA3Jmlt8LqRXNjPEiqXmYrx2ej0VRPAIAJ1MZgr9zE
axJ0BgbYzv7zBU5W0ZjCxVqHQMjHnP5i2DkQOjGMaVSe/bp8Nwe1dN1fX2fbhuEol8LXAPA8cb3o
jX9LIeH97yg6STwo8jOagapiYRLTTiyoE1HlUsqOWKFjld6JyG6MuGKNW4zt2laT9zwAmX133zXS
nt2XzMw1aE4CX2/u3EdEN+PRJansWbiRHnSgy/kCXSsfZSY4nhH+0fRGBTOmTjTVC9If2fASw80l
LxfEZL0GXCBSJeieo/eIgaFoxktO7q69PnxhSo3hbAQbAVj2jDDHzdHZgGXlKJCvZmN3DsmPFGhl
konLFhfwJSx8D4uOmLbGgvWT5nAJnHIu8/4Ozd/33TrVlN1QA5QucwqVmscLnYOHkC1ASMf6/2sQ
mUv/QW/kOK0Q8bBGB1xtUS3BQksHKsNyUd0JtCkRLXKZee1PAUhldGLSRDZWdqEZJcViJUyMIi+D
ofyXT5QSQKvZtl+E0rOSW67WIEN9gG2Zc5+Hrwx8XoyJBASWCq8+Sk7nE/285VmSnZm16Ys2OdJp
jkt670+wxbivUveIRsO+bYpKXMMecFLqaoc1z8LpbwXiM/uW6IFhvcdr4eEMx87FR4s2P124Kjmh
VtxNWsXygXHN4ekf52SKef5oKDyF2yy+GmhcQPnmdNd51kJgX0gFlobs9/DKLHFG/5JmJ3thXjM3
Z9QSuwLO974jbjigwL3SV5tMH3Cre7hDpChG2KPUGA3mwwbYu88uxQyOqfm7GoAKLBLAbK2wnlq9
rgHegISMCNFVlDMvJNSYfauQc5QIdWqYQ7iklORBhXvxt5BrKn6HDZbUeIXuoUovi8ei/Ks11nXE
ngwFOGfDB76Fc1yyOn+RSyJ1Vw5TmNKivD+eMXppQCKWq77sgCPIrlLSv0nOa1R2mYfp2YApvFsc
4eYE0ae6NElp3baEIYteNQrvhLMcqx0F43txFUHETEGLTQL0xyqkMFtaDoTtcyENog3wndq06tNI
ydNRXW695kI7MeHWGT2mX8Uvlx4IDlQ/s+ST3pp3uHLcIAjigrqzdgwKW/XlSLA0Q8Q44U6/o0dZ
K9ygTFBqb+YbJTaHdIjqI7lVg09SI9KuuW7Sc6I5l3iVfy0+bWNEdO9pVP24ZXkOvf6awQpZXjZs
g6HI++1ZhhzucT1swG/2j7LmKF9DaoKNJaE3IwXCTaO0qc28P/goI3zF6fCTHs0SdMLgvsiHsi6p
aNa61KpFAX3Qaf9bnYlw+z/T2M9c4Q7HIo+b+Hi9NJHdDvRnLfKdfl7bs8hONCH1uMvN2IMCvqbB
1WYW4citZO7tuaUqry2b4v06Gvwqqv2VbjWndGVo/ukOmbHBGefr3uLFppceMDGmC8HBoZhV//5h
OFRqNcPHpt16in/8MGCkP6ibd6Fqd8bylEQ7daB6MzXzBbtxCMqaV3/Rc0q0w/wtvC9yg5sgdo+N
TiC/RQ+bNd7Ui7F8AEPcnz6BQjVLZvyN9d8kpYC5ADloJbAOq3n4XTzd8VAlARcl1DRqGLoRfTCD
o2BmL9h9xYyCYCfB0HCyBSv64Ooz/ctrADqkmTvaCj3tO5OPA/c+H+C6uTLDKdBV8wbqfZqLRNjg
VJS+8gwcH/7ZBzzQGAYk7es2CIIK+asmCPu+DlL5kRdo3gJ4upQFpe0ice1wOXDO+iswrgyW/1Hx
Cv362uc+F7gTP+F4Up/uELlxeCwfHCnejzTLZwOJvwSVVYAwedBFYISIlumAjotW7LBTRzzCYM8R
ynCAP9PB5hqMKqiRV/r7tVvVfI0u8isEuX484qv6BiPXMDEVlHvADIy2sa57NWE9leBQAfBUx+tH
pcys0MbBwWzLYNsl9PIMzgzYRxBeWh37tR07Tiph6ExJwEMbIJvBzIjbpKkwXYDFb27CdzA5wVKO
UIaLOlNdyEgsSBbn43/n4jYLeUWH6TvkPk81Q8gn9qEuyy5GkMKvkl3WgNveCuYoLer9Cz8NqQDj
QZPqLsh+6QTYYyARDglwXaPN9bauMj3HWTi6dtndXd068a7MfckT5YZsdZ6m9BRKglqk3UAc5hDi
ycF0ZRqcgG1EIgc0xQTvfcGHhCxEir4TCLY44bMWRbdz/0rgkhiuvEg7ZEYoy7fpBP5oDcWMdPMG
2/kpmtd9udtk3AZL37nma1SqJ75KnsH/LYBi07MxcNSX/n3MM2keiEZyfANkXTDTH07Sc4JZTuy8
d6PCF7L2PkPoqASAABAjIJuMB8Nbr1fINqJo/Se1Lbo9CB81K2gZEoTzwGHRYrncQY9dMXGPu4NB
fWyeClHQNgVvcMhcU9GR2wQDMLonEs3PHpo5z0njiAzJSowQHLgcQegc9rxQ441Ra9GuhFyPQKeE
U8Zj13dBu3R75HvXJITPPdlP81R6i3zdA3QzoO1l4s2xBtzsJjo2GcpdjxagT9DaFPpJAvhmvBJV
ySv3x0YXKLKOwr0qKcMw6NbzSLbJ1H8/8YY6n2rAZSPttsBI60F8PC7dsQOyhKiIP1OOps3eacDM
Ob7wNmQOt8Jrv/Sv+YlfJUQFNiAfwO/UCMK59/SmqTBXMb8Ar3pC8dIjFolWQrXzXv+9dDlEf6/0
tn00iwTrpcoOSa1Se95ecxBIU5SS3QM9hEkfWFuWCDMuh6BfHKwXy35/rVO7g58CxOeZwGUOtee5
qZyF13IPR9+6R6NyxBnLBcqR8qOtLDbopGCCVD5H2u09t2A1d6G6W4zpZgHjVhKI3owDZUiQyUrY
OFHENlxlI57SYknDifJjWdrYeIFY/7GiBc2u0KfUCmNGImSF+p+EFXAQJlL0axmA2WoqbeZJ6jad
eayA6nwUH7q9hQpGNDoJNkEd70t36lBkadcJWAov98FXRR71uiv1f7CiXBnWzwzxegSL0P34bjZa
I113jtSA67OP/ZbOwBW4nnarhSglRQkBRl84wl8bus/xf3E1QpwX38XmkiK9YdDfx0cgiDpj+XM8
p9wHc9UWhnsd6ESQuwcg1nyUWwooeSIP46/XiNNNdKy8+yD62hfWs5lLNFMunNcnvQIAzPhKHD4p
i8Df7GjnPJPqSockJXl0sByI3Cssc/uQ6hd6NtnhXFkRiYGul2T15Jca+zUZFNtBSsq55S2dj+dM
NMbUZxpQhNGhsi8HEdSKOJCr4Y85K40o8vBVsDF2J9G9b6un7CAI7S3agriVLeT+5WEoaDx/WK9E
v9GGVzkvygP2X4XzhDypCq+zltAQsnY+4c4c0VRp+uTaaXgVXPwEq6tQaacMn/3iCR9n+zI8h/vX
B2RbJ2YmOno0uDEzOlOC8o5ur+7GATbWlnzTM/35NiF6qXmCiBo45Q63GQVfsa3WvthVJepJkV2r
LZt7CtziCduFUQWR2FAiDydvZiQi0QP5BOkqnc9k1BpDLovNpxsLVaM/KtbKwF04sGd5HX4FSaME
cTBNVl+NWQOCts5Vu9IObF6uJCBAoTV8hs5VvSlnk9Sh13oBNgFxrwMa4V5vh5brX+VopWol77zo
zC2kp3dFEFD6kFfe7Z8GuB3KwgQ8CF1jKHRKr+zfwDINalWI/qFWnkFlDoiLhoUlqpPl1WSoR6iL
GH997dSK/wbJ2+mw+F1kCr01i+RXLm0jzyJW8FZAsdT+SP7TV5c/qTDzFJEaaqppsaFS+bvYfpBv
1Rwf1d/NdRVcvbNXLFJO2U+tzI6bFUpXySyc+5vMCbWTik1EGvd6REgt2sJPmNdSKANsENDoC47o
13JYj63VWtcFYZjRl8X/1DDg3CC8wwFk+tbthvHI2dxhrmLJYfquyLkcvNkJEutd6d/hF/XDQyEH
RI9UqaZnnBnfVoV8+qufwNDRaDgeHngWivoZcouYJ5/GnJcckaL24ylhriMZnStYh6bF5e4LLfv6
pARTsoi0ayTzxOax9SLC7+Md2bEOakPck9Ipcrf2b/GLTwF40/r7KyO7xyTan8n/mAewQmZBtVtS
W1GrVliaaPS8CYW14gtzP7rYcxMSIvH6F2Z6N7yqYqquatFoShKQo7QH5z5KiGE1tvG1VtyRWO2e
xSEaMYYL1ncIuuLQ/wJWh37zSAmEuCoJ262+5/8ocuZZeWWKtU7FiwL1Tt57a3TJUH0u0Oml8Zsy
RlPxhlzGYkr+R/mfN70IEwJCWPJrXbMOFlnqBh2ZnhadoRGZ0vunECuceUxJ3A+/87yWyz+rnIlv
VMY5LEFJ1/fx1ePiB7JouyqWzPHxiKxFrAnNnJ+Ae/dOKShp6X5J2JMCu3CilplURBiLOgeep8An
scuZr6Rvwag2cdVfBlSW237DysXmwLNMja3geKOpk4IHD5BWsHOPp+mYxK984NI3yIEjR+7tghSB
q00Eg5H0UPy5FEN7iGHlKP0tEnnGmD+tztfO18pENR0yU3RIebVVPihIZw/u3wkSyYOvu/tFSo+4
RfvCQij/1hUfHnayJpkuvHsrbQe3b2MBYSE5qDim8Cok6mb4Aha+bi9w6iDowZqUsnpbYNexYJ0P
1pTwf0BDsAVwGfONKAii5Zb2LZ53F/PTvZZsD3XWKdQd1Jb+S2JVBXzqsy8oKK4UaCZzLYAprx7d
ioLprR4A0oYvTYuoYplkFPsEnPf5PWzpsmKbdupDyhHJW3ptg5g+ZcCgaH7gKkxk95hTusDJxfwk
TXI1qUwMeBHY4GINlPpaEMTjUbEhTxf8H9ADOaI9fsy+nPh4W9xubedH/Fs5wNmd+/E7bfvI09cv
KrbGr90u2Ty3bd/FNrfGglC5Jdxy5/WcCdvG4JR/rbH6njzManscZKUkWQbM2/na3MfJ6uhYxbRk
nzwy6Ci3ocbo2fLKdyMnD9mFqvLUL/hejX6aVtPz8BXspzCk1xbz0V3pLgGYQuWcTAFWaXur6Sim
ILn4ClUbDYIgl+Ua6kwODttcs3Wv4q1w2m3eQtkZXbMzwiC5MCg3UZm/Vn5PKXypdZtATJQMQjJ+
m9ahKl+/tIhwi/YWBWJ97aj6swQNDrhhLfWCgSBnZOciKtfOiVXQpk3TaiurVcG60o7dUUJsg/JO
ZrD7aDqAeyHlHgqy1fhQfnHjhMwmlTqFkuCBBe7SCCiPy5l/BfqTVAnNHJZaYte9Z104soLPp5eP
2MLdTMR3n4YtvUB9fWysn6AJcSlSYjXLliCouMjsZ4vZIXYUDyvJk3JjZp0/AVwTDsEGaTWZHXfX
76ssbdQjrxVUt7JRV1Fv/I/AyPoAm+EjqJcR4QaWSiDYiyBHjEedA+xdXsOUVFRCfvo7V2ToFj9x
uoFxLxwVxCv+UkSCvsg1J3uIaVA9xB06MDNZUOjSVdJGSltNgIUgmqXK1E8YBWH7UONfjQdfd9ze
Uas8Qk759pSXesyJ7bABxjcFWzQLfm7SWfFVUyAO9YCsElBopUs98YggtwEOZyGhiVdoStMgKUH4
M+uyIQ7/B+kXU+nywt+TRYfHVwvJMlcY7w7iGGaT64IQ/J1ByLXzEY+wXoydKH8R5xoEN6+fhkAn
BDvYyLzVRLuHe0RtM0xG37bjkSwCoK/gBVDZCmiqbiWrtLAywZIamjgad5IIoAjwiQtVEJl6G2vG
RcFnrPNhYZz4L7XZlPOzBWB2m60xEgBz+NoLPF+EFW1SFfDm7JtA2G40YVGOEU9OS216tsqKPLg7
hVCGkhq5mAhwKAz3taHQu76HXG4XEDbwEvAUPw7GkU7sQTIpwvjInWfg6hCmNtS3NKCPXJwyf2xf
OIcOsJpciX/vzGmQMsuz0cVNIL0/ILb8YEo3DWR82/Q/j71DpPyAiXFMehlIx756x1+deBFhR9de
88r6i1ohEKP+6UOtJFTPCXmewEWM24gC7daVLf2rbM8yMFnh0siBadWEroZDFvXILPwyA5A3O6v0
RYNMnVeZXcJiU0fZUOGSUPeMfqNoHHeofrAWWSe1BTMrrWaprEw0D6dOdauNS+Qj5hU3Ek/wYkwW
w9MTG/NSwxHugqWomJuAo4xo3y4siJJLS2orHnnDdfgVHlixTXeORm6KjyFFi28429AtDhITBJd6
ho7OKu5wIquopTKLZH6SU2JqPkJfnjqDUhLIN9wLcAIOYQNazEeDuECST32/3eIkP2H8jG29ZGYz
MaScYlUaxQ66WstxKxd0uJptxYlPP653lCMuKrL2uyfy3TANKVp3ONCg3BezEuv86H4CKTqqXfev
uJfGm1LY9kavnFsgcPVqOsgPG+pYSnDSgDb5TH8GQhsVMrj4mZd+piMandppWC7cRh1ZkOjQdoo8
puvCW8IsLmXPpb//0F0cmNDmPh4ePY6ePw5jCpwRV9YWFkZBG3VPtwAF9Q/XhaqapmqnCFLEQI8p
31C1jTGl8BiccqUUOyV0T/L04LS66fVBeIPptNr/TltRPEBMtP6izv8IjXoNNDfbXR2olmeCxXWh
i/VV0SpSRXWbgm8uLtE+6j03OByvgsKViyyg/GEcIqQWyuKb/qCiE8VjzrSXTSQCniFnsYe8NP5G
3WjpgwTjq1jwqE2rTkRiQCJuQJQkiOqqs7HhZsSwIRUmtb29UXITZuuHdNFhEcyn966iNkK1B+az
tkF1E8wrExOD1yvCaMzkhgXcDJwB5YGBexAmA9u1rWCmy4o7v1KycUehzt3ZynDdiJGiTQ9ccAcB
CFo9/t+/PGpudxvMytin9qvLY4ZTR5ocb8YK0TlQogNkmwCdULDbjv3+0umIBaRmuI73hsVJePIV
Ew5b/F1PnG8enwfI5J88C+sSLSiVWaGcUXGcqpCqaUJvlCuyccB4KUYyBxbDkKoPU5O9+YDd2qUX
rq7DWouWNQ2/sbbuZnwXb0dS2pAtOUKLKXV9tZ0duRm7RD50CPWC4LoOLtMr1xY/BLxUaRYyawUZ
N1OK1mWTeDOLkNIq3kGo0vZe3jfFg4URTG70zV9m9d02QvK8AadOYKV9x5CL4w9KBiaGt0FFApFo
bARih4hr0EwjvvnwLVxloeI2zB6hPIjLxJZ4Y+Vzafe8ReKHQE+fLJM+Vdz6KuOOVwbZKEkZWb2V
oWMHeBXi6TPTTugkEJoKMsc9cpnWQASZvrFw10pLA+2Ex6KHkqtM17JUlUdhYwLsRbNbFxVebIVL
9xuaqt7XPosz/jL+mGq9vepUStWdg9Tb/vgKjDGCd9PEexG88XN8F4H/JleGiK2kNxvICt565aK4
F5nThVDCIU9xig8xj6RqF7bN486XcMhy9Q4EzWio7tnJ++B+6Dt2nG9o7QIXqUinw/Bptf8Trr0P
1CfLP8GK12ZkRbCIXglN8JZUAOLNYr0IQ8N82lWY9DKHh5vhZHbyiA+XmBSBFvh7jLd9BIRlqWls
k6cvyFm5pjaztKjiSUwsmv8V58ZKUZunnJBDzVGlCSfL+KKKwsHzzy6uX6Yt7MtsmBdHQuA+JvnR
T8TCWa5tkyavQArnrKg4p3TW3J/NLfLObV/BG3ab/o9miFUprvscggus/f1lks8duXxzSK1l7WOX
tXL52HawYmTLYRAoz9p4xHNdr5xvl2lZwrgUsHPZFoKUWRU2M5GDPzVHW9+/d/EkiaYmW0cp8psT
qWIKDHeGabRfZ5C+YWaJi+sZOThJkeTP5wc53UyijCftkr8iogORtBaRqQh/F60/oCEZZcpqLald
TmSRggFr/rEiTlvAWNKQLTo9rw/CL3fOy/8VLOIkEKCs4Cm0T4UlsyMWjiqTxjGNO1hWbdmXwKid
Qf9VcPA9+MoBB3+UbV4kG4Vj5q/udwQxPdo1DTB620waLaIhjgXQh1fNq/IPwwl+j+x1pklywVPD
5GpNP6VSwnh77OBVHrzoqspo/EYte5u1ocOZVpgVMrH2KdV6svEq3QjvjYBOiPI7+03WpjDvCBMC
g7fEqxRJRVbRCW+z/6AV73spTDKoPRwMUr4BUse5TDp9R3O84vcUnAavmU3TnAFqEPA5qfpGMIZ7
82sRrXP1B9MLxZzcB1hokHhVZPvUR6AexZPxNoKH+k4fVrLB/SqEGM4c/GhMWstItJ6lEiwlF0/6
hwl34r+GChvXsrnab2VYSnQiVWFluNNk5aOFlnWxyKIV6Ue5XRbfRbDa5GlgyiWyFB6FWFt+zXak
YEHwkyt2Sj6D92o30QLK2b6Tvvst54qWJFTbFHXyQJ689qrOvfyuNTQNhQgNQ72CR0IFCNPjbbx/
edpo8660O5Nor4z741H8zxLhoRy+Oy+Pj6wiSYT2aGO2IyukbI9/L9YrOcQlarVf8SxJT0y4EEqz
JyGiDn9elWzueLASC1LwJ6zqhzO659iiOI1pNIyjb9Y34j7FN3y7gW+1YhYtRTzf6ac6+2HL49+m
jafTlgsQl3IdMnYuu4ZOJ1mjW2Bkz+VQQkWz4rwOk8QqyG/Kva61BeB3o60QfLxBcUf7msXfPzzO
LMXygANfL7ccUuCW8s7XmvxCWqY1S+FG7Sqw2q7Ci21SeYnij9352Qx0Xq7Pzkae9RamdwZmt1vV
VEhzFLNaKWGCQk1lhEo7xq6weAOdqb1bVbaIF6jqiFU/D91WIve2tYcRDu9sN1MMeXEfQXmNQvhF
TNq702QME1Z8+Mcai73CUnZujxFlX/1bj6IRmSIbN4wnaJwqifZctM0IdbfQj4lIo2F6+GiU06X2
5ZWpRrurWXyQNjYXourD0IQpl0GNAPXT+bNZVHx1ZiU4JAO5JUYGuiNXZJLqFKf80TUYWGzxWudX
7vGhTge6EziXnpLM78LZrPrHWWpuxlqV6k51bzZE156f6jfIoVZrwxfXbDmLVhtwWQgimBUpWJu+
8bTy4QPx12an4H3sLW4X8NqKk153iR9hoRrmJhJI2ByMgoB+V4dcHatB3TF6Nfmmfb+tlZRRMnzT
t3tx6rhfkLMjgESfBDLKwY0xR76OeaGnjurY6Ne0hznoAJlnpQ2TjMYaK+1DybAbFreqbUEI3gt8
CIOMCiythEMjWNiX5B4iOL70qfZRCJQ2hx5nDoi2ia5oBthlliyso1J2HUA/VaB1UUU1TIoVrhe9
uz56bVwI8X9ajq5cQCbV5Fed90s9RwcXFrmgBN6+bv9h5gruvZcX4E8vt1f0kJhBF+oHi7YmBtaG
aqxOWpeK5ZY7c7OQsbCS8O6ZQkWz7MRakNDDNRvpGMttG5IykwOaUXeSxXfsWDjwaOF2bkDJ0Mp4
Nqt6YiHxUC/1EQGya2hd57sHqGQi1z2z5WbvPs/VSPq0S+qK6S3HCTvDHHBbz2zdj0jEsh+324eW
pTQ0Qg8IGDLfDHNQ0xRQ3zPVA5Eq7NRlrq0wzesDgJqlwDLTFhgZAl84slCSccWZ+jpBPfWknrey
YJ0ihJRxLgaHSTQmFX8jH1dlXLclwsqE3ItlZ7QyiPyhkvbJz/aPJAR7Q/Xf2FV0/DtmsyWTcdbB
msZbQ7iPfICv7P6nQDhVdH8gwKEaGUtoU8BhZLNLLPoeKyMHKhRv9dS6YzJFojbjAN/SuMtEsUhw
Zu76z3exH9WqvnqIPxTmOtiA580Z7io78RgryKqm8bab5tMaN23TIX/15hPG0ov2lLta0NQtnUGW
OLNwgxrAyB9196Y3hIr/ACY400jL9r3RkHxem5dtGTCM2AOumPBZCYow/g+9gOo+mpo5XE16O5rL
WOwhhfvyKMy7H0LSoQPL+lWPCasJ1c1JvGmGC+5kBlSQ6dBJfqmoD+0IbgIVFO6FVPZaF4t4xzQ9
XLEZiq4hJ22cHASx
`pragma protect end_protected
