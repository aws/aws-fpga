// SHA: 43f4f449b937011c34848123159f70bd11b98098
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
ED9zJslU7vets1Xxou96qP07dsNGL3/HWUXHdZUc5Drn7ia2ERH1m6WxUcm+hBehe3ZCd1s4zP46
rM4rGjI19W1DsbRv7vedB8Pyd7Jvq956xeEGKnij1jBkTN5pCkHDaFIgCJddUlabyHsJ40XOKzPP
zCPG6h12nlCIqAmAmrm6RYPx4OXdlfgtneGIwssrJwt32EkMYMiK8IvdUoQOi6RVSU2qzowOVyG/
7/LNzKLzStT82mWyJA92lmzGk9yLPsZ/b6P5G+Ee/sCShaXZpvMC+YIO65B97XkowF3vX+aTdzwE
NB1hhSC5TA/Y1O93HaRKKEb0/BBv/RxHlPmE0g==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
KWnRg1ImeB5NFIbaX04JeMw10iOBKWz/mFdKpwUkInXDTdXau7CfeEW2k5nCWFgyDqyDGgoLf0cp
5nVQ37W9MoZxSMb9qkldHwkip43d1EkcgrCrBg7TOmc92juUhOrl11Z1E7VxanwpaCbO5xvtaRgG
Z6gS2gSAToSprsaRk3o=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
GxacmuYzlmBAGM3F/2aj1xefr5ifWQovzAx9hX4VJ6vqehd8+s7my49bAClqJmkTVaM9jhKo0KLT
TgPlDKzdNZ2/AGTbu4SRV2RFSdQgy2/rGbuL623MoB13rmd88SsDaYg+Rspw9frPfqqEHtGNj3+W
TuwSw0HzcBqk+Mz4q94=

`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
QN1prkvvRkuk7IjhEhfi0Rn3bLrWe3tXnwTwsicX4zP2GaMpBO7+b59cSrkvklU8zw9I1kDNmSbx
6qRjGYGtdw==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3504)
`pragma protect data_block
KEmB3uLa/kQpgB68vSJb/wZaeKpZe1guRoGvKIW3hPKoNqmXkOI1XaR6CNIfBHqIkcPndv/kIG9e
bkbA9cYxcCROEa64bUu5ELsMrDydcM/7qLajX5yiqyKxiR1twXEX+zOstp3/8EtXC/AeXE8VB257
p9epderBGbhQj0Y56knrxXSOAPvqBoGiX79ruVAkYnxdj73antVdilpKrnM52KNuOv2XSe8fc4fJ
hwA+2lmoJ52AXwiuh5K7p+O3H2LnTUpuTaZQEfkdCs2qHLV2MiuREUMO55Oz3YVDlflVjhUhbXxn
50HhROYn+zxdNFzTlUBY5sijGQGpe3+ZvuVn/Aog2JHxaDPiguCplxcO1K712DaaNqCRkWM6ezDh
DgfS8g0iksOv5jUVlFeQQIW8SLnAEzuO2KFHDnfNMpv5hs9uZXwlGjTGbrYGjRx16oKpzWtWcEP0
UMwn7Wr8aErm6kYp+Kn9RwOo8Po94a31Wn3h2mD46eg8Z8N7YYWdcjU78SoYhAWWmL6Y95umFZgj
lLVHfIio5uTFEoEu0qQZpfOwghgJv5n1lsVQniaESubdDx8Z6sWRU5tTMcHGNIL9qJUvtohKR1P+
vI/4tqI8jY9UtGF4tV0n2ybju7PWxU0fvklnvyiJK6LjWniXk/CAgISSFJhU+xG/i8vxo+P3UBlX
yzGdPbiUijmLhKdUv7ZmycAMi0jYL+ppv1dJfZ1nwDtW1MKUO7oxBP1wtOXfi5XVQBNlyvJNLfzf
vyLvaSnXWy4c1XHguMRyS2kaOFA1jQe9ZsjOXwe4S0/Xh2f5T0qxBMeEgejtod1Upek3uNZzamvK
Kmhe+nEfKXderX+2B7IXWjCT76yozadbjoQmVPcUZrHehjofWcAYlLt8YOjz3mbL+2aqyBHNjUEV
hVoQJqw22miaHSxE2iYQWFOhAu5K16bxKAqaVZuVDqy56TqPGypX4CTvhzaxdEuJYMkD0LKwF9IF
ZUGJBn64hA8532nVrGAiXeJU/hdf8l5+crV3J2UO0mF3jREyoIfn6/2AV22uyfkvhAyEVEpthW80
ImWi6EWpi3wntSSbCfPIspeIHd+VDK4/yKQDrSUJa5xYENib2XYoUNY632aVNN6+X7Ejpcueal3J
kOeXFQeI5Sps6W/BMOyuO2523XDLgwp9qxXt1rWW7l50E/TvEibp4c113QorWNzR6BFgj5t74j+N
RbByCaH6CyBDKPrg+SZ147MIOmkD+fEaSK81hHAxR2XSn+EMffHQq42s6K9TmJNbbYOlZqZ77iGA
6fIc2iMpaievR/7ovKLAvUQy5Qh9E723ZSzz4sE/u1g8gKZDtNHe1jfB4rgkfQhUfSvN6sboQfna
fOKehRULCTWd01DnvBBaEmuVdtR7UVqhRUcvH/YAcmtsHxNXMdc3vyg2DlvlOzJI9yYj4jSIUyEZ
dx+Go0R/z9cVXmUEvKSeFZGk8UedJZwy0dQutrg/9i1FDKqKq4dob9vULU+s7xL/KD9KuDOBUY+v
2djNxA/3Ay5FcQplM0u04FngJwz3+O9XJ2xLkYX78q3NaH0wrLa203Rqx7RAyYYpfSi3ODp1eW0Y
sp5gK5bfJSt57hFB+liSJQ1Y7zNxbQNn5KnTs1RRlEIcNi1phueRYVUgY5hTpJVx0eI8SGR/4Epj
MdGqq9Xodlb9KbG37gzkDTyIZnYSIwRxvf5gK/F+OC0IvKLDI/n7UwSmABbWputMpMzJAbfct8nB
PSA6At5bvq4iSPwHl/UrxXHgaHPj9yjtNoC/OKepPH78aI47nisbjF+/SeQQkTe3Vy2C8i4BUToM
8oj+XtPco4uUnhq2qGkyddxfK++hpIwKFzc3wyTlOXT+ApRAI9q1ZtcC37NfLcOfWaGwXBS4d2RZ
+y36SNwKV0u1K7IOGBtleJD0Y9BzuK83Xi1EUqvyFXfZMgQ+ugBnyFTQ72P69Nit+Hsc4uheI8a4
l1hPYjlBjkzARcs3kuXYKzvdMi8oiNiHqBjQDDLgbDCEcwI0K0FvzVkrirvPi03WP8AzRtb+r71v
uiecb5dQfbll6J1dREfIsCjo72qm4PeqkET06pWK/K/pkRHsDxyo53NZXNmskrs8bIMiv48xOFpj
Ztf6STFqMgL+d2YccehuYxNFpSeVsae68t0Opvd29QO7B03ERZGk4/Cy6RvC0znD0KgWP+tXu7l5
XFNDqcJgjbQ8qGP+ov/JrnIwpScqdYHBCIRzUpUQcxI7m74Q/dMfPwBxl2TznzYWfhx0W9azAwo1
WPfk1g4Hzdn+ZGd80NIJnJmTBA/6KLbcEJG8NEcJDSto7w5mWN4t5Qfgo1N++kG+Bql0YD+GPY+u
R3ScmiQ8VKQZ4t/Rg1JWxJZ76J+u35Siqe9jGET5DCI+B7jJMsLpm8dN2qxc9F0bd+BU1cWcF0na
OwSoUVBEJeF6rto3f5Rl9KKIM9lYS2h1uJePZoilfA6JfeNf5Jk9Q4eX7Kjc4uMQw71PfkKfz3Nz
u4H4RbSRCikty8JFRqyz/qkKp/Mc6Nol7B03mewdCe2B6j2J+jogpTg4leLmtbHGuI+uH13M6LGY
7dD/O+gRjF62xNEmI0LJZVrW2ebcE7FwE1jnu+d0nc3oFefOzKXJNJ4Y8PyvF6ECKjAusSqLmQ+/
mw8WNDwNiAwwJ2cFfx70t2ESr2CurCw3kgqrNkv4ctqjV1/lyVxDLF0wQmCn2/xAXM7ok5/XVHz4
7yCGQZj1g66+MuuIZZeD1eUNwijDZDM27lr+dOhxQZDELMG7nsRpgtBkALRW/MHRno3qWbLg4BeB
ttqkvF+vjFTRAX7IukspJXxDBXcSqGODVyx4Q/UDcRiGqjdi1/YenX6+6e/7UFb8a4WhzccWVEkw
cqp/CTb24GYy+dmftSqlMJjDhexa3rG34Xi0V04ZKpGZZBzOFs2JxaSUrouwXNpEKc/EHdzUUtey
34gtWyz7MVVoHnlj4ACouzC3FNrHCetsWhuzh7vqTzCKruxir3SIv4jiPP0A0LLLHiKvYtkuOFUj
3Oj4h4tZW5hoNyNJcIZTB9DRzQbqmvqF2DyOjpPnHX5GwtFIHDB01ACavTFyUADoozpdRd1+hd6X
pq+gtNkwEWcbwB4+boD7HuIJ3GyVV2fI/oC3KsdPI6N3AuWJq6B3KTOlyC1sN9Cnj8A5QSHHKoj5
SkiukB7Zc/8yd+Kt7jm4un7yooJ5OT0CBVhndiemjqWDcQ9lniFIGT9qmK2Pd29i7lAb7cmwn3Y+
oSnRv4f4cXXFgywxEEuDJ9dsmzbkLdMcnBmy89jSHcaP5Y6VefEBAA07K2vXvwm45jGZVA3R4WBh
5O1oy+X3+nzeXRk0tMQT8vUJZc6+3kSeYsNXWdBwjRHCthhoA6a1fnmNp7us59wbXWdB2mCnxLiR
2D0YSAUCfaQ/zb1QI9fj/egYe2RhR+lQ8q/aj4mAVV1zS5mmVtjSbjlKP52P9U6SYrtVe/WyDqlo
+VRJCBPZmDnxA1WWNPVC39utztgG1n8aQ9sp6YRwxVHHEKEbtYcFQ+9UCCY9ThUF2oNwW/SORVKF
SARFQ3NTclqbNTGIno2Ho/qRcbdmZxxQOnQ8LfoOq0TQnyJHEXJyB5MnLcZkPvPudIMVSEu76bqo
dosEeTpBwwumVtblXa7raFTgqPJX0ysqViRXAh/1PfQBT+sDQ1xmGA3Y1sCuTB2jEaS6RWjBIMZ6
kWxqncHFgyirSeXIGFvL7juq4XhHH6f+BW8Cmujf4tC4AX9Y4VFCst8/qDctgvGQDrCoBkTys48X
EFNmQIuMy5yXJwSPgVr5tV/131eCwZIPgC3reCdxCNfuCkhHMDpqU/ALPIDSPzxRIa/lM8pQhku+
DKQcRnXjDvEsXNJkZuHOkvjrJHgD+5eq0zGQ2Zf2cFDCf7FX420tberDqDM6uWskFORTaw85bXND
L506+qfJGwtHJOJQsLNhkXzUV2ZlK9IZ1ovhYHdtpacAdg1MgVkEdfFpCQjmgbQTtw8Jl/bRlKJK
YoEh96Af76aAvN9QazxsyS1wd/ZXc5JvIfdm1tMVdVDPt4ueiJ0OvC1kEsjRSsQBdjXejvETaX/2
N6dOSKC3chdyzUL+6Dzilz/cBW/s/QnLtczP713hmWcw9QiiLPBmsEIEnmyTEK71YLh4rpmEdPNX
7zwiXdK+PXsAxhh6u3It7wZhtY+1JzEpgxf6ucdAi8jD5WErdmczNFXhqMlZndr8rqKSitqtqNB8
DxZxC/4h4Fjy6eATmBT2WG1IpDxliUr758nQdVefQ4+dLXdI58VGKEdmZ3XSmbp7weJBbbkySpfr
SIJFTrsa+LZcSk2nNzxJWHlItOwC9Erk7QFNVKkuBMSftMYGhPboUk+Gxz8j9/CdW6JzMkQnkaNS
WjqqaLTp+cUm+F2r7NpYD1yOwWIyMiL3MJuGBrxo6b54jMA3XabFexikv1c0vyIm7QvAciosJQNU
o5Iyueoopa/aSqfwDq46j0yShUUoKUakn27XudzaPjaUCdApigucIK7ulG0wCoMT7giJsS457nJB
3dpf1Dm4Xc1TckrK+M4wqb2QtxL2ZAHot9oPnffZxbg+6/Y1rJm0ZZDtTsNTFoYdlmfuzk+cfcvx
0XmwGrTSNFPxozZwPeFpUWythTjk0wjlzQX6
`pragma protect end_protected
