// Amazon FPGA Hardware Development Kit
//
// Copyright 2016 Amazon.com, Inc. or its affiliates. All Rights Reserved.
//
// Licensed under the Amazon Software License (the "License"). You may not use
// this file except in compliance with the License. A copy of the License is
// located at
//
//    http://aws.amazon.com/asl/
//
// or in the "license" file accompanying this file. This file is distributed on
// an "AS IS" BASIS, WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, express or
// implied. See the License for the specific language governing permissions and
// limitations under the License.
// Restricted NDA Material
// =============================================================================

`ifdef ECC_DIRECT_EN
 `ifndef ECC_ADDR_HI
  `define ECC_ADDR_HI 5000
 `endif
 `ifndef ECC_ADDR_LO
  `define ECC_ADDR_LO 4000
 `endif
`endif

`ifdef RND_ECC_EN
 `ifndef RND_ECC_WEIGHT
   `define RND_ECC_WEIGHT 50
 `endif
`endif

module sh_ddr #( parameter DDR_A_PRESENT = 1,
                 parameter DDR_B_PRESENT = 1,
                 parameter DDR_D_PRESENT = 1,

                 //NOTE TO CL DEVELOPERS:
                 // The below two parameters should not be changed.
                 // Changing these parameters will cause place errors for DDR_A and DDR_D pins.
                 // When set to 1, they will ensure that DDR_A/D IO buffers are correctly instanced
                 parameter DDR_A_IO = 1,
                 parameter DDR_D_IO = 1

)
   (

   //---------------------------
   // Main clock/reset
   //---------------------------
   input clk,
   input rst_n,

   input stat_clk,                           //Stats interface clock
   input stat_rst_n,

   //--------------------------
   // DDR Physical Interface
   //--------------------------

// ------------------- DDR4 x72 RDIMM 2100 Interface A ----------------------------------
    input                CLK_300M_DIMM0_DP,
    input                CLK_300M_DIMM0_DN,
    output logic         M_A_ACT_N,
    output logic[16:0]   M_A_MA,
    output logic[1:0]    M_A_BA,
    output logic[1:0]    M_A_BG,
    output logic[0:0]    M_A_CKE,
    output logic[0:0]    M_A_ODT,
    output logic[0:0]    M_A_CS_N,
    output logic[0:0]    M_A_CLK_DN,
    output logic[0:0]    M_A_CLK_DP,
    output logic         M_A_PAR,
    inout  [63:0]        M_A_DQ,
    inout  [7:0]         M_A_ECC,
    inout  [17:0]        M_A_DQS_DP,
    inout  [17:0]        M_A_DQS_DN,
    output logic cl_RST_DIMM_A_N,

// ------------------- DDR4 x72 RDIMM 2100 Interface B ----------------------------------
    input                CLK_300M_DIMM1_DP,
    input                CLK_300M_DIMM1_DN,
    output logic         M_B_ACT_N,
    output logic[16:0]   M_B_MA,
    output logic[1:0]    M_B_BA,
    output logic[1:0]    M_B_BG,
    output logic[0:0]    M_B_CKE,
    output logic[0:0]    M_B_ODT,
    output logic[0:0]    M_B_CS_N,
    output logic[0:0]    M_B_CLK_DN,
    output logic[0:0]    M_B_CLK_DP,
    output logic         M_B_PAR,
    inout  [63:0]        M_B_DQ,
    inout  [7:0]         M_B_ECC,
    inout  [17:0]        M_B_DQS_DP,
    inout  [17:0]        M_B_DQS_DN,
    output logic cl_RST_DIMM_B_N,

// ------------------- DDR4 x72 RDIMM 2100 Interface D ----------------------------------
    input                CLK_300M_DIMM3_DP,
    input                CLK_300M_DIMM3_DN,
    output logic         M_D_ACT_N,
    output logic[16:0]   M_D_MA,
    output logic[1:0]    M_D_BA,
    output logic[1:0]    M_D_BG,
    output logic[0:0]    M_D_CKE,
    output logic[0:0]    M_D_ODT,
    output logic[0:0]    M_D_CS_N,
    output logic[0:0]    M_D_CLK_DN,
    output logic[0:0]    M_D_CLK_DP,
    output logic         M_D_PAR,
    inout  [63:0]        M_D_DQ,
    inout  [7:0]         M_D_ECC,
    inout  [17:0]        M_D_DQS_DP,
    inout  [17:0]        M_D_DQS_DN,
    output logic cl_RST_DIMM_D_N,


   //------------------------------------------------------
   // DDR-4 Interface from CL (AXI-4)
   //------------------------------------------------------
   input[15:0] cl_sh_ddr_awid[2:0],
   input[63:0] cl_sh_ddr_awaddr[2:0],
   input[7:0] cl_sh_ddr_awlen[2:0],
   input[2:0] cl_sh_ddr_awsize[2:0],
   input[1:0] cl_sh_ddr_awburst[2:0],        //Note only INCR/WRAP supported.  If un-supported mode on this signal, will default to INCR
   input      cl_sh_ddr_awuser[2:0],
   input cl_sh_ddr_awvalid[2:0],
   output logic[2:0] sh_cl_ddr_awready,

   input[15:0] cl_sh_ddr_wid[2:0],
   input[511:0] cl_sh_ddr_wdata[2:0],
   input[63:0] cl_sh_ddr_wstrb[2:0],
   input[2:0] cl_sh_ddr_wlast,
   input[2:0] cl_sh_ddr_wvalid,
   output logic[2:0] sh_cl_ddr_wready,

   output logic[15:0] sh_cl_ddr_bid[2:0],
   output logic[1:0] sh_cl_ddr_bresp[2:0],
   output logic[2:0] sh_cl_ddr_bvalid,
   input[2:0] cl_sh_ddr_bready,

   input[15:0] cl_sh_ddr_arid[2:0],
   input[63:0] cl_sh_ddr_araddr[2:0],
   input[7:0] cl_sh_ddr_arlen[2:0],
   input[2:0] cl_sh_ddr_arsize[2:0],
   input      cl_sh_ddr_aruser[2:0],
   input[1:0] cl_sh_ddr_arburst[2:0],     //Note only INCR/WRAP supported.  If un-supported mode on this signal, will default to INCR
   input[2:0] cl_sh_ddr_arvalid,
   output logic[2:0] sh_cl_ddr_arready,

   output logic[15:0] sh_cl_ddr_rid[2:0],
   output logic[511:0] sh_cl_ddr_rdata[2:0],
   output logic[1:0] sh_cl_ddr_rresp[2:0],
   output logic[2:0] sh_cl_ddr_rlast,
   output logic[2:0] sh_cl_ddr_rvalid,
   input[2:0] cl_sh_ddr_rready,

   output logic[2:0] sh_cl_ddr_is_ready,

   input[7:0] sh_ddr_stat_addr0,
   input sh_ddr_stat_wr0,
   input sh_ddr_stat_rd0,
   input[31:0] sh_ddr_stat_wdata0,

   output logic ddr_sh_stat_ack0,
   output logic[31:0] ddr_sh_stat_rdata0,
   output logic[7:0] ddr_sh_stat_int0,

   input[7:0] sh_ddr_stat_addr1,
   input sh_ddr_stat_wr1,
   input sh_ddr_stat_rd1,
   input[31:0] sh_ddr_stat_wdata1,

   output logic ddr_sh_stat_ack1,
   output logic[31:0] ddr_sh_stat_rdata1,
   output logic[7:0] ddr_sh_stat_int1,

   input[7:0] sh_ddr_stat_addr2,
   input sh_ddr_stat_wr2,
   input sh_ddr_stat_rd2,
   input[31:0] sh_ddr_stat_wdata2,

   output logic ddr_sh_stat_ack2,
   output logic[31:0] ddr_sh_stat_rdata2,
   output logic[7:0] ddr_sh_stat_int2



   );

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2020.1"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
S1nfxyo6VkjEyNmkUIW/n+NsteolI37Zh2912x01jnhIT5hQMQ3pZd60zvEUaeqwueyGdVJDxCxY
QTgnmNCP20I9AaWRyqtC52m7YXFRdvO72PYcxUdidBNVUoK2B4R4jEIcV9S+ZkmVX8i6C0w7GJNc
7VmWm1jW1RBBI1Kjt86xOwel1QkL1K37niJv0NBLxxk9XLFLmr6upLBSTjM9RsBIxWRC6AOzmH74
/pD/KApA71M1oO6eumHOCzDYMNqnhfUk5G4LJ+o+T6KnIo6UqH10xUx1QZa6wkhbzcAvUSWwIQHb
nFvn6QVPBbqsdxvAuaC7SRam9HpXVE8zE4FQTA==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
q8Mfn8DigAeTt9xIyuOacaf4k1h/M00961hget4VxBsr8+uxdx9RFpeBQBEbapjqiFMiF4ItKBY/
0KR564BStJiTnwPRprXpXkcB4GCMFlFD+IluF4alWFDVo57CA+XfRhoTPPD2pcvaIL2FPCxJpczk
vJ1tq3qz9p9eItypHBs=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
L8IWnxuT2pr9RequGy/0R9p22yuf627FbyJHHV5JuRCa8injC8lR4HeWv/GZi91T72GCapPFI4JB
tSfR9AOhKXMlNZRW06k5BVmHtxkNM9VlCW7lIS9bVRNGweQgFGIlpUjkpPnn/1k6HB/1Ok6YXu4G
NPCG59tU33gjQsxP9L0=

`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
n7ztbgP0tByYOb0u5aABK1Y86n65ueuTLZTOk+tQJWYuYBBOKPiaoKisi7VkeiJeERCfRjRlpAa6
wQfsY8CWeA==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 75568)
`pragma protect data_block
G0VI4zv//fiz0RkMtPrDU0kQVxYb5KBJdpedicaf6pW/9xkPV4XBmvzq3GbwJ0L8PYljqwL1v2RF
2oD1OUaPrE2h1BZ0MxqsU6mzUcb7UcDSOfzIzkXCzaSNOO5h1COKG5MsVj1ulsQQZdcEzUQs1PR4
F+mmgRmist1kUF7icvrz70lE+oAWxinf5C4OC8RtXfMuAGJ4iG9J3XBARhIwgWt8MDntzbGAuCo+
Z+sxowbi2lJsub1dIkbvEWxvMVfbDvrZ1TKj3/tHi4JrAJlYqoCWBfw5gmsiU/ZyRgYZ7XE95VFr
3Lz9I9fa+kRh0oz3nWh9R1ZmartZm9PPD4aSouk70RnMCERNpIft8Wsdh39gOeYhwsMg7xr++/WN
9bObWxDo6YuS/BmrY6li3GO6uaMZefEO0/uSEJE+j4+8Jw9nF/bLJY4d+hHKjxxkWaZxmc7gNhwY
X6d8PcBmC1y3+b0FT+7ZG76RDxFLpP+OgBlN5ADnc+nnigd21QSTT9Ns+51ltwiSgVyFDgTJgDse
alaIDW/ulmT7r+54Nkmid8K/J0rV0YrvhBcznyBKp3fDX5JT3M2IJ7oykuOsxL1wde9UklkaCmA7
cTT2NReBJC6vZq0+Oa8drj9l2M81EMSK9vRO8jvb1UF1YwT5xRSgxGdaSPW0JGmXgcxs4nX/j/sw
h09HPnHHmA7mU+1K4AAdmdpLFM9TAFsg/owdwa+qZc/d1U7WW/YRmIHtoom2tOfONRyoyovGseCW
KBzkMIkZYlFpcMwbQq/pcoPSumGzlAgiFYLr+OKpJdVfLnlhj8XC4zFQCpy0HxeNf+QD89j6k/Oa
hpP41rtM19wtaKoQTyT9on9diGymyzgppCWx1ufgDN5k1u3ss8xhK4mBbnqk0z/NgE8+vNM8gqOD
/P/RkWtH+mc5JdwkyFDDVLcI2g9IdOO8fq+ocpjWLbwh/FmETATZxpJPnAneMXGZuWMJcPpjjmoP
xBIYW46ct+0aQjBQhtf21ngLIYk8d8gMKHjJlbLjyk06zMx80hTLfoMjikV0pPW1nOrCsBvIK4kD
9u3jcP7lJQ5CcWtp4v4sK5KNWNjVKGTmXJCMWzXmoTpwgWdWh/G7kV5QZe83szyVUL/xZCUUI7sh
vq8aObha4vuFtRpv1PnC1uFSxoSKKyIjnBym90b+KNRWW8xvVRNZUR6o9/2wpTWgW07RgI2JIGfi
m5KRAfTRUkqjGRZgvPjnp8CbjluLhb2LzxWI5lZMTZsNFaKi2IRWYC2+Juqedm7wziji1u5n1vzh
L7zOADia3ClHrgQIms2wqtgGP16DhKJqt6Nt30I1gJXbbPKCvfLPStkJ2D/pqeDdHesBO6Fe6sHc
VUCgICip0SKIip/DAu68SCmdtX2UhAoZAv4VJjKP9lWA0oo7adq3ayJstoMRNpVM7j8OSuB0WQ84
dSWNnhX8GIsKKGoG0hhT/aMQfp3Sh2xRI2YsObgh4USywMHfjv7LkHqOa8KCi/PnbFWVx0fSat8l
5v837T3bCPUXdtW/C9x6pBwfgZR07kkrPxVLSEv0vmfBLVcSh31OBFKoyJKStGhyhAUAwQV+Wapc
94eWw2nn2QjSkQQUnvBiM8FEzbKI3174WWX20kR/SMVQkc7QBnfT631DHjLFxvRtU7U3W/zaMcG6
CF8SBo+M4UEnpqu3+g5CZPl/IW+KeKVx7W6SWebUPlPl517jgHlcB9EROL3JWL0Tysgy2X1Q3ldD
iOMv+9aA3YFIzhGcEdGCNzzw2YyBAmYPT1OXn4dkqd7roC5iI7bL0dU+E8Zmh/6B2gqBiEUVexRW
uWgm4+Lu7Ioi0SkaUSEeLZH+3Zd4MLRxts8i90m+26hCVipbvdwfLpJAobv2qc3eUm74GE0zcOQb
pxuklAeAXPlgx+yOE0aBUm6RBiK16z+meBmKOU5QKMbZK24ewVSZIESzNIZMY/blWVLBHg6U0NHq
71lzyNvmSPNtiHwGT4CEpRAAIh1M2xnXc30Y4yuV6dWoBV0Zhhed5gpEUm1uIwDfTJ1UWcYaCeF5
x2uv/662RGj46fEKsQuDB60Gkv4WBEaYbZHz6JLeoX1c/Gp/jU6FliFcHn7Zh9pGlWNwdUe392Jy
829kK1oGdsD9Qw8HFzh8ISSeqidWxQZ+UjvRmQiVxiEj2M6mfV3mioQJalYkAFiUgy5WWGz1j3GZ
NIm0QDzjS1GUnb7C3NZAnufkOoVMFiQWL1O9//vimbkFxeR6PzllQZW1x6Ot+KWSCorrgsF0FJ/R
V6L8dKLjilknfQJyA8gdcPE5/caLKDDzYd/1Ci0bjJ1JxG2klSf1pxLGF+KVaa9AmwVhvWUCrbVA
QxY6Gsp+fIVDhQ81KtxfmS21a8nsK9QRfX1T1BsOJy4sIZvKmIpJN+dC3h+56IIx4hHb7DVtWRDL
O7N6UIY/I7uY17GlURG2vg+wSEmivL8eorkpJJZOE83xDgyjG3z/n6i5JL5uqJovCVesJ87lHqZT
RxhqCdYWeOqZWxWa5zNTOo+CYla4ulTdiB2S07UKLElZWm+iW/bJn4mGzcmZNJiACjp/CUc2FqZm
9dQuHrIb2p6P7kni+I+D3LoMtc4Ho6uz4s4AWZsnoVUApVcuNKoCtznpx0VJzCJRVImQCNLH6ORE
lLbfsNTeQPj6gA4Ew5iQtk1y+iEOpyFOD0cuRkUQ6II6fhnJbZshqDTS4GjjOj6XIoNWVmS7hlM3
W6FNpLvMmPSF2AaUvVauNSUmivURi+fq+3uwgEKT1WT00BzLkb0B4v88I6+t8NIRhH5lYOJbz9CG
bhhO0O0O0zyL1KtaViBOhmlXsZ9nm0Mvns2JMbjaUXtbg20G4Ees5m4npoA34sFhJ2htwEBY+GnM
mVzuzMKYE6tjMAEfzSlrSK4M/Te6YT6Yz0QX1vfZ6kaKqSNXnlII6Ru/z9Y2Uju5+LkOiwGxKijj
lDqRrtWLNDbWq4V2t5PGfB0uXMH54cZSlYBXGt86gvp79zli4TLPSxjNKagnfQDBg1IhNXlQQjGN
Vk53Z3L4HMnjHTb5Iss3IP1PS5G9Hpx9iDgCceHidJGFjGto5Mq8k/D61oMyUznsshPZptCIEO8c
DKPwbmllOLtVL9aPURcHuAZnGRm/Y243zSIYJULB0e2U8zFpV2JX0Fv1Uk0wxRcVhi/29Lo6zkk0
WKyhzMohHUPGNaOmnXLO3B20x+Qbn2VU7kRk7fZM2hJrav/AoENoHsR10EER5xm2K0oRjb8BpqdB
qCf/Nu5rJm0usmD4bKanzc3n/OqIZCVnfPylmDIf6exzmhCcaxb8pDGwSS+M9HhgP6RZmV4O2Qii
crnfTKwrfOOEYMleMtN18aEvNQZp0qTukEPuqoyFUAfytv+bFR/H+6hJsCfz0ykWfj/pZHkzanDq
11WFfgibUPjfqZ0uujWXVHCSJHgiYvmWFKhgYpt7YCnyT97v+xOuQtYulI4s3tS5z49jFu2l1+JR
Zv4w7b8kClpu1RUX+gF+sM219LKb8+uvLOkrxgxz5cMLynpoT9Vt+vVFdfJ7a4py637Jt/jLUvJ5
GzMJ1vfTxk2ub9W32hOELixnx8EIRxuNN5+QsI+NsJhHqQottLZb8DFGocog1PDLPgJ9EGirsJAL
2NHA7HFHuYh/FFgSBDNhssMyfwxzTVtQBX/buX9AUEV9NyKm39TJ5J8tT7/aozHvBpnrCNsuFc2J
8Mhi6ShFaMUrmBeMk3fDH1LEnsr5L7TKscVczyphAk2wSxE5aWDhPdrBO7r6JLz4lzJughH+fNY2
yJ6NyXTja0wdpXBscT7KczyqVJMwXVAki03O2mwYfcWFnjp3Zlx/WNQmSRBrV3Mq3hjA6G0+sm8+
JAlJgOmwTDRbDjGqiO+RhNGkNDZmPWn2mombYsgfH4MTdQsjQLuSIq1tnwfUJIAxuqLE7Pwh1KiZ
K3+mLwtviiHc2D7chGeKGzkr6AbV33IKuR7clebwPh6rHBIJK21v7HTQknJiQdg/KdpR2SJFex9D
6bNvJJjrKIiX7xETTtaIzS9S9+rj2jB3elESvekJyIZYKDL7qOBoQ0YuwjNc7vW/yj73cT71xWE0
PYutQMYYgAWtf2kBdpdDcwIHP80tKtaRlD4felHT4pZDbV2HeEPvqwouDABSbdcQPyJXnGrcyW68
XWxo+dtv1mNw8Je87upyKGlMYaha34N0b1O8Z7rgiUR2fSS7roy6AHkLdyvvDWVxv1WwYGUyCpAm
+sa1e8yOwXU3TdHoavCDy5V19eWmhQpAAoybcWkjqO8sjp0uJrFWjSZowL5IutJJIbPjqFe9SC8A
M5M1bTHaJZWXf0dpm8qDwY0Vas4gmNux+SaBT83mQpZBg/qcc4nwrxWY7sO/+HIDM9iuEftV/Hkr
/yp9Fg40QcEBpY3pVBxTIkiflgfnt4LdNklccjUCVjMG6zqfr1X1QY/Jz8MVA+yLAN771eHtsZf8
Ff+CCUFBvhrUXQvJFWL2FX+Qf5cIZFIDn/8nBh3+MS78ABSqXjJ8DxhiOJtc9Rq/wuPhVOyu8zr4
TirRrNpk+xACKj1xY8PMVrXNwrrNsV2JaCLnBrapd/OkdWyO6csNOm+WsLWtRrPeBE9gGx7/EJcw
iXjbvO46ATjn4aij+xNHGN3j8pDYvjFGRfPu48lYADK/7ARhZ+2C7tV9SgLY1ert2RjKGbS2KsCE
/EvmB28Pqi9PDffAQxymGSUC+kdXLEfuM9kkeC84ZJFiRo2NP2UJxBjBJk6boZXGlZGmqFaU0MUN
uasPSvdfxt8wYHwW3yp7Vd6ZPQvpu4JmUQGdT4LNkgivh3kakNQjbkt6GFI8msDN8rnkxWIR+KUW
dyTZO53AR8T/MKlReazvUMtlbH/1n8fUjQVWsXY5d6He6Hh25dyAErm+RvddKcA/fl+u4OpjuYmh
RRAVukEM7YX/gdrI4xpAQSV6fcyaHZPIkJFIEelJ7d3N/RztCrYSrMWWkdiKL4+Hnz91bX9n+fAc
Pp3DfIr3sBX85I3RVzkhIs8O2cAPBZg0GFERt/TrldQA+zV+Rl+Ncr1Quxp4PyChVHz075/Rr+Ac
II1+69nDuglng4oSIPtd60E/W7ys9pTIoHYSSQoL7y8wMgfkfWdjGpCsSu228hr3K842g5aGqy2S
Z+8pGKd6ggH4cp4e8hi/VdQVWSRENGaoj1Jc1T7Sg/tNjO9HUbVNAu+P1XM9xbWONhvh9DznP/Iu
Rwt8I+tAirP1iRP93yMq0JiyFp8crMTqe6KCbUtSrgcDbfCGj4RPgfsji7WyVrNk/ONpTjh9IH/d
jQDfRVXvS6cVftYXPLATrmOLF7frXZIz0REGQp7XxBsDj0//h0AJuI4J+3A8KW2z6K+z3DlO52Fk
ywzeh+e3PuiOXUgJ8FeQopNUvPhqDJdYMVczMqU6QccJHPQLk1hEIlnop7NCh29x0z6vMwTQkQif
73CE3GQOqzVCjgV0uF6YgMdrwkENIyF7cQ/Zyitzets9bhgkYh2RPhT3y+s7CRB8NkAN8LmeVuZm
lxqzr4AUiIfwzVtTXFDhe11IyMUOO5vVZw1pyVrxLHDv9OcvLy+fBrKplEiqRW+hgvtb7PbtQzGM
VINgwYEDt1y9rxrX2vyW0gAERXY8IqmPzDeqS4UyIQ7sxV520LfvihK5oZkSMMkcBwUHWuKhzUKl
YlXbfnZ6NsHcuyDPmKfpfewmHD6ycERUYvqKVbpL4JHamiRISLaTJa42mBRpcM0bx5pnRrmQZ36i
MK9sFy/y6uQrjwE2f2xX1QR4Vj1pC8G8Z99hYGSGy6omnF/ndTGuE8OF5u7hfxFjPxnrfYa6sMa5
UmTeg+Rr5Psq1YNbvkbVHpiGf4SYOo4+z3JG5U0gNazMqyvxjCZOcHFm4Ja0xoFQzpxwa4kJQO/B
My6Scv7myEJNZ/Eq0mdXXPA88/VtGFHoxKnd3YqSfllC5q6t/aS49UdB2ieZ6yvwBnkeonhl3w4b
CifLrmsPlmq39DW6fXZVo9JpSyxMpvBFMhBU/A5XME09C1qFk3GDi+W0CgEFRKxugOH2cv+96iYP
CJvc+pKUfpQ83BUihxLo1WtfzR1dHdL34M80xDpjHCbWRnEZX/ViymtmwVcT65LLMV+whh2EMNfK
ZzGT+1lT9jlkqopMJndp2KuWYEHcd8bUW0bEVPz6XHqkuSTazch2+3dAFHB55icZHnDBfzoYOnNH
wZH4QWEUN20zBYIESxns++r+ElIv6xTHgi3/3ETou8qo+zl9rOOO+F62A6klRUTZdWg90Cl5wN2H
dF1Kf/pqcAuIBK96GWDA+db6lpmXGAcBT/DzthVzsNe06qNmY4DkthW3rcuI3/071muYHd5fetjB
RY7JLg+0pv/bZB7KEQswg/Cr2MTzLjhhDt1iaHLKB5FXSsNuexgfTCxgNRrLsRdN6KjKxnJp+3w6
jzmALLv6EdHCJu8rdX7Pvqy+Zr/SWtiAnraG/NAucPSltjB86KUm8F6KuUyoctmEqTpzlIHGsbRb
3PTG1FMrLHXfqT7nE+Dt3r/hRGRLKwREf03BrPlcMDNG0srPgd9RVJu3oHeGqZlzP80YA0I93n90
5SH1OYX6HpxSyuD1iF8Yok5m+43q2UFhCCobE0SFeVTOZlYVj8fbpbaEW4NE0LaU24dvl2PKb+8T
c+NT7Ps7mbPX+lTCotYBJ+CKGMXd3aKC8AbTZOaptdYe+9VaH03oCTgS+ll5l8e7CsClDksbt4QN
oLkH35Cqyw8XTLCknFf2uXT4XlKH62WMTlZcrw8nw39Xy5HcTHA52Twv8cwHuvx8WZY9qOwyzQLF
AqPdTXFBLejfpXMC4RdhY012DgPgF/APGEpR3IOHGLzTiil/DE7qvisYxrM9Koppctgp+TK3q0r5
zyqwGEM3luQmbL5ZnX/CdUDSRsE4lw1eKVKrMzPf0Wu9Vg3xGFOpg5Yx5owkqnQFLPEhJ1xV5II3
9NEu6UkkttYg4focAevIwhi5hQivTUszTmwAASWVsYAHAlAyDrqy2v97ZxnycXq3lmH1s/NtdQbE
2T2nFHOJYGolSUHf6eKiHAVfMczqGA8/D7I490q+XVWF3bYDTpK0dXt0dNhwNSgqDo+Uyq1whzrW
znAAxCYyJCFqilmKVE+IZEGyNev1mr3dVrhctfT9L0RDxv+o9WvJHyUJHllvQN+8+EBJTgFM9rjq
JLtU6kV+v5D+0gV05dwe6UveQADK4QKFdbTQ//AMFJMXWL8wChXkdXUdf5tMeofNS4RutYJPUfAP
5pj2+cmKpBjrZln8lxbW8Gd/tIMOMUM4JpClD3q++sf8kkPjr2oVwv02YZSzQV/LlR3nle1HMtP1
FiYte7bowxEbqAOBgr/COXJBj16/biqTQA83IyAbBFovVbBvhUDuiyoO6fNJOkj5DIRu5DZ/i0pO
rPTjwrrs3yZWI4tu+XwKXrCdi9uyiTh1Xl3OQMopDYxExRovt+qJPh7dk4G+6QYONaMO5Y/DO2ki
WZzSQy7c7LhUapod47C9OA9rj6pZHskFyfxNT3maSxbSrGZQnS5Qix21Jx6KGZRCvudtgkrx9ry/
V8hW8L8GjP69Txoa5z5w415hBReOpwJsZutIRCRIv7LZmoX6V+8EdTGhjN2edK8zuwjytEkPXTVk
tjxAndLrto8dlSdpV4iP5zZT630yIFycuxGKYpd5D5qfppbxOZDUj4MatOg7ulT3hwJx4rjmU2Xp
u1GxueqZZFku50C52ZLggBxp1kGZQaSKAIGikushsljUV1b3FO5jxlVnRqbWKK7RR98pdR377ZFW
kQUxdK0KcDRTxwmHEiQZbcVvZ4Y0bkQP1HYC7klkiEEl4yCa4ZEZUoAAvFXVcY0BRCBkSC9AkKwF
BnR8NA22ml0snMKnO3V1ag31lCYa9iHbw8oxXtFTXPbR22qzn8GWB1f7So8whn9JFk1j8Vkr0Ov5
Axukmx/5y+vDgJtLQdwOPqOFneqsjaxsn6JhTVeVEXhUytTAS5ixeASkJ+028rluoed5fQMZk7R6
D/LCdZp4O4VVE8sbaNy/Fz3CLpwfuMfaQcmis4gapKK9SXsc0qbomxre1QZ9AP7NEUPtQ438FRZ8
q6oTw1lPkOPDSMcd1CvKBGHCIT9urIB5YV3L/RGtXhHZRAMmZDs+bnhIqQmDVl42RTVXUUHFtFvP
sikL82qiWc/4GC41h8hswoO4+41MDyFOto4pNRVmxgvz9jWqZvSz2KvXSGvERnAR08XnLtndRVDh
7CbQwGcF+hJG+EH6sZJIVEyC3GENEP6+S8Mn15zl9dtRT5CuYoKUp5W6A2HcTaBFY7JZtrmIgfqD
gD5och9HsN4zmLkTZfC2I/u9iNlSMNEDfMXp2agDhpL0BMgLNoqoCelXoII+X00zBWC2SwVGHqjW
FLQxR+kaLheGHCAWu/uA2SB2X6HTH9zhwOVhp60e3Ujt3Xz1ZRmVQaMxdzgE8gr9GAGDVeYeaYJT
xYysJs3fQnFqMG3lkzgW9rkVnFs0+S/mH+/oXYNQLIQ06SY/EJQjyCOnrxMfVGJoNLL4AvYNscv7
RfH0rnbOHDXK8xzq2FcNsiY7JZ5gb+Z1pgjc1DO/5ajqwxgiwQkCh8FrZ2ZAkGXi2g4F9nhmOybE
LdEjF6aTAmtHIpgdKFdg2A+Vg9fv8iAs3u1kkNc/gHGaDvcGUSvoamgSo6k14Zr3r3zOEnGjr41V
4AHHM/2xLPwPk4ZU1aH1g7D2oXmVlTdTFZZ6KYfYIhkMlq5c/0IDNxI5Y3vkD5nxPlpXDwb8kxYJ
Tf9G3+jl1hoQLJTeQDAVXD57J2Q54jQQsQdV13mQ87les4Db49eOLB50y8UOr1uI8zjpYnTkA6QW
ftwg5Jmp+JvGgh885oNpacJtPRSLT+Vyzi1Y05Bo8yZByGaWVGeGyvh2SLClWKzQclGBY+fEDeqX
F10wNbRfNVDYCURKDuAVAioFQDpxXFfH6uZmx+Ke/uI3QEoALYnoKLZ5tWe6J0WghWNLzoyUn14h
JzsImcX1zZ8xlg60pg8H7XSgKcAW1VTOdxpuu8BoxpEMWIZgRUoCNZpxfgNAkMI+shEeChR6cxy+
utiIVo911awT+y5L5MQJqrjeDJy969uUjiCcCxf2GuUGc1N/CcX3ajscIy750yq0uy5U3B47Vjtj
Z8lg4JR+j/nZ/i798liooX7UaG7ReJg9at54vN3fOf5vTID9OjCf9AGSGJEYnaTrndPtGwehPSLy
tk/CWRR9AM3RSCBOA1kbRoOisNs5ZETX/4kHpnLun4tHjj9FupB/eV19KdTS3XQSp/ix1Vd7x3yo
/LdN9wxYLYO0aGMJMTZiuxxjGRr1rMFaJOlazArtNhmgFnVVbzWeYOTLYqkCez4M3LnzPVLX/bby
3rvFlRCDR8jyt/uvdgno0nhGcF0/y0BuQRmwBGArUuSZXkYmKhLg+dLeseLKywaxXvvR/0DYO6nq
OK7JMyZ4ifD4DohDNZGJe/F5fbEgGzw+IgVxGywd8Ds7j78M4okstnmNJyNysni4o2f+hj8kthwT
1RBwWJrTmD7IdI6oLjRIBqSIT0bammtUmA6PW/6Af8QgEC32DercOImd7fExesAtI3MbuVKpLG/b
P7U0Ay3x7mibgzXReAWhaDcYQUgAJoejrR7XCuQ4QagLxcpEn6K5L3Cfu1wt75a9KXHNnz2RwC6x
DZFsZm5pfZySKZvtjITL1VtQYiDBa9uXNlLmVdZMalkYQj7i3awlaJRRweZ2xddDtX1xRGiV8q4S
Nxim8guP/cXtRHak/8Gm483O0BNg2l0GIjMae5OYVNz3XT0rIIcuv2r9GomPRDPuUV4K8jbjaeeL
QIIlr1p5fP9ckznggOgW1gIeKOifE91+v3hmj8EgfAinL07MgCL69/dZooUfEhHA3ePqWvXZ/cJ5
1VcD42vyOBYrLolzrsMQWcqfeN0nwSdPxPWFCjwkdahMlVxf+3U9SV2jttdN8dF1bsC2lViVA7Ug
qWg2YW5ZYQJzn1M7PrK/ypOkiwApYGOwEsAZjXJLxBra53GZ3vrpr2s8vVUVBURgwtftHZ1pMTdK
ethavV/7T6uC3f/isAkOx6DKFDO3+A10O5YK94s+cazCkBl1tvRnH+mfOdBdKXrTOPJDMGguuzSv
dV/xcKGMKMDMl3Da9IabsLem/IxdOeRi/H+l0hn2a54z9YZbT8Bi//XbTwQMGoqgWQm3M9LolIKZ
x4our4dgUDxl/NXcBLhHpb5gpWWVgWunkcZ55LjIdW6+kIuPUYqA3Ov8r5HVGdWmQ/w6MDMA2CVw
I2yncHFtjnOGPjt190FH2PVnFpH+/LrtDZ/Q0M45TdZLAyvBd9HlzwX7xR+OGR8VNSKWj6mX0OV2
o86MdBLU3gFNATJtBNIZUsSe4vMJKYK5ib2Ju6XvCZcy8ZBnkJXz2JRh3zjyJ1IMHVPcBv8Saqxs
yjDs/6kQPis1Eowxo3sJClq6M2YDJ8QDml7NZZIplCmqxFv90lhAs+uJwCLA2qmtQ+BAll8cnUSH
lwUyqA1+twBFCR0V64ULpUOHvhrFH+roePobIHTJjiXEvcb3p+JWn1ULn7scx8BsOUyGjN63Jgg9
Q4GwBji/Yh2yIXYU+s9fh2BRW18xh+gkTcq2YjJY8MD9Edecq+Emtdc5aTFppD+9M9ygWnf/Mibg
JBX2jDfs1ixKIhyOkUpUSVIs0H/nfDmjzy6Ra60QWjDETzFkn6iPOUTFpjnmCnGZ5vBqTsNcH9NR
C31kOfzDkfuV0X09+KeG3UOchcFnQ6o6zFQxD9e4SllRTp9coKDeb1cB0JZvDKOsBkYbE3U55DG3
olSVGLFY0FLuqGorL3O7savdIdSRItzEEBQC4OnqyV8N08vxhUt0TkXj6nhffzZPyC2WzkbpE8w4
LZowXnd5/VwEqskwuWg1cEE6bNKkRe82jmvZ0WfNCwOXgowT8CXpkjM+DMqR+vEHEL7Wun1BGR+i
LDVBVcK3BtiW5m6XUgu7EZQWdt7hvPKn8HZlNNk5FRusyrwhkjtO739x1mec3EqeOBx2V6DZSk3n
at2FZrNfd3Ty/fnjHB+o6EwSBpFbKypNmeZk0eAsVQ+n7TS3FPmkyCOMAEsThjDxfsVOpSkX1B+7
hBYoc1rJTVpL6RSEn6QY5/4ff5ARDIShB3X0vPIZ2Sm04F/Wt68/nq16Y02IaOKW4sfGQAkWjMKa
Og59+tF7pzAJrRcBDUxQdDmr2RNlU6kVWHmc6fy6iBWF9AreVi83PHMmD55/phqdrB7EfyS6gvzG
QtR9Uq+7sNcddba99FgWZdbOOSXoJzHxkpVksVk0d1QmB27jdMvNyaK2lPIORQSNhiHGSHbX9Wz0
+VYztkvlZJbOngs3YiTXXs1pxwF7kPaKFayDfLzOhO4K/d3W43NGXavQrPBUuxPPrFZIKrqm9+94
y0g57vk1DTYvYo9EoYWP99FF8JIoMejGTuPTNfRf5u4ktL0HNkYkYLYoJkjv45EdGWaxh9Ta0yuO
XGlnDnbyPpYPG+NTN1lqsYKR+c2WrQQjVMWnyVpSeQtP1UW5uLHg71WxpbU22FJPJLLkfZN+glpX
1Pn6wAzGn4aa9olnqSDeyh1tb9GcmuAXi1NGFsHzUk/E/DwPvY4wNTrYl1eknVk180zpmyPy4qkZ
JfwGjMMu7b1swwt1hCW6bU7xhd2U5PQ+ylXJtcWKvalvhXpUhpaNQhp0JTayV9maiHrkG9u55MYD
MukpsRXdEvvDojtEVRlbLLWJYws+aaTJGjY0ddXXujYCVkdwr5reYagPhFDzKDYauhXIZ5enfHVm
DIZupmkBbZJWZfWuxEAcXNGEWPZUMDM6l2C0m47RayOjkOAzKhxVHY6s2vw/2nD6XeQaPI/9QrOi
apTh15kaEIuEowOzYeOMfanRBmn+TCx2ue8Y/4UcmBgN3f8S3eWr/A7demNjGYlomQCJML0rCPgr
FeFK5xnjmHxUDRxOFF6n6JXgJdUmX0Sdzozabk63FldTQLRPIOl/8tJAUyUmSedNOdrXuTb71/NF
01aQhf9k85tom2Oyxox1506DQLjOgkkM+NvxUOl6iTNjPe7ENXPHsIQem0pG3b+0wreGAYwoxe0F
UUCBPbfsxsj5qm3kYDGOY0MvFShARvXLq/g5cCwqTy/mMFOGqu0EdEfQHPLg5lsxgpCA4pckkdSo
T2U3E8h5GG5NgvKdMfH7jd2t5Q1Ks9ICgOZfR2PEoNkdtm4ONGZeOnH0WNEhFw7AdNbVrRjOwclh
4V1MpW2AvFxR0g2oXbR40pio6iAnb90YKrfrLmNwVwRIKXidM0vEhla7hfpz/5OdKUqduPg8J7nb
dbNNuXv/3k2hUDI32bzhjKp9qI3cD+wO5U86/6OVf2cd6CpZsFbC7mgcnX0EUdluR98wI0otpnkB
maZKaX8DYoT4gQvQ/UZIC0arJkFjmvcqTNe/ebAulPco95Rwi2qm3PiIWsb6qbl0l5b2a+ibLc2B
BNCXL2Y4mSYEHVbCuAq90hnW0csTvfEFlK8stpkbX9tQ1To8XVnyJx0J3Lh/pLpdT6ZYV+VscLze
3uTrhxNVcDy8CxITF7xw/SXFJB5NTq6adunMLkfjo+VFT7uGwgz8dWpo1ydAqJYgdzDS6VwakL9/
/N0Qlz4ydjJHUg500FVmy4XnVMO51Sx2ZR6sYj4yETc+sRF+T6JhMs7GF7RGcFH1DQB29MvCVgR5
0juxheBFZe4zkjdZdeW4BifiP5nLvhm7BTweK3fl+Z4cilfF3mrZlkkLrgV0o7l1eaDjIRDcbJD8
XvnTjKtwpu6nwMchMuA8Gb/Bi2Ki/srERthyz9HvES76r7xvFGo3kUE1TYX0pgrSBOommMdMYMVq
WV7n/afG4HzAycYhvEQpBU8NIDE8+GiPZk/hM/myJnpUvCRYR059cunoQI4X4udsCMbj1XmhBgho
CGxWQfhCkOtymkfPxRjFH5MvU9A6A9eIjaYrM2pELVqX9Svr0+8jleQg6kBaLCCGU2ANIUqRWH59
wj/o6jzVGZ6naH3QMgCLk7nKAh9HsQ75Lr60oCfRsy31bi/7esiUOkPq4u1H1hjEFo/vux3LLYtI
nnvfD02fZTWC8MATL6RSk7S1QhMGDYkq7LYWYYhRdHlbr/iNa/vAdnEiZFMUu7z+g39N9mTY7VCz
JFMdK9jPbwl79WZEEpnoF6KgFj4VldmMD7Vre3UI1VTeXpcHEZpe2A6YUROV3S8EtE30WGG25byX
BZ08qWtrT4ipn8rz4Wu6yv8UIx3VH5xWA6rX8FkBo/9aWCeDdPwqmzAs8Ar1hqBSBWhfUWSDebGc
k5NQdhf4u8mezx7tfLBiazgd2Wbfn7GFrHD9ErayJiTmF6l2sANO/6CGmmLCGMFdVBbjFOU1NKvm
RUwCXupOQ5KtvzLfLwsnBKyyoL3CF3HUExZHv0G0Ap68YHCKg5DOccccGlGYzRpvkJTiSqhT0pCJ
4WleRJgvc08OqoYOn6geX9RidFR3jv5QKLF+TDPVlC5yr2ea5ue4JriSbk+WQ/l9LeAsBynGb1HB
dZH6aAy0Bo+UJe26oRQW6kizz/aJuFPOL21cTgaJENzmykp7wpnpPDm7hTgwkI8VUyAgcIqdouqx
watFxng/gfCIPPPZ9gHKkcsZHFXnKaLpP4EUSJOfBey9WOD5ka9Tlbq/ba7AYFI0K4WGeXv+duTj
FUbUS+Govo/d0a0GIwlTZHTSBDeNS9xgSqgxJQZXCD8YzSQ83QuQuJbQXdX5aq+kcPm6bPeSIguL
nL2aeAoN1d+BdXbkV9z1wEkUq4+lutxM8WwwkorqUzK9swfW0YVNw1kqlHj1H12Rq1HQ9TcIWhid
8xLXkVw8J/b9kpQkAFzMG6Ofb9XeDIp/caWtcByW/7628myWmgkWDen3CdcXOXIYEW6JBTeVzvgy
5Irg5f38FSKuB9if/ZqxLj8uxqH+CHb02M0kddzb5fQGJ1bVNI+2D2hIzyF5yFLNqroUdvCgPL+P
5m8mGAScEmEZs77ukcgI0xFUqnMjJyQuVMRPcTwzfOxAOsDh6A8Wn3cklwJk2t+Btd6RwdMJr/TK
vNdhl8tiD0gV+cCd/k99kq3NGIkwVn9Y8Q8o6asXajTC1muZ3woouMsOZbn2gGtlIOyg812Uuk6V
dS6z+yDilRv8h4sKqV+6QrliMfVD6MYjVXTMDze8VZ/yRHKksONqoQUyfQCFX4vX9FtKG2OljyNo
6z35VW9uPg2czFOCco5ZJ3wKTdlz5/GgImjrJoESFMA6MS906EUY+9BIOUi9lKD0ju91Q0LOOS+l
3fnIQPVn9PW0Y+XQgkgbUdUU/zjZE1MZZYeWf+Dm16vQtijCHk5M8R9pEzQEHcgWcNo6zmFVg0Wu
rYlU5DHWI975Rf5jcCFQcf9k8RAyGs+cu3UJYBKdWIxCBUhBu8USoI9+fX26sl6LSxpnbS7sSgrH
bHLH3TtbRKTzD0/Q0SULq2vH2Wq7e1jd5zZO+MMtNP3LIX/PJuGjGtWUfX5d6A4GuwprXXIXqMyT
pNOOl53xaj9X3Cx47J/Z4tuE6S0X5gx+ancgzgaW+nXG8FywX0HkthsFqLgnBUF+96X4KRDSlt15
EBgecbvw/un2o5Xfe0heJ+uUae1JMpkD2DQfz0sNe4ppWx5Ws2+Rg99+HH5ufaUchkezvt98som4
sTJkOeqoews8OJApsyfJCaIrEhNruEJfbdj1KsEdoRbrGwvfy+ty0gTFPvWx28HirLzoVeft6eFO
fDZZTTBep9UIJMI0H1tf7QKnEBt/v1HeWN0ozZqkiz4q8zCp06QUswLmeLNfg+eBf3daE8eIgBwC
1fAPdJLlPAwozxQgZImCUsRsPJh5Kk2XiCBZf2fYYwogRNJvmKHjTvHewDeA8w9l6C++S2qeuAnV
Nq/I01KqcTv6tQsMzkxUxvfq3R0JrJdifK79ZLd1ph46hJv0XI2UwECdkBoZyqakKmtrCeYFZeYc
xFDk/l+o6U59GqBiMphKTRzE6qXNBzrqbHolCbnvD/SdeVStuA5aZ4IorqCk3aWUVZvkQHwXHSEL
8KdJskyLAIAFAn5IM5pqPDeUZTLsci41N1i5P5oXvj2+gb9pKBbFPuBTwEU2O81y2BnR0QuQAqfh
BC/YptEpI6RwVKt8czkgb6Nots67qcMJY0D44uHhnqgBdsR4vyUUr+PTuWqhTq2kRdS8GjZrWZse
qjoa2qR2AIeYUtjY2F0fT2xJD6mvgnnuPbgWRj7QnF7GvbH6bMaY+3AqnYHV1FWxHFp/5auANR5Q
jWvp+SMwia9NLNru/vPp8jPL4SM0a/NIG7QI/yR8nbv/Ljy1p/1imQs7PP/dA5DH6+fkxtfp1MB1
2hcWLpGoa0zByuGnfKuaEWYxd9TqmTvHvZtzwtPU0awHW0dr23/SMMcgX/GS5VgM3hjzJuZeNC21
FiCk8DehYPUs/pxdJC+RSykrm25V5LFObrxesr2KmcRcJZx3QofNBm2u1j5vGYDTC4zSj2gKRBE8
sNBGJ2l0NUsG742PY6u7GQVVSSDlwsUNceg6iFpJJvbINSF+dpFF2IK5FVMrvI6irShsG3eW4DDk
IQ6HRQ4HkhQxlYmX5sKsvpU6DqDu1AkLLxqaat162HG/qFdBcaJTZlzLQM11S24C24wLpAwvbAOL
/e9pZmWeYVKatgF5zBfIoBWUSA4wdaHK22H6/i05S3Qf3HA3z/e9kTM8RzD4HMg9ygrhnzP8FQJF
yK5HwINY4/oPnzpPXIhbiyz67B+2Ea990mQgtG2JEWPwc6nZr1GWDdR+2+v1og9+Gqps+QjlikXj
9gJj5PwJd24d5O1KKx5mWNQLxtvOt7MFTmJHWveos55H4SYzg4IA4zCLVRAWdP2JWp2+7lLejpqO
VzA6DgnOojM6Kga77opSPQDAMcwAtu89bgqcD+gR1EiefUWM8UZloYGKjqqd5LN0UClkUar6Ijyr
fmaJ8JWipycHhB94gRgYR+VI3O3dTrfuqYUYvIGmmY9BTqnLttePJd/AXMC6jU9A1jI3nO6Ea/OC
2S2LP76r9MkJofUCilkSysI4O89ZflHoCuvtWGtGwplFADWvw/8Kyz3n6kFsUJSLcDj5hhfgiJIb
JwV1qRHV8Ab8c8g2wyo6D8QuW0bDdjUNl9cmJkDf9vxv6D8XutEezkswCd0r/A/MsrvSnl4Iv67v
Cci1ciso6/SWCAgBN+TGj29lrVgP3q9NkndofeCQUaFjLQ9Py6K0NsH/Mh2ZbWQdeCz8ei5kONzf
UuuJzWs8N7VLJxIrLD4HMvpJvynZ4qAj2rFnZ+MJ0S8yA5XSTCnC5rfLbClUshCzna2IBbhGdcsX
Op7QPh3gBWlNSBv+xwbguZyAtZvLCVYCCRwV0Vs8LU+YbddqzekehjEboT5YhFjTY9hTTz/87LO0
T8jIezpp1lY9KNcgcSu6W7/kxgzsX5nhTimZBJEaVtjsUJEN8HZ91YGR/SSUwjoXc11e8t1XRB2G
HwPUqGreN07p2mi7mL08x59AWQU174zNfvdBwU/hUus0VUNB08Px+gbC1ZF1FJ+XahrA+WF+Unb+
zUCJJcZvU+wh/ZnFnoxLMr5bl9vob51RNrl9bxi1tax3anl2fxbJRDPsf1BMTkXWaY97GZXAPScq
hIgH/s3UTpdyL4VVJiRX8rNScpFM0lC8Gh1QWgDzuaRG+0ipA8aG8WFO4FE1TQCNa/6XSzpsUd2f
MtBPI1100pZ/lYhnZtoY6ONEcbsC2vnSV1sbSStdEyGsk9ae5q1l2sVGPvUR+mNAGkayVQpWqh8A
vMQJO9nrRETlQ9/3zb9P2U8akwqyqTTp/7pIEnmZsZXMYCBsHoZa1wJB/gaOJq+WMd7XXv3pMpH5
jnsagHOzWn+toYLWd1l/Clae0uCa0CHPv2nndal5ByQDN9NVydRHxbf3OKoNteGW6pmz1KwFEvVW
Bdg8uwOtkt7AGdtbIXEdXoHVnj5SeEkMYZXFyjYabvGVDxfB1Sye76qmqyaIjDO5Nuqoo2lZGnu8
Wo9nDQHElQ+o1JKosl54ZA+lDeuCCg4AHo0t/EZ7pjXZEsxXV8d8/yi0yMUq2vhfGPxQfNM+e9aG
s2SMptSnKQxcT3vhYDRcmIMq4Bvz/EdFzbF6r1l0+NASOfodhlunSIQ5jwKKItx4c63urA1MonU7
ZqWoyBFGho2XSdQqFx7CbsNbhaQaz2AZ9Yx/eCjV/7a6zqEiE653VoJvz7naMVOvhI17bXe+ZRui
vTz75XpOnTkOOmJYJNWid1mCQGhHlAE+paDj6jCR36ZyrtlTr10rKKRMAM2YxpeDpF9QWHaibFcZ
1/QSebdVvvBqIxi2kF0mfYvulAEy5bDEKnf0ugkGK+ropofXj7Z6t79rPmq1kojoJBJ1pmKN+KRd
ghDACPie9NSRKr2Snz7K9KOKT4yQpUn0oduM/Fc/6glAiAvd4/Ru72w+oMfIsxCz1IyZU2ncxPim
gTA4lgBfwx26wir0NCxMLKb5U+I0AAKK3BBgC6V3LH/LLnoxXQS8MyJhb4kXzEu+aCxzN1d0yLV+
0tGPCVOoVMWZBhfqa87l0y9kBECaCS1qSvl9JSaERx8Yu/Zvga3GjJ0wnRLh1uhVUSbpLZUysIBk
OlaLL93LnmyQwlRVvQtXxa14frqOKL0q6vZ9lI9YxeQbQ0Q9q2QEymftl/2RIrJ4j7V3i9z2AIvg
bLmOVcR1yV1hzlOX35pOeK6kXV0XJC6uK7xYwoPG3FJIoD7dHL4NdJuFy9OXHemNJTWSlMMjHeUW
Ow9YwibPUm+6UKPfJDZPtOysQXAKZ7nzCEIaIfZ1N3sGyiiQvND0YBUkrPJC4j67Vt3N03NM24XZ
V9V8rrK+Q7BGq8nn09BN0p/sSXagZi/ldkejcEKaqVJt78bT2MnTJgYQept9fgd07F66h4PN9GxI
KvTbRAE/k/V2nGLTo4e2l5zti7/D+8Zwo744YUpcQ+/hWappEpqoYW46lbsXGClhGkaDIJaYpGF3
/RjQ1xN4iFaDMOblEzqPrMicDjT02X2COaFHz60dbVo/Nmp/Ud3Xid9fBSwVeCGj21daIvadKAMs
fRgYQTLTSoKuRQzxcZgYQ4C5+lAm38GpF6ys9BUL0lWqqVYEBwcZHm4t+0vcx6YlutpB/WUlvClG
SOuvljjh3kR85k8KHSMJhP0R1UZ0U1ua5sbY3qbOriQY8AOD7ImObKGywi5+KnQL/I4uvmgiQHJp
H7hDL5oZCz5YbxKS0Sfm2fMAtMtYAzhmADkPi4SGDhXdLKylemmxRdoc+EQY1g35pfXMLAY0WOXL
qKFcv/kXiCA9AYETKzZabcIN5jCAtznzxFKbnJNSsr7DVwbBk3QrXj8vshM/I4US0A3SvywD6yQM
YumfslO4jSHPHVxTy5oUY2/4x2P6mIUiuIEPPLH12luswLc1aYO34Cua/Zu3co7NSBIPLK5D/LRI
jWGgVdJRsWC1iSoI7PiLL5FK+gerxSnuX68alnH1UmV5tC/zIVy5qk1x9oCXGnfLdFiJ9xBiu5uU
+eFomkd1SD1//jPjpfuauGsOA1mvCGaZUDOiw4W8pDuUJlos3io4MwTXJQ/4ZnZ8hNmbneAxmmea
CASy/X3x5zYBPc1m322gEm1If+QoYgozn4xl2X7Eu9DsQKSXJnUJqoneqKmyswnUVGF360WiOU/t
kxCP0NvGz3u+dBkRGDI0eLLdFJHaDBrTPtEYwy+AYUBGZfYT6gDQqU7q7C4YJfOuWQN/enngIcBa
+NvYPm4yiYaS4iwt6WGmSK0nbUKr/2uE7A5YjJF8fIBQV/vq1iR4z4UvGcXbA+fX5T2AIVrrMTw0
9pw3h2zRHhNm6SYMm6W9esUDXWXdcgCZKCOgQCI4BG+5l6YCWYdiO/hnvJEMy5ZHl78BO+hrg2Ly
N+tCWO3+ovJD22zVQCK7TNGr5J6XhsYjm2yP84+4hWiDEuywB2u6lZW+GArmhkb1HwcTpf8tpEAK
FHFsjzshpUDNI1ZjxCZqgYqofj5KRf36UemaaHlg/RUXVQXwFHrmQeOhuLswhSr654syaTFWDCKU
4fxn1cSUXXPCN0HGoJylDEBTCt4vHBwhn8dbQ8n8voLpn31+7YcPxRr23oE7Ty5v+cCFNBnkvryR
/4MrmSALLaFHMqmzbf8U7z/bgjvVB8Rub6Gj/lGjHacsXwIox+MmtlaO3cv5qa7QuyGXOeklfdkU
xUwOcP67kFom53ct6DrGw1G3KAluuIXH6mhCEFlZUBluL4iGDPgF4X96F3eKDPNuapZl6sH26q3s
j2qqSP3QdQOfiJfFXOkKLX9ZDw/830LnUwUlMfPAMdyvo7yY7AkVjfwReuw3zK/0PG9fCxb6zKba
8ovpwCBQqofeL6uWzklin7F8veKjrSVdGd2YPH3qnjlXq1jExLdWQUC7B0ZnVbjY7VEhiqdV3VPb
FfyQO4V82265SHCWOyLjMW/+iQMDnsALulCEW9yGDadrKpvTkyjm96ymvA8xbcDNwf4EAWIAnL8Q
qzuAstG/07x1X0J9dhtLUsDjn4rqw0ikZ8CUgoTAyxhLI634/FpEoHoKGbaCOHypjcy4CFzq/oT3
vEA2s1ruRXbDjD2pg2pCfVk98PxzLZSTF/dVxAL94+a9aYaiVmFP4zKnqHrj/1W+NODBpWdS8r09
1463Yn02vtjK7rnPumnYCT/Y/GrLzEloWXsh/lqdIrTUs/ZRvXHHvqluGdzccea8iw/pmgxhxfC+
7VqCmMAHaawBrI+B1uEmvsJbT0cJLw/ASvONKtMfMxCJ2rRU6qbg/Bu8BxSajnpFpydRrzlAMKzg
YXq+aV4ULmi8wsUFgBAQivH9KV2EpPi8IlaXL/cTYaAf+teSpe/8qkWSnxZR4TzZxHI8dZUBYjvH
iNqneUtyz616GNJspZMDX1u+OmXVj5UAhlMRTFwWzo3PSQTgzbSolGUyLb6KVczgI0IFiEdcA1En
vykAVm+sZtYtM3Ox7vo3pQmknDGB6HzOs37xZ/oP/vo6G8r9VeSMpwQOJ85tTbFZ1SUMwR/x8MjU
ni2fXgtSTKSpaKb70IHMfvS6yD6cVkehnetPFKU0CSmbr/NKzqDV/ZHUTTko623bOkI/HHSxbPGf
DYnN5ASY4NS2lSe0/ndAM7ZdvXR6wWFt121zCvvaiKDHoShN9Jdoy9Hsf7cZ9IThBD6z2CQq0P8i
BZC/kOqdy/ByZVS5i2q4AJMnkM3gpoaN25XbKef6KQSA6JHUVzRLjeYlf0eA/Rz0XVqgoPh7AReh
sFae8C2waepCJfscK9aQgBlklAAcFbuqcN4+69sLIjy1X5nbY0bmG3qSl+6XHy81y8EFcBtbkD7M
erziR8YTdguZqyWdE15ewpGxRwi9/2S31+ennWkQi1H9ULFJSmPUsGI70/3FfjDIcAn+/WqbRldj
n2CSNAFfdF2AQKux3ur5avtag24I097nK5Cs3E4yxVmxQPCHAS9+aoQ6ws1Lh4fy21sVla7KQ/tm
vzHMqeosNa9JKkL/QeqLPZNLdKL6SjEBC5GXcXnV6ulyYAjSS0xtRDHrKlzbvEMn7pPPp2bh+TwW
u92HIXKiRlu7lhhtGs33uRvddLZOiB4zj3uMEEIh8x84MMPG5tUrSS8kdv2TtvIQSUflQhVQs4HF
vqWk3jHKqSoYDpDynWiqjW1CY56xmIsi64WgO94peeDGtMvNIR0udynZKTPG8rbZL8s3r8jzp59k
VBCDPJMJItmRCwumhoe+y2XVzuIMSpZp86fPsAKWR4MjsIdjUpwrW5z/5Gd46poMAUYxXQt9wZIS
25KTp/rOc8b36fE/EglcqUjq5Irg0uq4M8FvJrJlQf169JQZs13Oc3g0/L+3iSxHWAl5wJtVEY7C
Io1QrmqStROj2UdsqjD4HrZ0oVGa/oHYTPsla/y19yXruN1gbuy9Px8HpfS+5oNuMK8mX47uVNwi
DhQZQt1Wl8ThSKrefZ0DM47l2wl9IZOcIsBVPlEwwTlK+L3l9IMSyyJgUEudvKoK4DvMioBH98M4
3giuLboAGdLKUyiLAqWEOMOB7UnznQ5ZbhVdaIZVlfPbOK/f2wPTvpV8aZYLa/zZs+MAVzvEzlfu
b7+n2E65Zwy1VVCu1zMZW9Wzq8u+6De/OYa7IA1tY9lJ6VnOiiSSkwM4vK43vnGek+0P7r4Yj4E8
bGoB6L7zcnz7zdAcVEv1SSl/Uzzdw6HIoFXFEasOtQ4grSIY1iSnL1RNJzRidjIm6E7yspC1GyGA
vSeJzFlqe542apY2WTCTOAne/gkgEHi94oUwNPICv9VsmQhY25gkCsE9eUWxmk9jdgeRP490AOAz
ij9i415PwPfixJfSpMkzHyzG9YD0UZLpcYwT8iRUrA6bQHE+T81Q800wtYZWipb3LUkh40A7bR9C
80r/H9BWUDmQykvyv88ce0JyWT3r5k54FDYfbweYntWwXMJiNxeN9AxZjft9KBGTVssXqWpG0i/2
KE8RC7nIIGybXaHTD8oqmzun3uD8O22288Z2HEyaXmJVi7mo2+Yos1ljyx2bBvWDYyR5a3WDNiZO
pcw//31LTwuVuqLE5jmNQp7Zy8KuDVwR7Nch7a4S/h1/80o2Cos0UqHREAevQ4H5eOKD8e03i/+q
ntfY/fbV+nPmxtQeWHTBIBJGnuAzm+I4Feqrh1s1x0zGrHKk8Ce4NKcQDLUnDs9EPybnY5LXt/Ue
c5W92WV06ulDRuD3y+xgkzB3jUzUXIrQHB0ySL5J0+Sq83XBDbbRzNH5nGvfJqll/5XtXlqXjIFi
ldy27gRXZTbhK3wd8+7UYJrTBZESAOSpZh4n09l34UwW/24oVAbHauAWyMqqBYXHISYESQXF+gCB
3DshR+Sjh7pAzHkeMD2VBXHv8/ofCivxxIOnR0OeMZAThJ2FX73elicFeA2IemKLIPgUgBtUdkpO
CFrvRsmx7yZLqLhCi+jSDjKs9gEnSyaR8pbnAFpmJ/TvlF+Nr8KKUTxcBMHaDgUTMJa88vamI/t2
9xKR802zn/rdQHGXvldKTE2BA6jmE/DK2Ia7yWbOuodARFfWUua7JPXnlhsKfF3vjWm5KtmvV2HE
svMOWddgLYP+Gr07mcAlzT/iGXtit5BoHFDRs2MS92+yI/LoCLl7b8GBiAUtuI+6Sp/A0BL75x5U
hGMkRsC6eYj+5s5gvXJLiEnOupOP5ZzClyCXAw1oG3ySKPWfIl2gZKs2qBDy9hdEy7uNW4dcpA2v
Nuw0TNgdV8BnI5O7S0cKg9iBPH2Vlcw/nPg7sXs3Z/f6FmPaSGMrAOLgdfDlFq/lBmBHsu1w6Pyz
17DYxr10mu5vv+Zo9zb0zST4ht1VWiO6PHUqdR7PCk1umtBuFOQ9gOJRFtvOp3AFF58zxd59koP5
Xdoz4FRnbzazdZaGigJlCscaQJmieK7+rUPO8X8fq6UUArc8yT9Lm/XsrS1iMAJFlN9H2d9QooSX
oyb+ucJ5aezPFi5tCb6SfxGW4p0fLprBLcDEoySnuYoV85Zyd2SoJ1TSduvIePjOEuDBTcjg0qDv
tqCPKSc3iuHfAHXafYptyg7tB4UG8vhfTWBuqBa05Z1WZrtyop2B1Th1WxywzdojD9yaVtyl9rsi
Kpbam4qQPghLG5hSxVT3Weuc3udZGb7JT+nJhhYJ1/iOihd4Ep3VTDTMxyBwTFzyV6/tr/WCHZ6p
OpL6qEMT8xbO80ZLw5Sc8DwYXzZ1zlmhHNb+/AdW3zx/wvkfESqUMLKExPDwPNzWQJal1NRvgzCX
j3D6twVcF0eIRdS5uyJFbGfE8GJrtLK5fTJEnAg1Q4eFVF3KOyQEuWaImUwwxJfp5OOXTy/fdpMh
5Id1pmR4rxACoSfjwxGZFy0EcRBU/IH5Dxb8N/53dsbHisJSA9DWPijfZPz7jELyTLHpTAR2cdN+
7aNO0WDrwZDh3guY7KsaDeFIyrsgHiBsQKOOtmGDF67GvqdGEpQv6py5fRTTPiw8RVdLK2jOYb4c
UET0GUHey0r7MVVoGdNIXyaelRtrVeWQlhtRpPjzE+QrVcZiq9BEWT+GAsUlQAD0zAG1vq4+AkJa
0jhlw8Aqwp5jw6PjNeiPfzHf2WIjIZDvJrQJo2n/TrkbJ5Wjvpg+byk1rUKzq3/LjOJWpeaUtigg
pOusrGBCTJaJaOruPByEIktHlZcqkTseYPfajylNv2jpbK2egk3DZjZEjAmSflqGuBRQ+4VFGi9e
HTHQ8JtG8woSd1tdVnM5q6an/ai13Tk8c5Q6vfzG0hijcebCI+bfoRr9wZFLEWokHlmtcUwhcFsy
iv6j9T+K6kKjEzizVlBiDR9mErhnhVmLr7Lzy/c5kCxjJ3JgV6UDpHEaQXWnT+jxQ4iH6cL7vHCu
KVMYpxlFAJhP4ZvktqhPyQXsuiie6e6LPeHDgYTFNZw2zzEJcz5lU6vloPmZ8H5AtCdr7Ipn6z6b
/bQIYVmoMJ+Ukg86R6E/iIErf19gSSqdkIAIt4sXot/BEPtxAHvdz5a6/LnpL/VBBVaQM3x3nZt/
7n0ueAcP9yHjrU3BzK9zzMPqbfEP0iCkcXja3VO3NgJ2JNWHIJHEizFew81ZaCnTajVsRqF3ew6j
ykKbVkAomSPNIUFJKMEfSCHBg5Pr8bQocmajD7yuujdweZKEdAVTR4okTSly1+L9tMJi/gRQavaO
idV+PCl0vare6Tmig8ow9OArwOwueCceqCx79DTzL5N5FdtkMaZMr7uxF0jb2WXGtpTr7G2nJvjg
gEi+fSzHzVrFD/g4fr5LzYp1Z3dReJCr8KxoEZK/o/e7XarSVnKp+cjBEkF+Cl9m58fRivNkP2FG
OOHUS39am2Ip0sFfwvj5tRtuFMHEo0164cK86pxbek83hPzVXPyzVh+mvUL1/wtGgzePiXphuIfs
Ltj0pD9qNN5CWH7n3J/yfDpj+SAvC0qPvqD1/TIUkfyuXY4kOpmw4iPTjwIxmRul4yugdmqXb/nT
Yo4NqSa0qoCBW3iCAb2oT8AzGGPsKSzR0RjqJLlAkoHnbTtc29VjO4qEU9DQEzEXxnZmqa0LkwjT
PjQPdaEaYa18Ql/NnGagMj/Hi2NyfoAlthF6McVQEeemO1Zht83pwpd/cs3GEYBn0jrwHbLSo4xu
HeeqDmwn1MMc0JL8d57FqMAyPBOxIKiV+mKeEm0yVHk6u3ifs0r8FDZSQCcJPOiG33kWVbv0Eo3Y
sgLNIxPdYMiZdj7t34Hj3ZefHCEUxLkQcDmZm8HRTd2kwPy2lr+7VckUxcB/0xC63TDvZNxbfU+o
0axSJvNGxvX9nC9tYI/korXocFnLfJkVBSX+7IBPihZwaU5noyS7XVbEi/mZolXjW4efzYQiPsI6
nJG/o7IeiWcSJnKPEyQqyQUFaQVNy1p8oayFPLHsMspbIZ94SBp55DTVBgG908NHZXWbpEEwwyAG
KHoVxG0wCPWXIR7Xwy4/SycsNJQOYQZ6BuzJ8Q7Tk2gBmZ3cC0uLB6JIsKeUkdhoQaLA8Kt+5mTU
djZNWbNI66rtEg9ekhV1pqOi1DAF7mUQ2eq68zqNAS5BS2B9x+dpl1hwYxzNTC/yFWm2id6F3i7o
Mg36bZ+ho7LrJYiFT9ORLGeNv3SfWXBBTCz/6SgHzhvfs0ERdTT31MJem7MeselDHuUvYN0Ibohv
8UgCtSaLRL3CzsHvpexy3uROvsrCi1h7I079F+gOJf+a+aTDSfyWs5NA6PBfU7VCKd5T35/8l9nj
C4pTSJLzr3+XixN81n85iIfbs+nR+0DhCoMORCh0VpPcESUqqiyj296673QtcV+6Tok1oBsYyeZe
u6iZejklxAerp4xeLObTjiR1n7SxhI1pIwonIJXzMnTaRgriuUUii3nC/lZuTb0oU5x3D8YOiegr
shM1xZHo99gOJ+QYcwuKcNuwxdplfGTeW/j5egePg1qSh2nlzl33qtZwFm537paUdvJki34hcXfz
ktxZImOb/FWZOVNRcpCAgi8Z7cq0ZXVENsE2V4Xn/vMJHwtOgHhax+qy+Zp6ak6ZtTLuKQK/Lmur
03cUiF0l1Xc2nTEMDfHPVcDM8Jjh5OLg7pbshHkWgQpSbJqmQvuukCGdc/8gaoIUcZ9fJPzf3ZYW
Pk+/HYbGJMwzPnYAofDgBQKtu3JBfHDWAtwf0geiNX0uG/zj273FP8ZWQNaHBG+ZTgrJ44cGS6Uv
mH2beuubV8Ri6MpWtTd05SdUCG8PGdeMLCH1jOarpmqXaxcda5AVEWJPZ5cJ2d+sNyOdx5gn0HGZ
4Jb5weF1c3v5E8rokhbRqtpXSIci2vornYKB8bvCn6uGvR/1lu/DZXRsTqFvGtYGZHsKtCX+cThi
XpqixXGK9YDShwT0tnnEsYrcgwBgmb9aDhU3dWDUVKaQ3T/q/1db1K8eGLPuejf5eNwmg1F5qsUG
0TRcEtvXA0iIJPxSAFq2HNZ/5bWpG8iKgsoM+xJDqPR/sUDVxhpyB0TiUQz91JIxe5xI+OyIGiE2
Xa5liSni4B0NvmzuYfl+k/R+Xv9YhGmWzaCfVZeIH9psYlDYJiEkSu+TrRTZNBzPDBpDgx7A6K3Y
vijTLqWHbxru3tTuNnur3nnSHaoy6b+XHeKd5hEs3/jNQoFcfMNAjeouX8Z5LPHUTUQeaZZZxRWW
0BfNMUND4sYgWw3iQeDA+x3BL95el6DK/O1SjNI0rCb3hKXS+45qWjfnmdhKkcUXZwyDzxAvzIkQ
3egg0MESbE42/jW+ptbUL+6yLy3t2AhD1X02kA96Lt5fiFPQKW3zaQWKD7S3dRPZtOlNHJ0CxAz6
ehGLFbWd9CC5MmrS1kRzUOPj3hL9rqXPmEn+n8mfzf8oW1xXhIIQqMuxXh1tHZZCZsIECM5prR+l
w5UBjIjReLWAOoOPLAma40t6yBN+jiNqswarNCf697HaD775ymm5u7d9vg5yP28mTmM1jCtgpHE3
AjllfqkjTuE0sedj7AYaXfd+UHhHqdAspkdFQJY/T7CcR5mvmPciWau9AB7WmvJwcG7zhXLLo5rX
t8O0xXNyCKRitdRXXUzAmrpDeUKz+486M+ruUJabiNwAwhpcehopQbikJavWpshMxZL68VDih2BL
J4/jrv/evfakYMtWmH3m+9BQ4Y7lz1kMA8gTxG9RphSIR1WN5pvEds3IaFBiiRb6+ZbE06+Ls6hd
PFK9088lUM/rhXm233G5c2XvgwOGNkThSXfa0V2Cnsqd6hr23f4cg21mt/HEe4y6Of6IwWOQ1d5l
OjE58xcLAuyAczwLIorZ+r+s/2zmPrD0AzP17/E5BeHLuJPvkEkNv+r9lwqmK1rT1DF8QMIBo0sx
OOhXdxaDtVXjqQFtBkMKMxaSUuV89E9wRQmBh0UZ8OS2wxIatNorpiNkGc3wK1fcwiSCL2mgWkC7
GLphzOti+U7gC0XNOHNgdGp/mm6KPzAOqcsaI1hl6nfMjYm8Eg0fqt+95LqCpaqyFYjNZKIvd7Gq
ODjaBRbaEz5nnlkdsg8fVD3uD2tFbxWmBcECq8lM8xMIU3IJfomrGzxixYAFE0HlR7b91VvzHc61
pSDCXbcXP2162W1a2BsmR7GVuvdWHCfUbHXTrRxWc/1l5zFZiFeMgSa122RGdZbt+KwHwIr29NuJ
mCRKOTXe0SU5007M1wmqDD7uHRGJo2s0iAp8etCypLDCPuNOzbn3/Irfg35RflMglToACv7yDVGU
IENeZEeKCSKFhp66ZiAFjGHn22Ml6csPHD0zVMGbI/43bPSKXXpi4KUn8CEGpCtb9k/NUgqDQouT
qX+vzxdCG/ZtdC+pXffVhcp/6SasXCkBYDkv2EXmq1/1/F4U4Htcs2arr/3FmjXeUac1UN05O9qP
4ZbjAwmVJsBTEIP1usxL0xUO0Zi/QRRS33CjQEqzuQ+u7ukIv/5GR0dwambyxLz4RViOINjAVxiR
bfdG1RQyhUeOvT+nKLXjlE6KF9ZX69jFsbpmHZtH0lHdO98KpViuqisVE6O0BZC36/1WoGk0ZWWj
SYqhBS6fcVPmr7D1KpK4VWVPT2DNCpve0BYtZ7WiWm1tyjDu7lRiImE7BGjqvWJKenaZqq15qOoz
mnV/tK5qBfpsJxlJnioUhmyMMrz6NMkj1gJdTuaskBZ0fZ4JJR7/Jx/DsJKRs3k7fgH2sRAJsU/q
PsFoHPOtgrshEkhwUl8Isyi7ZLAkYQmA1xMVs1PN5jIc9CnV3Op3XheYHCaRtsyB+SKVSUsLQR4q
zva5kh6SRLUZmATY0OWm30ruIP+fMgpEM9qCy2cg2tSKJT/fM68q5a3yIC8LqMVA2MBprw7217kC
l0zoKJzSb++w+u11JWgp/fQDPnK83lpjYqOBvkU2ncY566vwvtv9JTBYYFfRHHuGTSI089W/rXgv
g04iZHJg5mWQxvb12ptOAPkJik/Nt5vjNIj9E9atvQTHw38xoKAc25CeJnYdwMd4zAgpeWivamjM
moJq+hFS6Ir0N9R39W4K6D16x9yUvIKyZzMLbHXuDy4BfZOHDRUJeXFPHmrfKAmy171fl2UgihIo
iFQJpehP3xbqRISSl5i6tsABiwWISJy6554SQ0+HQ/EdpgjFuxurOQ8vw/kPt6BBaR4CxWXM/23t
OH0VOtrivU877vCj9etvHBxMr6CO84fQp1JzWgLWLJks/1Wypb7wNcTZ7eVlxaE5kTnlnOPbjWHv
C9+SDA8i+/kKBltDlSTsXwuXIp9l5+kER/XLb0dsjqZBSThK3ZvcXggKx7bkbt3QRt7+Q32l8OOP
bUIOfqPJOLhSg9umQczMgAJxCR+CSPqzVCp4fGesDhCw4rTd8GnCiTmCKjHQBeVhIOO8/rTz++RM
Tlm2fKtFD1uFfvujgcde9g6CrnPCBk1IRtLyyuF+H/w4baYyzIX0vMTUk3r3gljq9mhfSuGHPHOI
AOab1iqFqc7vQ0uzVNJ88ztdkgAd4o9gK0HGfNAHA370ql2KXXi9dcYf9xmdozDSNcVZXnvWwmtl
AM4rIAGx+GBdm0srlQ1O/xG1HFDS+ez0+P3/n2RMCgkVhcsMj3KnJWZ+plJJlP5d7Cm4XOEBMOo2
p9vEB/NaiyXFZBjUXReLusDo4TeFPAzG4/6OM/9kn/HjTimw/g8eaZrDivLqSY8Rs/VEoKgqh4uX
zD+AW5UaMWAf/NOEx1QWLdLSR4EWaYlulgNynmWNpemSEWz7Czwv9tkUeEDDncKzz4UcDprCqZmf
Cq0EHV/U1iAy4s5ELe+9PtVbTHtNPweckuYB7stp7AKdJk7R99W/dqDnFmXVN8guDhkWP1IHZiYF
ffGrt+j9HukVTO/vOGq2T5MyfPFdwKcoMmBaK2jK9YQ3mqfbu6Vke/WFXUNA3hFl93/1ZHxBPy9i
a5nDtpGp7YP8vmWDqj6a9RA9HYEoWdVvVy1konoJBvPB69kI91IkISIlCqc8pPhXVou7YX4TWOYM
K6SINbmAcZ3SygC/MSal7SCSnlvDYxNb3rhDdRALrjg9iraYaAYoiwNe3+SeN+ADDlxOQCjW5Ie5
AGxSH0x1ZKHupxll8Q8N2qsbnRTwzAqAudSW7HL+71H8NUr4UP3UVBL0Bg7s/z8HNp2lBlmSpHR/
yZ1LJPlv8a4eeobzY1HO5HtK4bH7kjA/mC1WD+Q6j2+D6FqV77X1MRVcHgWYMyKeF2+8UOSwXAJW
BFCxbyZcHc6K7bHf/RwPL9DsFKh+NbobcNf0SYMSctx5CPhyc/wYvxzCnaxsEI4oh4xgxKyAOhA9
+0H/o87CaIzBjONNkVvPYouUzL3i58nvoNc59bezR80mLjuz3u67jqQnaFSegMGpaABJszmQflcT
l8fxkrQFFWdn3SSoU39mSZNkiVDxxbDg69Lg+15+EGsa6puG4+jH3LaDsSqPbukzLdHoJEwo+1BP
MNxvMgoyGvFlz0YD5IO3U/7NTL2K4kHrQdIn5PU8C9Emv3SmrKhviNJzAuUSladtVLzQzXpi3E7F
BuRUF36Jln4fGpwChD039QSwfBY4x/LRbpYTUd8yfode3Ckd5rcKQIgHm7sUhcQfjJjjZCCOhTGo
nzObh/z1lr8Gpe881BR3HNOt3EnMU5io2dJL2sv4yS0M3/+nYGm9XSW9COq8tDKnRA2b8UcrSyW0
mW1OkyDxvEDgqEdqM3wA7E9lYF8t5fkK39g9wKiyVoHcI47a0OpZ19d+5vHjOCMRjUH+B9raDyb4
lDJYKsksVS5H7bHP+/bDWCnwR7mdboD/7t7QYkyrGyNoSZ1l5JWIDIzeEge2gs+L3x1g1uFt8wYl
78i8Xxh4X80yvy7idVf92r9PQuOI9AnZxP+wpc/zc97z7+gmJnPWzzsLgyJ6XJLnGV4fB97qhUZ/
B1BXbnTL/v5rRczhCye8K7tq9z41jzEM56zUnndOJHERLopY1fH0DxJPbBU8twyrN+iIMpzt8Ql9
PIzDTfScsNRn4pFobbM0emvbfv/2u5HBNYLYOj7ctCBw7GBv1t5QVxjep14LxxLzj4Ji2aNELGhs
4pmk9W5qMpzVSPNSlpeqdOzGyqz/EpTsofSewX0nTL726a/C5Q8KAGm9WqpeM3yLT/v7wMqpSw0Q
rVADt/R8F3Ou4+8FEbcP8GzIkcKoSfhbTyJMyel73UCVy3hMJSiiFWlMhrlBan3Pl01nfEdXyBdK
v6qPrtcuI4hTAxN1xjRWg2iqHJXFfKOdGN0Ivh4QbasquEYxxAuRobzYzddH8ceC7bNzySeJl6v/
ljUGwl5OSdYa5sqEvx/4nd7hsjDNMeawGfkKoa3Liq0EQv80mXvJrnEWEyO74dQNi0xuTTFtT3cc
nHeQ02U70P3sh1qVjobUcV2DawOUvMFq9fqyjAa3lSt6Be+n5NPdNAhTwh4M+CfEiLZYjJbEtmNp
D8HxfyMD3f6ZBVkuv7+k67ImZ+pXX/FQKqT/6Wlq8QjwFeaCP4qU640S6Sg50slB0Yj0Xb8PMTWf
aQtJnNTf2bTzl7unX4eS4f/5qK90WCWYhMzsEbP2ksyLoOoiu3pV2qw+9DAS/7wht9Jx6ABEKfb+
fYVUts1fiwIBPSFf38xxrzjJqe3mTRVt/PDTrKi/VfdWGuzLAjcvl15TRmYpSoSA7Zn0EbfFo1AQ
6oOqXTAl5YthmiSZROBF+JCLS1Jg1IamFQps8d2KlYAM8yY9TrUrG77iSvndQDXxLm+f8j91XZ6w
zR4WapAMytRxcm+3PYW4c9jTD6LSu66WoFkm0mvN295KsKpDoPW4E/9gqO/HV+8zNrrFMvNVl2iE
t2yDqMGiG45rM6cC8JL6V8nn8yQYrZSV0xHAR8Q98qGilNJK/Z/yd22j3/5KUT62NP71eMia5b8U
mtk8EQsrsp9IEEu/uMNuXcaxJQ0y4BEze4EzFi1wABcaVLmxvDTMNPEatYakKO2ZPlaszpMm9Zgn
FX1d2HCEFBJiDtrY3OTdokfOjx2vP0oOO+AF4M531QdF9qN2XbIfqQcn7n9sG+oBSpT8JiAWgAyB
TF5rxagWBS3ThZ85OdD05UtcwDCO+CKID1OwpJ4AoL46uFoVqr3W9zE/k9i5Jt8G58DLrraN5uJH
lETg6kYdn2Vae3D6SeaDvf5S9AWqgHl9GrzsieiyJdgYddx7N6OP9OHFZ048vHVY5dIjx5CzEbsJ
QN7Q6BAyMHOPWZvbYxVC36ekvJ18QnOp9T7s7D1R15JNoaxwza29j65hD0pN4gkpGkF6q4HVcBYR
4qrkXyFusT3rQ8uYKgqGsu/7S9rs0v+Nmw3QS+DB0aFvTwwWEx6DVecmpjWf9CXmEPWzfixdAM/6
TTiPb2QAaws9kaAOHEJaKejNAcGQQdm/07Hf7qv9by4xdpo+XTFbVPz13/nLmY6JGue2d8OvX5oF
zWA6KUKiU8q8WoAsCobM6hOrJ8OEdb8l45O6jabGX029NxvF2OYXuxeikltuxP2ADMmab7WjXqVr
efHhfxuX7/+KHsx//EzFagqphBxeLtNUIPweBJXwqdRM6IOs0e8HzzT/84Fi5eTV0pu3Oc9MO4Tn
N5M/kGuAeb+II1HxdR6NmJnQOgSpw5cToOfjB6YFeP2oNyD4V5iWOCV6hp51FwDc5nJKPoKyuZc4
yuKUG7F6+oPd6zRx90huGDqUe9paOlnGHEELzR0c88tPz29dNt2NNnP7dzkP8Y2kd3G3iJP+R+sE
8fwUba68qmniB7SHk0LFKiZYmXyMocGyG5byL52r+LfIT4pukNWLTW37VYk7FokdW67lWi4KEzIc
ZqkfW47GrFX7k6cGpOenAqrtBD7uWZCUJF3ydr/grAvUNegSjSYIb550Frr67ug8T4JvH6NIlQ7R
Gk6FvzKwIaIZal3Aq9mwxMYuVfmHbA0Vz2AOfcG3HvhT7JPuTlu8T6p5P4cqkhhGhRZyiL+Plf/k
cPm/qQITs2a9LjnXHjkER8xexRtLUyq7geUw7/e/S201T286jITffoFhoSCCZqRmqihEjyjuM42P
OLrU3nn4YXM04IVP/7GjZTQigqrpJ6izXfZsk0z7iVxCTtgW47nzqqFBs0mVVojz948QUCt6a+bL
QglSZ2WjITDjvM5gWtgNJYc/xL4oyErwqF6YjvfmMdhypZHWA6JA3O0xaC0rL8RIMUyuu2j4C9R1
diwtNluKSX/xVkPwU5Uq3ynBOs0q/+zMPsMRqCA9qrPytCsKoY4PqNbSvsIDmfhFR8pSzIpSL5fV
op2PAD7uzs94JXJYOv4FtjipbjtLrmS0IfoU4DHEzyZ7FqwT+u/qRykSDK+fhu/mmYPGgH3D+MXw
F4/5Qf5UUPWjiEqOpirl7YhzOAIw9Uu49HhbCY0fI0AlzSKZcuyD3MnfJ8DIZjbAof5Ga7zsvGQ9
H0zFgdUfej5BKXM+yZpAG96Zs350R/QMAxa7a3bYcyZWkLPh+YHRhIn3EH50YMMyxt1a/ACGKbCb
5JKIGqQbtFxrH1oqw8dzsYj7AIs6f8mQoomAK6rGflnF6Y37mlfcKmN21nNQEqFf3Y2Op1WOBV9U
TTOES6Red3X8E234iZbBhEGnp4AwbNKi5jRQFpkgbCH0ek/R//s+GLR0yv3eu2NN2YZ2W+4xPS55
sNylRoGIeodbbU+6Nk2Dji1kkyex6POcH9uC3aMf6JaSFpOXlBoTSVBVzl4NsxeJ7NA28a7ICXWS
a89NwUPaM+pkYG6WqUbO11IVKm4+P0ItZtaYDpWpURFDjcZIpKf6SnpK3b/W6uowueMV5pdKmxl7
/9U88y5GvFsXgIbPG+dDkI4qiAAKeMAmBlVnd8RYcsUlXNN8bwyVVHU4/MwQLdjpVCcKFBAkmcXs
XiF7/uJbyNz6Si4JJI1L/HkNpMFWvjA0PpqlUzjCCUJvIU5w1UTaRfpw5xamy5JGxCDsgIb1WjaW
XuMm+WEW7XnCqbI0mEST1vtin1wW53k6xQazDvZENI0ZiasaXSMusFKII3G+SR58Fw3xiXBGogLe
nAi4vXYLgE9eH1U84XWwqXUk+m3tgBMta0y9/LgI1nOGPkTGMC1jcdg6CykbhG/CcDpiGcuYmXr7
TDLAEc5+MgTPj3VFTvw5dLmo4wLyc4piockJl/b0Iwq5Ng5C1Gu/bec86vX8lZoyR/47jIbz5FzR
qCIHNs3zmhdyCL+7QwkgaS7zPuq8kdavONrJCk4R2ubTfTjpsNiygWh8DIKUTY/9/z20xCaDIAhu
7JvxNwRF49g51a/mg0KoiJme6fdatjgA98hYbTQuv6tVYGikFltrt4b6eU2Q4eS/CR/lw55n6SLn
YWOImYJYgXjN6LOx/ChVePfKwlJQ/7KRZZYTeDHBwN07JVKATFQ+9HBIPh00ADO2ZJbVVF0e8QXc
O5XCrC25zIsldVzu6j0Id4Oz8EPbt+wPevKrvfBqdiIxvH9rf4D++/YHL0PjOQ34ErbV5HS41ag1
JUdJb8YPjVAuYNfKcG4YsXT5ByDCryGmMsX5cZWpVMSCUA77zRa/502Dr6iO1YVVveUbxkyqsWUu
NxE7UOIglrPzOVdGUgfd2k2RsNi2Ke+Ue9mQ8Re7FvZyOIyzCyTHm3qAFNkAhUaMCfwJL3THwDV5
o8+T+gIB9kLbPAVSe3HrfTZcIGYvHBuWeo5Y4CS7Do4eioDRVifJ2sJZ8W8erhCIBa50crdjCf7H
UPtg0eLu5ayfJOmTmQlDRoEmrnl/WgeP8W73KGqOEAvbr4iKcD7HaOsyjiRICD5w4v8fYxvj/med
swYQ/LPQFAuQR2HM/r9t/mNRMRno+GTJ+0l9CEy/7fPf++V5fkQgIupaBK0c9VKcdW4m1WIJJJHp
YDaoDFCblLaDpbhep/1xG8y1J1Ew9I52+HN5g171WFHWAV9VwGFGV+NzKLF3Czq4qTEzJPaKrubu
0fJxF4Ljygb36ija4Vj+f9HeWwXnWlzDAZFdNfuQa1QcTkQDkWleddUjpNh/6HGrqcWOSQW0BO2U
MBUQFSGzBUfSWiQ3/lGnu5QQ83j9bb83u2IzGKtgX0xx2aXdmSS41IRyLVRShbOGf9WQv4G65sVo
Sh99bVHVBHVFkk3A4JFY9sYQCovNRphqm+bfzH6VcmF7n9vN6uCrUmjTrogR0pb2fwsUojzTubiA
FbuH1zXdshXjLat9zvQ9rtHxcijz+EibxIhKTLzXtSjNPozVC5bPx+mr5xXPLdrL49o8WSXjjCw6
dARkbLyoEWzxXL2moo/gEsKDk6L9NviBMujKYv8GAkheiu2dspmWAlxTzQjk4kUnqIC0XxBPALe4
PHDce/70NQ/RggqaInzc4w6I3jC40R0Rlu3pEk4VI2MEi2v3uIDW5F7yFSPlAgOyf8qWilByS99M
b6S4bIWAxqmTFNP8etfyjzYPEp4DuAdyPwaS7bDNQApCSyheZzf5FY3OTzVygTrtwUQbx/hDRKiB
/9SGj0TxF2oBoq4CnqBnwoFBU0Mj5BE3KC31kcTmAVYMqlyGH5WmeFD294mhEuVQSoZk1dR+JPHI
e9Dt6UDdxgIaGlVNhAE/M1iNPQ7dfIhtY+JkxeNxXr2+nTcW/bz90LJzm4pwO3T/VcNzLATWlJGk
Po9TaNAQl15TerUEr91BXAu/Bwv7Zjq4s1OxxpgeCUzdSB1tFnvmhienWTJzxzY7L2z6gi6cU4g1
s2g/0VoiiFMIttllx3C0ceDsFaks0FUmQu5qJwVMRxprPO2Gzd890rM8o561FC6UCh0yjmlPAT0k
B3nEZVzd+zRjcdkbG8mSlYuOPT33bXK9GUuFH8UdRq0d/CYycqU1PGYFdSZKc6cXeMaCv2CDF1rx
nTKtyRDob23zLq50xYg+KazT+INahhhbP4QqmgKGVCZg7Bf8nKDpnp4jc2KRCXQMn/j6bsYXkJcS
a7CRkeri9btB7mtm4Y5UGhFGY/bwwWrvbKWPO9vL51QMNxGdhtSVQ/aurLosqv8qJrWvuIJtEVdI
kwNM977dV2VpjIbciXfKGOu6yV9Zqynq1vB/ahieATHMrEdlWzA0fyMTGrOnPGSricY0/zJwO/RW
7mxMw/OOwkvkrENluu+MmYsnNtsck039Q4DPoicuTxwfwcD1QDPOaPap4in07xnYs/qGh8kajvRL
FF/H1IJypuctrosv7874UvSZLt/hi5ia6awOXTRbi/ygjMEpT0jQ9kQPrk4Nq+FCUfVCfAZbMy6F
hW2Tbbc90m3kpTWFRr+IvgMnhbCrvJv0EjUQ018XPKqzbct5pp/4fMmV/dWW09MiLi3ues5nN4y6
vilfziCz6yabfZ1C/ebiNy36DagJtUAT3SEAIXjpnpVLCEbIoPeVH0Td4cfVyOwrFbCyf14Em+r7
iztM9Ey6a4ECGtJrWL0G1/PjX3ZUw7Y9FFwVOuF1GMP9RUtHvk7WeHb/eReJ/vBJuynpwMsp4J9p
KX52gJXMXvtLgWdI4tj4j9+NNeWBfe6EQ6Zp61X71YQ/VRK4KkjWiqlYEzG/t59ekSwpH+tEKSjF
QYPm4X26YHdMa+C45Frc30AxqV843nJjT2WqJwkJaYnCvRr8ZK69D2gZOu3ryoPb2BCXAQjdeRKT
14BvOIM++ayb1kW35T2ntZ6vsawUbYDlxKkBrqzP8cATp7jXTLly+LFP7Ugv3BX1GQZ0F68vaveh
40CUEBseHxwVqfkstXCwiNMrYq8Hkd4XwN/KcaTpzPRa+iixoWVP861egXQF47hvEYBtnkcRekW8
Qz/VU5AEzgQy35yuGkBrsSw1iS70Rq/StUQLpNmII0tgPMnIaAZ89zcubAf03fxIHc6WZuyPwORQ
5rTVSwuZUkxNO626dMdtuDAQrpGGUbiBAh1cYZiomlkRcVdZy+0OTafhfmWLfWikmNdcHBDOrPF2
E8Vvf8H5eQdPzZYMY7z1f3Jji8+1yAdbrnlgAmxUJR1FQKXMcAViO865BEGSZOAJL3YhBqwRmWij
Bp4jF91NqufPK/7VkpINV2LdueXonPhfnDgdX4ZLbu7kcAtUgO2gVgbV2GbZg4eEE24LIAIPJPuy
Chzw2WI8aADk1RWZuY142L7v7C8wNto+6XQHTWNuQAB6Vur6cH4oHXdvT2NfWXdav6jyWxSU+Fwl
lq/acn2ei2igihE+BAaLrsMCE9dLw8jYkslIcCBjNID2J/rLRz0kZwLvF5t9JyPnrlu25fp3sV1j
l5QYDkSGfNgaGMbCQTHUjcDY3OB0NXuSOAzkuUG8n2dhWZIdvyx8sVBQGU14oYBEEJbOt9IhdOYP
PDD6J0DUtzUlwPMOul4ZTSXGbycuq79auKF6S6q1ojarhPDPsTIOKpDxfaBck13EOsSAHUz8mwKx
/3UbXvjTeI8VJNuJVycr//qsCHMxtHDbnjMDJP34SEkBX4idXWPnZQBC1gN0oJTLRCNmdXRaqhv3
ayIBQaB+u7XoTQhjoodXq8RzYLLYpzzptU8MbC1wEloSOXZZAQjZ6ylXqZnyBg6ttQ6cXG1p+ppx
S38gJj5dPV3c/o6RGc0vblaxNls4ZqYWHd4SIg7VGalKRZCLwFxNEXb/QAuYDmMY0O2ceETxo1v1
3i5U3/L1Z70VpeYWSfqEQIptE+tAjbSTuFrKzecgYqficUad8MK8yws2JFmHzb4YrJ0qt/NKje8u
3qJdzSFIq0kdHK/0cAfshtBoymKocDX/vEe4nOIXjvIG24UmIJp0UpeZYjwaDxQ01rxqdZfisdhq
IFGvB3q0H5o1souyqMTrBfAJEXBeyQtmHyLPR4LX0/ON7DJ1MO3r4DpgUVnowmnTOsJxTIG3AeD4
yDQdJA80rrwzY6lS1ymmtMFB2WvLrcaNOjdPYGeFMu8NO6ckGGsoGJO0DDm5f94U4KkmRPVZ1WXd
Tdq6eYX1cu/YF+Y4elatwrA6EJZnTMbDag4/NKR7Dqli9JUCNwmBWAxMO1LWRd+LQLrBM3uzjFJA
38xcXx+QT/zxRmWHGQKYZV8hF8okknGAeq4CnC+nJdFlaaUPranUws9qbIq6FWs9TLovKCejF2Wo
W2A3RV8rPcYwCicPbwgNQt0YNqluh8lUzLRnsizeZ5+a7Rdat9/UFptqC3W3GSb54cyQ3vf599cR
w9ThY3805aoTFDi42OhKvW/4pJgepEKvFixdwYQgkPykhk9vqXOmfcGV0FMcelI2SNowUIFSwPHK
kvyU4NB2GNGjB/gEwcYi6fuAlcf+/XEvcsWYj5zECqA+yLn6wDKRlObM3QrfmYBxGfQO8vMNfiMR
Ayy30Fk9itbwCbT4rfilIgJcbenviVFRKISqHGtT7UafqcTQsxVjJoqfryeA8PlzKcDhnMQxHpgz
gBy30pz0EoM1nMQYa00OqkCI8EFTW0zg86xd2Xn6EzAoiJyK2hnOxemQlhlupmTjaIsLeie+g4qF
O5C/is4/LYWjxC7wQ2SfUOf9m0f+saU4oqwckwTNM4VME9937oLSDF3fFzXUFXXHri4ChbwxGFMa
YJlsku/sg+dAMWTEMQMl2ntSP3fFsQrj6hpP36Y3V3F9P05Y3wODE7dRnpTMw1pv+Mu49hw48zmq
2szXeZ6MFLJ8hNjH5dVWpFpayuIAi/SPsyqgp3Sz1CtCjOy/fXt4pBnO7AJ1tAKQSia6g4fJ+Kdp
cDMlsZ/zen7+Cm55QJAdYfdd8i3YFbe/5tZkTZhMP7MyLckAv4XurVnKy6FabA68JReOOkUbNmBg
DOPRABUCBnD+wbUbsdPP/YXIrH/8DGynnGBLyuFD0/aQ/DMS2ZJqNPbhVrTZTRUl/oaS35EGDXgI
mWXOWpLbA8CUvWYW7ate4SGqoTyKniH6GwWHv11EK/nScSukM3KY673yWEDBK18kqnCv5BiG2AIQ
xoHUJxUkEnBTA1DsT3fphqEOoKBwUx1OwnDavQkgW82S5sXOFpOzsxvyFegFcd8+0JSFsjNk7amD
IE7M4Py7SNB2iLY7ybMt08mPoMLAFekz3GXkrNhOvKwaQLvow+WI6rXlLpGK43V3bbYNmei0nEY/
+i6trZzX1IDTHRODJ9sG2Kf6PlehxyseYtDAcw6Q9aryR2iIqCZEkOweCLDqGxVpTyZ7vfX+MuCW
4kBc9jc98FdfWKdGhHlshCGKS881GKGIAoyY4Myx9awEi/UQtWCa2eo/wNcymlbUAZxwgYynwD9p
RcyLiLVq5Ay72/jsGv4ULs7Rk3wywT/mKtHjL19MxPFHdSqnmkFujgySlwNZA+5yRPHiarfr5v7y
mvc8EG+dUD9jxw2+NG/GdFq112+3y1gdV+bpgQkcvoaAXUbFa11bv6w/LIdMy9MR0ZXhVjPtDLm2
/ZTS3vXaOTg+9UK0zWoyP6TTgH8QgeOU64rXSKhoFB+EX7nHJ3mfCNwwkmVp+dBmLU8jhrM+Afgu
rJAT0HtmF/+d15c6bmwBoVmRbR0iwH4tdrsmlqo6ws6tFPSpPJ7G194WZ0yjk4q+svM1HQwyy2BG
egmIxnS4e5+j8JSCB2KK/d8mvL5u98Gy2ps7GxF6Sf+0WzNjwf3pFC3egnbg6xt4MRgjlwpm1qBI
6sExNsGGYzV763Z/C60myXTQdCTZfARYiuW6rAx4hwI2Efhhcw/roOhaEmMrL0XmTki5fjNMiB7p
CEWGhnz6Qbv/J0ky2mHqXgovm8ex/aduHw2V31N8oUeQ8B/hC7N7TnDaP1z3g2R4yAJq3WrOinUr
xM/3Xr0TrKahILHcJkdoIerVD1OYcvgbW0kyz3/WQOsPZgKqqIeUPYaYSMuUuYGuo5UWQei44EJK
GvY6pKH5/k5eNTpnHOI6SXuLyn1YrxVVonbEnF+Vyl8Om8QjYKV5d7kRl9M6+GruUND2IBtiZi6D
BDjnqvxEcnTDeKe8uZkpEmWu60JoxVgUhvYQobmRriwa5R4r8cqSlKkMNUsKxQYjZWf44Ec2wtWz
sBI6BJvfQFi3OE1IBusDTqoN9hKQ4Qcbm7LbT4KSiNqZsAiW7ZiPbSZHSFG16T2mB97lBlskTrRd
wCn6TQPqgcAX+OVNvAUdSZbwHWZwI/BlwDpbgmHSg+l/3wEUMBv4DgkBgktNvSPLBXf6n2G3oCet
IWAIFQVZOxHI2RTR2a9kTQbZ8bil3GXX0Te0s9BaVt7bFOyOI5JOI6jVGEZDV16+MxADjtQQ+/f/
EB6cxzjxEGnjjdn1RQV1GLmIySBoM+PiEqvqV7IAKXWOM+gIhRrTA89IVtHzRvnLYFLTgjq1LN+M
LB2HYP0CWTEiOuwqX14ywNZaPGWsrWbC8AVsyh+S3TkHZdE7JxiPp5oO55WjlI3A9Aevn96MPF6v
hltVLOcakya+EYvfeH/YAiU5ukFzDTy92SBB/7sGtLK7PV8FgSosbKbc6gD6hjdvzsx8q3riYPqS
wBP2lNEjvDBU0lAimMSyqzP+s6uGGAyTP+ezIJHq6iWrybzjDs5xjhLE/Ll+VDZ0M7xaL8eQSb+6
vIv9llffu66aUPPRETLtVp/+PZUmr0oBOFSuwnDZDZrAqSAbbl5yQ7jKt2szxoYADbRLDDGW7HAx
nYWj6379NwsZTzhF5jv6XOoKsvqMxr3OjSBr2gh/bqPa3Vp3ojJyV0qohIfBbb4loh9ILJrjBDvX
C8mDRFHaoJqNTcsBQBKyhvPYoBoCt7/eOBBi5vZlkC6Rf6p0uNHMnio5xhzHmJnvbDjHE1K0gOVK
u0bz5b3I4i9ayFZl5NHnONwDbbuszOdVDFfHHWNs6kIpYp9eFkB6tiYGu9hcaVc00wBQifmkzi23
xSqzGdy9cegr+66JqCGYiZ/V5xggtjEbZPozeVHJDIj/mcovTiGyXrEecPVyE4gpVraToumZ+vwo
qQXIggQQ0d4Tbb+kY6QWHKGjTq9X1Omh8b54n+v2W4JNAOPbflfw78cebxyLw+CgLYeMnpP4YGo3
Wj05yCotDvrvLFHyf5kP4NONjgk9j2p7bZhvGg8ifcTpTlP0RCmB8A43wAHL3i3LhaHEb5/TtH7q
0xa4VkeeQwFSR+mkB3YGp2ye6ya0sqlCUI6zOeJgcFVy01EhHlFpazomMQxKccH3oV0safwbe2bv
zV/6DMcQij+lf1frYavig0bj4HD/e5XfrTLRLHTwLNmUtdZiLGZOQ+5+wGzfDxctOep6B+cwn8fH
Od5s4QUaDiZXsGJelLn7JVLI8e4M6iHVb/j11OWLLITFpyTwTqZHJsh7jBMiY7WhNVy9LjGR615T
0oNElSkmYbMCy8srwkRouiAV0u4TRKeDI3Gvbj1qU06L2Z2ukZJHb1xEwg4vwBEa2FKA0b4G1mjy
qjyH5HztQvcqq/kKNqFcFP2fyMylF3ybmsc96zrMS4tJ8mqIjHpX/U7WiYLagRLZjKxv3GAH8r2N
lOnQbqdKBuWwpEWyz2qx9toZiKEdE2lBXWmpbAnhvzXauCTLWPb4j0qBthMQUkZTcmnNiqjptY0o
03LYhSsjUjxbkwwcNTP1iAt2hC/fIr0rbiVizj/nY/c1cybFTZffGXCAYuy5ha9dT5qSgaztdRMm
/a4tyB+gbjzOwhZCEpO5AsUVmlQl3pFs9VysdvmK87pIO/hOH4Gzw3RQgNPLL354DtQoAq5nMa7b
/8LbD4z4kBdSfydTkglxMyHOpDMnEbpaT3ysEYCFf3whijncLUoBWm2j6m5Tc9U7UmLq1bcoY4fA
bKl2Z0oVtUIsqInmVk6ELmNpiXzReYJaQnGc3j6w978g64CWxSeOdJxSBkEgGxnpKfXE4XbngmzS
2xzDZoyA5XHTyLaVt0YqMOIGlpAC/PQ2r2SmQfCVTuTSYpoS7jGIOPoGWsStRj6jaz1l0xjQvtzT
sLBRCtN+uLyE+MWuobeibPZNeKr55RdCaCqR/qZgjfbshro8yWVQ6JBjjwsiNhjaGNoeHE2F3BiQ
8vG2jXtTwgRD1CCDtWJQW2hw0YmMSyBOBXk2b6XuIxdMfM81IbQ+6w3is8WiZXB23LnPkw9c8Dxy
54JPMlF2gWvPeHfy6oEpl/iyTnZnY/dAtO/dq5LVsTKKp2Y8AKHRoo1d3H5Z5uzKAVnenNUBeih0
H4ZNM5DWUngKo+KaGutDwRt/0vFe2r5bgVSBNJU4XKrnJrok4lEmDlIhkzt1VxNJoZQu8crLrGmI
TccXBVvmSivUL1RPaos2X5/sFswbB1fJr6XDP+W0ifUo/7dB0Z8BMdSzRVj+J8Xa10pNIy5+D93l
ED0UJqGwpG8qWlg0NUC1rFYO64oYb3yp82pv/R3R3Zn4h4IZ2DhD3VOJyAxgcCJizFVcaIY01D1y
rsorUV0EtlUIy9XKltTW5deo6TnHvci3YMiXMJ/Q3R7Aggss8i0AN1VoaqL/F87IMPDNZIxD8FnR
QAXLL6CJu/JZFfBkh8pzMlNOc4bOVDwksrBfspd+j7E7QZehls8nhiZ5zMOlp3OzOF/s6uAGDIFo
BQ96zNsFT9IUCV1ZINMNWjbAJ7TLgCRHrIYTq4iexcIFHoNGJbcU2cLtgSinft3CVvUCIBDs6ZcP
EzoayF0Zl2BCqyqvBwtDwebkH11sEPUcJ3EtsDDa1s8KCMfxPA4WFfGBAWCr4YHkowqxLyH0mTIt
NpVsNtm6BohG/TnW0U4ZkqgoA184hProfFRTbB+uti08tn9g0zdzh0B3V3CQq2adfdCwDLyXkuXJ
VrPtNTe2d/jA7rITNnHDX3EsrEJepVaqhSKzx7j75Xs0FncCtCSrM2rYnYNz3dXxiONXlzOHVyIy
ptFKB1JSfvIaRnkyJAx7nO7XLz9z+/srV6oyQNG+JpMmb2+1PSj+FzVQLuLCned1vAypt/e7uw/Y
QEdKlXfK3fiDivQ6WLZDKpIml8yOYW5xc4gl3l+YRDA/LruKZPmMzramlvWguiTdfeVpmqIsYCno
3LiDl0OlsLcj/NDdCbOSDn0ybeEnPjKWM3wvjOaKi58O2XPK6z06I/2cgDze7QTT6BomDGS33JQE
397J3O1Teep/czMT6w1hTptFe/Z1JOoqkMbzik4JiyHQl/KsijQ/zP2qNqCPk2LWdbURwVU3nwOW
7lqqmcO8sPSuoYWbGyNkKPgNt8l6ceI3g7LUMvy/iZifsOcggh67Ybsmi6p6Q79wfQadAg4qBR4R
yIJ1SQ4YUB4LJ4IXORzvo+qYqLSl+6FH2yP7SFCUQr3/KZDPASk8w8Xb7xkYW7gupa+fHoAXmrok
naaSD1jCqtaVMn4rkCMYJzoZGwOOy4Z3RBgWyGfnu8H3JQQGqYbOeD/lWCeJT3zNjFZhGeRtV8sL
PhUtyr/AvmmjabWRBLvSVVwSzsznYZl1PnYEhLn0O5uqW1VopnVuo1bAj0tn3RsNkK1jaxTBkG5z
TdLUSgIq7hJcJKrAYKhRaSMg/Xtpecno8bKiD+2eP1mch9l1QWAoMkUJnhzkwIg/E+S6HUjlY4Dq
m6bBak4RM2Os1xNy2mnPZVPRUf2Lh+s26cndn+lAnq8UPh4UkQPVoTX21GTy8OnG4sq6EFEbWJOa
UE/DMkVSBTTS8uXukbviqWHVctp5L4YAhc8jVPsB9KeBTrmQVgwc9YNmUFlu62ogHow9GtAgMzCf
GVmeKJpv2Xg5cGQ0fi3A448ftQisYKfHeJq9O3ov4whY1d+4dAlzcN6HOO23rsaYQdsUbKVSS4Cs
4nJ3k74aZuITLOWTyZUCcNP2xRiCLUc8La2WEYsEORWOA53Je/Yq+hXn7DrW4EKCnjUW1uFgXL7b
5vWdFnRC42o72SJprmOef2YQ8qyE9F6fldt7jbAB0MsmcpB1fvhAR95ouQ+0xNh5N0nOMCpO+N/8
zZcOzRZmVl36Hqo9WrLclMZnPUQCBDI62T6nxIg7kwRfRM1LBwoD/XpCbwQRIqV5PFrPoAWAK4+9
RnSEMyjM7YUxdTyGl3FHSXUjbE+CG50/JUg14W/UH75MjKiBHCJ/Y9gNuQXu7AQA0yui+0U8RBJm
gStwUqlQkBCRIqFPjlDGKkhPMdl1l2+9dNJbovLBdOV8SlDD3/Raoil4j+T97tX6Uj39bNYbxtjk
nVxvftLEpTinHUqBmawcwtAhssqitLS7Z1N179ZcbXnijLzXxfRDQb0FTw2N2n4nslG2o5uiTZVy
DHIFCG54Tz/3jF/3wpsyqKE4w6ick6WkBvbVSvrj5bdDuTLtNKcxy/mNFUcfO6pmtN8l1V8jFUaj
jb8UP1gm9lm62VbTadZTCbPntsyJRSWmksQCIFOeXfiCP5gXxV50Azb9F46xq/BBFjYAh5z5Xn3K
VwHM2dFDAzAL0d6noeRd0moa08+O5UszeU/9EYg1ddIwzS0tQy7rmvmAkQ98rLOB9rzjxujBoXOb
d/QetY8wmTsZ5Bq7uZvJvxbzfJql2UViCQGMM90pEeiqEeR/5NGoH4fHP0t9Aq02KD98S610Ip/l
VjoyQKZwqFAo8L7z47idfkj9DqlUtsNl1s8cMR8yWg+eS0N5K767t4aTL620hqXO+Ccs/fF5lF+K
+mG9RK/PdyHLUBHMqDsmqROwoV2SHo/nlomeglIBYHRavV1qG0HjYVr9L47OPLw92koipJSvVHDb
SF+B7t1aESJHH+sOs/743WEJc+Sz4q6nr06LrMEwswweOAyWeCBcc3ISTY/2mgkvQalHBwBBT8ls
+6rEQ/epI4AXh/XwowXx9/Jc9q/PPbBPZNlEZt8nOZ/Q27S7Kl+F97Bjc9VXRfhqQjH5nd9FB2Ok
iALAJ9EILVZspAJFimz+0KpvafuNq35sB3f0pafYqCRUJk3n1qwYbKSHbDfBoJMQ93ghZ3EFYfC4
d3yCfUd8qN33FeCyphwKd0s7SjFdpQ0O/ANx3bDrEzGeaMOg6fZ509FvLmnoof4IptYXzG5q0ynf
JacxyMjPBYeCiEOLPP3jps5Sle3bq4s3nhI/uWclANR1mIqlxrCfGELaHaHhqbcc261yImnks0yB
7W20E91xle0PpvRvTJmLMzFOhkcC66aorJOzhYDz7IJhTLbzx1ItvYIW7785gEaEUuxGMTohBsEj
UPb2dKNAPDS3amxbmHGm1lPIAUhfHo602SNz3gUb5OqmvNL6Kdbl76n8CdqOFH48W7WI2ZqpsO1B
7XYqkO3qQ0Sd3KtU0/pI4BYhy1qaugdSv+iRZUlY+CPDuwrXIeM9rZtWbrBF+y07PbEEPT54Zfll
L3eNB53PZkqtS4yv6YQ2f7F7/npiscdUYSf5Ijbf3pWka924W6M7sUBg8G9OE+8+cucZxspraGXR
7o0+qS7TBYCPLovkJrzsof0cDZfrKq736EuDnYWZIYu8/B1pm2R28oWU2UUfv/6V0P/9ob04NqP7
V7eRHNaj6IS/V6uL8wdwD8ocJZBLoJ4hiqXqsMhNUeVhS3zj3F7TE851RpijvQY/1afb+UBRW6bm
l/Se/koUWR0A1o+sN8fPVdXXoGR8rGAcmv+XJ9GGr2RXD0AGQKxBHqgwZAr5halijmC4XASaKfj2
dRlYv9V8h3iFRsL5LRrGpFCypC/R+hHy65/AqyMHfB9EyKggQqeBnfZfgf/4l3hZp4i3y8Oo+bh+
MOZwx8qCt4DsP4wq1MZWWM0Le5fBegLQO4DOXrhuCl5FqLr9QN0U0VEy/cwZ0HsOPED14Y9CCmm2
9AnEG2n5eRECrtk7+hvP+LZNYYrOE2sa7JVpLjYunlMXlQcVzTxgwOkEIjqwOmsDRkVW+e6P0Wmq
ukIV+shlv0+xwHWprjY8sxyzyioTmBXY23gaI/I8F8unKUb5im1VdVjIXypXXP/+xSYrTtCKbASW
4mUMJi0UZaLzMsLDtzxdu++idk+MSrxPWF9fIhOLAhX+cGwnih4KlnP8EJ4ulzYsyUcho10IB8EN
81D5+h5dIKNEFtH0i2noQBeEnIuQ8XM2NuZ3tf65e/Us37K8/myzjzvVv9rebzUlE9BVDfNGCzcQ
WH+zVpkkJU73yvk788iGbLmZtBZZdLGJQqvYfrRNVR2Kd+8qKihkIUtrK+lATF8O8mAmgBRbbtRH
oeYwrs3J3RdYhEvVMsiuGi3KBcZCcFCfKpTEWqCIHhmbr7ALsLO66ETiHLG1U8p3hd2SVHzWz80k
thOjYkU+S9Ia4hsYj1FewHVqID74lBoAPKo8p6vw+F7NfxCBWsnlDSMhXTmpDjrI3HUZGl+sVbZe
25CMY9bzKjBI+9Wxv/Z4umX2cZls8I7pHRUZee5mNXd9PfQnX2DoBn3gBS3o0ITwePcyWYCtwl3M
AgUmDY7mMXmPsxVooLtWZ2rrWSfRQ9OHvmtOx0K23bG2ewqRQxWD5h70jLJ6VYLxaiTzH0i1NwF5
6qouX9+BSYK5nKA8NBMNAzh6tI5/MI0eDHuoaTawcqK+Z5thWhfUKvo3rlzWmu0zUQPfTr8svTyu
dmezTTQP0fRRbYOZt6S2Thw7aLERd9pgBsHikDLkmSCLTJfl9jKLXtzrmLNyIF0XE027UPCXd6h7
8AT9Q0drEEmtLTaRL0y0tL4qoeqfK5kPLVpwmQUMw8P6K238I/mqG2y7Xlx1zMC7+N0H+/qL3MYB
6HMIDaarTpGZ5J8mipT1krN9OPm0W4zb9enG6lNQdybUU0W9YLOe9sCYerRqFk2EG2mrDhrVi1jn
y7mb/iKqvA0M8opujUzzfkoGg5TEvPkvWT6RfVd5KO6gyMKX4asZFfr7Hkb3ZOOCMcnvrQMFu2DU
XgZMMjB1nB3aFWlhv5I8A2FfdDyZ7LTZe8VLDAKcPEWre7rDoJpkV6lMfvvMlWLUKuaDxndFFC8D
vVKZORPX6E9N7PjD6Dc7DfYGBluM1U5f6fIXhwuqRIpW5oFXEZP/TC8uQVgyOYpRsSduR8ry05gd
gEW7mhSskcjxOCs/2fWq2BKhpChzk+k28jOYvgRV7dhWSPIWWrMkR55yZtl636F/3RqDuEHq9wnz
EJq2rGUvZP2EItSqfSGIbm3LbY6cNjfIzRwdIcyaG44lHMK9ctfjlhV3zIPbIHeUNT7dYuHhqPxi
XDCUsZ7rZfWxGin0kBZz2d8W/rpyHsI4w5adImq5k6V3melZaPKOVEzAdMKj9VJAFseVK3+DsL+D
PpzYUw78WFxvXLkMQcl/JtCNhRTdKyOqYw3HI30WYnKEsnW+wVbfjtmIMuXtjLZWCMpGnBOvOHXw
4SKqZw/b19o3Yel8RuaFHOVZeq4IP68E5hqwPPJSvc6by3H2xLpSZPcX8hI2mg25bCh8CDBN5uDF
JQJIzu2vJb6Ziv20mLqZ8uUXb7KqEJYKajXH5a/wnafev+s60d2X3x3YW6UBg6kU3YQ5ZQ94FMeo
rD0QI9+W9wtRSbu41A9S30mV2IxhN3p8j1VxGDDcvuVCdnkeErr96pYT1Gc0IhrWTxY2+54KHH/K
TUrYTLEE2U7k35tCgfEgrEisbST1Cl8QNib3YhI0EJwu39cL7zVe4d1ArH2Wl1E+0E0QxWC2ntrJ
yxgc+IZE3soXnfjIF63BPEWAdXQd7jlfvGWKbhs3RwVc6ePAANVVl9+kQRh5YsAhzfCzJblh6z10
IlvjTM3gkoqgDqVJDLD2orBbO4AqXuf6iunTDbG9QWOBUpDKyqsoeiCg1l+Ko9FiTlzR+WtZD3Hk
54YFi5crgjneXuTYd8OSkur4GX0YSqIxpWTfuOiKUDg3nym0697oytGCBDbL47ezq/ct7z9LWtAQ
JxplnW/HTJR3OASxr6Up8W2SUNqRDY83+ShwpEL3BYfqLae42/MkxXAI3BQ2roqjOUgsGMii6HzY
Z7M51Latcl0LPxGaURb4LF9jl9ChZjJznK6yek/cSobuoYuTjcR4VrC+p01OaIRGtogj7/OgdoE2
S/Tz21IL9KzLqyH7D5ZgkL6NtL3UFaK3KlFew3idWe8pKJBD/wnm36/lXrT51WaU6QVgqdlc8EZN
oWXsPDzLhKk4d+6Uykj5bXHRNX6ZfzJLufonrK/BcSi9zILOUsPNAaAiiAHi7x8BuoiMI1ft92Ex
KMz0EQXgzVCtCJ0RKiGO+E/VR3ryrdWanTXUdLz4Fkphhv4C16TT8yvN+UBb5YnfobbQXh3yICHA
tY4pfOSswhCvBZNyAheUAjMM8kR3XSk0RVb5B4/XdPTMWJHWB9e8Da+MLpRf/AMaANhYy6Cy7fCN
gxFY3Rbo6jYOfIhs7qeuQHYntiMg8FEEe2JIqx/0jwdPi6ApFzrFfK1D/LzU/Jv6sJG/R8A6pcI0
tOyJEUSm73PzKRq+NIcB/pbQIuJBBJWihvzsHjnxlMccb4ctV60u5EeB24CplNqjGGW4hXe1kE73
hKEtiIN3T4UEiHspGZEGJLYQCoFSkmmzg2Xg4D0vD5xk0EJ6guXTI1DVlk3j642ae0pI3FeueFBA
dmDT/hdwNLL/kxlT4KSzei+tMO1E6D/T4SzGCSw861COiHsibpC9t5aj/UEUylktsl3erwihlqIm
tkY4XFFClz1dlJWN0jC8/19f06DyjIRYnjOajELrAziE6UvLVLJyvKm/RJwvyOz6uiGrAuAFoObB
1p3DrgcNpFAngXhOOy0xMX1+Yb8cj6gmI3Kfc8h/fFDqafRY3f8cU7tUQHG8FXR3NWg5Wp2s5xVe
P4LfguEKkOfB9SXLzYH5wR6J/e42YgfHol1whNYPOspx89eKGu3qiQBAoty7xH70j/Qd5EPcweay
x0fXPVseNIm/BDhzzctQloQIW8FCDbewksOZOO27sCjuIBSwPX2IITau8e7OkJlHVAx+eWb6M84B
YhhK/4on3y9R1p48cJbG27TtRoeNExh7Rd944zoykrVQboqttXiavWTOxobJU6y17DRFHy0kA2RA
V7wq9zJPZGJoh01o82686uFh5pCXJDxppIl/bGd7TxQt2wq4Fl7W4hxiR+r/I8ysfPnCR51prTHF
w8XqdvQaBh6nMVA1gQvzlvPMYtvvH5tB0nhgzDSSV9wvRhyKtL6Bf/CAGrERrJm5XmBRhhFbMLxA
XpTDgaKBpRI163D71ncuiOTmP1JXlCkSJ+j1mGXNBdALN0gHbHucp3eMF2fjfodhyf9rGwql2TI/
1P7vKnQEnJiPHG9WoWMCApHuuVR50eahFjxRsFoRtmtQh+ANf5y6n4z9RgGwaSwlo1hi3Qr/XPnz
CenHQh59K+aS6yPsSrfQDsXWb6Z3EG8kkDNj2bFeZGQb/8ZeRyUdrNG21aWFb2NZwdR9ouA+rdRx
KSK6CQUimBMAizWBJosrKvwxfCobxrVcBztlUnmpEBQuq0U0fNKfxKEiW2vWsfQl048PddISl/iF
HuT7EKvChtC+1M1Htc5fhE9WPwKYPy6tMYyqZc+3ty2fG51JbHXk7DTfp34TlSsp597yckVkGw8y
A5vazu7B3zJ9ugb6GFIfmUq/RW04GZxLrfXMx5pRhUp76Z2GzVNEAnGrPq3a1xxmvaWpdUzaZWVA
q3rhitOycmdisknwblkdIplgo7o4ToeJWYK9rdlhsd1Te+x+Mk9JjylIei7qIzA0SYjlv24Ts6Bt
ySMKCOGjtU3Os0y4tJ6iFBjT5nFlWZCzo5dVEacxlrrNAGFiF+SwDr2WtK/vjTMEZ2tCgSdk/Hiu
Qpq3d2QUPdNQUwrdRvvugiXU5ViyC8Qi14wBe9ur2+71JIBqvdTKG7WJa0JaGCOUSEkSEUIWdZiB
Z9sUT9XQ5HX0NrW3NCxiaVrfr/o7hAUiv++pXqA710mqsQ3zyUzErhSv6j7mmW/7fdMNkNoLPH9h
6PWJuCBbDgwLF9qhBrW/mXl8TKR0ra1jDGMEfLGUqbWsngf0zQSXwdQT+6hgwBy2tjIE2RmwewaA
z9DX2htTskx5/MuPMfOTi08PEGNR1f0mHWV6K9fSRt9YMbWCe9m446xUba3Kilrv70d2xm4JLeOv
lL6umGfhY7etf30BRKhDgoBo4dDRjfsH9B8TvBcCi1Nx2yfmYTZXi+w26iItwwenJ6sgGCfaJb9S
UqFUDZl4BmlQGUY1oTCXud7Q8YtGz1gcFKJweWLVenn5dYc/XalpVYz11Tj7+RN8SG/CKEViK7rx
6n3cjomRUoLqeB0A34J/mj0/sJMZ1kSyU0kbBXAa0oyYOEaCxvjn+pkkr18oLMPcOAbnRa8VDAMO
Fo2IxvC+fPR8zQtN9wB04DKNt2aM1hkFm7hDuwZz93dXeHm0Q3B+w244xyI6kQ7PC2MQcUdkV7a+
Unfz94xa4ym11l2hdKwYEYfHsqRi7WD7evV3egc5V0ew7ai+cb1zJSqcTp3fblzx4zFOTb1y5lRu
/ZRWfaoC7GssB5SKEdlfmhIFdANZ22z333zWFbYQs5QTXdHoewn+RLwe5Vzu+2b+jzrR+oT6rbVs
WNUYYLiqcaAYBB8X4HOq/rCt89BN20vgFGEwTiphirOvVFVUVFr2Ji1Cv1dGGeXZdX73y1k/Xijs
PvjvweJgAzpIAULN03UUxymHCjx7UiP5UTENIuD6uN6AxBjMzdAE3c7/Mu6Oj2moiIh4WxDgvvhM
csEcWG1H9g0/YZ7LxXIvpSZCxfbf6v9W126RY9TJ5woQsm6cQHtkuYDT3toGv27S4RJy3ZNgoQ8k
lrOcvdeskd3ULPWRU6vf2h6kpg7zHBMlG66ZvDA3a3nEjTOZPUeKfJBddK5eCwCeHNRPmDdDgpp8
hMy0fivoVchYnMuBW6Wa1VD62etSuqfdVSuReQTs3efgaOC+LSvGTaX9898VJgb6C0h6qTZfFG21
LWGYw5UqbOAn6X/Feuga56/aWC8CL83+gaqr9eOZqM14weg/2QgdU21iWyR3UDut4rbfD2HNjQLP
WsM4AY08fiOwLp69JyavGc8yytGf3jgq/ALlaycnxObVTrJKT+rojBhN6aDaILSaFbsfP8GVmIIJ
9bEvL9V1UkKIQg/dQ4FIo+1TZkbCbxHRafFEgTWadNNvtmJbrGl7/2AAOEYPhys4cqLmd4zUEk0U
kMxpPQ8LMEVjewJIV5O8aGU9HTyvNrnDGJ6nQRGEp2c83lzBY1gyFzAo2g6tXM0Wot3XEZWIQt5w
Jwvxf7RhVqy7p5OHBKYrHmQXMFMF0FHfLaqtuNqf1u9iRr6jrVqXUDrlFLNGtMBqF1gWKmymMnso
yYkwbeiL5/a+ug975s5nRrwX68O/DgS+yXVG3Pr/tEBDb1Whu+53jIPKKfbiFxewYEqr427I3vvR
yFHKRv6yG3sErBl/dGtpxS1a/BiKr3o53sXPAjAFF8OdyJMNxNrT0O7/vu/y4x72KmWkjBH6tUgs
tUca6b/kRgow/SccTmyAE4QH9kTYBUxlqvgHzTrRwaXkM41mJpaJ6nY0Fytx/Lo2c1L7p45jk55i
d7z/QEe1wBJ+6W7vm2/sGgYPp/Z6qy/vvVlbh6KBoYNGzkTFYO821kHn+w7+T1vgHuhB9HmbFY+O
5qkxi/zdljh0LGRbKPQyTo2exjXXm+85rmFKTW+uZcN9t4BIJfA0RiYkOmRihIzKuRFzIWX2MU19
c4zZ9wOYrbS4jogW/eQW4nz0si0W4cQ4OTD3nrqvQtHTYENStk8Aeokwjhtsqs+C039pir0MH3XH
QG+iCJ2UeUbXft8OWkLjQiIZNehTA5E0hA8g1uVpfV7ea6NEbzzusxF/vv9nQnSxG/PWX1YZx5Em
HgfiajIxF+DHX141z0s0O6Nv2+Bp4k4JVS3CF36I6x3dm2RoVzBgChvGYpKa+2gt3t//svQUKUoZ
jpa+9CzLP1KNBtzZCILiBn4Jiovk/vnSHPTam6kmkqpNw8EC2XE0/CKnUU1YiiFqHulOjiqfEUE9
CteJ6o6bIJ77TtYqn2h0h1sSOt48/pjpcOFl39ognlDkEkYlkJOyeA54OWGOKWAIUH4yMyFKIl1U
nqhlJx9yIngjgzW903+kEpzDmTTqqxuepIQJwV+ua4701aejKatnmpIdVjJJvNYY8T5tts7wrVwf
QsObWvP+qVaFLPqyGa38XaD53ErXcDiW6VLPXTdY/cMjC3IXdOQIJlPm1cCJaUgWGoRs7n8Q0zrm
kpoKfwTGTYjjY3gBVVIbk8Xsju5wQonTUEi/YGuJU08G6gMm45G+Sq0FM6utRGfD+tM3o+VC+BDC
jsrBbz+6PC8YWpvSUI6VvsFzoV/aHkSsrmyW9PO9Q1E/Gqge6L2VB+UwMsBSt/3Yv+JuC0+rQ1WS
bUz8grRuqwO1vFSk0VI7u/8AXU3HaEgEgc+7zDI9GqGyKUkHQ7ZoBm/uzqT0n4bxTig2oZ9MN6sk
xonixmV2ULSEtD2XaH0tCzBVhItyJD7mRMJa3Og40R4/Oj4VPKXO/Fb4IwQG2TaU5sFRcSGvJInU
S3AI6Ef0HY2CDJ6vF3/450F/+0MyHUWpOktWStF8X5UT0pQqBx8lnesIf3Yor2lOzEJzy+EFZ1F7
X4792AvSj8dOa0bDVLQZuZyi8qmCDIOUt5oMUc6zLkssAdQFR/YdG68oOCgShOTCkJST4ST3f4wM
oHzyZ4O/NJd1+fSNAPsFZIWtArAfV4jfjTJKkt/9AlzIkyTK9b8Pyx1bliX12y20s/OEhGFpjAl0
JNYM+XaJWCHOa7+WIDSJHGCK1+UkaU7R4GWLY9tiCLUqSjM5pC6lSVeAgcmQGQYmZ1bBy03++sz3
beqI+sl1z+kDtdI2jsF8FmoE0Ni/3fRupnCocj69qjB7p9Nx7347UqnQht7fYfxfjQor8tOy53Xh
lK8KHmPVRPvgPKWjV6OFs5Cfi5GVcIOwc7WpFqlfkblNYUtQtJx6oWQqf7+J/sqV1cS+NQ/9squj
uKdn0pcoRnyoN0yUkE/WBJzf+KpaVysTizzkK1eE4iQtHVIRtbS7yE1onZc3qldDhnmTWJiBiZlX
X33dd6WLxEJEIU9Upp9PzH8OtyY/O47Uq/aV7G4zZnbiZkoMQAPXdGfnBwCBtK33BuXw83yZirwG
P2VD5SS3dr5Ts/Ts+sYKvq7/7CnIkxJbjd3rxyM6WKRoOOA3ljikpqvjVIOeJByzrXN+U/c4TJ+z
ftnyz8FHRrvyxz4e2BRoRpU1Oi0dZoaaaYpg63nfMTQZwfTTSjCX3NfbLyZDrkGV/hs5ABl9Hu/1
csd7Yrg+ewBebfQoaxJtmX1fURvnMbgouqV2ofIMTTfQZVcemaH4PWRJYXlizLB1MXs/00keEpXG
QMa/BM19UVe/rqpNNpoO1zibqgdUQvkV1M7fb4lJmNnYP+89/4RM8s44u1TL9dpL06zm3TpCZfup
GMSEISBF+QqVYZnuxQ1BTJMmK2gmXdFqiN8w/bzZufTSQ60wGWlCuqha1GBjmnbXGhm5QnZbCRB0
zKlv0W/QwP3P4teAp9yEwV9MBpusUgp+xDc47oDUN7TPCrDbtB8w1AtR4awX0+TqfmQ7yM00sqyF
h5Fg9Ip0iYQmAoDSa8waDxQI2PatYc5nK/VkCOs7AA7OT8GyC9ctiDt50mfWQSHyeNj0oCx256NN
ZtjhDslnhAsn6l9fi/TR41sKCrN6o3CSo/8iaIRraFpbHo+07U5MQTXbg+v7VwmAo8rA6iM9942q
WIFU5TZ2sEZPYFOk/FxBKpUdsVDVPqD7YGRtx06z04t/+P27g1wiMzI5dYFTrM8wGKbfuT/k6/82
iQLUOoL8DXlltkhpqKJlrjnUpaZhwejAM6noheCZYNu5k3BNAUf+FJL40RQegtkz7xJd9hLCmkaj
JRS23qn8PJWWPyyUaSyKiqmAMtTxZaR/avjFYRVJU1Y3SowBObhnPwlLW5mtqDc+qKZ1lTBvqAyY
4VqvJ/5EarWYJxP7F7SHHV0A7BRETSQl8Bb/esEEU8qx2m1GzhLUA5KOmnSyAPjdLK0pY+c1aUXf
Ywc8RBCrJv5svJFVpTturoUpsdIUMZTUUB6S2l45bMpgpGzOKydV9Nwlc+lZLBBuVFuuWcvN6qZz
RTwO72KPMT/EIjPOQOXZlwi6sW58qjaYILJgfbApeSjUtyxdx0pcBoMFgrXdQysq7v8taKDu5sdL
q3Y/eXbPpI48s25LHVRo+GWI+M/P1ORMWYFGDPsTrXP0RF+e4QuCDtqIm1ewEbE0+3w92THozZQv
hmVCoppSFYeH+sgC7sXebPMGScapwmFlLbRXXr8XPwWKrslQyQHmO3EvfZwj9bGANzEZ8SIQyNEQ
JUmk0uYAON7gaY0erukNl5rrjACU1PMoeT/am4dwNtV8WfV2w8UJWzSox9va9d81Ehl8jtXKlwia
IQyDfquTe6QM9Y/x5XlFioXLJzhj6oisJXnBis3R8W0rF5cc7S0wPqolh10PPC+ePT7kIqCfkYrw
7a4A9PpykbPYvxpSFQ18LsI+Dc1iuPiIi/a5PESoqXwImSm9n1cRMOEpVr7H99PB8JA9F4S+m+u1
fZTm4a2lU3XqjRJVbqw5A9alaZ2e9u+4XHwebhzoT9+KnfsHSALtRPxSbcmke/KFZcmXl65fDL7+
BRUdyghDjHu5c1iDDDqxDQoKjaVPIK+IY5i7dLVzorIvpAFIgWjg8da3b0S+UCulXbNhixfQNZMO
4uURkYmca9oOJuwYNNoWl2NhJc6L2nwY4bYGBuQpTx3Zgk9xvKRS01sI4z8Y7bCjlZtheorXWAfa
6SB4fmKUAAsZbaJCgIUuBrtqDl0jmrTI4ENlffvHEHi0Kz4yIBrJfHxk4UQnzwrf1nd+flSWksAj
SJDtKiS56xy1JDEgLqrQxeiU9GVe2tFji+38eUnb/XJQT/mPlqorZltXtzxaKo/kYTTdhS1XFOgp
DgejYZ8tDrL4b8K0pMOhU5mWcldi8cwggp2Tpx/xUVDE7ppNByxTDKIrhUnzC6vgoDVFUzvH1JD9
0rCd4JhYI9TiHIs0eX5FtF2EOtAKraAPnlukoEIqj6Etif6ZTSuOXxnsOxWqwlkvvfLo6U7pC4Fh
JFNz/IzTDuYo6Xdbea4k4X+yk1UHemvyHADP7Rri2I+P/0EVhtXkRVRFP5F+RUcgl0OiLS+jG1/O
RwgTjn+PBjGOID9nAll94NaEwgUGiWpOysyzfrXjteY/773LgXn5P4a8ENq1sdzDmfiZoZD5AtFe
7vS95e7CyyHjabsldxLtAJR50Co/DieOHESIQJCTQluc+vTD600IsQgVtjfMrfme6U2pA45Nk1xL
fJmcEWq4OrxMyRxWLqwSRkq7zDotrbZuQF1715AXDAzm3iPhduNTR0BzbQdrGP1Ie4FbqTgM0FAE
/+FmgmRo/ya51ynQfSNw1xWp0ImPhxnuyiy7Myl+t9b+h0F5UQZyK9XYpV5nWKuioo8igJlNg3JB
NhlYwqwO5AcCv9/DKCni7PS+J534Xjf7RX3kbdJZuacidcAgHqaXdWH7sep3vCrioqUGoTQaPSDW
nwf+75/AYHp0ICp/y9d41QDElkdmB3usfXvpbd1XGDi93BYSFaJ8aZEbsJ0XIu7RNYfp8fcRIZM4
2Wtffe3bFmV/FS3TGGmDFfUZwAS2lufso7wzh9htMu2SBIfO+WN5IvoanZL0zAUa6+GT14ZESJRW
M/S1BmKLDVLi32zhgWv/9mVfjxy5V/eYWhC38Ya8tYTXgiM33b2Uyto456amLNsYRWtMdDdc4hiB
z4hP3kdftPiG854N9LtdTa+1KrC5aO8+qN9H19m6A5Mv/ZSpn0evFLdYxZaqcg23N2B2OTfra6ej
BjGKn34Kqg9HKgLorO151jRC28eYHNZbQT3HWJ7UAickfBFkCQIIWHOenuLC9g6lGL4toaVkXcZo
CHzYtWaphcZssDOAL4p8T2jTiP2m481aW6wsI7IXKE8mRbbPaIT21SwVGHgNq3mieGvk6/TrKtnZ
ksD5fFXZancPMYpRqYgIus0EiR9KtBAhO6/IUXjZoV8tGv9yZbWK7Qux5VrUdJVV3g2TGlvRI4zb
goQPsMt9Qs4zjiY8XuGjI9uM19OzO/O8EhWPcWvzPzjqns1hv7DLDI/m5pEdNHA0pbI7P1im36Mw
aFPHmjN0jZ/dfX3KP9Z5VGXSbvisdSA6Q3qA2wYh/BWEGgdLU50yi+Z0Dn6bMzydR5q2RCYUq4iB
ZJNQ66JeqKeQNNadrjYyZ1PQ2sWudUo1X4RVFrUkiPmGby5fIDpOpXYqneLIBfC8UyBcGn14deTu
o7kB3wHktVIzX4qxcCxTr9LmOdCII9yJMfmRfDWkNSj7sFiPDVjShamAEOQT3oifnoqMd9xDx2PI
cZFHGR//JT+JJ/PYUSnFjGK77yGUHhWh6fJGNA0LNcDIxAAdgT3Zfox62nO0zqMqm4JavVFpOdWq
pHKi8A5XiTfQddTy3P/DKpBtSiI5RROqAP7LacQ5e55ByUL/Lz4biHzNyYijChA/x02oyAOUTguz
v5jueuusttfb5J8paP2AO7/tfbaHKP0sA3wAkG1tudalZD+oDPySpuplaiKs/bSz1pYvDywTgfr8
sfUFSNuDwh1zug6MEzuYWjOZoTs7v51/qTXFZeH+DFwy5ayXl9hr0/U9hUDeaEr63CPBCwqS6DpF
C1GlP8fB6gfl4JYHMNd0EtmoeVdk0aFeR4bA/Kdm0QzofzLEBiGGF+hUfEaqxINJdeQRM0afFfVq
+sGPK4WZz/3HXUFliRkcbsz/++v49agT7b+OdCo9uIvlkgE1hWE89n8A/zjKYPohVI4/CyidzT6A
Pab6vlSrwgjwCgIOHRExwgsHi45nSjIS9OyQkSPCWllcj+is/7N3J2jfNwiHe6I9hFpBN3vNRHVb
ofn2QI0h4fwa4G30+1jZasa65jUn6CTt227QQhxdxdpB1JQCgAmp3nRN6lD36ti3KHr8ZZ4kSEVI
ViVRuaIlxSo/itbt9B+YZotY4gIl/vAo5eUsldv8tbFgYCzKFmMaUT4GzuiFwM7ufXS3GuoTa+6r
hTSGzzHTAX11Bbifss3Ewn2u4FcRsErTPb3symsjsG1/1hR2A5IPE/CAv8YomYbJzyqiODOyZpee
DK+JqhXX9SGJRTC1la56O9kODatC5q/rTbvgq8re6zskMTwwiT4zP70gS7e1lhMQ1b4vBiZpEVu9
d6+lPTWtlbRF42AmXdgN/xNZcVJve43dQjRNrhtToDuNnZ1ki8G9V25yxRFIMO+p611YelpvNick
tMdsGBUifSrJ+9m5AJa+YdtK2RJYNhKoCU0N/6nvegqCiHy2DtDtU2MuTbzx6y3MdqpEUWt0W927
mp93lzn9itVNFPJYnTAqkpoOjZ9SgYlDfvvjhyZV7v5ZAFpqdq4pQ0RBIV6Upjz/rPAFXeeuAotv
/lftVV43JqwNUuwxYkb3gWkjtXyr+gBGyLWi2qtFrN0a1+Go/lgppw03dhyNbEZ6YLVRS4s9JDVV
WRAVIOP3EmlT5aosBHRtgZEadVwFzmlNDVc/PGHSaJHiyR7hN7gzlGssnbi/ebdCsd+x5GJWs7nU
xHtcW8JUn6cyH8df97VPHIwUrcOPWbyDd8xyz3Jn9s8Jaj5lE4iJCDt34mftBYD/MR3Rllzvy3OP
5LS88pKnz+8x8XCpDjN01TM4ZKYGcAWPuU2616x3+/QwSdav336nEgtlBPYFrd6yTvb3RsPLhgMB
Iz6299ZilBtaygJEWgdSGxd839YpTIL7W29G6BrYCXlx0l2r2AgHRcAMFdq5XuLx6E/v+qQrxsuD
MCQH8LUrMkGB0HBj/fLwdkSzGPasQZXeDDwHRveLJX5R7pW81rAqwzb1DU9fZBIzy1+cmHY1ij56
mXVJJJ4VozCtfDBrxloj12GjH6nyQISCzRY/uKUmyT6We3/ECMPLHKXu7yl90DR6E/b2PbJOktr/
ADqT0bpQqYEE1mFK3xxtw+rwChtI35WnM78QLNPQvOpwfqJRDDO4Cgqdj3KB5iXcogjVYCOF8Qsr
PrzoXrvtuNIM2Qz5J5XxcjVSCFr29fu/mzyTGcJqUULt51THoMqyapFjVc/y1L/xoZSbnbfbWpij
btiKzmSi/XG41snL8H4vhtqbgGl3Pq0WizORysjV6VcsrULmaisqnPJb4PgIBuXlgS5aGQGJfvpC
x4Naapml0qVmdzrvy1uHGfLKTX1oi9DzaGLdXA5iafizp9EF2fwEVIIeEUEymxZlP7hqqaR76eeJ
m2rz/33yzrkxoZcmz9f2xvD7gLoHTutBUtV3+VS3L0x5FKwZEnGFJRLJTXWoAuRy+qu22SfSssRI
/w0poTve330DFHcV3bLyL/dXheZDsvQ2SGB+bGj6OQ2EDT99ZXQZvozMpTI89i028LuyZnqHfnhZ
mF2rsXzQ3lISrot/OC2PuNwKHZXO51nnMj2he5zPIzP8dGZx5jeUsMptcIg5wGxOqkHra71gy7Zd
2LEr3P5z19JMC/Hg9HCRyH76lrhcQQVWuUV0ToowHhqFK7kBr/NdoipfA71wiqO2BBb4E7/kc13Q
jGmavr3rnGmDFRCEP0/0jhJL3ekpyFdp7BsJforrMz5SuQiwsvQCXTnfDl362XB88sdpzNMtrUbD
Kr+p008/0BS0HS7XXOuJvwj9oAHFoWwyZwLoS+KS/ipcsEaE1juGJwlgbJ8Bu7DodIHhAxh3uKT7
cDH/Bk4MNxRNy076h3f+m/hLMPbemyhMnbDN/l/bQ0wzvs7AP77QPlJP7yudeXcI+AfqjOjtRL4F
H+4XP3aP13NjKhEoqlRx4Id8ppFM0Crp3O8hITSkxZ06ZTAoO4wF+q1p6uQ3SLLo9duo3wgBINo9
8Bqe7o7G64xVcASPdoo9UqiM+xlW5sSdGEA7ecnCAwQpK7NjeQkw/BLC0tWHjy63bFAa+vkay1Y2
+K3NUkHe9wO59m1Ma08nIsbBw6AGu/bxfORukj8SADZtaiVZsuiayFeMVu0WJRG/NMAhWS6wNzWh
nMUT1ozTySuMDAsiSWrRlZYgWZhDI3oXRxwZilLPJhGmj+50dcrOHkMbxFk/V+ZaBJS8xrFUeypA
AehdzLCndrLMpegTNA0UPoXXDLQ4HYRqU3iSro3kl/3ei80T9pAO3uGrADcNEpT2rGbtzmxgVgGt
72boYxpK2vjTr2CY1lkwbP4SDpoc5fINoxdPJ+hTMPXHCHlYC/XmS8yhSQr7Bbb/teNZFmmkDH/z
UnPx6wYmasjpACTrKZIMJpgAnFw607TaiFhBFQPrk2LytsK+agsmF6PETFpAkGgVg2q/tnW+Do+s
7gEhngEiCZ47syNO48KCWCWPy6XhHWbN6cpspwvDbi8zhYbciFrWLUN2mOF8MBsKXxt3VijA0w/c
q0KW30vFE0a+UIwaTEBQBRdO10CS/4rPv8zB0Ad3P3TiRuowfsoQC2ypSXEElzHp0OlwmugED4dv
Fpo7jbKdwU5WKXcTSiXYTkFxG5mN1kQetCfX4MpUTa7Q/aU2CgKqgn4EMhfV0DcHOotXKArEG6eO
eorfLtI4b90mwKM7Ci+RKxNg9bgiIt9XR4GZgPK8sLQe3f7p9r+BYkwxm8epejGHylgwPMkPkzxl
nhDiRW+8sTfFAJ2sni7LyeVOIAiWJFdVT0FhCgqsoskBlQQgT6WRETAQB7jn2PMXISQNQN/5pI8F
GrDHV4mGfeXo4phJvO9Rpp/Jnk0gdA13cM3kPARgUAuHw/XDh6X8+wF0fYrhOzPPeAh90sBHz+k5
F+FNSQEzyU83oayc5qJVLflx1Us47zF6/IxuI+qn1BG8YHyCSSTsKbSZvKVTXDmDugRxFAfVtl+G
YOq/VnFCLSHsbUCMj/iyx2AA+1G7Oh56c8pMsJFadKeOiV09/vCYZvUPmRU6Pymz6emkMcsPQIip
Euf8xxuKuPkURqyT2pCR7zP8iTeTSdeSjw8BLdHOloUt0teFVgoNwmcRN5acAUXbrErEB7sgjtHH
G0deMAd4ddTW/Cqc8NF4WTM5Tsw/a+LjzmoqsGBh05EXgM/zq6QvQRwDoI/GigzPeNTdhFJ8IKVk
8+Ll52lWVQ5A9kWXOAR2hvqAUfWXUD4JqM3xsn742QDj5MbhkfUDN02cYMii1qpjz7fBFk3EVCH1
PwIuLobqeuoAZZJkNvlG2wBzpOU8AV12ZYDips7o+jn8LqcdQXJC6QdkRqqjRodpFIbaaNe8EmFA
UTssU6KD0UZwohd9DT7VZ0cwCz0/5rnouMz8wEoMZmUbqPXKV0lL0PVMPwANAp+UWC2g8MoUJpME
6DFxI3yCL4K2COkqm7teB1YS5goWkqd4t8L2tKpOh4c34L7k75Dtvao4cm9wPWJ6xkiXECxHHjrE
23vHBggpIQ17zuRDqth7wqzS+DFPuSXxOYp91r+Lezdg5JiA3+3Ixiot45lvLDSDuIJKEXYKgdeD
nZ106cJAcENaxgKt9VG/3iRRl5NXjTrsCwqqvZbYRtgcXIfRngJj+gStiYJ9neXzbRC/iQtNh+YC
RsT3S9BsitKByTeMq9DDk9+Iir5im82tM0/KymoqHi58Yl8k/ETZY07XrnhHoa/dKey4F35e8kHX
A2vtQNtHnh8Y4/ZT5u0/8xCu6swTlcybP7CuGjvANTPv80tMvHg/H8GXYtDxvdupJarSEROs1Fyj
acOqCzHUZJ8d7X0zfTxXYaFm1bBOy5CcBrs0Hudpf9EZMt3NJsJ9bjRoWBUHG6u+LpZVc4aO/9Tn
Oha7AuCbgHVKJmtLyabjTE1e70fTtDuaAq0e/XojcoCZOLXXPcXsUlLXJpctD1efJYSuvK7h9NvI
ojvR4/tgLb0uMf4ePlR4d6vDt8p7MgPJKmfhZIRiF7MiKWfvIKzZzDJGTqPSJQxT3Sb1kP1mXFT9
Fwp5e3SDkm12FQFluBam2z6b5mJvCMuU9ahDNDH3jfkEku4cYpinbW1B6EaNRgJh2QsiGNrYL6b7
MPcC7BEKyNVR2zcuPfKIxKvxc6FKjMdhWoJTeCp+6qJT7xByRtk4+t9RpSZnGMinxXAtiRWFE1Yx
EauN9smc3F6+Xi6LAFkud6G4Sf0tdhKnvJn/tTi4n8Mbe2IrVOu7VB4KAw6xGI0txBb8tfBxdKn3
U5WgG25ZsW1RxYnktcLvbxE/DhcYq0Q5F1SAnmOB//x6SnpQ8JqbXrydsmHJW8Hg/ywNnkPKBOg0
ynh6TaTWSdnIjK4bECqug90ss8lXLAJ4Iu8jcYWq5G10fPEIIp4yBrlIFLmdtOHOSv1/Ft0unkmr
4Uo7+YWw7GUoQMo8WoBgpyh/N+Ft+IajI3L/2PmHB+iHsZKo6spHm3WtEvzuIUcdfpKfN+OaoYDN
jW74LRE2ObrLX3wT5U/l00hnBgCeAKSid+VklVzwe2Efc8e12+FcYkMLol99vCDHCEEsrRolQjf8
gJqkb+soHhYm7VcQVP+sWjp25XHaMnLMb5x+V8kHAmlIRk21JmwpI1So252Xz+XgCJFOFZwkSWSQ
Do8JpB+1uXPASJhcZo8KmbGCJItukLEpZ7p7Ss/9IZSxTVLzPVg256whNpa/goMnS4ghM1o76y5r
KHw+U67N7ETUpR8Fw5/W3kpXpRTOu2taAy5GNuO31UNT1Svgtfips9k09xLuhHA5sM+DMMd/6UOs
gNkblOWLC/AjF1daRTrOphdnNwFBt15CpEg1EeRJX0ZF/xdClKtWhhOhlVrWtRA4KLbe5VNsZP7F
Rl0iV7mTWAxjRLo7Od/1FlWJ/b0oM9W3lv4u3iU3n3CgaI18YTUyPhH4FJXh6OboBeBhcvR+1RbD
nRFNXwZlT2lauhU+aNnjepUd3gLtknFwUDulsd0jM0jpPdFXXTG2PKOqQotOg48D510G9nqL5Mpt
ekxzcGs3L9Rc/TVAjj6ytbiJbgPAwjUTRInG4/4s8TdDpMvA815Qu5wbbwB3O+1qfoJCMiQOutD0
XJbJryyWJMV0DIiiF5U9kKp+UcOuWiT8SOEBJ+pgDzJ1xBfJFPBSCi25XlxwCRMQvUWws1hX8G1H
wqe68PRpzOXLQ/McwjQ6fAXMU1hHFcg/YFOzdBb/nqA3w+2YB1feMRuNNVG4dGyEjOsYuNz8SaXX
4Fnjl2JnQnrul6Nfgv69S8gtFfFASlggtiSFKuQFh5Ix1v9SvqKVgpicn+3XqvHH3hiCNVdKyAvl
ygg6E6U503PAdfmIpcIaiq8ERNY9NhbnxmqCEcn/13tfhGCuC+RSZBrhG6y/uLcErNP7diceufT/
FZwzt6sY5MajSK/eR+7Ey7ArJ8Ab8qrMqFuDcTpcl99LGbqBw7eT4Xep3ZtjEm0xutaDBHpmfthp
nUkwQq3XO0it2vyn4OMDZ7CtnSF/7j3S8ETmrjEm5Q0ziVxg0qYtQIsqZQi+7VJnScMGp7SVzd7C
lFcJqDmYM2ZMUNz4dsX8i3AK51+5UMjX1On7tErNjdd8gXbi3cLgf0PD8xwKBKfLh49AQ9e55WF6
0WpBv0gd3cHqwwRONwo/t4c9J0V9RV8PpVyvWVMUINyI6Uuw+a7RLXlM5A6uk+35JSf++xjY7dYg
O9xpEunpbkr+to8x3EbtQ/C1LK75oMha4tSn2QoIaPpQVDr5ulwC1v3XEbSO/4ZL3dLihX7wY7Ve
/4aDv4oeI7+QOlASjJBoELlU7v8vhKcSHwOkPRvB8oc8qIQYA2p3tpvQTagL0DSJ+YRUmQNLqCh0
iKSXYjDTa+Gh58vywsgFEaA4mxu6P+5Bu6VMXmFIWzlSR2B9m6r8bkSHnOHANz//xUMPigzHeV3b
pmidcOkjVCQ19vxULDlOaZqMWfGnq9DTz2tScqh4Zjb1JEMeSf5edchc2qr6NiYXV1/T1kbSrfFT
smpgv+m7CVQRo5PtWOPEfF4WWlFI7InUML+lH/1whgrXe0khQC6TH8wQhu5CKJUAAqWFUFdY6Sf7
v7zUOINxUmTkyJBbNeaaqM6SxfFoNX4lIQkFm0lvhZYsg81WJoPfHmwzAr/7lAbBZIynrEWEWNCz
KJLBGno79v2CfSGARJN6OtvGMt7iPZ1vbW/QjIJelQqzjaXfRtm8+i052pY9QsUjN0YKFViSWhVW
0ZwnV0ogNdSU8k8O4GKaWdSZ1oRRP+9qUja5ro0nsC61pAF+1zzPPBYJGbarIR+RIZR2pr+ipxHU
NqUNecLE3qdNEWm30f53o+v/ssmc+Y15FjdTVibebo7hEoWKcAGg+kYwd82NmO0nvsR+vKIO+EQP
bkwetVjI44EAHATFU44GD/6nIvNdYndBljmnrVGIIFtDVMJvFfbnV54Y0B8+w7sLCrR7eMWtReHc
uKZhK2LlQdTKMlvHJGmq8lwReU12uhivkDq1wk5mI4t+r+s56Wqs+pPnfLSzRd5JSrCcLi7qPEAH
NLw9FdSEufAVBDPweayQNzq9uRgCUCpNpGOF7f2dPBvx44mOCSSSh82Yde8Vr0Furgc2clr9BPGS
NyQSP5oD23jm7ISsJtuhNT+1yhuh8wPnpIUJ5+z35Tf4fVckC+Ww3cs3D7DCA8U2VtG4V9WnLZC9
GmiexvqCN9pufYNO9XgHo2Ntn9kGuYOoE0JOf5oZrHIrWKRC0xKlwPoArKXytH9svWZ/NSCDnuta
j+mW9GR6thF0/yDfVUExunBEigNVzel0Vh0EE0Ak9ecwwoop9wNJeLnln5p/U6KjzKYTT8Ysm4V7
EVnLzgM/OIYFdupVN7D5grGTueziZ/+dzSrIPj5OEPbTdQzeWAplNPc6B35qUrZ7aTCOvEArjDiy
3edARuYVnT0zyhUPTZCGL0PiYmdU84vY9F7HRoFzknYY2/gkltn7W80f+O32nsq7GYlAn8mGNHB/
u1if/hrZyYSZsgkc8KoWDCgqed2Bg17fuLw5mi4yNUQV0spms29jrJyezymq9UCL8rLhKxSK4pKz
0ZeOpS9sIXupi4R5s5FcfwmtNj309I6YwiFsOHwmGzfG17XTywxqq7/Szn5Z/TYjPoHw7eVmFYKR
eo6C9ltFmEAjd5rWRrVfXL00TPCrT5CA3zpTIC9Cz6Bglg+D3RBQ62nDefZIq5YScNBufUc8QdJl
tlN3AMFtFU8Ns3/VgC3MARvq1Dylcpccfuo9qYtE25w2Tpa+0jfbHVnjN/IUx9eWFxOZeEpRLvNQ
aOzomZZV8KAVZEJTKmzYqTcin6uul+rISC08pbmxLxrGTRXgJXbCytS+3oLKpY+szX9P2WBTB+95
0jHelHaGOEfyKBd3kEj1E5td50hPiO9ioVSMkJm4BMJ87fR97n7jWvRNEc3hxczlnBHfMeDNIoFw
FRFBCyHhE4FaqgejWUi+A+4dqVR+eeURe15+raW2nnScRe2yeEd/V+9iEgFX2vYS88XOluGu7b19
AJuRky93wd9a7ppqP+InSdKB+M+3hmj3jzC3FPI0SlcdnPofMiJx3w/AizvsbKMRBk7ii8HQqE4d
nqgpG417G+LuYxGioPYNpJFawwEHLY1gOUxEfynnj8JZ3tTBpHZArJyyxXbELbUQTIJnK3ReE8ue
IPP+x3OFSLqBWi2eDJgDtlyyPFt8JO+nBjIg15a2PSCH3HHkQZuIVVvDdn9DFX8Lr7JDkYOg30Hn
Wfm+Te3bTJ64TLD9Zld6owxPLtvFxdDQU0Se/aoTva7ZNOP375WccQ87LgHZdyKodmlvKwRHm5ad
zq2QNiVIFCRlyPwrmNrpNhK4L+y5iun8F8NdB9TmoPPlrZlFCc4+RjqZ919u7zv4XNWqncMAd8F4
anqMRxUWcaZ9FzFwgt+xNOc3oZ2q443tJVcJBkZbXI0KjUYgQVPAyE+gQzgOlUTGTrpjtEW+AW+5
I1zC2vbcKBgKEQqGcN8GURXufx+cEMHOsIDC7D8AT6lM+vkJkiXyYzqNMXxfTc98amyEnVw1KLCx
OnjHhe0U+8d87S9M7nxnzmx7hmNaBJ9W6tKSQn3csmMbTMO6SYxvbVk1mCMo/Wye+ubHAqMer9Hv
LqzarXLKOb6/UrolhmGp4tWkJLeCFYtaUnAVYlE7w5MtYWvdNUm6ZiFGslH6BosdLkiFF1pJeQZN
GwPaXIRK6Wlu1nkEo541C/KCTg3HWQeTo5ntprAoVQ7Za+U7sGZmbxM4hQs02hbNcYOFD5bGt0QI
FPdYlmDHljzdY7XYgILJPm5TkUovsBm2vJ3P6KpqyA0x2BpLFvcUuLHos9w4iCmYhoUsmJqO+dP3
lPY9DzhUunjbwxfS+TB9boXur1jjDbxYIDdsHHHBpWHVrj92a9XZsyyOmaB9IiByV6XfcGiuaxEh
3hz1Ql8Rltu8nm1vzUwkspUXgfwB2w4TbD06QkZbCdvYZyjl8ej4skYZzVDk4nsmoAUtHzbBj2fC
BgT2+Ay9oiL2PcpRa2PNrpztwikg9RSXh7yfMELeC8QlEY4qv2CXCLenrQU8oFycFmjSzw6PVpGD
7Nc4FQQzhQRxukPsosftuS+pu/cOFetbf7Be0r+lVyuk569EE0cGfXFBzmq1qo94cBInNzyzTSdq
Kz2j9gLNxQjdw/7D4ERFOGa3z4loUFIaFthLSKVZ+85s8x6nQM6QWMqrT8efBZFtwXstFxkbWPys
FiH/dK9RyDoX4dKwIf+x9BgwzcNeGWrCC8DsRGDegBXjthBzq7ihEpNAAnHPpxcYQxmXL6uvtFCB
rM7WsRh3jR3T8jy+PNE/qLlf/5bDeVh2gH+5Og3VNe5bjExc7aRI/4DuJFD+10wgRd0Tw4WGoAWv
EbPmAb2rudAXeQP/+zXohJu8YLMm9UYIx78KY/e4TPzrGwPd1SrYmPlrAnsyNg5jYF6XPGaQ9dZG
0V/myi3Jmh0HonRXQrvREfqlYx0Asw6CmovQeR2dmJDAyXcD5NWNkGDq5s4Waeq3rNMczLvFmTTz
RQKXHpvb2SNi+dBhFUD1rY7Xeja9FIkYrsC77UCYMH0wWBpDGkvu24wRdtyg0qI2jT6Bc1zwL8wv
8X38Wp6fmoWbyHgItC//FMUKr/OnN8uQpmMpDcGWKQApL6RRaSNGNzuRjQlBWKu8PKpwcbRqqET5
ujWC/svPwUkULB1h6VbVEV4vkSF6oQ5BezTRt0Pto1j+N6PcTuvfFM5aiyQ5UwMnc/Jw3NarkUZ1
t7O+PIb6zTUvXIZytU70ZfxEPPMo4EYpK8UrWWBblnEr/TanP/5GE/0nL8JpjSXSm3NxMSEA1dax
HNrpkhSJCbxe9GJwFlmoiEFFBvWI5fqZPxoqz6urjhXt3X3IkdeQ9ynHpabAcGgh2z793xpo2YUE
FZVdKxlShYqMD0qa004Q6/P0C7Q7aQ19b5sC/7vlXPEx7RNrbws6GEEoMpL0AU2Jwec9ec/YLiDD
iWJwIc3moty9PHITRsT1CjGmb+nMoSgM7gO8a1Iv/IbQyoSVXHlPBFx4YehRSj7XgW091tnjiKPx
6tFHclyX7zpdUSnilhiJAEJKQhf0JrWsntv7uLysvAxHqloaNPp/r19j73NrEM/OQbx8DICpT7dk
bpKRMZqY6hoG1WimgbYKd4AVSQcaj8Y1cg7W8eZUaJXYjRR3S80gBzGu7mvvDrdjNnuorx6ozTO/
NLv5SChXNOHEqKHDBclE3Nrul98OambXCEDCOaJqwroyErzvfa0v8vYMlNqQry0DXRWDshGnRKx+
+FKhJ6IMVMJ8YvlBdz3N4yCoKqSTsNdkH/10uVQk/kGlXw6hfz8NmQugikUq4hvLRJfxOWJkJCgx
37Rb7Zbaiu5y6ru3HwEGwdfsBWJjJg/jF8zdS3nCQ/aPpe+kHTgrUaSxSmSEMWS02tVxJ+JQ9fGs
s5nEbZZ7e+BebgJ951X5osRVd2RjkPvv1vZjgagqybC3aOW+zCag/XAexEKtXCe39ig4F/Egr30W
cI1j/XuN/GZ8AZW+RO8ZvkKPtdtRrUdSZd6sGHyW1ABAK40QatpHlTZRsGdfrgJl3ibr6CHuWFmj
GekDtskOq4g8kG/WVeUSuvHrKI9K4u9wPcsCbyFLvifUAgLTJ0sq8XeBZDhzQ0XuYKHwDwYKdkHt
47i+cwH1J9f8TJW2NVraodfia7jd4qWH9bdCW0agg6NLsbK3BPmokZRTwgKYvrvneWtdkYGLjcDg
CQR9UJQ85gMMFS7UHzfXQm8wCP1Lap3UqrUXb6zoxBN85VI7EDDgMFjr5BE9WhYwM60y40EX+8lC
6UBE7oOCOJRu4Y6jiJZz9eEOowt+TOqfUyd02mFn3xK30k2XRIaX0tYZubsyy7bYjJLjAWQCcMt/
WHfRdoFuoz8fuD8LDEK5Wz2XOTfz7u74i/H0H0zENliPUERce2jJ1AonjI0l66wxVr6FI983wDE3
1TF3sZRHPhzXXY++gzXjzHrdaObVLI6KIIexenlgrDIdPA9yGGRSdNES6mrKt8+IP0BWUhzQPCRM
UTu3N0CcEK4WsgbBGDx0hRVe41EFlbw8u93IyHApdL2FxhOBeZ6Ddhv3gemOFvgQeOodJJCNIk2E
gIQ4lRK5jSlhvhQ3PAMRFaxW2YAXgqydfFLIsHCcEfOwzGzgyh8j034BBdgRJ3Xffp2CtvwoY8Qv
YZ/h5fq9kRCyCi8uRtGl4aGYbwcpQlFSR3LbQrBZhVR0bCr6mXpRn0a+Wo03PbLRhgof3l/kp538
XhQzTXe8pJkSYhM0cgoUPe5ziehfVwyIwltnP9Lj4OPZd02HjelRLdKs0Vfp+tS53XzxOht3c2/G
ZqmheBDoapuu1QZE2nk/W6O4YoINMH2YsUqhMrmOGIdIKwOE1PsDjg8khs0HghfJ7TmtL8/TRr3U
HUDpSc23ewCgKSXtvqmRhHZulF7Arb1QhyJ5mvXGt/m/R/veQ1oDvqW0ckthV+Yf86SqaZoiiVQk
ccIaI2XbdHNTEgjZFru5zwDONCbSKcTDLdEUYar3Frz/J/bXgDFgM2j3ndLRdLtIOWNkQBmxw4qI
1TTP67CLY4lS+0OA4dqOUDAYR4illEbOdfoH8+x+mw2F3upyynsD4HQf52JZSaCaHEldP4/sZu4X
8zdSFiOaLLIX2RrFIJZg8fy1GCNm/EsS6KWlOur3LY1/pP3flD92gn60zDxRoIr7qUIN110VsFCC
OSupzbkEeY9JzdZW4c8G3DXExztl/wb/zOoHdtBFRNxtVGkiAvdEDwIs6Ktn5SyxFBJRMtSQDX5g
Xcy5xQtlatobSKRNPOVoZQ3rveF0dGsh0cPn/bGz793Wh9djsSUUW1CBB/K7VgDF6o5HF5EvpNmR
1LT5ywAzRcwYMS1jFJboOdrVmUl3V7wZdTvO/+zbyh4Lc3TYsuwxxdVq1okOPZxA8rn5GFuSduHP
HOIf/LA16BtEaK5CkTjk2WsX0NGKCpo3KnvANCdzdxemJLJh8gSE7fuz+rYGmeYQMLr3Ihhp2PSS
+6+1VzthgAb0nSe5z7oRYwj2eYJ4BuYu/bGUHWWz1jUA6TOdygezRGCoot5+6u8e/Za8Ml1B1quS
F9l3Tw8p2PMY7QvSkfZ2HsCdWs4fE+2hpULwi2EVeROflyyyk8C/XnNk2ASCM/d/PW2bocVLi+ax
MnGZrDz+mEh+G2jx9ncP0n9WvU2X7DGj8VuZVwh288KRWYUTTQ4g3DwrIlwV5jq55eTTFoH2DbDr
vazdsFDy4SCXl3O6QsUUQrZ/Y8GRX3WHlCRRQgRI8VNFrVsHgpIrfRZS4Ba0bHPz5Wa0b8YeHvf+
EgfXiiP3N1wXlRd8iprNSk3Jw/z6GuthDv5C7PZAzU3TTIf37g3MmNT/Q3JXLYRKNJ2K09uPfOXr
ldQvbV3xpMD7VOx+C41gq1f9fOWfui4/K87scQowT+vgz5HUAz3bLztVMo0LoTMNLv/TjbFXRoZ7
FSQtGLlwd5GS/+bqLUTBe0EJ1RECfeU4qzNN66qegstF25+NCNe7Q7YHDSn+eQb2MfMVpSs5UtqH
ZHFeTLRtYY6fzBtGFTcxROY3y8AHyzdjZUJIN7SKOtQT5JxkJK1AKboyqG9WG9F7pUMC1uTMk7kt
9bpqRfcQKAJH8xcQPPmMYfNVCZr6NHR3aGWrQFC+bvY5WiVT2ui+OEQsknE4Q1CV2Niu745eUff8
/S4vsb3Wdnbv03IFWTj0mY7yFmU/hBxwPFQeJvT75exDTPWOtmWC26en3jTMYfAANKTE/jVzRItd
FfmhZrPjruJ5nT/yH0NHG3IH7n+cHwrlECjK+G+vK85gHeOSgORLFmMqYRaR9WSAROqrbPOve6LF
ILCg8mA3qfiDqaadmVOYfaiGgBo6C4x9DLHJpu+nCJA6QoqV7cKaGmWv5cy/hmkr8EjhmJbvxtKY
iLJt1O0q5jLyERoPEqt7H9GkmAGihMopsmLrX5VBlrFDkU/kagky9CIwRO1wHUMegbfksAeiwCsk
/8CqW3xHkwQikhKuFnbITEFOpmrjJmaLyINTWEULaTZZD3lEEYg8aE+JZEcIl716wBE7lKh7HQ4v
9FD/L5/EtR1yQGfzlWkMLf03pqw60qMNhglalV1MeO/WqTmIuRzOyY4M+Z0/6tHtJSNfkRI2wasv
k2SZsKuoWEk+AiobZl3BL/deAgYcuH3cftAhKLAccZroyZwppxTfNy4/xa3noYcwz542LdAcl9Pd
219LIIjGqNif2M9u1MpmSPqNeo6q1ZTtldnnQJq5SamCjhhIEZtxGdfd7sVrMun/pP+gGQK8M4pj
atuwHHUtSjRG0Q9ObLiG94iLCuVAyHUB1I2wzcT7C4UJUms7fiycHcTsq3K2TNDGpLpjnOB9HKDP
efr2aifll/4iFnqAL7cZXk+2acA2taTbUJ7+0S2k2MHM7SJDWBdF3zHQMpM/1H7Tg6O0CoEyyrn3
4MvDLQ2bteq47s/+2RlnAVqdljku3ko28PB5I2dDxo45XquulOju81emkLsUDTWxcVD201Nf0uRu
SIUpF/q1m4s3tTa6XDIoFCDo2jktK7Q+6kyjPR+QkXbTIpj4ttEPDFcomLupUe6F+v0aYmpl2S/X
u6XTUp5swyF3e8KGWBTO0mJh64uWaeNwNDfUAR9OmdaY1aWJh+3dMNVQAwLX/HsoGxwd+ilnYHoL
4sfiC4kQ7O/lapLFnp44KhTa3GrzQ+WZ+HwlMxUBbu2AYsLHUfuBnoM/q8Au2PWgsTFmBoIra10d
ojlOBKidOevVXSNjzjxsbdP9kkrfU2SMd2F3+/WpsrgqT490THNZFtISNt27DioYTXx1UfwHJCIT
ejNbiGeeRigR2UpjaKdIZcsZZ4sUyLkFSE5c6Ap6TFO1w3spmXnKpqBGeDGB+L7wf0t8g0C29XcM
K1n98k0HlukhqhIvAc5c0B7HVUwDopT640io632QQh2GGdfuy9wy07IBzRMqnsN3iTEHR13xAXRZ
DC3zXnEnMzlDBsBKYVV9OPXf7JauTJ0A3dbeICZ92DYwXPyqBIYHOlSX+Y8rox637nuM0DA4446q
yZN2xDqIRergstPih6zmmDcK50a10/3icJqbJ6sCerQZPhyHcK7zw0dPCT3ouAYuQzOKOZOXe4so
ab9dCX/cAlT9E/6kO2ohCeiO1p1DTFNVjv9722iUkNxwKijI9C/4xCIJhsOLMblUCPx4imFVGkhW
0P+2xRc/AUYNLSoJyCp0xZQAkes1kfos6bJUPsBOuOahGM1h7nD+7AhLGMU0o1RZ4Spzz4H7MGC2
psT0mNgCZhCrevtx7TY3hMoUrL2N8bpvdYA6f6E5HQLwwLE6PnzdE7rt88ZxsuUvLaUEJkBh+6fc
ccF9qK9m2SXC5JKQ99fPwN0I1i1yV9NbPC4yqbk8yzc5CKfc84oKg4bbAky4+32kYtDBrbtaEnb1
JU5f3L09c8sOxjGeNbDiiBMG2Q31wyG+4JRKPWjCCbIBv5lzgDONAdeq//pC/hLwmOU5TxdsNQZZ
oBI0X7+KEGOQo3rW9FposD8Bj2YhhG8clnw5hekOtlNtq/y3zf30SGn4ynAhgFgLUbISb/Ufiafi
mFy+VyQTBX90bkpP4XlXZMK5GJNlGhrTyHRrV8OBAgE6iw3CSfYNxeKZObvF7JuglTqsgo6I3+K6
5tEncC9C1y01bKZf2JLVALMDE/gw7M74uW+0LJ3+nnZKym2sFJnQRUL9wbjotXFuF5T5Qp6/9wGI
qE4miNRmQDPP1d5iAjr7WmyJYmSx3dsLSdLO7TES8zR3heEVkco7CwCkQk7s8VPDNnqmyy5ZrkLU
+po0ORhSTUBc1KUWShN5DY/eDeeOS8Vd2Eu9svR0Zxp24vjKnK1Ht+NhkAo9GswgHoy6pZVKmxUb
YrAw/d+9XSm3/IEATr/cqOoZwjwRtzkvU/kfJBrb+4Hc3EKNU9lPcSNLEUy38/QS8bUNdeWawZEg
ja2nyMtKexshqk3csub2JvvC+BDFQcoVeSNsotY5SXdCKSl12uuOAwncPAwE5qJYqVdcP3I04TQC
u7wklBgGU69sTR03xCz6f1aCTwkkVjUhXR4eC6i5l+I62OU2r5eElFGFsyqBXb8LFhAZUiT7YdxN
RR1I4ZWgLKHsqHEUBoq06xLldWn217shj6VMcdRwR+liHnGEv6hiU5UkTed5s6ZYlH7/XbeHZpOa
056RtUlIadMg3yHe9YRjLtHY2GjhBMPncDOW/0d/Xu+ADNinxROumNbZUETXWcGlMMvkJgPa/rKF
7tHosDBhSvZuqmfofNS23rR33iMuXMj6HH7v0FC0YVs6r3xPM/9esLvWKUOrPDdbLpj6wR9l3ZVg
WS9ucXJUV3yhkKW+ypEK/LwFSbuzVzI3kv8sBLnrKHK1P3ZCMLJzxj+0XA26voO5kRZakMpp1UnO
dBBc/qbNObRp+n9UVZI67xWIudVUzNqfdS3GEYU4VFKI6xoB2iE0VQ1i5Wb54uAnrcs5CXkvru/d
JgEj8ysDi7Dg57X9p2LL57xbkvmt2FZSCDbDnu1HlugClv1MVK/Tc19mTacr+ek+P8ufFxvSVJ/G
d2GwYbapkuDjVuwf4mkJ0ILwrW4OZDoktpa6ulWudMEHed1cjUDICKZwczIkCwV/IYP3HNMiPmMK
k1g1Ic1Pi4SsexGGxkb2MsMDJ32IUHHrJPhptfEjlCYVqKdKakUBcZDNzPRfpkqi4+s5bT+B+azy
VavUxYLG7KqbErYTlkXknsvcVz17RHCMr77vC3gSnDZS1KhFW3RVUVEGPPTrKikGG6/Xx75LV4I9
jSWzjLzi37eDn82jXiNgKHMmvu5SLpsm3iu735sKkzjDtbLMe63E+Q+R+WLRUCP6fPR4bclYQlJf
Oh2PLvCI+LlYeV+uet5HeUWWRBFgL60PxnbBR3pi5p1hyfEGtFKV8fR6A5WUCXNOnVksIXZj2d9s
Tw+V+Nv2QyNDlVCNN/ciSS0QeBblGulJiCFIUUUiyF+V3gECckBG9ONqbFYh9TFxArr3Hmkf+mrE
k6sr/4axmenIca5nIHseZfffdsCSD9NwINzUlvcMJTWjrdrCaVK49gFEEgxJU6fDd2s7ePOpVDoG
fRpADJEVBzZN0eskeQG562sAHrxC552SJDuXGt+/1s0TqjZseNcSTQIUAKI95zz1F/5GdtNBRr1e
bjPNWJBaFlFXBKIcyEJBw8W1n7A2UIbMAxrnIXkXe9eSBaMKryJaWbc14yXmHurEQbK3FITIJ3E1
olnpRYaMxEtuM7RljNOzccthmS8pG2ExA6NWInj5NFij1ZYnB4NMA5ruUfjBKfnRoeKfs7v3OQ6r
PTsw21QqkEk1s4xFURKgzZjy0xLTaMLcB8TbZWkDm8eYowecNLZDwi4HofTjG0FUOI658RG8EsaO
9cq/WPU0aDh4wwfE2ppx/iE0Cg2ldyJ3xgaBRryivnzIMTRPS+S3AbSoL6t2hM9LD+GokfB5Ebz4
oQdE4/gMwyi/IDKVdOnmGXh5zDJzDCO17ghmVFivwLn3WPKSz5snCC3kkYCrNItYseX5ER1Viro/
6KppRbp73Ygc2Xx+KpmuLGzjMoIisb4s7q6G31yh/LcRNRUnWEMlHSmtUm7Y6po+J1OMpS9qOLUG
gQgewgMuZsTwA6HOFQ/z+qX2N5eOGDWFtkwHznF7a+60Cs9tW7+9EuyEDMYL0HY6Pb6+PAV8dH86
vVqfKnqX2+U2qLdObQ/Eac/G3il9kA4OwRdN1hbcNxCz9kxv1GSJLDHVr72kZWHjG460EE54gce6
nj2lHCs6PgsQloEGl/fchYdHaVWK/inQ4Ury8h6/rxK2Pu4AY6QaXW16maiTDTVMFbfUkLzJe1xt
rAFLRIkqJothuqfCdxQU78/mrGklTmeKoaEhM+2Xulc7RN+FjwJwaZVoEQB2GooHK9kejVgBL2aU
0C22reF2JGn9RKO2ABaXmMXx/np2Uhey2Hz3zvY909+ouTAfoG2plvQ3Umxo71IyiTndafIZ62fl
Lj/43GGIp1CLj7nSNbvLTB85fWyz4gX2qJOUZ/OqTrNeZzNv6nZBnvQYuqtEtg1ndMuokfxSIAuy
/uBw3GlEQUs1dXDNPlm78bo3whhZdmL0RKuUygREFlpGydo86F7MynW6aVgY/8en0FNDep/Tbczi
y4tRb6kD+7kg9tCMCDo4AV4ZQmUh1uKHIvc16/3OmpjSI1dIpOmMt9QTT1iJVhKpr54+tng6Y6rH
t5DzgCbF1tE8lKxMr+OaFxe5o1zShhxIjdxAULA0mn7k/DGKqPf69xZCdFistOJTi/r21/vo3DBF
qmFreYtzsK5aACzfOjHzB5R9cLaBodBxzyatOiru90siw7S2EAxAk4l+xBKWllQ2ckWKPILzMTpv
9oy2bZHQdPVzZjqF3filSdPTwLU6ekxw4jZ71N4+GcC0wHVz4+2X8nVIbFBXy8D2/fmFKdoGFzLh
t1RGqkXlf5O5tG8zMa3rZ7UsPQ2f14h88H2VtKsAVww3MVgNjKRB4yMaCP1JWC9o3hOsOxTehuwR
ArbiJoOtljszq+2F/P3vN7vpwnCQxAakupSCnzsk+J9gIO8AHfq7cP+/ccyYhNLv+ewBY1qEeCbP
sBi7DWhKOAjF+B3GPK1r/J6Sh9sDuvTjN56iuX6nsUBx4wzu9LFSffPi+GV0P1HHaSo5L0ZtAms0
MGTmOaA91mhZOODHGRUZ+jRBcKBlHjVvNk3zMAuIa3iGVqyOt9F3sMpQUFt64eOaYcOUy8tisQGu
28YXHqH7rrhLn119Mjzc5KrN9QNrShORcoYtWw5YLqtCFFx1OKdr5vu9MDliDliiQTSLrJaTWVZs
d5JUUhB5Sxks/oeHKts4H1TlnfAomr1LtxYQ08oceTYYakdSU1fSLz9rjmtMZ7ZrfoBHDf9jfNED
m9sEjBP88R6eTPR0m14xgxV8+VGho6uZ0ubEdffXd0zAsYxznl+M2R2bZhU47CAW/vckJPzoA7OZ
jZODamDRy3hwgan0h74Ljr5ArVSMEMgk3E6WAM2mnH2/eeicCmPwa7Mq+7qOZ+4c5W56UudUorko
OEF96zK6+inhh/hBPxPJ1w3YjqPHx+iaqRwbVJC+sBHqc8HY1Ef9YhhL6SWhxJLabAhsGswWSadM
ofittcYKXVlQnuhUg8BGUCCSG5X/o+XPHv78TLE26knxso6YMut8yZ/oqhM6oiV+M3LOcJiqO9P/
qcuDDGWkdLkAfqsyZO/vlPO97wWhNxtqRxwRk9oYydPXL1qQkF3eT+QgCVAcw8MoQGCvDhnwk28N
TAkRcARotZIpSsqMQyJfqU+MgukTr1uFfwLzBGTKchLHBXp7t4dM3xgtoHX6UfxSjJynNO1bEPAk
h6hJL04z7orQ4i8VHMI7NtNgq9d8czzDTls7xXBQJbpvHRWS+fj7PNPBCvW9N0hodJctv7pSYpCL
HeE5SmT1lpps7Pmr+bKmkNyLGo/7AGPzxGU2FL80s6xZZNmcU51KaUuAU+j/Iu8gg0h2KgevZJoD
uREcBP99t/uGEtRIaMzxaQJLAm9Tlkgra0sIYRNmOxU8F/Fthx6/F3zAgulOcVZZJ/fH4BRpbKpa
+Rz6lmZQIxO/Z4SKUtJEZd+xhmELxKdNiFUAmPJObxUKQLsN6SfyfLN2n7SWfV7mKjupN/8zsG0X
WZGknfCaOvpcj+msrNK+nWX8GN0vr7oQNAFtDamif4XJWscLcWL93yIwAL/cOE6RJKZmm3spBI5i
AsksDaHO2i2tp55Hin4haB7zPALrnLWpIeh3qul5/TliGNwiNK/ZuvnMsIcYrMGo4pf+V2uH3CDs
Im+ZRi3t7eVZaphPqta6Iegm0MvFYxZz7gIg4by6QJZ5BMO8wLS+fxs1YcI4pb9qau3507qpxyxF
zN3jjVd0oFdd8hyG+h76kcoY3ZVVT6AoOLkFpyWqDbkXmsFnqgre1f9FF8jGHaL23V71PSTJN5nG
3NQViOQZGJdu3g5sch8mJYzxqPf9+oxRKP3VKufIc02kc39i+/Bc00teW9MoZuZYXcqZjvPX4kLE
IUvjOBEsM+zP7I00QarkY20i+mAVq5mMo9XWltyWJ7OqeeWue2ZUOTmFimJAh4DEIu2dIa0amVDe
QB4Zhmgnalw+L97dy9cfgsJM4KcKaObhBWFX5Y8LL0xh+hbpHOFolVW+g23RZtw9Xn6sd3uXM25K
8Vr49lmPW/BmidMxGLo7owhp0RhdkIfGSjVabEn7cRxKj/2LxkGZpcR9ec1qTubLpfHGjA/Csmou
EWQlipI20kMLjRfCb2aLpVB8a0m68y9WvavUFsXJQnOq0ZW5T/p56UszC+Qin3LjyDk7Yay8egYX
xWPUvWt/XQU7eYh1AlGu/d4HOmS4Ta7qgUo9Pab2s3/IMJf49K61gqfMeNtOf07JwjQGsW6fyY/Q
F47obgA2gg4iShxA1iMJ8nXPqkL9wwyoeNO85sSGlsTKsJHonx1OtDuu42jlCdFw5pkhjJppUvZp
C77YoxgDyURxw4TFV3iyAMMOCz5PQ41OX6lF7IiA3CKRkVQnYUd7J57a7doN2iiEzAR4cct7CyKg
hlzevB53W+8Q0eQcmFhFDZ55vOzhvN30B8fCD/Gwn7F13NUsvlqGf8G1HLw3bWQvOkYRS9Xj8ove
TqXCsciPBM/4tEFrKjioSoSU2kUe4GHO5bb7SVkcYfka6wRtrJkhLBRDRhWkwLd8WO2mZVUNCxj2
H0xfnkWJbuaWMVNj1gMEJVq15reXTZmVwkjtJtOOxFqWnwgO8qclpIktgg8OEHcN2sxRfHLD8jT2
7su/rKevxQLYQryuaWPGsfwtqHoewxnojQ3Oj8jP7YL6mfkucOKTvJ6I9FmFvXkp8XhhkOT/4UwV
WYTht4BaPJ1qnj3oIeJxtSreqbjcYGtpHUuOKuOc//gktrxeSZvYwMHFUOTPgx9kJKcIuhopMzvv
5dKktTn/DN7na/nQ+YPiys3OphjwVXk8s2AVouOFLuHuFJkyHMsBBBVQJAwvw1+pGdiFWcni71Vz
lErstOK5e/0qsMbIya4VLISGcIyr15VPVZJqLJ6itFZjYmzfqrNEgXhuRyMkC/kzm/eBpdrak951
SoOnb3HlayIhiqUxUREIj6edcplUEqdvsLi2PzJ+xIkbOA9o7zw23aeE1z+n+OAfg6i8og9ti0hx
2g8sdpSRdF2TckPJTdsCrTm8sDa8dPIwOG4jSJP3/MoPfG1mTjVDRHl712T77yQ5d29lPkWRXWqU
BVR01fhyoTYcnkNG3khciqwBix7rmDlJseHYr6BvjRIYhzWMBqgVvPpjXL8sSghANsrvWoZMLz3L
RMWZLPhRUrnWCOsbJFGUqWP0F6SQkztxLXs3Knr4CRijbUWdSB3L1pxOv0LFrDkiMjWkPDPu99Y6
rNBzS9wIjQ27hdfySo8uSyQBntcwztaDCTSwM/hqYyQNelPQIt3MC0lULOkUT8VJSELZ6RC08mDp
es6cVpL/AezC2nn2RTJhcS6x8ZPvaoUnLecp/5KGkX+cBLcwiR4uadgSZFniPrCG1Lon7YQm2Rxb
GjnkhLAZvIz4QVulEbGah7z40Y+FH29z73Zo6eNBrEJ0R14CZNAr6wFeX45dvYUAxHgVtE8cltnN
Eur320EElGnOP6NTmxY0yuGcmaiC4W+vwjs2Y6CVtfdseu6/QWUAyfDFt+yKwCunaXEgUlblIsjA
aWuLPG1fxlrYJGbNcgotWI3Wrn4f633ZYYe+45hjiZBXjz8k44SrJDK8pr7ngkRsU1M6cOUskVIP
U03XXZqrtVZ1qMlm/Qs+j7bwqzKFv6WUWd55MG5z6auy5U4zxI4UNuXzC7QqypYhKerg/qZjZfOg
WF43klBJ+1VMidIsOmJGh/i1LRvVe2l8lPMgJUuqNOmIVUhky0glSnmbVdX93v2ixEis//HtSWUD
N3qtxfzWRP69BFex7rfwnsb2B03IeNUSK/a/q+3CmBIa0Zesga0rrLHwz5qIezRKp5iaYFVEJ978
kb4Cgv4sNSpRTbrSgJhP07FiKIXXPhmPcl/TpIWFVXIBnG1YadQCAZLXnmjiBBj46DGc64D7Fgv2
c7OaMlgij3l75YrO34X6HCNLg/t07FC0mEaKaAfLQszGJw/14ykJixoMosDIOt9w5zhapIJCIU2O
XcSaaw0f4pvsG7ut1bF/Jt/4K7/ewWkR2XKsRtn1G0xDcfBDZ3IWA8/4pZGg8ejNwuRI2YoWvak1
oP8EiSCNxQntbY7gnH7swmAojUt1eCIYxBzS+98QjpKtCpro7SyVSsG1pqDKO/1mItEClTq6SXgl
hB72qwxnkCcfipNeXa3DrqIs/i2KkrwDSDTQXtyB0rk2usfD3itxHExnsD3EIe881+KMwp+WN7hI
wwV6ekpzZOwt4fq+j8UorqptNVZK8gK0jyCSS9WE5nlSnRLhm449cFYMDf2yUirzPGK7gSCG1dfW
gM/A3xB3hqScC7jGK0ulNyUCcGDOjKgvhivCflGhCotNHkcCGuHSHxvYdxs4+RkDGYF/tFJ2dv4H
Paub9VhOfQlTzgNxpPht43CR+UTynpB7d6IK1NL3fjpHhhoFimR7b7mky9Tme0o9tnETQjBIWfjK
PqbJn8UlttTgJbX2MXb/Thcsjdd8sR2l+LamaaNtSzXrYlGCGmjK99MkdAKT7rJZeLqwaHMVg2SH
WMU1OP++6boiEcPfyQ0feM7OFjK5R3/Td34DCs5ORn03DIwZqyD1VYcy9cDT6bmxxp8ghQTMmj46
Gc7qEgd87AxsbKp18Dw2ADW7AznY8s+ce7SQ7Me/rtnee4PrSosythGt63vYj+P86Pyg2n43btAs
5hipBzCZYWdkWqjHASlyLhBP+dKD/4e6JSmDstyfW1SjQo65GaFC06LJLQ0Sn4jBJH+VXmTQAVhb
ePemwoPQoqKyS91qUJ6tfd2u3bP27YFm3X4hzXNyZL4yTEh4BbdxPQksLyLmVW9hTO7NTO9LmDrs
3iMHQW7bZ/iIerr4+nWO+oQ0wujN6FK/lTOMxWT0Rk5+nNpdRY7R1pKhoUpBg/ySjf3SVdQ+LIHc
cKIUjxtF4m25kD9FtjK6CryUfQIhEhSQKuxGq7jbBB4SG1+pWb90m9IVsIIVmQ5t9CYh8ZSvm1qH
1Z9kWoo4ItzcjMoiPB9m2YcyzHvNgeCTVg/R39ctUVVHv5FaRYXm9QGZNOYmfZBwO1aRago2oM4v
9YrsM2Mwa88wvPnXvjpk0iAeTtfhRpSsdnNS4rWC4yteiTr7ZhbBCp/h9Jgmx3L+NmmAqc7l5xKX
QwWA5Eomzg56JQ1ylaGkLS6TPKmWsHMjMBqtCWoi866Vq4s6MJWNhAO+uZU60FZ174nPzST7CM2X
cgKIqPpDmOfddY/3TK3fVaSULGgEOe6nQbbxwi2Yp10ONw5dk8Gx9YIwai/s+mKy2BHtvI96F1sC
/JJQRxDsOleE5+FgxFtExos76Mxpw1nVJ1/vTSPD5n7ktE1FahLgOoz6kIlaFgJTLQa8+/09wSu8
D3t9RPQNqsloHt5RF5EwboOTNufqv9DvZvi9SF1Zjt4+a2l5Wlu3HFSnkRyb7pu55Q5D40TlPEM4
gWCGyPuO0yxjUnUVnx5fL5mZpm7zeQlqpf9X/LZbvj6VZFCnPT8Fk+2eqhvQtiZ2g9jakVY3LFNj
8sAmDobGTYYl1HSweZUJkUNMugOiiPVDO8YZ4Wv/ZnjviwSHZlI6JCo6Bk1Z2ubjbpCZnAu3iP/C
fbpKmsy7+E6j7riLfgQpSozLFYZnSi2Sogn0/bVApK3NibxMMb71KZ9fNAfIraq/Eme1Ke6tBn0Z
PS7D4lrFts8mxPEjhX4SVYPRKlaIW0988LI6jzaM50w7aeanwobdVyxl13/XM4Y1TAkJ9NUqkmTx
2PfZbTayIHsvMk+I7REPZ78IKaCIRJJoynvpQsO9cJd3RBQACwMDqXfje+vLF2Ricn1sfCE5U2Y+
M0fkhYQh4x/6KypiVbwBFyt4bLXp/0c+y1MmK6S7gWm7EwizR1Mr7fY7N847kZZ0vv7VWnVaVpjA
3k8VPu1cvuHo+RG/vAnvyeYnf/x3hPgFSfBKhFnL+JDsk4KYxnqRohmcLjDMigkRA7oV4VzF1Q0u
UfNy2uLW9hFJFYkqlSn2jNNTsquh5O6FIZlsmxDI+ndSmtnmxTqWYJ3DOL4OwFha5tZ0DkLjJfMA
4NAxPXorytFevR8132fMWMXEZtQXc8GT+Z265myjKBanxcQgNh7TgPg9X2+vG/28EUTS8AEzuCyw
VpOu2AtB1+DRialalZQHS7WOkzYJ+03Zz2N3jga8EOpiqTLrBP2ltXnlAQtUYWgb3pKzJK4jQo6x
QHZKuOkO12tB3RtxTv9zv5ReuiCPL5U6yNpp+j8mkanH17IvpH82daVozQaBibJ6DGiZOSjKggZd
qjz5inkRAyvuMImTvILTDDl/yFg4UGqrbkZvLG/VOmhRODQN5gKKzr4NRg/RTzxtnOF+78DDhNlI
xUwpn/vKITqktK922dDRylZKScfkfPTr3IefJXmw9qjhoq1VJkgwcm7ukULrpQqABXQdmZdC67zS
3p7DVzDY/cDGqyy7I8dCHKzFc6jjPzZD2L2mC3D6s8QLSHGPb3yLlAo+jBpVsJ25cnupX7WyBCpN
kkvWuF3Cc23jeIPIs0CrWFiQwX/MG1tfYCJUSj+kJThple1hYIVw5tp2QzpQH74xOxV50DE+guK0
YMHDLyKe/kBmWX7/mc8ktrQUv5jJUnoBZvBFOjz3EXmQSNDQbKqjKAIIEIbZr4dM5Q8BihT5WXMa
lT099vbWPMyyfLkaICfnwqABNuB6YHPJxJJ9mvDo8/XWWiQ9zwEmA1HclXah9Ehaz/PixQ/74hqh
nEwx6fv4j6Nbvav2ISZNplCtwDltxjECgNeD8icsBP1DmREjak6a1ZhYgwjj2fA+NE5a7Y1pb6Le
TZOl4h5v5lmcIGuEG3I6RVYNRNIEwPY4k89uVZaCz+1cSyfZd+9Wrgiwa57rXsCVFsezx4MVLelV
zZJoVAt0wUIlAxJDaCCITvVeP2tZKRIOPChh2pmPhXACNzQMYqd2ctIF96mMcrNg9b2nmg4VSYmA
3yAJhHD6ZQTiYf1MT5nNAPX00wx/x32MsxmfU35etx4vVouY3cZCTC47fITOkQ3OBW7XBbtQHAgh
jgbTtOdPpUKhn7DcdVOLfQMeU1BwL8fwKvA3YuzkXR04+vE0UC6yYXHy4HpEqpYbB0QH6BXTJEEG
313+HYKnoMDmD1QnF8eqJ9ZoULqI0QDgePl/8x7cMvsNct/aF5pfvydVx8G8oSQhIVhu790amPVJ
ZfgaHRciKXyyALY7pxBcCRQOdojZXleHH2WllPyqRYLNJXb3iqp48D+NiCIDCs/w3GBWrXMYBLuG
b56VAOnGS/vauD1hX/pOerSf/326D6YOs5GMluIzMSLz2Z6WY2G99mbo/DaPGSTcShwU5EnhNSQe
QmlIX13fFxB4NDtxhpn+2uM/P22JIvR4p0fFVIQ1fHMK8c5/BgiLo/3+JX7sYHpr1dS4cein6RMw
VMt0y9xJU0YkOwDic2LGQiMJABIDisDUrw7eZZUYUIfeLt9FFiB/9ZfRClCpxwMmLDc7OxFNKkQf
S7p542cgT0EgsZ7W9J0w+LCL02dB6a0y5VgcHO6sjevsSS/5kp3BMhFqb40Pk73VW7+LpmtU6A+e
Zs0dXBhM3m4IWnRCfRRQhB6Ajntb/nO9FGgf8AC4OWSTH1JFQiKlbzZ+ZSvm+P5812fwsEotKEB9
iB6l5sepKYc3UgBMa5GpxnCFSBP0v5YkTNQKJRjqURwBpiLo1s49beji9LnvP9i6EYeL/VBcGZJP
oLbOfBptXOTZutRiEPCd1cyMjXjpTyLCC5MP7qkaol26xFzEsS3WqPdDlf1cvc9mV/2X6RqE4t5i
8DwIdQrF3cFfJV1DsQD2PYyROdIo/zcQBO4400zq4BYYEi2Z8lHpjiF82H1M3A1ipeD4m9ogFgaC
cg2yrOVJ1pwzbZYpYxwOn5LTQa24Tu6HAZ6lHTN0OUBxjCr/UiD7GLo30HohRY2N3c3r5pTXrhwy
081W2f7rGSUsrTvJidKx35W/FXR/8X/1PdCJfLYEkWZU5lr1voMkhZB+GX+sUkBxOws0rww9sBcp
Vi3ecRl8qX9xpRnotu4do823l9uGr3kqivQakLYKhMIyfAhLiVx4NSpPNTz2GAPvJ5gawoXhvEPg
iT7WXlNOQX1uzrPev4ImiwyFinfbmutK/N/iAkUYJToSQc6bIhkboUMNHynveVfZMj9QIpJ3YPJj
mKST9SnMDzT6VQkeKcMA47o3+bM24UBz+X8QhIJmJ27spQZ7x/9QYtsfOJnZdcdJCsn5ItdK2gOj
TqdKDKn0vcY1cx2nvEDxMwMjVCvzDWmOvEm0crgLrrOCUs4MsVuWxGrI5kCrA5qetf0Rk60+CjQ0
cFYSkPiqmakKCXDYe+egLmsUA/ieLnWLSPLLK73O4HJXH/OSIfRh4b3JMmgPbfeDNNxf9kjFyZ1O
Mw6MqS1stSbjZJ2zgibIRKK4iq+reLZNRwrPdyB+jmlrDkMN44pQ3PHphw4rcxIWGDyEdvaBtxYK
kZpOcQqWSo4gcHmDSl1uLiKfkVxV08FexHrWGFq0N5K5ZCUHvKuJbRtBUR3eYHlAnI7Wd4PkCCnk
T2IfEFuXhdVO1cWZsMpYHDkT14I9mKL8PE+fZEsl1i1BvGFj/ks8KrdUMmcQG7NwJuhip/1t7KXq
m4Rx/1pzscoIH1gbgh46Hm7X6fwG8Y8xfm/Az44ZOlPFcs4X5YuAFdsBhXDLe7uuwQ45ct42m3Ta
+DapBZnXsuU3dJO62MUW3KIpuddlWgYDv+DMFuHb/daH3+YmOqjkEMyauMHCJem1+A9KaD+U0oUB
4MGcQy16EDXmhF7FSvHwRwifQNXTIQtKasZyygAyC4YU9KlWjt2NH6gNGYsh+OBMoQ7Cfwrhb0OT
5mNqF1fmDEDwNIID+Ma8se38/bhp78maeFwhCHQJAdSEjbDMQOGN5/Stap67gwfsVkeGSVPYD1H1
SG0HqgIzz5a+fV46XXddy+HG8LkpTeAMOgTUbXLFKIAd6NmpMA6XHoEn/3wibtr9v834fzf7vfAW
z56Sjwc2miyMEKgrPyJoKDckA4Pr6X2rgaN4DqVPpYPMtvjpnvoWm2/8pZJY3afYbPBqq1ZlsITT
ijCRsylv/jn3UPZv6Zq+z+JLzfGM77p5smiUAZKBgj9sn7TkKV8UbWJNh38jFkCj5kpmCMYAV45K
Mx3R0xb+LDMIUD/7su7W3y3LoLotKMYoyhgz93yIl/0i6WNYLvEd6o5htVe1YVLUadURYyWsSjs6
p8jYzQhPl0ALi4ZcT0w4MKx1RhKiSOJdEsd5cXjj6/DxhWYA6yw/J9ckJzFnu4ng05RShkhlj5UD
TYOWQvO/qP3eFBjOkgBekyleNIMv9fUIONklTUyqPEjEFKTPLHf2vKvI2zq9UwJA483JWaJsTe48
QfDkb3E9tgqnwqwp4HbSmquFy1lgoIhps31lJZd5wZsuQK/R2LevvOLTBVT3Fl8Qj+uX22z4sZnP
amxJq5H7Oiu14dd0eT74n2QM4kMmjfRXT6NEL5o+wcycEEfVxsYSqbOSuvr0Yhs8wwBW+KV2uqWy
0sAn2BIvO+SRjhkB/ebqclYZZUPnATnr1leD8Mp4MmDQdSmdi+TrPEM3nzx4VRjHKPwPhovrV+s5
eOGjKi+z9suJRdeVUNWu0xGXTypJFtA6CGA46G9oyrBiVhKtDaDJq3JlYKoi5KDdDUl7TZcIM7BA
RWVXp3hO7ViJukGwPBEA86SGaRxwTCfJKYmsYEdrGgJeBKvaNcCgpWtwxPxVE2KFIy3mQRT+gS8M
JO6tuk13CGnKo3NoMxsomdkvQsGKmRMAAzbCLSqx0HRrZGP1nyxhdsmyYO3DK277esr4gpblFN+Q
wolMYufHZWVDRv+nqYZIee++xkVOomhBKt9GAdFLAuoruF1n4W/4HkW2SNM82D7lamnhHLVa53zQ
SRIScCzLV6jzfHdpmxAr8NfmaIHpbSRYfuvXMUtg14qWjwPPg0YGpQaArhi29U2X23REvfvxJOgN
oKkCuLXIK2WpBw9rYe8sxXmlsNxWJfCqebnhnNp2QwPsIDgSAPvwsUmZJJqxnL7uNE3zL986nP2q
Qu7vqSnGN8Q6jdCNvVdAXL3J2SldmLsqWHxklrB7+/VXq6tzlkU83BPmJz9SAAUfzCNv8Guwqxx3
AzxDN1G7eu2Gvwgbq9PToGQ9nRK4A/E9cvherhUL8WTnSLgIzaxcMDo7Kyvu6/4RezyVOrIh4IoR
JuTdxMSXVubROyV0Z8wa/Txvw5oeiiVhbUSo2HMdGvSBHcNCQlrwVsaMZm+mPkcvZzarf/JOpDJo
Xp03564KdhTD0rFCanXxv+B0x/8spIJaX+ugW5JaF+oM//BKuw8BfR8Bkn6C7iFmIz0/SLJ00oiK
M47WGKlhQprti74LX2QkraAi4RAYUY+7gjqhPA/otwIiSOPpy0gQcct6Q42LxKX7wL66lrPlCO5K
WCS8knXvsoj4kT3mBjUNZjdrPGt+yxY/RQ3sdcifG6x2vWq+qK4sjKfdzFuij3IiODRqv3SCX8pg
bUxOPfh92yaDWaMeoxuO/iDxlDZlTUCMCLCw9b2kZXOB9Cpkf4reiqgWz/rB7Xnhw/pDqnuM8R2e
6jgTR+n+2U5ri7+XzTDPjAp7VHLEF2TVocFyQXUdS7Aa7P66E2uHIp611bniurtxKsqBacefzJRV
JAGB+hsdfU37wxCTfYaSoAU1d+IZauoF0yMLSKRZpLiIF2/VHLVMOp/pqEAaZYW1kTya+lPUbeqR
4uSFF6Jny4vokrKKgLs9GNlNIzzGn7TR3btCFs2aTImCxHlf4TidMZfOVdyk18mWmxH0YXLWSybc
NMLSLgENvISDWe4UE2jFwbdl+4QkHGrCBnMe7+1l/WGbSWGrtYb+eRf7puWef/dZdkH51IfVy3gL
GJ+4ygZ8K1yEZKDl2KP893cH9WcOX3fYNOX0sRLWD0zNtYzbmmibfcU2WPXtbssX3HGt+stDBLVc
8a3ez1Jl89FWjWp5wBsEU+kq1yuMNoU3F/LUrFOnRSkuzbT/lLBfg5b4j3NEEzNOYVB+O2iF7f5h
8vnRgs/Pil0fZOWNKLtbSo2Ek1VnQjoT9LiRrGPHTExQkVPPVq5zBdEjle8JxaWFzIfmu4Cis8b+
KvWbpiCaO879xygGSe8QjBPYMfI0bcqpLvqLePoQNbwl+Crc3nfKEcnZlfnEZiTLhYSDuxs/uuTQ
8nRbT5nw3xYoMj/cXO1Y5JfidXzleNQRKNH503LuRpQ8SqP+4G6d3klAm/2SsoY1HC5ymAQtCgXN
7UDz02xLRH/NmVFKR9ggzBhS489U44obXle+5PtPCvj5LcJkqkFqvrwTyfGt1mRtr90bySxnyxXq
wLKw3G9/20Ww6ApcIdJ6rBDO2YKhY7IRKY4uqj5quiWe3z4Gb20jmnGERBqA9to9P+45WVpKyD31
0hIkioovlNjNobf3QS1axXrNmTVunCqcmpX16rrb1L25vsSqVtJpuWFidXoHNr1TqkATL6+8h14A
lQctsf2+cY+AXoNuiT2hW0FKC1TQP239vAwozQxxQNE2Sp2HipXVuh2Iejnr6oO3qv7DrnOkAoaQ
Aoswi382Xgl7ca3bS97ZKtxYqexXkq2H02Bg0OoMAh5bxxp2iTK4IcmGvY6DARBtewI29uPfmy25
vO73JBHMtXxoomTHu177L5KMbX2d4zEQ8/3DFbsLrsryFvFxdpuBaRCvnpbei9jIzmJU9x1n5Yjv
/Ef4SvE5Q0UM9x5L6N0crBWA9tGdLSRWHqTh5Da+zd+BMatuSsIPde7JyBUQUisB8q1BPBEutfot
VPqMKTJJIiuDPiyCkCCgb3oCeg15ctPbEZheGlVGfSfqICcPhzwDtCx6inRMthbVYzuF+kf94prI
5yU4YygWon0C7S4N57tg+c3yjzMxvVT88QFPjUYA5xpYyvrQcj1G9qJQGRiSnYuFIS2VPA8wt2Xi
flxRQjOZ72DHoxxp+dtO+RreUZ+mYHADVi6Vjgbq0HVgSWhUs0ET8eZJXZHxviy2lxhjEncRB207
X7V85r97xZDO/81y+5g7qto86lj1boyxifQXcMPYvqA2kg/jj436FyobU0YcCRsBFENDC6PJ2otP
m0aoUhzoC4nt4Re148iELa3siOsH3rXQ5Pe/sFw5A8LR5o+2PdKOlBZX3A4LAq/cUDk7o4HDQu4N
YDmL+6kp1LHelJw6NwFnGqvozD4shgZt/kaZhCIZ8nf2nqd4/T3BgRY4nFFfreVLDPj+zRHwsEXk
QS9fKTEcac3DX40MaT8xGv06l5kAkUuEGs53bNA3oyq03RmLJh9OlCqBg/bZhRmvLtTs3mGvgBi8
tZEHxz8WmrzvuYctvNm+j24/zkLBYYE6iUYEBqmZDZApEX82QwtwbqtNrOFK2feQLWCLqSW0/G2m
/BBzNfn/4JRWsbX5Ys99Bsc9qYrRA5r1YojbT19P973v3pTvMRAy1dVp/k2AXaQkYGwCM0HbOUVj
NRhCDKKld1GbV4k1M91m0uhg3nKQIWuQHl9hsvEESlZLsbteheEZdceaLgqLBkwz4L8tgL6bMfwN
yh3ANdo3ieXUFGWLxZpWvHBO3sPCWwVg22Cu5w+fN1O5VTFG2laTArRqimhEX9LVA3hawQLEd9QY
jFPxmSeDKugQ18t9oA2AG/ThWqzw8K1vBVwu4dEvQ1UwPt4FNN7NHn3PJ8k/uSOs688gIOQNE4qt
k2q/UjUEGU8wAPsfpMCFThn5eJRCquGKzPdYh+i18wXuCF9LTSpolQ17UGsaL+2xWKhZi3l09H+r
vrsBP7uuQyzXplvZWJfT4oldQ2AjV4AvXSfhY76Npuf+Pc5RStExmjeLafb5K8mOfAdKd7jP0aeD
xGagZN1ZJn/UU8g5MCbCQ2Fww1sX/w/LCyHebfKQ1+bgRbmYe4UvKM14Tx7pY8RD6Pb8+cmDeQaJ
5A27NimFdG+VLSIB96MPQ+vOipRJAm2PFQGIYA8hhjXQMGdyD37rUOw6OMVrpSKgp2bK2vq0GGSx
hdHbxVUdptEQtgGXCr1VoCJoRnQ1wlJG/1Kqu//+VcAAg/s3d1zAJauwh1gtq2d9SQBlHP2n0iCi
QOtR5SppMOOFC4/K8LB1nv9qtaXmuejiIKHnW4hJAwUnLscXWEZ1ZZGErEt/bOZALQs0s7Ivl/Qa
AT9H7KmTaiheJ2kgwiGJVok9E+5pOQay4PuGp2oyZLmTI9flrKEtLdyDfwLgB+cUOcx8jzAE8wkS
RG1WWA0FH8Fr/FyNIhQEDZTVADX6XbmoicULR2WHMFaYpv24LQASzO/d5TkOTGkk/Yak3Dxuam3o
9YoTRhARAlBsPiT1jO12RqpROqwotk6NoAfQA0OoOT+hO/9XTYDnOxSwqVp/UH8nrs0iRENE3eg5
nnzVhGNbRcnabdkU2t5KgFCG8wdeQt+b6iuOP0pXoE5fcpOWi9C1imWKzi+QbtEZy1P+UWB5v0W7
DfSqyw4TaNz9nq36oPnIz/mPo4CNRH06QJszKSuta4XRMPI7tdu9+3s9F1k9P1JuUbuAzSzVjmLD
1wZ0XRus9Nu+2TYcqX3rjR9ZOWy/UGLHaAsaIEmE8/EYuweQv9ur/6lsR0+9SDaS64zK3jcq6NfP
XsdoGt1CK9YMzNNsSbgQ1FZUkZpISIjMWXDE7BLXBlXwg54B2EEuBPLxChVIuL96rKFZgUtE03aB
5r5ADUD6cMTYJEvq6LNOwDaJTaNnT6i7gz3ln6JZsOFIPhlP3rXlBv05jMpEYjx72YkRLIDf0U1D
tK7ptVUuUwGIfTNckReDHCMw+3IRYQ+oOgGEOtO/gbxQZpb8AafROD7aYeDla2E91yCqTCxv9mby
rYrJrb/eULQeE3q/VN+QBEcf/CV8ygwF6nx+zg4qLJJpyDTboBGBzMMe/lqmf1N8YIql1CbUMofY
Ih/WxMkyUzXS7KVdsqg/eOm8sziGWC9Ku0TFQbxO/fSDyP1V/EFMDX220+p35kV4IBEvUqAVa3DA
NqZEsFMoGiNuu3bMLZuj6Yd3fEuSsyi2HA5JYbYhIqSXtwH+TxbJfLz+ZWadpTiQMU/ScbtrzZrE
RRKd+kipt9sJLTYRdKVdttxNUSsYzhcWXHm3UR+y28KwEYPd6nCnil6xn5sc5OLp0zZOeLOcKam1
LkvhgyaDVBZspFjwrJ9B7Pk6mfDNi8IIPGGMSJh597y06tlhWM9iu7AEzyl+dzVcHTTAIuiNOUMk
2GeNArG//hmO/6HLYbeOEF2hy8amcKgJCk3qTcjTfbOEPbsDKKBfCOb9jky9t26zjRmznDOxTfEy
3OzO24WsQP1GdTbQ1aIACydgwo7fiJOvL32/MEGPpUiWEB+izyHFv5dB9JV9g+dFkOItowX5s6Wf
1a2IhLSgnXPHElDO86mPWANPveVbzw67dNh8Whm2xiYnFJJBPz4mTNinVoQnY2H+fIOUDxIvZrmR
PqUFp7Dfzlwf/cZKyT0tFr80NarH3fW3473xQ9Azoh2GN6qdc1nNNIKA37RtQGzxtwTeEH9D7qv5
GTZUBDyDQXvwz1cg/fjrLT3UGuqxmkcHSC1xjT4III/6cV4bizXYy0a8L5sS6SZU9UeTcin2/U/L
wWcr/5kUYP4eaG65xmFvJpkE+26x0xBBTQnw5lNF9tVnWqlaTgYQhqjt6d6pdjVRHb51ywLeeX1I
rWaR22DwWOcL63W59Z9jzhccnvpS7/V5Hrv0rS3hlDMfOimjo4SAJWK6k0kBs7B29wBsWhb6Z8bR
o+vgiAMV3fbgMOoXuICQiWtMOaU3OGFpeuVaxORSmaXY31tln6RzOtBD/mkFrFvaxSnZkZ1ulOLX
SAWLYquk81ihDBpZTyFrJmBFeY/7koqGC3ndArAya/t6UX5V3gbFqQ0RBBuTfgmnab235a0OpuR0
MehcpjHQp3mGG6C8yZJMg2TOGh2PpSzJ0djC4nPkK+Jf9LQCC0ZUUkqwnl0K3k5Yd8vgc2m+exun
S8rTpEr7ANeZCYSx8CzTQFEy78paWlNLRiBYN0cpFSIpjlxT9Ub7mU2ib5jiBL72QtwAdfn6nY0S
5hoVYCurgONzs+lGqOBsmKhmipxIrztzAFCPwFABsGayLhWbvfDyaZ2qaiS+zOVHeCf3EJzUBXPu
Aq/GsqGWpn7/lT0INwTKw6y4eMbqQj/0fN5WbHCrFWJ+DvIZYpuWCjiViNiMCkZOSwGxKdRAuxTB
NKOJu71/aUAXkYlSMBAyg9R5xKqp5jNEov/FsVMpnmtllKLlZN+l5M4QraIvTLoWyacECRuzyuiY
TV0JneBix4CELGWeWrw1DZtfhGrDoqDU2WACp7HFh1QdZekDR3dOjKQxC0ICjxdFHdGo94Tm4jl3
kxua8eCKlYzq9KtzIPzXeP5VEGaFGJ6kMnUgajx3QjjFuXerCwj9mN0RYWfJCEJ5Ta3z4Cw0Z/zE
TO+TeHyux3wuGzva6w3jiTTGxlZihF+O/hntJBrMabHJfQkobBWfMStw01mch8nFPFkDVMJF1THW
GoM8lOhYK3SyVrs60E0HKf39A1mPX6i9nlYpNDJF7ik/SDywIE51SMBkpWdo+bVSXNTVQEgzSWiP
6GqqrS9rNYti/05IqkdHk3mk8IxmwuWVvF9osd5ix5aqAFT0mhaFAq4tSajD6kcTspjQ+s/fJ4IC
+XlGQ5QKKB9PQdQ8eARz8fGEjsnIqjwC7VDUyuNyi5ItIEDMTyOR5mM3HVA+qGZ16/iOouNENCBd
cPei+WWJYdWzHb6FkMYvFgz+hwwFE4UAo2Pu/4mhbpQQ4lDHrg/wdgIemjDh//Ys+AiCM0LFYSDk
xPQPIrenR2TYK3JBtEPUc75Q3d5Uy2X5z89ps5DXjv9STA0JdkVc3byrf6cEm8J4XLczttPb/hvc
YiFaB4EWIfjCiBgR7FVMEQ1kX4vqqNL8+E/z4yFGMdEC22qu7WLydKWj+E1IRfixVOAtq0OG8Nmu
bcuqaj7zc9RXwtK7w8JmoMCuF6H4sK8o0LKpgTsazJlpPY8M0yvZ1189JlVdSmJK4BVqRj/zYFvA
TLTyPkVdBO3uPKWdXnlve4Ai84vnxNudgAORdsIY8hTnNLhC5z+oQ7mnvV9+OH6lIH9V1U+Ha3+W
Exs3y5WJg8BX/XkUVVl+HgYJw/++7kQILYuosRpsrzXrHueEGuICqpfYl1UBJANvfPyNd+c7BUGY
6kowrvKLu61tPHFaKf0iEuChR2Db/LJgdYUU1OAl1bRNy/Zi1f6+Oc371DrWIsj45djhSLo0fNwb
klFWtaWLSSv6GgPhWH80BycqQ2ZHvQytW2uh6A97laFftXuKeIn90F7P4UD58BW+10li5AHngo6Q
x0Sv4k1w533gV/ztayp1xVNqFyMFs0z6H6dVF5ua252ie8ies0/PlNEGSgrxJU7y3/LAa2LUszos
4VcY7ebzOo20SmY0Uzh9RdPDVHNXe3lv1CIEJG/qy1ZFDZMAbFQgdibXG0qBxT6qbsMTCWGIZtAW
EumNQoHRy1Vg4qD5t759sV49TB+AEIuWaZrAS/+mjSrKI/7Y/Kc4H/TbrHSOfCKnqKvyaS8OlKNo
Y6khdm1qb53eB84llcF70NuxB2oVa2xaVKlHgAyV7AfQbYPCeR8shqHlEx7CX6TDBu7ecw/THxDh
tHesdVkEczTqffsujgAt4DJk3mend3ZPtTCRnxkCB0L8TWWgXex8R+TOlO8504lJmBaxLemvNvd4
TQ4GzEc2Z6DZauBu8lqqwpKdLijVS9Ogyop818R0eUNBZ2Dum1XtozN0O/iVNJ4qTwDJGnDXXhdu
6p5F3X+Sx316+CQ2TF3F3fuhlOq67mF9av8Qoqh6Ck2BXr7wODAckWoHEzok8qf0sh3u+ayFKPrK
0uRXaBVDLYnTEqhBhk7yek0+cEajXkCv1IPt9ne6Tfm9WKkGt4kIzFZ1Vzb0gLE5h0ZaauzNweld
WVb80soyNJYgaSSO2v9nMjXMBMboRyOJIU60BzUNyFo8G8Gpb+Bb9OsC/rH8IM/w1R0MXVCi8N3s
3jgSYUGpWx0G6dD2f14TFSzaGisEiGHQ7Se19Kt8xksL2i7kggY7ok1htuLDKFfSDsP9dPcLhqwB
xHg13pPUPhzLWb5RE5/O96Hb9E8Qm/6pNrQ2Mg1lqukHg5th3csefPD9Z7Nb+UF4eNSlHqeXSy0b
9OL3qYAUGKS1060U3Tvs7DaTES89ah8MjpCGU0iBYL5V17FDICQFelHGHJSIw9MBSBY/pwxGC2s1
WMAU7xss9yXaiuUiHMAwi3e/ys18W2/8gQftNzmsJ7FqkklVVtu+q3vF0ZcZLDY6xNNh0Pixjq2K
dFq8vx9TQ/pNCvGHpPmG7ZXCmoAR84A1ls2XO03kOzRkrxXimPAFWP3RmSE7pBbHKnlHLMBgL/xY
M1THtiMrqEpmum2sIPIjvbga2Xc5guxFyOugtdGuSfa/mZUW2039psn4/iI+2TkNrUPrBF/MXPbQ
klJNY0AmQ1vRdF028aknaPTLS5iKB9zTt5LMWrCq2bRBVhfVrG55sBqc/3WbBa0Fijnx6bxU04wq
YXGqtvJ7mb2bjCFi+n4OJPpiE2ksv92EYTuZ5i5fpIGF5id3g2aBpaPffjl+pcs8t1Di0aK/9EWu
ZXdMgjnxrDeT28/rmrhrDlBUhAscacMe+CibkzXwt8SbQuL5qpI5WWPfN1bllLCM1qvIoEdU8Akf
XPQOwvN7VbEhy8XX0wxBS2EdikhDFcS8JIigy/tBT6heRcleSGODgaHrM6ylbvc3KiyWSQuSlvvF
LHCTytIM+zFYkzY48k+LVqBo7TaZpnXmrhtlurWDr0cZrUOwIBtzs5JRWn9PaFxkaBIyHrk5AE8Y
VNAXWcL5vpjQpCaLMETAoAGaADI4SbmH7t41aiehD78SNjU6wr9VBfQk/3DK2uD0Y1YxiDBDMSkA
Dx9KbWBQGj9gXLVZPlA++IbtHnCgyUCO2nliZQ0yP0ctkP6/onsHIbo/eAtiwksJcqacpKunI5S4
8tZzWVvtdMzhuSGVfhbOcuq89P0kndr+y/OXy/j+2O5xK5LjNBbcYxXPZiWAhhuB6k6PaUVutgl8
DttvPwUgec6tf96KBlGgmfbD9Ybxs/IgVQf56SYgTJ/t0JSTNqC65+AZjaocW/ojnRGKVX1eriPi
S+5jm7AV52bDcFooHLuWygBl874NEsKZN1XDP0G4kbpzNHH6a8hTta1GQBB+kdDBuaSUh1FquKHx
LZVHDf1PJ8SMk319LVd0sR0GrGKO1BApxIL2NT48B68GL+d99ne2aTgBf5sbEE6gCGcKcwo/l6li
BnkT/0PdL2FZX3V9frwEVH0gcolHugBUpQXolqew9hpiq+SdJ5lNYm97CMuRkvYR//8Y5mrNhWlt
IDTFkSPe8lcgXYz/hC2eobfDEMnbi3WCN9KmbSR9YThYCSijBq+cTgg4/qPI/opw3E43/aLez2Dp
pGb+uVR5ROfjFZ+t/bCKk1iPhuhBXMkNC1uZaJQv5Jk8cdpwpdRgMnc3kLHpNje53h6i0I5ri3AJ
ZVR0Y7oUCpax7kmbWKGfp5hI1/37wUnctPTDujKFKinXK9biiAplRMYt6UdnI56FH4tPvBuxVzfx
Mg3lO0wdxPx57r2aq/5QJw0kEJecxT2QfRFXRz9MJhO3StjArJAIa5MJkly59xqRDAppAXWewzSq
uX+n+CUb4ZSQbgunQKbOas1zuk9m+kCHcgy/EnUb8QZYrQFNV7FT4iAT7mk0I/ojFd3ibSFsJyLU
1UQN9HaskmX1QirOoIEbkI+rz1bANTF/5gmeu89R0B+STXXRlwNucqZ+NR2pOW77yCnEaEExank4
C0fD3wQxdEOz8ORliOwP2WlpjMm2SqyCiNOcaKPj8xYXce1hPzwwBmxT8CZFozvcs72talaTVN0n
qjj/D4sGkj/MgwEUurwXL2hAChX9EselzZXpdT70OXFg5ImhaA6F55qA/3pQpZiPhZS3q+64WGBI
pbQze2QMxN6vgzOzDmNMTutzAd1xaLv/ZIRyYrxDWVMYQPyzT7b5YD5XrJEFPmAGfhxB7s/moJWu
4xY6Ks/sFpQgry91/6Hpg3JSx1gHQ2ZGESTh17yNO4Zdg/7PzYWb9lGbr7YT+LgwJ09p5G0CLphL
utLJwnO546toOVERFa1Kx+QMCHB2JGNLFjhDrTdaAd0nX0JxSOxFvb44NugQaVfm3qws05smmCUT
c7dBi7rSoRTFyk/CxOZuFxl3i74kFPuZQ9CaARLSe0dJ5Ym7+C3zAHnfuF8OkaUllw9g4HXFI09v
QzGc+D19kiwGTIL7oEj0VX336E0f87vNNM2Pm/yBOUTG8tiLbGf3jnDaSyh7EcwtRyZv9OVJzFlc
teJMRnySE+QZPNl5tJUcZNGHCRccq8NMPRwTclWzeXbzXiPUYoI0CGvhxQkkjCoYtB+qyK4Zwkic
2hhXO1lXqsGTTxb+Iy4M3jno1ZaMXgLn5sL66/oPD+c1FwmP7L6lIo5/T+cYH61gy/repRJb/Tyr
1KgmVM9gao2AtWmmRT0FgAvTZ43WtN0RPfRTJZgKG+mprv2j3I31lLNkZZuAEfCAWkFTorZpsy4F
gcyXPl9GawrZRvh/rZOy+AAJKpvOHU1pCK52IFPuF7PyWtOpsfH/3G/7cKyN0jXHt9n/ptXczp4W
sOrS2aFUN2c2NKa3F+RGl7ILKngLM51G/L4k1tJoHdsr3VkYllwrlaRfVbMqSGkuyoWXg5QIyooF
K9R2eOcVf91MVFv5aGVU9nXzzFByVRl91RAlSrcHtJ6db4g/Pvs7GPnWsUVgjJFqTsQl3/XJ/3I9
RCqQt8pwacJonZFZkUVbWHbLu1DfW9dwOxdGV9J9t+/BgSdEKZ2HbAlZCUDPaNFD52y/tIpr/89Y
vkmTBucZX0DPaHAKPrnDoD3XY+32M5htkonZ0kfC/o12EBjxjMJ+j7U5pWnYrN944tM34FNRrR8O
R2A0k47Z/5/6ckBVONw7X7F4iB9CPRDX6T5rdgLyIMpWcwIb5PIzgTlxeMTWUD1GD9x1LzZXcDdL
WdYJEJgcq2sopOHKHLBQhE7jacfHGtuIkKja8zs61GiDxrprtSKagywAzCbI/mvyWsWl0gjnWVdB
DxKHvJy2LwG8p9VCRnPfxpknz06Lo/Rhr78Rb8KIRHEtfaoP77OJO0thq0VImCQWnfHCZXMIO15x
iTL6NgZAuaRhFAKztQEl+6HTl9VdM73LrPzPHX9XFyQXu10BXcdca29Kwxiy0bF9RA6O5VV2D/mJ
NJI0JxtAcmqOn2vY7l1Wh8H9FhnHvbSViqvlmLzpOVHQTgkuNIVK47E8n7Iw0PFeddchplTezfF/
aAXF8oc99RfUW8yLzh2gkMSuwzTwrjHYT/pbVIm3iP5NGOYK+L3yB9eWVxsk2og6+0eCdlQnPbtU
346yGJmb9D+4KwdPXSGulFAwGg0Eq0p6+1y/dk0tmP8wllUprQFRuzTd3fLCUJDzrdciqO250v5t
BoTZOZ3hGdpbhrLd4xwS8n7SqJeWUHo5Lu/26GgmPdg6OElo1wU872nV3ndR8oHwaMJRlDVyvWC1
/hd/2+/OX22trltwdtBiZoC1CEnVT9DiWvN7rrygeUZUCtkjgHhn7i625/Jgj47Ku93SCH7dH72N
cauSGLChkntSXBH0AJyD/aM3dE8oC4aixnlM++o0QhtkIs4zj87jiEBDTSjPUPO8ohXLlqGGDo19
S9ysxToxHnEVRuYpvC/uIeVAOSX71EvyQC9pMax3gdXwKOQtoDXf3rvCX6BE6AHKE2HcekKhRw19
5LzjMK8yplSaNsKlcjUnL922UjRDfBiGqc8AicOFYPLgQoXqepOvSLa1irOR+eOd1pZKuv1R3xpq
WlGJyqc06vK8oaKPAsN5TFOE/0XtiqwRya6AtzayIDAE/1BgkRL/VWkVH9oOmQeRxVlxSmPijvfn
1RQb74QxU11ft+pEjn1YtHqvHDmHHsKIZY1piRNHQ2Pxv411jrMrurIqAvprvDP7vAwi9yGUEfBY
jiHMq4aZ60tl6CfrbOvjv3mDxrCOBI73cVVEo+5u6y9Ea7NhVwxQGKA/CjWYH90giyJjAiOsItU5
BsyTwX5xhb42EOOp8wpE521wA9GUD4+Zjz9cztahbJ3+6PHAxCpXqVC4WOSsnSFbK01zHFobHrBr
84IG0qgQx2KoqoqIutvTxJBo5R/PyVqwPQIJxPzoiLXVKI4t56P8XlVmsPo/5J+CpKtyoKok0Xu7
dxKK3iXejG4bWheqXkh0x4rUshfXBntmwc18KXbJY3g1Hh7/IA3gS+9rG5swzyuWdtd3RkWmk0CK
M3hIdH40OsIkckcoUGABtqTY2J+6AGbrp+SbGlfNkDtWQEjT4KUujjgap+zDPlpUTpzzpH8TOctC
5rOjQgZHYdAjfuVXqoNhnG89KtRCIg45sp+Lj5oCVl6/qjAGOnjs/uit5e0fcAgytv9EatZhlDdW
7/kZwyF2S3hbxiIn4DqWOMVI3pNMlgmy2C6++d0eAEgDUrtpGIxJ5a6+ijbV4JDUTRaIzxGPek3V
MAR44PJfONZfgjEDbv1q86BA/2Ze/oUkMMkCg9BEatNubP4i5XHvdI0XDZpBgo1tBqGKbLZGL8+f
n6iyImvupoUoPmrJGiiF5+5gCajONZcIU3A71o6mKTf0VYlIXIuxBZ6+SJWbe7RFk5GLJgRSy42+
m+S6qOsEQNp/9VOrLumqEjdb8023xDJ0B1brN3T5GudWMvV+mV1CsJ8EGb6xxhcvB43uViVRxrIQ
rxN8WWahOLxN5hlfDO09edghZhekYlQjQwJPZOlSnZLY1pPx0z/hnI7dI10NARpA1eiPk4FVe2SS
TGN5aVLds2OlA2leQJ4wvZ43EfI4hTDuMEo/Ws6Zer937wfl0E/UurUmMIWXH1bPzRLENGyzwPcS
+sRolQRZ7P8GyyogWxFXUf/m98oer8NcF8d7Tq4LuU6WlF7ofqfaeIilVwxgCr1gq75WDxc/mLBM
rKCS0PidZ0xzR79SAJZl9Oo7hw90wG6p0Ur2Gxin885NcFGyn/Zo3GhGsEAd0O2/7QyXIe+iq5ty
JyGNXQXto6F/jDuQ4Z6KbBP4PaqSG8LGud43ZuU9tSKLzyXDeb5S0DqXBKskzAx7Fo21jPc4XF9z
HOj9r4xTTQPyoUjO1kLn0BVOJ9cGoLgLY3wynEL1Xz4BJ2oTQivRwZNuIRYFN8BjaPfWb7fWAEMb
ovmEE3b4FvmQvMObEasYx5tImv+lWqxTlZwEHAfTylmDVtOhOgkMsCGYqkf6KptlphhwR4A5gEs/
87W3LS24sz8VEGhIjWIWcl4NuYyGzd9mpkn612MZffYx+UwUkGLsdkzB5ZgVvI1Mmkn3ngU6Q1P6
oTCK+SCcUuI9BZKjgatW4Gx5mg2DubdWxmg8MMh0Z4NiIUbbB0ZuSLKMHvbkCDK6IbYZ0b3diN0J
BU1IxU0fUr1HGjc7rOkbCLE/p3P/7znhE0of61qMkigM9V1AvlIOFC91Yf+f1E9G8qJjBCZ5/P36
Kf3mBOZvUcGxIkTfEhEYDBmM8vyHSieek2A4laYZL/Oiz2En/cAkvtL5/F5CRxsMWiN0mguO5OAZ
eixZVGl89SQdzLJlzNnychBXhKq5J10467lA6BREj6hWC0ddw0blDLu2DaUM9Str7h3VxvFRdegX
ZwgsGioTN8KZ3twLAE6IXusyhqLZJfIU5Sav6zmvFD0SXkeMhvXTQIkTMhVPoJ3ujkOl3vXy3Mtd
4jkkZHC+2ia6T2EBephYsI3SxwCi2nFlGg9eFY6fXk7fYy34/eK3fJtNa1wRDnlcjtG9DmauTADF
bZ3uNHmQwiYqcPq5OU/a3aAUfTlfGxMVmFz5/wglT6zeYFXcs4MdyyjSSbUUmYGV2ovOqBmFkQmB
We66VYm4x3RVRrl2cA8x5XbI60Kr+4etlqCoTNUbvIU8Pu5Eu2cpbGj+iHxK8waS4SOCWFBnCjD4
+W7BUjefu1Y5hZUUUwnO9b1/BTtj6XE29+pWsJJQDcEdBX121izB7Fnw7tp7VZlVNRm2ogxSgBTU
f1NGorRqA1RJI0DLMRXagp1w59N/fCf+cqCUeXtnBCz/HgZY8qUAuhJZyXG/LbAS57XyM1UOKRyl
fi9e4LhkBkJu4rpt32alD/tpxwAZMruacVA1O2uR2kIE92OtNB/0HV5meVPrsjmN+h+PeFTuGYmE
hkismABwAFdKfwS115eDz7E6NUmi1z1ogUUCs5Hhjkb7eFB1kb2/j3iTqzyr0x6ld8lW4MmMRuH7
HyLOgGodtH0xCCAT+iM/doPl0omxp93JP4RqEbNbaMnokQX0yGJNYA/tweCzOdHqGrJrFj1LEMl7
zTGmtCDaHGQg4t9gpuuHAnhPy1fLpvrI+mqlD2KnbeNswSkiY9o2Q1DQSQQh/WIPowayCHkPw9ik
P4OZn54vM6vxtiVhndMwpIiaqmW+holwKkclzdQ2P1HV9DcteKie8Vtd+TTxW+9sDBbiVKiO/8jS
EnK3zpr8v9SAE6Jr8BPGHbfGyF6SIyOzCd0lLhcEXxIFpMKBzGUBC99bE9QAr3O8YDzPGYQeDiwC
v5L40B35JQhVklBURyA2S7dm9haCSIhd0k7E9ChAtBseXZLelKpzAUDZ7JmyMA42hGzXWJkMR/FL
7Q7Oi38398coeQcto0C7BCwPwfCLV6/kqs+0ZcbLOKRuoI/5Z0ySHdV22erA8iFviJNxoaUqMPcJ
A7XaiheD+Ogo2hAVJNEw+9VOXx/2I6kWOwL8N9rX1WyUFoqCkuzFWUlLcx54i5trVi+X2ZJn69X2
SaVPVIvrc2q7NLa2PolVCPPfDQ6ZABiLEEdKdgReDhZeC1tiV2SjJ4L3F6+vM5uK7rSRGjFNjtLd
NogCmptweTdnmHgwW+o0xkzyjrn3BISu7w7ixNWQe9g6JOGxgbnNMtcU1/oLUXUNE3xFdIsZjoIc
JVzqKif8yqZhilgVfpB5D/Rm5EnPRXFT0TFghx9Yhtpl7BqwJsdVKPTMeutC0E1DuqwQY7lOStC7
acPbYBdhqhotWFWRfN5FXs1L56dE0ttLlzSypj3GSED09JYW/dRWXmV0hU/JXydhcvnIsix9p+Mw
9YGNMxvfyYOow305a3wEP6AFk5HMohBDgsy9mVU37uhqZxHn1kNWQgZsA1eBGRxhkd3LDz4kbNNo
hQTwlSjGYrQwIeCV1HrnV5pkSzpaFgspcb9bDQkkh8ozY7HdAHcUd1HYtKYCdgd7V4yZq60GyOhK
LTFAhb8F+3j6A4m77cUVdGHWi8OAvvk4rCTXi59zPGMyKgL9+RpZiXY5Vizmcmkqa2im+J5+s883
ZsIRZIFNYo+DTG7nPYHSJDchMr/aM0ni9tfnkYiNjxSNsvvuFeLQrJJUI5D90ak2sXTQuI6mBpKQ
/OGeM6HVDugemHb96BWwdZ+0E5/jNOp+5KklvNoiYZnyKr9q9G58ge7Vt8EFQrs/OkC+5c3uifBi
YrEOSyCA4gFxlQwQuNnZlU9gSsn1TQ6NQ6VSNWpG7A0pnJjUYOKW5/6NH8JUGT719lSCdDwGVJOF
pDpndRRvLNER/V/hExS+3G/ncbh605ffHm+hgilpTsdIuOiVkr7nncXkWrXAQxfCkgahZRnRkJMr
ZYsc9aTOzaWX+mUaC3DRIcrppXKxN1ARO9mBMzXHCUyZp6TIb2zAbUmBhGwAoTUb8VygJk0bOuJp
FWROltJVMyV9HsZ1WUN1K877fv+T6tI+QHLekSBOgbTaQws4XUtqDL8GKXVmQcjFlsxauphpnduh
w7epgFrjF1Po/ZFQO+O70pvd5tppKd7zUME9LCw5xb5IvcqNpQKSSJZ+TDhEY3xB3VsTrOkNtnr+
Qk5gmhtLW/S6o61bunhp1Zb93ytMXPS91kK/MQb5ZvJYUqWeDU1coMz/OAEcCzgEJXxDjBC2MzSq
VHNE/DGfA6NYcUbogwYEVUGc+RSfKJd+eWnTFQaJekDLmLDQJYT020CUHB1TBEw3QnlpxDsBbvIN
DyzPcJdcG/n4x7tpnrnWi/9UoBLCHx8veoe99vhz3vatLHnMUSHYxHi2BVhiFM/hj+8ATrranDdj
IWAlSswg9S7bG/pSjp2w5Fcc1bzTCXwxI5tVeVm/bjjpTl3Go3VVYiK5lSLhuEYVdhXNqbfK5oV7
/Z9h1h8J2Vmfie5RRsccFWzMbuy8VAiWOAMons0epjVjtZbWUoUB35PG44wL8pR8JEPxQDRNOrDk
Uq/qmHGM1Iz1LBMAzCFoW2cZAEli+f3yAhEzdxMFj96i1z+0S4am8MMljKf2jqb7dEIqUnf6+rOQ
kY50zQsPWeV3HdUDSeIPwpIzQdCj5FxzMDN9WnYApNHwSFFGYFDhd7tU7QXb6N+L7v9Xy9Fa3Ts5
IGnnZWaeY8w2nS8Hlxu5P3cNLHWk26eTwpZIoFPzfmxbeAalegHEbbTU98dG5IakY0iJE69u7B4A
yz4+AFSOwigDS5VvYWeynU5feD/uFpHw4XJ1tjr4js1/Zk385MH8/l5co0KTsg89bQUfnymNeO3i
Mu1hAyHccm5YHZufxJ/Njl6ClDLQygXklLjRV6kbrSWVAUAbiW6tMWfUi9zN1fdxcjq0nyqtmJL6
yixH83+7gTvIhc8AtvVFT0sdzQT4gYqvhDAI4/oEzRfjNRKJOSzxaE+qKx1aX+84HnY4ra/WtjXW
OsRVfB3xkIwSMZ7gx4OCLahw86+GY8+NjsrSeiTkky6+Bxl12c91ftg1GnHL7eidVWVgII4sEMYZ
Ow8Tf5d6UtUM6wekwvCpwAW+Gi9aLmwsYff0q+8KUhQMJq5DxSOuswbdtTyHfqQVbMrAULlITCgL
D8bcrBNiIcfDWJdQzyAqON7weLEB4JIfr/PRQA4tycDptOzty1uBorrsYmB6tIdod/RB9yTB1W3q
wWcfnDQRs2YJHznQo9YfFieu8ChMKSqcXN9Y5e+eC5BSXAi4w7ucrbZfB2HuhjqM9WOaKu4sOKZf
ABzThQMMqcagMtEht9eBfKHLf9odDeTN/oZEV8YS/Vqq7nO3+hke7wUIy9TC1mL2SA4EAklhn1Ds
iwHL6MDeN7EZ/c6bo6arsCRo3QBp8cCfbaKp4F8FcB5FxEGOjBChaiogKc0NDQ8b3u/RH3jbXptG
T0EPN96APHmR6NMzXSxVmB7AVQ9AFdVvkQXm1d55rcYE5fXSUYRSprO5N6FZAa0iWwigXM7fxFEN
ugExse+SF+wiEwExhTazupr6t0aNfsYlEYrFStqXrVE6BTGjD4d9aFcmeCQk/SBaLCkRJqpCjEZc
p5AfJgSCPlOW9We9etLLARiQpmlRlmWq/KKGRqL1pjNheh/+L0hlbnZcSpFLRbVJr1fStcPnzNLl
qoZ8Uz0o5fMqvD1Wmyr58Oj7U5gb3U8I6lKTiuCr7qx3wvny+ZvUrGa2keR+Dfei630tW+8844la
ylHCJFOBXUGOVQpDLmZVnBDo+SLtmw17Alkh+I++IATGB8m7DFKAyhst8coB1Fvp0bNVZcerszc2
TEXGrzIsKsJ1NfBsvqXjux23Ls3cEnViwdLL7sL81QpujDaDyqR8AE5119mntMhCC7Kx3GbhDMlV
3yBXHqPNLBkb486o+88OoM6q1RREHmXlwafZebcq9DS0W8AvJcMmCdE12H141kmO6hTR7VpCkRoZ
+BOnjl4b58P6g2j0eWI8vhXSl/rmp9e7+CmfmGPP1zmGpvPyGZds2dmzXgL4f3/HgqgfkV6n9fuv
nc5S0wvh3GzOs4r3Yew6Yt/Xoeys8gK3uOr+deYI7kgXRzO2BjYoOCfyq+59pIRwh4NMGi+topAu
0HXexW5XXEOwsXMhhBClMVkL3K97O7knZSL3KK8EInzQw4WHH34rtbNFNpkrSrTnLxjfd/cwIyaJ
ievX9ycjVKyZLAd0qrB869nRVjqUvoZKdLKUA487aBSIgI8Iwg+g/gkmYO7+cu3f1w3j9D7rITqG
Oc4Y1aZWnqmuAHnKLOkZG2qAvud9pJME0upIa9c7xBHWdFSXS4AMTObUo8lMIm8RNuDzCVywhZGb
mwtULjeobTfRnaLPjtPpfYVPFvXP+l4ehyhktStwZ2h62E1vVgxNP3ziJ7kkk1BoT+pptRWy3AJv
Kf9cjHfIxT9mST2fBRB+KBYssdb3y7G2UQdRmtawa9zGOWRlXalnwtS0jLDLdtFGHmATJlK4S5EK
AKkQQ9aByrpsmHWemytYhLMCKsO2VqiHvOXwWSlwlw+FBe2HdMiM+HzKO4YlsfCzEeSqffBXAqHo
sGG+Pttuopo0cgi0oOIBaBHg35IYi5j2eSmEokguMBntYyFnLmk1pUGwElmPuuy/hMWbxChmV6DD
gEXGPsLjb1tsFrzeq4gghckBjo0kxx6yjq48flOrfcgXpcuZ9XxR8v51DKbWkpXmJepLbMM7fmKF
dmV4UWt64u5/7MEV46zOHT4AKsEULoBgAebH9No53ETh+SJ1ozGf3Xv3TWfgV+8hsNrYhKAeLxGP
t/XkPSit83uoVFAKXSKhmGd19uZbfFhLX+SBgbpTlG4/Xe/5dqhgSvR96FQrqmku1l1sVTwdrJDV
BlqV0D2o7PCDGWVngRoGE8FzYFuLMV43prMv0EUk1WDXkR/BPdsMIAv/ov/JrIyj9BrhotTVAtNZ
6GgRMjhzk63jT0L88YY2XlVQhlpNRRU04Iux4+T6bF4t7mw4MAUUHnsb+HcOJnEeR5RI+XFwbVdr
LOQ4hPNYgRg53L3I2N/K82vnk5SB7WKl6LpxnsJkL63RSpXQudoQ8cPB8TgywbgJcl8yzQ8QsAOE
mtLLadolcXTWUhg/UinzzlLhhUec/FYHPonK5NGC927qq7p31HyeENrwZf6TCnMBD0FXenQ6uMZ0
TwKRyInusPfUNGZzvR1ADUSFv6OjfR7WOg81dkPpdxaHraJCm+CPGSm19/b/3lOeeV/pHEBn/qA7
3hMC/r1ZO+cwa1U8s1iAmNI/JKNSwnMPVFtaQbaoEc7PS3YpCk08Q6mADIXy7ka1hpFnIPFjrulN
k5OkzDt+ycrubeThCvhwQg0zJ5ktI3KLTUUHZYu3cWnZUu34idt+BTiAIjR/g2tcpuqce1DvoUiG
UV2BbFisTQp9KjTM/IiLnvbgQ4j4tCWif3oDuk2QkKX6oKtDzPraU4jXLNkrPbD0MWVcXTow2i9Y
lwr9xcx56VB8QNVrXGU/ULGtn+VfSDuLObYq2r9CtAf4n6AjzAIQV6It9I3IEYRPv1Z65uy6bjFT
ciztACOyhy4jMUm03RtPLh+j9GsB8NF+TTZzSdTh16M0BQ0iTts1ojH9QjD2fi3F7kUAakQTTvu/
gMVHUPFBvhqi27k7FSfGqTJdxXHF/LcrIttH7JvMi76dN+3roUi8+ryd5SBAwTZfZeh6ebQZaKk8
xt94eRKg/+AuqQ24Kwsk1ivV+aabULdyfQFKtqTi+dGSH3mXAdPmjOM3IT4BbGtyBQpewQZd3KKn
2djIPY/UAfp6dej+CjgdYWgFXnrmHfp1jlXPQuUvki6rMRLpL6AzNGfyxw==
`pragma protect end_protected
endmodule
