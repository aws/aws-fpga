`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2024.1"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2023_11", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
OCYOVRDiQ0PRLh53jjE5hOV9QIwYIMRuQmQz+AxH0I08pPxHoNv7VXKLphlUnKboY9gJ2aR4bdkU
U6NrXISEfZExzQmXi/HrXwJRYQ38b/xTFm9U3pJRVnm10Pb+2nRMZzGTrVGK2bHzKe5m7sEnd4Ck
cbNFyvLsLx41OH+shnVKrZdWvQvyLxE1lrFIKyyCO1IgGScFSuuCzsnddZsi1jNaRE4rVZFYdF7t
gPRhdJuTnX9xwQZ5Apw5dhZhpK1y+njO2VLCE/Rx/CFAM/anLyVc2VqGkQhUHFxxOiyMqHeIWuBq
WrC3Bq4QF2VhKY676y4/vzbNmbad3pH7Wee97A==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
E++ENnp/xsbGu5w0Dy0rDXAhiQOR6lFVKGv4RtcMtxPdFHL0G7wZKLLZbgAPKhCv4l45PPH8buWK
Pv88n0dgaFp11bT11yibvwol2MYv07cie4lSAUs6z7sTBMhOJ20delOT7H/OmsAQKGShrQpicAtW
SEn+4yVUC2Oo9a3vrWY=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
E3VI1XnOysIc6I7W4w28bby0F/2Blv676OCmQdvM5NlAZInWM+o3syjpPf9hQRd1tup2MMQLkdit
7Kg66wyroUDz4ZPbFjMbl1n0MCCZCcHKtjYXqd5+wTN/0ZqzC5hROZSkxAi1CJnN3K+0+oF68Odl
2epLkPmBzCbkLdVJ6J0=

`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
ppY+e42LXakuw1nzOzUPpTQTND9ShoEm6qKzHUGx/qGah81Gdqq8FZN7aF07KTmx7Jw4axRP6kTs
xRbz9Ku7kw==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3136)
`pragma protect data_block
8RsmBRSg70zL6vRlrQaBsayFTQY8Yrb7FiWtZQ7CnXrPA61VrQdyGcTkILpl3R8f2PRKCNXiVblP
RMMBo8wnwQThZ+/l1w5kJQB622dbezXn8QgwL9vkOkJi3Oy9L2uDEkt/2fGbIayBjflevaIIByu5
VpDcyhhsz7w7t5mRI1VDGv+5PuJ2EGTOFuKydXNQE0GgYDnBin4hDy2+iwvuKZMkAC3L/qIZeeXX
lRvvBm/ny+P9t+Np78j90r1kDuOnV9M6eA7y1+i6sxuYfPe1whgDxAHLGyGA1BtwmHTiUac5t+ej
Bo4tILfwZKYN65ZEgGhBOI/nIY1mXt046UIwhgkEA4r96Nv46K5N4SDMH4rDuU+xXyZt2O0OJzbk
8c1U8C1UxNWI7rtrNXHAn1/X2QAhIChCPNndQywaJ/qMOdXp9Cd+cqr/YF0m2hcX31b2NkLJ7ZyW
QG8MNoETZ6anv9qZtSJ8gErnbuF474/wuvRUQ+lB8lGMejoCFUoB0syCvrwVfuQfYfQ1hyKqdH44
SraMQTIBfJ5mBlCCC9LsvsxjF9Ael1SbgFoh9n/zA/3/69qC+AAyFI1AsXp6Ywm9rxTK5xT5j8wh
v/OIVQs7/H7jeY3oX4zEGehxN2cwkZN3Zlt70hqzVojZOK0lkQCDoYUEyaqblMvEE5o19ufLJF07
Z+COSHsnWwsVFPqgheQZTNR8Vcrmtv6j285qBFGqprQg9/ALZVYibEAUjM7Vo8sYKtRQfbqtEJuQ
x/XKle8xuJPNZcD2R3B6yd1vWHxWyC3SUvec4lO2kmG3Psb3nZPp2fhK/EdcDJRo4OI+Kc791Rmr
Hb1ULeb4BU2iqxIj4it8RB3i+yH6um9X5tfnIl7760Q916n6eN0bL6V5neW4xS0yNrHUTwLkmYCu
Ry2ozJL9rHdv9+laYVhs0gO0qeO1ohOLxX3Vtq9amOlhmP6EXfx7P58kiBjAk8ZU7nYWdhrmsEln
XLPXeY/b+rVD29wr1DvnjyI4KQcRYwWxEhuaT8n4LnhcVYqhpKTsoJIuTIGJzZVmF19mPCCEO63z
GvA97tsSu9tzeCb27EbE0fZ3BdiCAb4nkG+g9Qprx53cpualE26i0uDtgFgP8YOtTu3N8Sv17Wib
47nDaq1PNr64i3+RbBWTBrd1UNTRoQqKDi2ame4bhzB6Z2/5YIk4Lz3rV453UpG6gkGUZVU5jVEe
3u4sO3p3Tf5Fhi8vFc85Z8873old35/pjkyYutxCp/fyhbFuWf08nZ2pns4UnemFEmU/Jse13Rqe
mAxnc+CwW3fS9gQhJOC9pKlT8EJep+/s/+aHxzskCkPbTao9aUOwXxX9Df/aj8YdZdViHdOXKgq4
nIU1DWn2KJ/LaCu3JvA0Km/MF7noCMamHq2sgpxls87XFWx5lGPcrScUDX6EEs9SzXI1+aZdKR7N
jyURx6Y+moJEbG7ErGwJChPnHqnHS9eQDa2h3UG60E50HclACIhYfAc0GAwr9/6oHSyC5wueWoCY
43ctHT/BXrkyZRheHAVn52oDAyfIXlV7H3Qb2/h6pyIq3KNHbOEir5cKxFgLAHD/y9hG3mG3JbA9
rLXH5t/2CJODl1WpZl+XsXNCcuTkbc70FQvlNqT+kp/DjXnq68luYlKapfARlui6QtgAa3akdceB
25U8Pt6OFDFfMpENP/+u0VHTL2xEIaiXeXlC7ZyLuHamb4muaF1LEMl5xnKwIl2fkmVCP25fPUcz
7e3KlNd2zEfy4Kkyvqu+c5YAFRV3jdSWvgbokKGinKKfTgwZ5gCBvquLPBFMAmbI/jhdSFPslDdN
WBe1cOhu0xVa6tbHBKthMIIMSJ5A4OpPlWp+Z1vfNsrpagbhGXeYdGwT/pPAG8C+xFtZn4FoQebC
Wm8IxfBVwPK6JwiSTwbXaH8T0tW1AeTuu8sICnT9kKPMQQ1l8BwHHUG1Bq0GO6D1NCoWH7qeiCVL
yZNHSr8QPIT6AleJerQCQHSxiffoGIwefcCoq8ZyoW6o8XJsIS6ESB3Bv/xXgoM6/E2GJvkT+inL
1Ex7Vyi33fs8j9f4H/lr4uT2kTBWxzibzIk5rWlGhndyIqaT58CGYwPiicNZD771PZ0Y6DwiN0zJ
B44gl78x9kUX601yjbOQb3T0XaAwdbXiogGRxtA1wmzoL8GkLT6pWX2UBbJNG3fjTJXkE0lcaSKz
klIBe8sKOg5YxfMogTS0lQMh3+rCjAkiOdpoQxxIBj8U+bO6gebkdKiVbH9A4DUQLpufvDpbdnXM
AqU3DdKfE0m2ZgS4YnN7UusXbsVU7JF1hTxMKgXLePYAtR9HTRbr2vvERSb80LVONMtCy4D/9FzU
VvqJjRpSwBzdyiROjSfhubZZTXI5enA4NP6kDE88DTJnuovBvwAdzs1fPjJZc/RZAG4ba0s/iZgG
E2PHWiRKkOQVSSItOqacVGZ9TZ8e+xytnaVskUCWic1BZHHViKfc8OGF7rE3VuwDE2WlCudjUpxA
RpVgehwKt6a4a7YPxKY3rbEAbAewjMmIkrkN/xS0AF6PCibUnLRHzbNpRpXPPNmY26O7UT/8nzPV
8JmLyYolJdM3el8JHNARMhMUeNdU5ihTEkSbVS3S9aVLQgxk4YDuQU1Z2DD4hEjxrGQaTdNMoOQe
ZHJDnF+UzHDzbFyTVx36iI3c98OIjZq0LNWlFApL0R+ovfS3C8iXNSHImil9kaCAJpwdwd1UgVQ3
jTwQpX7WELxuzc7a3Fe2c9sk4aWV+rYsQqBRchg9bzCHmoE3NlqRs+hasSbYXadi6z+HXzUw4s4j
rO6GYGqNNAQjTUQL8BrfuaQLgX4I6SgGCN4Zene02Gfr9yrH4rDH+nUac+eDPtOeO6z4bsS/VFWj
2X/48RaXv/g7qP6N8h6qYapp5KdlDXCNNrYZxJzNzFQy8QFt5zWptp1TbrXP6/MhyhVKqsh6R7De
lqfPjm8io7DxE93N38WfO/YlQtL9CGiTss3VP66Ch/uEwSkKg9me7DsmqTTzEOiAzJNj0J6jU8oj
X7a1jUao2yRwF3D+wzjqpC/0smamoUg5K7sF0BVv0oWcqUxQ0DnkEIzKq1iP0Z1RR6Up1YaXm4P7
LqKkA8i5DsrMZ2cCzaEzSyNO9rnexqWLdAtSPGKE5suFSVS8ni+wTo+wMXMicmfzV6gAwUmjpip9
GfWBGNIoE63ZLXpg9YuclHogp8PtYy/HGYgPKCBgQxut6rXerWX3QZ64mK4DwerlRUeJxRG8UfY7
FE3z/gpJlcVucibEf2PhUA6YlD+FbDyj52ZPPj9tVgd5aLo/bKLFI2zNjC5eZ6cnOtzUiwS8eihY
IRHaA0C6yvd46wU0JWfYyfaPrCjlRp4Ln9GJV1eWuvI3WiAxAdtt1ev1PLjcsm6SIiLyLdTd0fxY
lBCmZOp5U2fpXmbc/6ZKkQjJD6wiq2d4zrVuFL6YGhgqnEMjWTUld3facgTotxnhlYPwm6PLkd4o
IHV+cvl22P5FiaTihk5U+5fcXmTlldpplJADh5yGS8hEbj4j8mqe+KXJNrzWlhELbDvKVpBMaftd
vCgyxRCMy9MejJqnsw/a/k2QXJdF4DvboR9XVmhNTEFcU7WNaaCQ4WSgjjSnRizOq2Fy3std5T/J
u1eym5sbmCLNbBeFcTZgNJkSD4Id+X+bHhugWgDdPQsCzso5LIm+353er3GTFaEs8eptJ3h3+Ce/
8xGGv4PSlRUqUeuT7c9B5lc/qzzO0YLCApqBwQ+B/xOkUeyWw+rEVe85qlH2TQePygl+C1qVtU/z
n/ASqMpcmHH64AP69VzMNf3b0SWh9GTRw+NVJspBHqvjga6JNF1rN7tj6n0Er+VCCova3r6NTYZX
H+sdxylLFi+j1shKeUsoWd0w+kKbTq6ENgbUeT5o5plAVONlzbfwntTxXznObpmvP1D7GD1CJ+pg
44dPmDMRCSH73TNBUbJPm6lQAzxVpEyJ3n/kpMIVDFer/BtH16n4qC9xBwI2elxvp2Q8e1Sa6YDy
wlKIK7B0g9PzlGZQxwntxhpEJxTNgjMv9h7IMdUpzA9kIVlUvs3kOx2mcOfxFF5AJytvPmB0QWx9
k/plcuaaHiIJSApNAZhPTLs3/4hUxrrumdkm0g1qnsyhl0V/Q3WQE79FiJ/xYZuOzIWZzZgbvhjU
FA==
`pragma protect end_protected
