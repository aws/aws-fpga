// =============================================================================
// Copyright 2016 Amazon.com, Inc. or its affiliates.
// All Rights Reserved Worldwide.
// Amazon Confidential information
// Restricted NDA Material
// =============================================================================

//--------------------------------------------------------------------------------
// Stats interface registers
//Register MAP
// 0x00 - GPIO 0 - read/write scratchpad
// 0x04 - GPIO 1 - read/write scratchpad
// 0x08 - DDR is ready status (bit 0)
// 0x0c - DDR reset (bit 0).  Set to drive reset to the DDR core.
// 0x10 - AXI Address - AXI Address for accessing DDR core (refer to Xilinx DDR specification - pg150)
// 0x14 - AXI Data - AXI Data access for accessing DDR core.  Read or write this register
//                   to read or write the Xilinx DDR controller registers.
// 0x20 - Write Words Low - Stats, number of words written (512-bit words).  Write to clear.  note is 64-bit counter
// 0x24 - Write Words High - Note can write either register to clear entire 64-bits
// 0x28 - Read Words Low - Stats, number of read words writen (512-bit words).  Write to clear
// 0x2c - Read Words High
//
// Interrupt Status0 - bit0: AXI-Lite interrupt from DDR core (refer to Xilinx DDR specification - pg150)


//--------------------------------------------------------------------------------

module sh_ddr #( parameter NUM_DDR = 3)
   (

   //---------------------------
   // Main clock/reset
   //---------------------------
   input clk,
   input rst_n,

   //--------------------------
   // DDR Physical Interface
   //--------------------------

// ------------------- DDR4 x72 RDIMM 2100 Interface A ----------------------------------
    input                CLK_300M_DIMM0_DP,
    input                CLK_300M_DIMM0_DN,
    output logic         M_A_ACT_N,
    output logic[16:0]   M_A_MA,
    output logic[1:0]    M_A_BA,
    output logic[1:0]    M_A_BG,
    output logic[0:0]    M_A_CKE,
    output logic[0:0]    M_A_ODT,
    output logic[0:0]    M_A_CS_N,
    output logic[0:0]    M_A_CLK_DN,
    output logic[0:0]    M_A_CLK_DP,
    output logic         RST_DIMM_A_N,
    output logic         M_A_PAR,
    inout  [63:0]        M_A_DQ,
    inout  [7:0]         M_A_ECC,
    inout  [17:0]        M_A_DQS_DP,
    inout  [17:0]        M_A_DQS_DN,

// ------------------- DDR4 x72 RDIMM 2100 Interface B ----------------------------------
    input                CLK_300M_DIMM1_DP,
    input                CLK_300M_DIMM1_DN,
    output logic         M_B_ACT_N,
    output logic[16:0]   M_B_MA,
    output logic[1:0]    M_B_BA,
    output logic[1:0]    M_B_BG,
    output logic[0:0]    M_B_CKE,
    output logic[0:0]    M_B_ODT,
    output logic[0:0]    M_B_CS_N,
    output logic[0:0]    M_B_CLK_DN,
    output logic[0:0]    M_B_CLK_DP,
    output logic         RST_DIMM_B_N,
    output logic         M_B_PAR,
    inout  [63:0]        M_B_DQ,
    inout  [7:0]         M_B_ECC,
    inout  [17:0]        M_B_DQS_DP,
    inout  [17:0]        M_B_DQS_DN,

// ------------------- DDR4 x72 RDIMM 2100 Interface C ----------------------------------
    input                CLK_300M_DIMM2_DP,
    input                CLK_300M_DIMM2_DN,
    output logic         M_C_ACT_N,
    output logic[16:0]   M_C_MA,
    output logic[1:0]    M_C_BA,
    output logic[1:0]    M_C_BG,
    output logic[0:0]    M_C_CKE,
    output logic[0:0]    M_C_ODT,
    output logic[0:0]    M_C_CS_N,
    output logic[0:0]    M_C_CLK_DN,
    output logic[0:0]    M_C_CLK_DP,
    output logic         RST_DIMM_C_N,
    output logic         M_C_PAR,
    inout  [63:0]        M_C_DQ,
    inout  [7:0]         M_C_ECC,
    inout  [17:0]        M_C_DQS_DP,
    inout  [17:0]        M_C_DQS_DN,

// ------------------- DDR4 x72 RDIMM 2100 Interface D ----------------------------------
    input                CLK_300M_DIMM3_DP,
    input                CLK_300M_DIMM3_DN,
    output logic         M_D_ACT_N,
    output logic[16:0]   M_D_MA,
    output logic[1:0]    M_D_BA,
    output logic[1:0]    M_D_BG,
    output logic[0:0]    M_D_CKE,
    output logic[0:0]    M_D_ODT,
    output logic[0:0]    M_D_CS_N,
    output logic[0:0]    M_D_CLK_DN,
    output logic[0:0]    M_D_CLK_DP,
    output logic         RST_DIMM_D_N,
    output logic         M_D_PAR,
    inout  [63:0]        M_D_DQ,
    inout  [7:0]         M_D_ECC,
    inout  [17:0]        M_D_DQS_DP,
    inout  [17:0]        M_D_DQS_DN,


   //------------------------------------------------------
   // DDR-4 Interface from CL (AXI-4)
   //------------------------------------------------------
   input[5:0] cl_sh_ddr_awid[NUM_DDR-1:0],
   input[63:0] cl_sh_ddr_awaddr[NUM_DDR-1:0],
   input[7:0] cl_sh_ddr_awlen[NUM_DDR-1:0],
   //input[10:0] cl_sh_ddr_awuser[NUM_DDR-1:0],
   input cl_sh_ddr_awvalid[NUM_DDR-1:0],
   output logic[NUM_DDR-1:0] sh_cl_ddr_awready,

   input[5:0] cl_sh_ddr_wid[NUM_DDR-1:0],
   input[511:0] cl_sh_ddr_wdata[NUM_DDR-1:0],
   input[63:0] cl_sh_ddr_wstrb[NUM_DDR-1:0],
   input[NUM_DDR-1:0] cl_sh_ddr_wlast,
   input[NUM_DDR-1:0] cl_sh_ddr_wvalid,
   output logic[NUM_DDR-1:0] sh_cl_ddr_wready,

   output logic[5:0] sh_cl_ddr_bid[NUM_DDR-1:0],
   output logic[1:0] sh_cl_ddr_bresp[NUM_DDR-1:0],
   output logic[NUM_DDR-1:0] sh_cl_ddr_bvalid,
   input[NUM_DDR-1:0] cl_sh_ddr_bready,

   input[5:0] cl_sh_ddr_arid[NUM_DDR-1:0],
   input[63:0] cl_sh_ddr_araddr[NUM_DDR-1:0],
   input[7:0] cl_sh_ddr_arlen[NUM_DDR-1:0],
   //input[10:0] cl_sh_ddr_aruser[NUM_DDR-1:0],
   input[NUM_DDR-1:0] cl_sh_ddr_arvalid,
   output logic[NUM_DDR-1:0] sh_cl_ddr_arready,

   output logic[5:0] sh_cl_ddr_rid[NUM_DDR-1:0],
   output logic[511:0] sh_cl_ddr_rdata[NUM_DDR-1:0],
   output logic[1:0] sh_cl_ddr_rresp[NUM_DDR-1:0],
   output logic[NUM_DDR-1:0] sh_cl_ddr_rlast,
   output logic[NUM_DDR-1:0] sh_cl_ddr_rvalid,
   input[NUM_DDR-1:0] cl_sh_ddr_rready,

   output logic[NUM_DDR-1:0] sh_cl_ddr_is_ready,

   input[7:0] sh_ddr_stat_addr[2:0],
   input[2:0] sh_ddr_stat_wr,
   input[2:0] sh_ddr_stat_rd,
   input[31:0] sh_ddr_stat_wdata[2:0],

   output logic[2:0] ddr_sh_stat_ack,
   output logic[31:0] ddr_sh_stat_rdata[2:0],
   output logic[7:0] ddr_sh_stat_int[2:0]
   );


`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
ACNU0P+gXXJrQHX6Amxx7lYUS2MmDZ1qYmPpOCHTv0sw6RphHiBCBEEKcttn4rITDBMpORGq4gbK
PSdcjlGQj/bpYp5DwaKw2qA6iSXNGahu8dE75l01vh8Wwrc0a1sIrNXjJ1pKrgaM0Qe+ByTmHIb+
vL3LxEaB2mbthnoouDooesdeWfCRF75+4dec13bFJTJE8aHptAduTQOxZXc308jc2L11Q92herLF
DY2LixriFXj9WZHtNoHAHYSdND0Z7P8Kpozdvy8tcLtpMxcufZwRsw95/bDPewblJEU+jQ7pTRFQ
1LgreSXuPtK0uTsBEm5csF0bQR7ZFpF8pc0ZCA==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
rLRjwE7cuboHu4Qqus1M69UVjTiCN1BBFZb1Qttx7/ojZf52x9LwkabUhNlg5cGckYXWOiM9eakz
O1c6tmfo3/mYjopYGBmufc6YVNNsTO1iNPBG4ffZcUZdghnS60M5lKQsFi8tnup0Cl98dx//W7Ox
FwXefa5DF7J3Pdlf41w=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
R9Jl7U2on9I1qh4ImD3MCBMDMQ/1pOEIA4ka/SWXbi/tGTQCv4/5515v2+oRWl/ulj/uCbbBRLDd
8dsNICxOZjfHWLn2gQE74+XcJCm6NTGUTOwTHyWn/mXAig4TOdCQabmIcEJnNYRBvKeuV+YavHgY
3QIJtsdbuPru68G3r6U=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 35024)
`pragma protect data_block
Scy0Jzl5gMw0z+0B8NgJiDHMwO0g6fFPdg+2dxEkYE+rsQj+f7c+xoh+HLESEA2Y+9nKbCqViJQV
RkSrI9hHN6OCa4jFmU1PRf+o2KCbfUcwys4HskquU/6ahQWwK/kcKnKncxcxXefkP5YLrt2C8Oyd
oSyO5VwO/ToMPiZJO2Q8EEsEhKY8dG0dJV7RVtxVycuusmvqOdpSo3naEnAGC6+b64qCVg/bdPCK
baMup9ShqtN9KGel4+3fX+orNqJQRZffkPFTLFMFkqw5WEgOkR7Y9fJXr72aVDMbgdV37CHbxbIH
IpZ1k60JFk4LrjYI/5AblJ+7JTbv9Lm2P6XI1+amoKZLvE6pU6sdNpv8tKDcbKaXo4JOCLUnzYHk
eckmGvHnY/+eVSmpIc7rV2dz9VFvjPClIHibQPx0VhjOgPGuo49z2stS4Ey2KwznyLjuseOQxn2w
BjVxkHckywPnP5QfTS6ptmYDcDnWI3MMF/06fTLLwzjnJx/3csf5ieKUoco7g/cJKY7had6kjTzT
Vf2CJPVeJvxGQemch3ufExn3JgeK97CeZPIH8ItmunSH2cxZtwDjEMzNVGi8ZLr1X43LXac8967f
GdW0VofYjlDAjf7j34dCjbu9vkXuCotgKuzYY+Dc/22n3pqhiN6dvT5V2kQWRYPHsl84bw93J/UQ
B6WVFeThn8szFiPqMJX2Ywhyx7qr3Wx+oQHKB4Qc323UefXslEOnteWW0YsOsUxQofPY0uRdM7UO
8Aa4/oX1zCwdYyUd/o6BGjXu+d6ljWu/km/5HPTFz2EvMFyEHGKtmhh/Uyc03pKIhx10WR9L1uot
kqEeugByrzauWvyLb/lHVw4GtpV5vKShlOgoAiKtIKy42pb+cDxZFtuCrp9iLlret6nHlGH9WhGl
/IJ3FAWKIBZf7+3OGbo7YxS7t/KHm4N3450IEHWlOjOFNiF10pzvitOvoU5Wy1yzsko13ZhMrNSB
Mo+/HYs63GB6zNohhti2j745nhp3AOfY3LbqJzJRii2CxzslIjacxhBXNeFTqit0YFFOCCISmPdY
5UnUtz1O4ryJr49Ya6Q4pjTPUuh/YpFt+GhfTGLHaf526hjQAtRNOuQSbZgeyQscluYBmS6veXjN
iwM9lAePK/eoINbBJaoeVbiLBdwUTEl6vdsYEVVGJb6q47wJi54w5xl/Jm7eF/ilqvxsAL0ogLC/
jNDwhFSdBzu8lkOo1AxY4AkUvmNF0iEz8jQ9LQuhpcBPGB8MPrOCOFANukrdMpuyUuX47++oP5ba
5iWJWhdjxfNAuEG1h9lVzxqRrwtDR37TEQDe/zROSgCicOFqenxYCrsqLtKeZBXd1q1DCIo4FL20
4FS1qTSLVSRBcxZ0DZekrBh6XGjJnTIEajijYl/D0qZ3G6ONC1RYiTh6AgQNBkC0Mv4vYAVlzNOC
JssLj+Un5hy5EABl+a2zXviLvzc08ema2Ulepp0iaXqYxSgmqJ2EgYkcZQRYtAD1b6I0DVk2v2yi
aap23CKWeCZJOht2y/6z1gtj4h6tV6KD2T41HM89yRhS1UdssnoZd8po/o2wc5RUH/lmxkfkj0f9
YQaCBCmKbHOUVDNmtcUrWURN/iWIdGNU9UE+DVVW3wID/hsvdwBYK/RHBn7HKr2O+Gx3Jb+++pyf
uE0dzdFfqY3Q/XmlJXx+jQyAKBm7F4dzZLqRpk1GfIXWUxNq5dAr/H+340V8BxlUPP74yilIC3GC
z8wRU5qaSI4/SHqUnpLU5RcNfhWxlZ6GTbi+SZ0Y6onMtO4WNLO8bbMK352nDQKrbglk9rdkdcbp
WSDBQB0TI44+fXg5kns+tuS+QhgLBLF7eUcA8uPs1NoTRD58G1Py+ieK2LzkhBC5bfzUUfGV9yvs
XVxB7zk3SJ3hCg2yHrs8iN0+CjPpxjwhu3kpQ9oXz35vSTRzF0pLkJKDpzbm79+F3gNRCLuk9Z4l
4l0FfjTqZATYEZmGepdhKsZOPuyPGwD84JgYuj5T3Z0JICiZeGS+xC7Beaikc0lEb74bXJtvKuIQ
KPzGwGUUnNQXIXQ0eaSo/D15tYafK6PciF+24QiHFoXDcX6ODYnWs7GTV0a1Sbj8iywr93SpiChr
GcmYWUxRKQ0S6SWguZk9kQWu0zSq41wEAhCA4l320mT+UMF2Gkl86aMK4u1etstT+2dRRppuEg5v
pdZnXpVKoSJs2/Jg/ghsgzEjUenKwLP7IwZCWtey3SaDlqVmS7c496pSDGhuyhyhT8SAdqBgWvtt
AV7KvHHLo8kaCTfaeQR4epocTVle52YZbXG6f54stmjKeX60WuLByoIixqIhyg4pTxHa/VKh1GUi
6YT5dhIdgTlmDEQBWsdHZf9p+ylpI7V/t3tj5vL6/lu7C8l8IR/S59CvZdmbAw/2l5X4hMdoC+e5
4p7GQB69ckXWZLsH1uNDVE1z+oV09kLI6rqW461TOt1tl3DYH7by7CX+/+eFQpeIzvgqhLVVw1So
B02g2xRPN4zcul0TOIeenpcwWVroRM4zvepQKIfFu38PGCXZxdc+2d9pifVFu39HG7lToLKPQnIZ
c50elKisHey5ihKMxQlkLJrCn/pR2U0jQtQohTBu8KebM+TAa0i7bUoYl1XBnMUS//kL7h5zn4Bq
ZLBdNGGxXgRgWPRjCvueHQiZrfahKzFeSuu+HmmZGSInSz9IbRKuIJCSsi/4hpxqzVb7hUA7tp1J
UoJgj6jniRAwI0170PayJk6Q3RaCPRvs02GOM3s9s7kGJJAABq9QpYUnWElgPtyBZ4Hrwm7C7CFX
ZiyEJJ6KVVLbLh7XmsKZL0DSx+p5lLd7nPZqaA2QOCN6tan+/UYN9w5/xJkLc/HcnHz+t/t2p/Mb
TtLgBp4Dea1G4w45x1FNMwszoKkjrQpiHfpRM6roMztAGBHouWgR+ajp0I+exFtnSdDNbK2whQ3O
9WrbwJGx73TSG0xTFACVPrT/Vt1XZtKYR+T6+6USnQs5xOjOjvwhxwVu6bOdsZlzXEEW2edP9hpD
DjEf8KPhT4YBiqJuSn3BQNOez3frw0U5CP1+shXGz5FyDWq9fplwTmHlRBEBHrZ59AjhXhEvDdnT
Inqugggr3xh6R7HLKhIxUe1ygoHmlaR43aTqMEZ493DyhR9aDlGJd75zIlFpEfgAr4ZQyjDoRMBP
jVLwGZuIzJYauhoYZ291afaHWo6V3Gx8UpiItnWaRWjmaTySM0j1IJuhw3/KzwxXbH7HzzLjXib3
qIUAFytfQcn+PZ7snA0B45zLNvsA1HlQzq46EFnsXTeORCb87BHZqkWmgXmd+0Xe+7jw122vFatz
JGEMgBgYnvU2iH3Y+KCnyE58sUBr00MTCijbSoH4ln/sMWfozde2oV69uNOdT0Y0HPyGjCbL0CwA
4Djp8gpag1z5m5EdT+eFex1L5mHr2ahNgqXQrhVAvB9yaEIXF2YzVyNDpUuL9pPFHlpM04v/IO2I
LqUEsfc8yqDCgFbLtb+aycJmzcYFR3mUJIOmJb6j26N57jPP6CqLbG2dj0y7z1lNMwL9j345tdKp
U2hqWXtCHb2gpREP6tLi4VMPx6rBvHxGoFDtvY3CTDWCM/7Djh1CrVn4QNqvxF2N01Pss0isn/wY
vQHZPi6rUHCt2UQbGXbk90N0FkR/5QsoUdxc8TI7fPTiTu4HZ6+PkmYTHn8kbZA4f4bq28rhyhLR
LWmWTvdzE7shs7usG/jeb5zZdci6Eqp7EjSuxH8e0KsnlFm1XqCfr8EyYVjAiHJG+Is+lg8XvlNr
yTT2cnC6eLXV/si3+SlxmtAxGLlJX+xUT8PZlICnAgrl+d7Ri8ZccNd1LUQRn72SCDTbE5Dsuz49
iBSmRJ3XXGVO8dWV77PST6pTJzSWRNqaOb1iydwcaT5t6MByPGHHJ2xI8MLytJhcamBC395OsbOA
Bo+BblclunC7tm05eqPGFg7kM4Zy7RE/wnle+yu8JbfKE/t8DXF1DD2qutxM12UZp0sRvGFfbO/K
ymbasz2u6ibDbO1wP/Co3/YbmF+rwLPWm1MHG+MIC4DsbtuNzxdCi1ea0gemYKlrZa/3/37qixnE
QmNfk3Dk8aMsmqQhNYt2XrR4SHL+8obkSeFZeUFlI3rH4tfX2VOrcN2wBaXNQr0Fx0qUF7aHUoOj
3ECY5N1PZSyI5r13zvjkykJK+CxNGFuv4NiFvBpRCYr6NuB1wxcUjxrQsGK2g2+Ppg5PPzAMLWv4
FyGPTxxDSU8ex5oUJ09VTmWSDmn8s6CTDHb/7y5bLo55VjFXMVPnAhp9nB447ww64Upa/e6i3VV2
nyAEcaihzU7J5lTMZI7u7RmfU9bClXTC1tjJfUx3QKzA4lPsWE9iygVT3OiUeDdEVWn7Bd89Z60v
TSXUe7pzZd3OF0kTW9F54RCQ5/Se+LggkE9F6hSsk376xfio5PRC2b/6UU5EqX4m70fptBrvjpu0
Z41eLcshJDFaTBOFCEdy2grVcgdZhOxUjKE/G20Glyj4pYqIE/zUVTXJRLztfCHW7mXiOtYYAFoJ
UBn/bcOVGzcViZ0SNuzxA8MJjQNDXlvefK2HCx2Gi44M0RP8N+IeTwEt0A0/FVz+ei7PRxSJX9R3
AZgdxK5i58IteDq7pCpfrpbAvZpP2n7AN0P24taAoAey/PC5cyrNheWgmB/a/7vegXK3ls1pPaeo
tjtH9ibBIxfKRPKDOsW3fwFNF+9Mx6dyqXdhTx2oCTbKS2V/LINEJarxSLAlvBsQFx1oNfBr0rWJ
wv+VKXNgCpWhluBkEa3rZ3I/6Ep6sDLbuINuRBnqim9PLbbjogbzddCM8Q979rNmFsNmn+UDR52x
Xi5HhpJkRQDhs6teYVsbBs7BZ1sNoKz1/BQi+OS23NRf3guqXkK+I898KMP7K0y8sFxcFqX+o76J
GDXP2QeCaBDQWM51EOVQEab5TNxUTOAzalDfTl54nKvN/rsYzwOOeTvN0a9fNykMg3Ge08fTiohC
ES4jsbGry544YmHKFF2vDYpUcKqYjHpHIWplqjgWJb4XcVh4Oa8P10GH0zOwX1V99ejrgLp+5G+P
Eievow9lRqT5zLh19yBzlwcp9GJzgBxpEQW0Mae4eGl26cBbA0MhmPmrkFmGT5dnSEM59Tu6RwOC
JdGt4qKnMnW4GmIp0hCI1twlEI44EQd1a3jp4p0nfeIyt24YmNwv/Oaz3ZROWh8BMMfbP5A6GFwc
xcijrdzEZ5JXprXsQIsYvZejZZMlPvMRtYNQ01hRMItoHXX42KvqseShYfqnabIki7VMSHPqtYSP
k36I27HAdc5wYgKu1yefwno96HbMzvoHHTBOjMxAye61D4Je0WuW24Xgz8Bs8X+Ybbr2BQ5bfexo
+XoqwTJXVAQi9QeYvG54NOMpxG5YYwoQoauuJYAr7r6pjKiiW345/shjCCZxjWBUgzzCSSz8EzIN
UtjDeltukacYOpkWl4/5UJEs4YoXM7cV6IqeS3iGvRcFEXBHoh6mIDfIUDzTWXLFSOuMJvYGyI5r
YtoMAR34HKKAoZuiAQUCVlGSBzbfeyyaZF6Q91YEKwWwd/PErAT+etOpyYIPSNda7Id4yjpJe3O4
J/32mb47t+zMXDjaVhFSL4l88cWLjTUo1sd+295veV1kN0nNEeja44imZbMRgrsjJHQLw/v8Na80
EfiUJ2u0o//asMaChhdGo/gkCS6kowoWU7clgGFDSz00fqsnmMkLiQG/91tvMq5sOIslGXnz2C6W
EA1lmXeUSyiwnF6su4kjMj68BQPBv9Rnx7ksbfT2mOWOltOTgVFoPbhDw1Gb8ixVVIQFctP1YBGo
OccHKp2qMC/3yBkeXLv16U6oyAXxIwtyFVFuV3BOScmyoyxsK1SdWO2sND0tc3+1wM/kBOT8CDgF
9pyNmOKwwRnDV+LN7CLrMRH8s0AuPXsnDwkrsRH56q2nAE46DS1I9MYh2dfX5SPDaNQvKkH683g2
q4eGLS2mdQCBy2s0V2/YduuSqP615QuVx2ImTmToOWB4dcxZR+kcMafMmIo8hj52En378YevQ25H
P5nq7BBZo1yMd04ydjOHo4/HiUbw4EQBnxvVZjY4Dyg6Pia/jVfu8VzWbL+BB08+TZofXn0VFSlj
b2LC5TEFMCP1okV0doXCsR2p6+3Yg+dEyu8T4RYWynDQWzBk35fHoQPU3aFiaapkcYjjHO+jAvnn
+02alhoNpw6i6EA+yZNS9bYGdwdNUSLRQnyrZ6oRR9luk+r5FnFiqmIFM5g/372iK4oOmEZh6Kxh
spcuaTF3e2bVMNBcSvlrp4FoN4GrBbgMUOKI5OiwyPCn/lDpmXw+H8bd03kUDIRLp6j8P0rWSPVH
qPhK3JiyRSo+ZjwedsSF+G+wKf9FLGfbUaqxcsksjyrvRiH2uKqavrNrizc4geuJ1zr6acMDPydc
YMA5Ul4PEAShWQAcYnyej+9adMTospEu8qtsznZc6gE8g3pFoNeW3jS/RC9dNMMyzS0ampluxPlk
IPJq3Ojf0/jjyiw61nnTvPPonQ7zcjhGu5nhXAkFr9OJoOuZ52lBU4LsGKNr9lZ+WHl+QBzs1SDI
S8qt/AKzDg/J5CIpjZecrYa50+Ms5ZrGA+mwf0zMYc0M+68GVLybHCNKKsyAOUOX9RNBzwhhkJbo
/1TWHROtrIuOzy37NHoSrjztjVbskdM8eLHeYM+dsC3d90GsF0MbBBVV4O0DEK47N3hYQ+nGgJIS
gvxhR7BSUPIWgOzKIAnZfcvCTrZVMnntfEdXjs8qaXhzKLV6kFlK9mqI5ceJU2e5WMLlM+PxrOX+
ma3EPdOYMKZ7YzA00WMf8zUmYP+QKXxI/FroifGfbFMjHADKNuCfhczfTeXM9kWHryQpqhcQaFqs
3x9QHyxJghrFbgCjxzB1zYq0Yc0xgc5DIzOERHyqHO8pSu9/EKIGuflPiblPXkpsDGXRF9dOfdBf
ZyzqU9+A8ye/gBQcGCV0H8e3fG6tZm+ZWDL33iKLFELwkMpRZxxrKCfk6+0x2tVESQz+uND0HVHc
BH/PyAH9Tgpf9h660M40gGYxsd/5fG0glfX/Vbd8VB5gPfn7qdZAOx8fUSQIrG8kLQ+yTUofU8nf
lTMlcgqu/ZaM3bX7VKPkh2ZQ4Salu/5h9PyDFVdfBNtd7UIDG/fsvBW08fXg8lZJs4T8a1CDUSII
G2ef/Xc6Q5ntCM9zU8/dfRR8FF4ICAcm0s9l0t54uZLQCFCnrcTW7oMrWZajO6iBBfrpRS9O769z
P25RdxICteKeOrIlyZoOBaBZ/OIWVBI+XR6zbTphsPwvn0S2nTXgMx0PJB+4sTmL1G9T0w7wRqsC
nomobLupDcVv3CeJdfHiBCmWWR+v1LrNLk8EAxP6VmTag5hjrX/m6BapE6klt9lsKrBFuwKb6xWD
dl2egxTYQFETX5wV4YHu02/FjbuM8LhoUVGxtUCJNNgIXsz/jod1vXhE03cSR1znTCb5YxvYgS+p
rke+/YOvK2/WYUJy5lnHY89YE+o8HNCBbsJriFp5CEZzm9C43kXwqCH3Lc+je8qFOUYEpOntHmWP
UMSUQvoEG/us3mNSNjmQC36NdsNdi+4RjEVWoN5DRuaveobfmjLuQN6xTrOxm9XRE4BpVYVkefSs
vQS5aNvY7I3c3KLsaqm9onhpp5lYmJ91yLLMz8KM3+214VsLLSL6e32ElHQNEmWac6R11ZDXHzmE
/KgvtOZDpjjW10b62UOKkk0+wNnW93/d8KXJw5RRP8SzeAy41m4SY+2EukuQgQbJ0t41VlP8QSBg
Fr2CfLxzEfyVyi3AfjO3WHTOeuSMY+Fc254my/D86aRWqENfKJ+o8JPoddgKuawhIgZlUkEaZQwn
lJqXo+sqvKwNKOmPj5gj0nw97biq5S3SPzX+h3Ma005zK1wOBbe6kvg91K2KM2crrdVs5BcHCvLA
iqEnb+G2MkLXY2ToI/8F8d+v7Hc2JkQPAX53UZD7XrK9ukxZp0SSJrsB4Dr/3SBWoBt8+FQH2es6
nOSZLdIvS1tPUMITvUBAXOToyFCfJ9xg6v4WibWazM3u02W6OLzHublvciDBJGje+kR+Fjh2qYHR
2KQPHirHd9EkpTYdJ8k0fNeedNG32z71l/Ua8StRqi6Sw2iYRKVtJsr3paKRIzfbjkhVk+R4FtR3
HhPP/fertNApQNF/yGq1xSTTDGDXWjcMYXF+6lCldva6WNH0jL9bjZjrASxcd5x2SeEHfFARSFRc
QQXcadVVBCuTz33zcom6YFyCNxfvUVQ6+XZf1LAYMxWpw6uDw54thZDiLtqfaoIjb7e6bo6L4qii
wJf4knKZINXbHin9s2Hd66ylMkIBiaRzQ0EHOvaanEbddB2ewcgbttKZQ4GnKECFYY309yway1wS
u7fM4hIeFxBhrtj7kiYJXvVDyk3l8N80Uyv2adX0vNgC/gE2t+K9AgPzgKi4LPrIoW34XeeNWX6P
xc8AVAwtbLQ+CS2DaUV22VeiNKJypOobNYKBiLfF+fSb0ACNsaG73+1CAmOyLQU3f8GRQsFCNx1Q
GdLGUY3+GnPQMzcV5YV4zleMu48WXWkdBW6sd3wBqE/p+SR6G35ZbGc3gPBfSWSVcHtEN/zi3YSv
hWukTq9X52vIE0Pn9Oeexzse/eEmoe25Ir9I+egTdBWDOdmEY2Fyotz2N85prwQDMUkjtLrhPALb
/JcAWdbl4vaw5KB4zS0ivGlT0Ikv4cn4yTcs1jc1sCK75Bi61BfEHqgy8tMi+nPvtW6WR5HP6ZoF
I6CRgnCsEnng9160HmOpzobyP8iZf71uw5Z1pSWDp4I4lEVK6/1ei1AbN744CFz0j0GZml5YG8Gd
PMznkRHb5fQHIde3FuI1ZWLVDPdT0cPVyET+GAEnoEOI+dCTBYnTIkOrD2JgKcBQ/lW/8xNYsfIJ
vAUQ5G6RMEVbyXlr2lt66yepTvhz+4ZyFV0FyL0wLOO6chJUpBXy+/WyUt22H3OQRzW5a5G7lHlL
WwlWAHAfoStthZS9G1Hl1VP1Y4e9faqaSZAMzBKHJwh1bGu7zbbn6UGjLXVA2L9yUHI5vHbVpFdR
9ft0XrVMXci7qSsJWBWJw0bZu9g4a7y1cUGigZYjp/ihDO/k21ugLs5iiquxseMPWUvrCHm3Ztr/
llaQ7NV8VuG3pufeSUOimljpJIOWdAPG0pGqnRazCMq9bht9PWEjLR6cB/4dAz1emvVNiS8jFBlf
M2QmItlxLatenmVmKnz3oyV76dhXesGOyNZ/eOGdP3hf1+7ofW7cf/nWexTdsKQIRtdi6kygcAzC
/Q3Utma2RrcPGP5RCm/EoHbMxOVmGaWm5jOCDP2LsQ8eave8c0LBlze5zs+gG9g6HXOtGMYDk7Pm
2PjISMaN16TNuUNUuv3f+BrHosMIsT9pVbV1fLvq4v/tst32m7fRI6IPy5x0URukdEb43+7nR1ch
xWC+CRvGzwGF7+twGR+SJ4PfaYDVuETKGzv1+UJFAqiB5uazZPjidC0faLIqaLAMwoucXfre4wo7
q3qu5XrHAnLFAcPOd1pCMZSHf1KmvbZL9Qt2nlfLcGUSRyEaRQWNMrLqBVSf99VApEhOUkPSmR6N
d/0U0Epwadb63pHAlihnku48PXo8Kv4wDu/uNw/h8T2tCB81Q8bU6JHrow9JIAD4OW4np6Eui0a4
dr91Toyk+K8ZJrMpDxr0aPvHobWwaTdTDbWm+pUF7/G1hgQyu9UeC/8vg6MlbRHnm3JIHNlHWmOv
Uup+98vqF5MtL9g0CHW3nFe/F4wUqKE8Jbi6IcV797CPCDdBPQL6By7yhSAxmE4RsjXJYOcH/UVe
V1res/iR7Quhr2rsogqgZbhW83l7VV63DZqFhOEnS5gWMz47USLL/kBKoRhfmyjT5UE+lpAgi0hT
yF6D/fLPNCZcxeNf36k7bvyRpair7oxJ7e9NaMkFXJh+RIHBy5Cxo0oPV0veB/oCD9/urK6LX6i2
fWw1a37kZdFagqVi3KO+aec70CYCaztGaE55FgWdiBheF1d6whRFHvHe8ANFqghayuJ1+Kl6KxxP
Ano9DY5zFGLVEMm2N0n/WmumDObsZc23aLQ3RgoMPguA1MCzz8LaRC7Hzi1Vl6eq7Uz7WGSZ+7+v
YDnNqUeK72vzfIt5/Yi7LSBJm/MddFHbbdixq9GBA+cNvIOLyKGMuv+E11/EzFB0geREoDS7sW4x
YmoqCG+9riACKjKJaJuTwlPuTW9JDaSDiXdte5pMthBSljcfJQ093ugKNG1bYlnjTTGhgjRy02a5
HC3mXbQMQEUxDay7QtLOEDEMO0fC6uYHLv21lSfI2Nyy4/r3e5C1nRPPn6ukaDfCZ0Jg7zLXPyQ1
ytCPzOuSAjKAXKAG7CU0tONQy5TUE/ShvUli076nufLHkE+0H6VcR85L9WjqzHCDIuSOKUWCEFXr
KScZIsbz6qbMco4rd6ML5p/z+qafHxiPGOUl4lA30kQsdYDQTVREwcIS8VDJ0cSwxCSB2dx4i14n
Aldoq3VlHMs1t2BHWzZ4r8BB/m9/BEIDPl0uBcjAtERqjFGZ4YS7A05kpPm3Huuu5NND5xNdSZhs
8ZUFeXrXl2OB//Or3YWBKKRxw75kP9XKcSD53NGVJDG6elFmCmvkCXtSwF32TOZirFafhl9uOYBj
5N1fktZ2rNmlvKi1T+8+DjgLkybReNO14gLm73NznOZpwZydqvXoYX3SNN8s7s11/+XwHmaLz3O/
yg5371YkyynzhkUAfNgKpcrZzHSnga73ek9BbmCsKNZkTpBXKzdxV1VyX0d0C3azh+Hlro3dgzTm
ypMZHyNFlqZjNWMQPSzZE/97CpXPcYocOLsYiU9W7HQZnmfCGyjo/NEe8QLHk6BiVXTjVzlZeaaV
HyXvf6N9+S8w2jgR0yxZlZWozxG5lpojGMNkn0IA2NW5DiX2U2+4II7vFvd58gSN9++mAQM+hYQE
u2987Rtf80q4NqlSXqbjZmfZLq3WfJWAaZlUnBa4ASIgyH9KQ+uhdp/av3NOL9Y1rM/NjACcKei/
b9uOwxGpEigsBpJdrdglQ/pSlM4Y5CWh+zub0pm5SLwvxaA4rTwUQdTB730vidoyILbKnyUupBz8
MzsvuaWCW/OHetdVAoM4XMXhBLvu5sijkNo84Ho8mRlh11luulQM/TrQq84omdeLkj+bFvjuO2jZ
Dols59aXhQW9fJSrBgDU8ZOGEQOdsA4rwAJo8p7PuS43ZYVnHyzvYPD9c/ThQwpS0MFoE4NNeKK2
ISd/3m0jtDajbDfhbAYo1mXo5gDD35NTBNB8lbGiIPfqVeSz6bSRu/ZtaSuqh2K1oKN67LISXD/S
aEB736LEPcLEdKPVrVYwmXcb1/ucfFBT4266AmFg5qRgaH/0Ljj3I3RENCkU2ud87dTo9UictUnP
+te37S+xmJHHs9sHNUzAQCJeo3wfWeeKJry1yNlRRwipza/+qbywMaXNiIMWEMW3xMuDX++oRTql
Fc+WcDb/qwWl22oLSojcKPmGkZTsNR4pomR+6f/DZYSbz/EEJjLtIXuROza4Kt/bF2VbYt/vagzY
0gMF/q9hfxpevZgGrRhEmfkjgFCjZdRBYTi7ZcrAerDMBlAevOk0hxX6Fo5QEjdII9h8qnSXZ01n
r/lmX0L80rQ07otiuTXkBcm+l/m2e+mB9ylPtMXrCgETbhR1Don+2RpRUN1GmAYEyBiGFpYEQfgr
kgVeKDjIgoYE4Y8hjBWBBkLYVSAnFrqwlOPL+oto2rkX6OA8oFOcsFefQuBDDDHXkGDynS529Am1
nXqmh+kh/ooLc6IjaqPCO/mzr/eqDtVabfr7mpOyGDHdiu66yeIFEQ5MBL/iEP+tuxgdSGhdADNH
xEPDFtmdq5B3ZH5FkisEHflPNQRiCZ5x88omUaCVVN6wDteJ/f+sbaBflTshNJ5vBsxh4VxNV787
QC6M0OOMC+1Y/2BeszwxZro7ZFyt+3S9ZEbM56uCFW9UHU+6VvRBTJeElrtLFsCZu31rWbm6TvUP
I6u2uY6tYZnDb7ACbo4uPlEZjYJlXR0xoeYWwUYVaTzZRd3UH0M/+aUTcNs7MrJPtNeqBuGJ29Tf
nxaciz6uxIRYQCia9fDnHLc5q4BPTriDwhVvam6e2BJ7gyS1lAAwNaOkNxv6OU8yKnEyMmPCWCAX
EK+g4Zx+y6N18WyGmXJJPMevyYlftDjhkNqhvrtIqqaPWyT2MsRVeJvzp7T0wDjVdfYvFeaucyDv
keNSPnCFSFdxDsEtlkzdC7qF2oQFE+bO+pL0pmIvSaFQoyYAnsgSm3/xhbevC3DIDbT0XSb3W/ex
PuOAvFB0cEXzer3PRBoO829uYTLbsOlruNWSbiB7X1WQIa7/SfQrGt0hOXIP1SFHm1RQEsFwXosp
zj8Ic9pYk6y4AIC9lJ27e2oJHIGqeY5HiRU6u6LzGrp5WKETYU8jBYDUFPrBGqOR6yP5UJK468IO
IkLIoSGzMD6f8ctgm36lTDix1bYb/+Iq1wYd33zMNo8Qh89s+r+KkW2QvVUfy4j1I+JB0D8/t9Yt
CJvJlDUSEzWu4c+1KX9EcpyQFVDZl1ZofIddHP1NYlDEI15go6JDQCimUU/jZy85VGDH1YzCpmuS
hAkXO27WjfowGmEhpeQ1V1+BpxG2Fzi3sHomukNbtBdHRhTvg+m7xjAxes+FrZFnRmDf22KVTqCM
sx1v8gouhys7NGzYMaZfXcfmyN8WpF89nWbt/TzFEFEfMq5pHwZ4msZtzDqMqCXnJyjYJ2/iGx35
YzM3ugIiYp2ashOMKMY8Lyr3Ye682KkQ3tp0DWZ0T397T5SC+L3CIPu0T0IDOJni7OKUvmf1v+3L
Z6+GgYfr4BWaj3xSQTo4wKqXG9PJ6YF4qKfEB92quzv4+Bc4XslTSEGtIwCKzyEDbcbGYWpdY5Qj
sh3r3N3tsuu6TTq8RM7KqLWhm/GbyTh76TTupRokWrQVxC662IBPvOscKjWM7W1u6ezhILaNvgeB
eZsWJUViTo7Ml6w60v7xNEoBHs5iRxPSoAgZx12fo0nhlyXAnJJrPecSB/lOCeDoAMyA1qUYwdKZ
KrWF3z3qpOSjywiaN22F4jb7FPETo49kgDd9RgjOijluV2FfdsK5Wo50MqfNDDjCqieuir0wE8lv
wbPSGosN31NzTioz+6WEyGLlpHfk3uA9PURPZ9JggrsEK7BbWVlyKSVoO7YF4cVrc4YNjeXitXT3
5xfmA/RIdFSI80t0feFwPbn4QE+shnv9fWeuhDREQosUXKS2VkyiERPiHmIDTbSQjh4+MwASEZyd
qgZKAB2R/bnM8MkPxFavr55Ss9bHb6qLNn19xMpU3CP6did5twNv33vjN20aqo2yR02nbBrpqIJu
cmD0fmMDZK+eM0TG/kFs2KHdgQSyi3RLOz8wQvdwoH70gbb6aeV94Tm/TCMZkJeAF7gMzzJ01eyp
ugPnJJjQj2tYitCk9d/y0HeMN0MAgmmCblNZb6TQ3q94bUQ64yCr1VHYESzdAxc4hpRluN+FifVK
nyz06inTHLozN862gsddjcV5NpgUzMGiEaadQNe6nl+dlZDVgTeeoTegHr+IFs99uOH5MyxZzye6
V+DDJRpUaDKiPcATqAakvSQxksBgcAOeP3oXeUaVW/58nKdS7ngrwEYWsXKLp/yfCSmVrFRCTGqX
OZzPP+Uz3Pyz97WKDYGlMPHNrQvA81wK6hyrXWBFzyYC4Cjz14fzWd94K8c/AkfAypp1eanROu1y
qoAkQO35nuo4GDDrfnYDpp1mlPXdXjUKT9INknde6tkkhgO9QtulQtWdiSzRDl7SNPQ5GQchZZzh
o4FeBu2/HYjxewp0p8/uKp9Tt5QRhwMOl3eajtRCGcAWn8NMKXhGPgwNLorwVWszbA3xq6EKeaSp
lL61Y4M8un/SUNJbAHZyBViG9d6Rmk/ccPw1dMDEZSS24Deix/12S/+nuyLwamFpLET9yTZU+ncb
ccfySsXCmuk6yb9pcLYD4Qwj8AhwdGtQiRCqyiqy8WBce5vEhZpmnh3A+oIXqy7k6Oag968H+PD2
0sGW7w5f5gRTWXayrpXA/+S4Wj/4vVS4MZJldzYYCuZERzLSbBRwqFWpWQwq3CP0Tf+kGwYhIuAU
LP8ue4A4JxV6xJg1QYQTXcZoRJupxmtjEls3Gq5lb0RX+B/IoHkaFedReM8+TLjDWTWN6xZugnZ/
6nXImvSL9uxt2TTHQ2TgAp5BKuJqC+XoqqPgVJSFYAfuPZDFkqGPte5+q/7MBI8umKZTuqNTxsr/
dMt5AKjJlBO2Z+zEUeL1Ya9RF6GcZaXc2ZUrcCAm8TR5DyPZLJQ/r7Hw/buO+zTxnoY+kLrBdS8U
r5a2SJQP9m3EIH3/X5wiqR6RH85FiEmWW3r3D6rIB9nwZAZnOXSbb5nHxM06VgIOAMnPgRX7O3sE
r76yQIGnMIBA+HXk+oZUQnzl03jIcYygnwPducnswCMOOSf2fCR8OeaSIZqjUTgoavKz9NGmfGen
3r9yTfBHzHgymPvUntjiPuwJ7oFFGrnTiGyXRHwYWzdfyuiD426DvcbBhWVSPcFVkO6GO52qhSR+
8z6YQTTCByd7nbgGhOnI8uByisyFtzsVD6AIdwrCRlMicf5n0DT7cD57eNDl9Y5Of/4Zw7HnKkK7
Tp9sR0xwcFZzfOBwKM/g0d/RpjvQdEDvau16SVVaLbqMrrHS9WEEvCxSV/bmPFWlkPsaJIV+ue5d
9AEekHnf399DUmv408MvWiFTf2ZER3f/gpPeUZhIyHKSNfwSVBYQWGpgsEtOWm4j3ZJ8SvFVvJL0
kYj1o/IlB2PMGg+omJ1tapYXAMDyASAbRgUOWpU+pR6/7AZG4kFwvarrocqOueoAEcjRjw1LMHiq
BebQ3iQkAxozHggCtWaWgx1j3gfJqDl9DbG4rkAQ3YvPRykROjUNsujHDqJtFtVBqrRJbZmzzzlN
ZWkpmx5aUpa7akc5P1m1Nl1F1ANmuJwTmYeQckyTfuwNOrS4VRt9hyhiThn8v5KuHL4IcMA01P9a
fG/bP3s2OTZ2fAuAqLbkeq+DUq1mKJD3XVykFtq6PZF6nqmXDTSNEF/8PPmNOaDr6wS/OO8+/q91
d+zd8QMKR7dsvd7sa19RhOhgOawmUUOB/EKglpeL8307DEQzkLHriipyGmfvKuz2JY0CD/11Bm4X
n0qRe77GQoiUI6C81KbCjYRQKSwFIWCAdIYmkKrGQ4z2k9JvC1i3ucwOqxKnUZUcgLTYw6bPAVma
0Xfbdot3er1TFuPx2yoxTeYIpbnXpHB3iB1PGaq8EnCkj3lUz2NIOVofsXGcf1cRIXukYF0Flyq9
VLwj2F5tqsIuhtXAh3PS7sFe0wrgJq7AKTKh2Z2b5GxU3UbGZEPan4qUIIJH+bku2x2KSE4LddM0
wIMa6lCFyehJNIJfeJpPK0/BnauJNGNys6N11i0lbxnsimIBa47H7scvxlo1E32MlBuvE8ekk/Mi
3wbMIZ27B2+RmjHpCEqI8r98RMxaUxVhyvhEXJY7T4fNyYOlgprDHWkq43pmMB/W1KW1FsZ62Fl8
S+EH4vB3wiMxbhjwuTDmd0dlKP+VN6Jopg66D8sX7qiUxCQ1voWNQkjj8pi7U7WwoqHUSUKJEoU+
D2VR90MnZhWvadztqbSruGVNEk2iTBT3vlR4KOAUVecauyw/jS4ceGVpQ7EHJ2g2CB6zRbTJedEQ
bzG8JGDkCX59pti5QJJ69rVUts90xu0isJeVGafO7ypZdNkLXnxp4gDy1NZmJR0k50IM1rrW+RSL
IKmx4cmUMF5fQNK3sJBip0ko7bYoRxOsu18Iy5kbqqJvwyqDNBcyz8lSFnzGAz8cFwCcGzHoKrEt
MKczy1FB+5Sh61PwArxMpqtNFqgfFohkRIlW39gEn/tTHPhjoJFjKBjtu+M/zaMPfu6Ha3aCpgGb
SrKdclQkoL0JtJAFqVkbS//+NyxYFbkGIq/w53TBo3AgW1PUOUfWuKLWggplaJRX4Qqz6Lbqf87N
xN08L1QmwdUPuNJnQ3o/hqLmlU35pkHxPpQePtseLsJ1LjiXqSoAqJNnsfbVXJGaXu3PHxb3zLNM
Q0S+2UjpupyhSJBEvQa/zObU3nCq5nHsXvaA3ZPdcxsxvg/xJH9+RCkN0jV03NxQrMFY1LaxYaNE
0BXZinQXuV9uh9KJKBHDAPWyPwutVerP8dxNUQuQtAfufS5bGEedTZJPqGaCp0w4Hth46RZRo1Xn
en/m9gQsXU2nMAFlolHAIk9WzjM4o10Vnj1t2mUDHkETWexMtVbNQICLruWMYgz5j4+0iZCG62eo
8QEQvvub6Dc349fnrg3s9JoY4KHRcZ+nO0q5Zw+az+1OhHCiIi23kpPM8vuiHhManEWh5dUicKY1
tQsjGI3I37hVLRtqC5WdUvKye5kzcsDnaMasLJuip92DYNGlrkcKa15+nt/tG8UMOKZW4TUlQSDO
vWFPJCausmm0Cejv2knZOK6JRncp8vgMgo3GKFrD7GHFHcbo9aezP5vh5oFNP9NdS6Yuv6mhhRBr
bts9+aympF9BMxTIvKmpei4vcaU8z400doYDJ4OXrLkhETSs59Ypu3TIOQ50ITWQ/aMuxsURlb7l
IKBt3Exjj65L6nHjzMO+dd7ocihT5XQofxjTOQhi9V33YKIZAqH7i2QOg593FXgv7t0tb6l/dw/g
vEXVV8RQgBvBp/4M4RYi4Wik6Y5G9nNAbov9jK1rBP1oS4ZFlIl7X3zw8fIqkavL4AiJ0q9cyuDF
A+JlOTXh35NlwzWfGP25CFt8Bfb7GpUKHd7bRkmQaSlN+soWujbcAcpy4eYNxBnFZOScvCplKSMa
f1VD7jG0UTHO5WG/9R6o+tcRnAu8tglxJC7m0gWh/3x6kFkYJgphdnZ+xYLmCDWkCh6zIZOugGSV
S/DoYWLvdE2oq+Kp19VDPNwUbgCCdSdUB6L+5Ym+cu8BqFrIUZN+MmhkMkEAis23TPvRLKgdWAyI
jkSUEpcOX+eM2o0uf2uoLb4Y8w/+Fq8YukecqUXqm8lpMvvD4CHeR9LbfnMz4uXADQXV8ZrqFkoj
2kyBqFYa9/qKnCYM4pZkYYG4NB5QR8IBAn2OIi2J1vCY2jmWEuYx4tegcOmb6bUa/duhEC1W4JXd
FKqQuwnuXehWplthOojDLNtBK47IQyGf9EpOHVkiPWm7dnbI0sKCRUB2WHIS+FLnC7QirmFdx0j3
Jicr0FV+YczUQqzKxyw8KutQ+zHFf6sINW0n//GVHgYov2MMYOHepATOv7Anzm2n+33C8za+jKvQ
hzyAQKQuXHU7R5y/uRhUTFNbQ+Ybce+/Qbe9JeRXFHeL7ZjPN+sVP6HwRGO7PaKn5CTzOucRsrSV
QdYBGOvYf1M7WO5OvkShOeb3CEhjmk+Pd90xouzXnLn8Cq7voUW/dYbAVPltDtu8BMBPQou2bMrs
M6cQbpIYXqmO8Q9UbQB65aWK96qdRJGj46bT50JD8w37CD6cw0c10b7Qe72ztWJdiXJ0KornSb47
hej7ejsq/bvWHD4ZvETNzybAVbRmqRk688rEDYRl2YspjxQFgKp7pKIWP3Hjpis4La2rxxFGecos
dfR+C8EguukWu/9rHR2xGP8nXFXhEwGC8hOeD5x1Nn7k6gt5BcivUHTYCTlBNawqwETO+DxUOHFl
2v93kJW8P8gY6fIqhJipvoOAt+QNh58SPF4ABj3GSPOOu3NjpPWYng+efdMKLNkssgdwVJeh7kgb
UhVS9SEQjMnzjz6y/3Fx35z72NqPm2y2ezQh8KEnArz9FiH5FPkJpyfieJRaToP+wbv9sfJ08BOm
twPxw2gLrgB4x00BPVHWpBfoIgOEUUUza+08OiGmRhluLZLQDaGtIs4GopJbeKE+AyQYCHK5SXsw
FASIMKVRoR1t+wPoP8tfkB1LcnWpNSEMJQ2OjIgXDjASaPOd1Zjzw72f7MhKQx6Ri3qUImyhUQrp
QZynvZfCpTVaCx7lCuWLBNej+A6GBmZfMm+/0UNp52zgFyF4xiWJCTEY5gdHpOhkJcdTCQl2NzBH
e82jBJCQCDOlqj/qiL3qlLiCzr6BRH+3zA4P8j7eFdAz5lt66KGNcqbvQ1qA0VbeE0EuHWMbjWba
dD1ht1Z5BCTZ1LDQ1J6HpzIZUOSPbzD0ey47uQ++wGz3lUQn77YlE0MsLvSlT2vhhkWI8ZbEa5Bp
3ILXtE7T2DnqQO+ET+Eva9wCDfhWSJGBkjxvEt38O/j67XaQVdWH827bI+Ei5YhfqseJzhgRNheg
70AmnKYWxKaCFKV/WPj7uYHlQsTEb5MoM5IachQIZc7jZgn0C412rLHfzvQtIDxyvNIdnIfAv4YV
5JjnAT9yd8kRJqaXcsF6viCYOOweRfWLiionU3nIL6NRX0YREbtB2E1jeVzauwYDqtfOBWwXUC48
qAguFwFmmwhZCcUWprnKgg5Y/NREHb98YQQU9XTQGnrYs6YekwWk+bMcsH3GUIsWlmaDKH9LGrbP
h/HgtZhOn9XnSsKFMv5lCfB5+0R/uMLct+5AQurIMeXyg1Z1REQEuhvfnTngC2EkBzYPecHBROll
kjcbxMRcxIA00O6wrH+lyANKaJPh3+hcleFcZDmusuAo3bFb5/1jsRjqbtmb4CPmhKed3JGHybJS
zpggm5d6HEmLjmar0OjVkJVbT88VX/lpxaKmK7CEZPaNHZSL/TFP4nDdiOIZrFX1VnbrPAO3HHwN
fJguT/sPizvyRWC+hO9jZwFsxvvtiQsU1JqP7Sm15fW04WBal1kkskXjEu+QPR24wN+ELxlPJQB8
1uobijqzUm22nMiH4Em+xh2Bn7SUtV3NrShhHTU/K90XVFwI2aGNlMq4SI9JED1L2PIlxWWUdHrF
CMsVhmJ2nfqux1TuF5rWeJax5FH5GghTZAfcmse87pfnZOO02WTPnSc4W3O/p5J+GnOOvctgtv1k
KKomwVvKAK2pAPN38Cv89PPbHSJ9NLPc8jNzbY5TmjFiK6wQXGS4/rIbF53Sn2qjOLXbS1ZZE9FP
yCm7CKo7RPBVQXxvuNivno7gXLtMLgOk5+bC3p9eJHy6/ayNwg8eeuwJ5dQBqil8bqChBIMeQ1sp
capgk57+kQbsnhgO38w+nYlkoHuCK46SefstQEUvs2PVYz+veqfNuwyX9csmsAgolLuIEJRaict9
8zHE0od2jxfa67O+ZKrijYjgZon9tKQe2tUvNKpFL1kC3LatER7vytTqsTOZMHLV5mgLmYzqefe6
pbcfyCc6DlMJ5ymg1CT2i/GqjnNs7LQVXYqwVQq7cY8YWr0GLhjgkyB6H6bcxQ2552EkhUIXv/h0
ht9xQIhYzfFV+1/38+rQPnf99/Bq0BLCYl8uUiUs5KC7mBmAVjdPiJMekwgV/S3X7e5eVxnDFoQV
Bv/5tv0oj6Ws6UiwsYDlB7nGl6tYPInfsg1JKNonIzVStbJc6428tZqq8U0exgI8ua3oLBUOasNa
hLrn7By8sZR6VV3elTPj1lPLReFG/6RCMHBqd5ra6R6eIFkz7l4IIhg3P5Np5ag4SJggQQjib6st
LimQ787IBfFg8/Uk7X7TZPEdgYPeSkRHQdU5wvAGpivqpYAAblHrTakHgKEVfeKPJIO5qOUUYAux
RVcnXfyOkm5g2j/jDTXPLPwTSgyMyHuTxSS59a0ymSVBAPnLgzU+yfIaZlaIQfor5PyuKHP/Jlm4
NykvxISxTDNjA6NbO2KnUM6Wtpgi2j7C9EfGvV5j8THJwLppeRQdCQGms/5s8KmwU3Gxv4I1xsZi
bVbVSllNZHmab+vMhocyQFTQDE7Nmn4/jmeO4aOEwJSXnz2nvQL3gqKuho8O2o82j+4romWyzQZR
ysl0us+JxTYZ7ISCBWaF9srS8EO+WpT74OCjqN3SgRlfEWJRcZhQODdfUzFGVbpBiMIi+b74rV+o
3hcXNJdKBaKr2tRwTpXhuPmysBOBkUK01chUhMzrwue0ySv884lCEk86+BXnPazrf3HJnzeaap5R
QdT1rCj0Wiwc6S2khyiTUmo1rk3GV710ttDlRNDCNXMbSGHcAqazaVl0MVOnOYDRzHZfO2oNLCkd
afcZnvPv/SRWEEop1aHWLRqAuTtwzdfu7M6keaDf+PSxM54WE7o8h70Xy+2v/msQ20X2dwqFIHit
1hfiRc7voCl8jYnPl4q1Y36KSrLVFGTbSdB1yeYr7jup8UWnXKyTYiLhgMi8ZNlKsdaGQdQETX50
7ucCRSYUcaK0GCQBo7Afulv5/GTK32Zoq0+nxvrZdPf5ksxj8dz3WhU213dYLeGp8KLD+0U3b7wU
PCwE1tBAcZjSQkNReO0RMPO4NeyVjLk1sxfzRGgoX65Quxks6D89lI53b8OPjesLJH/Mqrio1FsW
bMX6qp0NMjb53puE0ri05bt8cb7U0Ip8ZnbgoXBNjZKI7/e4fEiSCYiLUmiQrw6be0A2+ZiEfBiR
YPqMgzXRHGfZBui1nO5MVNLpUbAXh0MDe/P6jmfW3U+biWnAGi/o987RH/N71+rM+fSTt7/tKGUU
MTqR7Rt31LnvEyOWTDkaYocUrZ5+NXsaAVWvYUdJBEKmRnWgw5KUtccRqSw1bwAu9PfFvColT+5W
mI6AX4Gze2BSopbRQNVecoJ0fsZ5wW3QB1iRNb0RxQwYGYjeh68pnbJAfrWqpovjUqwPXmBjIlhy
9Fdt75SG576gWNcvkk9qhnaVWtFEWsyIZ5jHhs/Xk5UtvkimPV/PYHySCwTE5Z8ILuqCJH6IN6XA
aez1l8wajCn5q4CU9vJ17//UNALFR864RRhf6XhdUHYLaJoZiALBD54pArOcqEPoHpvGcO5DBNs+
zpZ5uKAi+1LJiGXUsJW58t7w6FGq1421YgMwB4r7z1gkGy0i/B8mbxMjuNiKHttxQnLz4do1s2U3
3JqzbjGGzx0liUZ2EXGE25BY3yNmC0KigwMVvNHvHm3CA+vBT7TKNoWailrUTPBSQo04pNl+Q4i5
rPMJ6q0SfS/qbsEwKuLQQ9f9GNh9yTfmI8ksvxpcHxJKHmyVC9IbzbBNjwIOX91GMa1EfpuQHEna
TT30t7f9umuK4S3Yn4LHPWmvrvX8gBmG74YAGjmUMdgV4Z78yXZNcAgyV+OoXUUN2pm2Ds8vOCNt
KsdbNEekdf27WYyVRrXbhFsECLkJ7cstzp8j37sI2SaCyPjN496LqdvLI8ohv6Vi+T2AI5z3mr1z
wH7o4gDnDYvarj9hNEic+3+zc/BHNnPRevmYVd8SFH0Ije37Mq8EsBheuso/e4x5WhLM0EmqHaal
v/etPfFMa3k5WXNRMwpaUBpP1fMvFrq/EKVsq1zgffXj/BhDbSTtLrXQzIrSfSx4pBkKs83s+8Mj
88vOVhIy+S2rwTziJJAxQN+9+7jh6tnQF7+jUZyUkaEOwc75szoCU5fSRa7svQpY8AobrmpjxY1a
R5iMWK7iG97vo8u1RQIoDHN+drvujkG9NZY2R35ltEbuxmnkNPGN61zg8CX9C57ANOXpGhBBAy6A
rIl62fVNuWRvUpxUCnCTZx5btWCJNMbfGqO6CmdC5IlHdV+DCeg5fyZNVI5kgCqg8pKTf76Ta9iy
F3eLu/5VeqwslMVp3rDY9N8TmrXD/zpLWlluN/Ytqu3SZaCxu3LIDGUHV7g/Sb+S4YrJEX/pJScc
38HBNr7eZr2uoTwLfst1pbLIM+CcTcuV17OXFZGqDnn/g39vLoQVxmpXLJCx+WksuilIQUFTWTTa
U5WniY3cWoyw3QxKQVTZMq5vLxV/DLQgFLZFbd6Moh67gIif4Xbxvoar4dXupcrteSXYnOne63/y
da9Czp0m3aKGt0QNl4gTIQZIGvLUdSVrWhvld0EpuylbeN/QEQSCYQ3Tp1TnY/AQZvsV74e1lmJq
uuSOGFRT1o6gV6jx7lxQfcEBrDgf2xmW2YsSSMXXnOvuRmvjKmP5GEqyr9DmMWKpht4hqTdLDkJu
9Ez56P0RZTjg7nMN7pLHLb/oDGNplUJwM8uyZxjeiRYFEeJDW2xks3HS1r165IoECZU7UAHlO/u3
NhopuXViHzamvDiLTtmT0pNe4FXiilVqJyZSAZsZ9aWWmk/VuCOMesEIp7J70Q64DugjKJ7/rNtg
SpIx/IWAPwp+0v4hxq96DF5tFpfnyf0WjGRTr47wr+UShUcVqzaEqptKvV8E3zTACxbdfciDl4jo
rB4G7al6Db96O6C7EY0YQXBGBwObA+GiHiQzbh0EMsALsv3d6GvwXrpO3fUK0k4hUuLXTnS5d6No
PdCTp3DX+fI4bA/EUNEkObkoiT0FNf9GmCHqv2yhAFzP2jWUBCpXCyvN+VOYwXrB0TmCucSEXC0p
YFSOgnxFDCmG4U5OTnCiZcqahjtkYaKk9RKQUiY+N5x35x0a7fFxY79IVjxEoyd0djjGbG07cM+v
rupnHuXjyZW3H5mlPbKLC/S4mQyNU8zHlrOgeVLKOThezfVsVPwEyNVf93dFCchQD8kqI1V/WrSM
jL2l+5RCzmVRP9f9oqjfVJH2nwXRlODCK/J2yTF/KZNcCgWUrYOCDcbUrzwHbOcWLAf/Vxa6kwEd
0R3dzxXm8IahX+5+MaHwoa7yORkephCu0ZUVVz6V39WtaLqfIGHlc6CcvsX4SkcVQV6XWB2H9mk/
e8pz3GWNuDpWBgDvu7xmOT+lTzURbQNhX0tdL4xjDWXkes7pTNAgGrMTePJk79ugftkHa9uAUgDl
c+F/0vmjoESsuTLo+/Vw8mMBuPJyClaa8Cjhxq/4b1Z/hoicCPbfgjE0Bnh4L4sCULChv86A6M1s
axwXsdKxQ5nr8hIla/MRf7vICwdiHlmKSqM3VhQbGKO2PQW+Omq2BVpjhq7B7WeDTcRye6JcyKHE
TwEFrsv8xoqqBn5zV/Hg2RXLMmSBbc4tSGn3e4tVhIo5DtX3AbGdFT2jSSEDFrqFG/PpAJisiuyH
1dBnyJAcx32peJ7ZlufKGK3DPQqV11gtEF1AYDZUqSZxEapb6nac+fmPUbT9g6L5iNB4D85mwiOO
E8xEKUm4nCQgW1NGpB8OmFyoG+7DzVLQGHYRQCLP0UTVUUFItH+qbJEbIoN6xwvwM87Uor/JgbB6
55RmPNimQeZxheTJvweEnUxJ28w1bVPTLJPvFoflohC4dRKxIEsblKK9Jpd1N95C1P/y7N0Bfak6
bEF8jgVUYRZWpyS6Cf726eovmP1B0NbVoHvVjRlM/kuZiSuFpT5WrPxrZ2fuUJ2L7KMF0tJ97XmN
+bM/DQKuYnZXTnQAuzMu/LZTn6HbEvDSjYiuqKE0kzKVN00AietU5PcA/Yt8oZOW8odasHKGnTQO
rDZMqP5EkWePxLNnadc2qZgiBm5UV8P69dXRle6A9cu+kyD7VpsgZs9oRJYbl3nAuTMxeCV4+jqW
XDLiuCpJoraDjzQzAgdTBJN9dgR7IuenWzHUsFt6vVFppOaijdEEIajUNteboXV9w9x0O2STH6AF
j/dUNlWsm4NpCc7U5HVjSi2k9vO2WCiX3nDxZVUTALoZ8A/j9aWdx07iWnH++xspTNMt0jPk4FqY
MF91jRDmgNaKPl/ps79f6oM7dUjOPJYfOzvrzNXAVJpZ/2UsqT8qf2PA+EBr7P4TbKL29pDS6nMJ
i4Hetav1cA4goGXZa3N0U1X9hrrtgUXzZVQMG1MNc5rQgxHVP9VzAnbtXVOztY6RHKe0wSXCE1Lh
fKcKPXkaif3uTFbpSxe/Fs1RKvFtcwplQhp6UbFjvp+XVbYZ8jQ2X68NZ6H1Ob/hJ0eIl4aADEin
su3IWRS9tutZ8axG4k8tP+w/L3zBRsePkeKPCNAQiR1sqj74PkDZUFmb6+lCURZQIyfmh6ZZCrQi
UkdpZ46N+k/3Qf8CD7VMUcwOnW27D9gpybKpkaushsb3DBdus2PJ1lgRnU4mukNI2Cx3ihGoUw+Q
LE5oSqf2nKxp1GmGEhLHjMQfoEunxcjf0BBI11OH5e6RHiY80s9cSj3ukrS8AqYr1H0qWU8bYXRu
4aeIDc67crpabUDPa44Z9gnEDaGNdNKl8LPJRshw7bVwm223IyBE6Tit/pjwUYX+wcvTlug4nuHj
bz6KvFhFrpBPW+/RYjNcSW2gFcu2tJsuYrapmMR1/5GLa8PyYV2Hd4evzzTAJT1BMeuQPMi66PNO
Iw2rbIIIMM/fztRTfCWPh49fdhpV1g6xHzRBBiwO7WGgwUpxCfIVWG3UQr9MhX93OI6rZ4EkMxia
qWxoqNL5VzQkFntP57+vBX2VpAMqdclRfmgZvpwxc/iQBtVACE5s32z/fnIUE8B5s2GZLIT73h4I
NsZNndqyULkTIOZgGKgMjBlS10I2ssdtSfapbuf/GE98nWsytNSmh/03pDVa7Z17f+lhfG6gqKy8
wt0ZjN9lFMinqGfZyHdwVWnFRpexMAvriowCQZCZvdKniS1C68ma9WOYVfSpO7WgbLH09DCit1ps
ypBA0ycfyu8GBW7DkSFUAjTbwoANxZT0bYOdEj67ulgqagATKkUO2pGIgsazymyqcS25EOxhz5f1
DaWvOTh2VnqFVm02bb8S1ES5HXke4vNSSuNrU/6HiodbcQkSI08UZDqddQYmGCrE7KA8ReTHUYuB
AQAl5QjplnmsRPiVElF1hCJ/0j9a4dNCVfR2/bzWdBopKBA9u22+Qt6lyWCNfAej0kaxFQXE5cRz
cKYdPOwBePlxT+ewtwjTLt7p4yw7bVceyWxeIx1B8aA/SjfT5rdNoTj51Hh5qe3d5K/yeeYoM5dk
qfInIh3dst+6AtJjszZGtWkr5t0QXdynn9F/wkhhqjtCX8H4Rqos1foEfHuQaClcGsU6VDa5cMNF
2vfDwgsb3gABgZZvUxzKb6oY+uyx4AH/4XMtQVzRRMy+lthUdgKrpLkMhzaisagLaEdGrHGknjpd
zxOXiocByygRFvcXrSkUzVzQx1bt8RObq0ch9Iao73vc8OR90PO87FCX7fmhs8MIKnF1bzlkYmU9
QdrbHPheHeFBlKSf+Kr+Z2F4gMWS7lelxPZAPduTsy/Jvze62CWTnEn/TF0rt9/ugBq33MNkvndb
7AV/j7Kl0X0W7VVRkkeUEypMLwT7ZE0ETM55yh4OvBxc8ABaZUvt22Qpp3Ewdn5p6/1Y6ZFOSiZo
BApRl9uLWoC+TvdP85qnLrC5X8XzrhgV96i3v5SGlVb5PLN59Snx2HLkVAa4yics27Qky04bnQj8
zJfVMiFWs0/OMxQufd1z2c7232rYzJFMAb/UtPdxxBagiwzyPfjNlJjTTkxNwh/O0RD16FyV4mWr
QKzyir5/KEYpQQsb0Gg/WmDSLCJw4ghN1XSM6M9vdh8DsaTzV/QNwbbE0JFmQXACwcbtrTD6cweI
7oYa/xbvK8ik91jLLkQt3YsOJ94cHcduQ1zoCgSVyqmy+nGG0s2xz0Omdv+V2bXgGU8IqZMwnfTv
qv7m4wvb+VVxivV45PZy+SBZDKb93Lk0gjDtnzoAWlOcvUwDxRT6wVjYpKhPdd9EtJhfEJ29lCan
lTGqHY9ujog8cIMeG4cT0twH2MSTwQLbbL4LAArlWeLia52Gr5t62wCOfMB/tDRAe6Eb5p1KYPXP
2Tkx9KXFpkhizNhHLUD2y606ULVgM6jnW0I4MxnEpW8YicaZm1FTGV8PHP9cN+wXCXMAWD10nIFc
YojGfUrRs4C7NIPLqsuLdkidps7sn2UZE/Vv3qr/g+NGlOxvN7Vtk2PjkRAz3yKL40a8XWRFF+13
4cY6jVRB8wf3MJ18jf6Vnvm3ePysjHYocdLpFPy/eOzgvYHxLT7xRgDjKXY1PR3HXWqjPnABXnqm
vZqJC35GYxprseyDdXL48b57Ea+ua0Dhk/40zBM+7JLkeej0zJ5rcT7f8YF8OoerURb/SfF90dQh
ZniRvB2aSkTNBzKKsE4P0J0lx0bTKwc4HzhYHLegnf1BtWyKnrhOpTuy4QmkLlmX0yYBxhkmRq+S
VGh9PUPjq3fAOv9jHl8YZwGhfWqy6hxcHXSlQGyaqEX54nij7ukmBCxY+edZIYqv0XgIE24i4yOF
oO0/B87wqXNfa9aTMR2bISw+joLVkARgkU14e3ty4aTbsLka8vVUiFqJA9DT9ClfxkdgWzSrz3AP
EG5uHkCkQU0H0KREK35wtcyMKpzqgBBkJ52NIcwug2DxujW9ycZtkPHICOjvnwf236eyqzuvbmgS
ncOTVFOjbQl8nuXBKNGolgaUk684kltidpEHZ9ki3sNBluNNqB4zU/s8z71BoeRxSLeWC45RSQ7L
oPMKDkhjBzyWe9e8FcXKyCA7QbuZ8msAR5t/Oa53xtCyMJiEXIkLDkDFZCf7O6xUFSNTKJbt5Lo/
O0VNOYX0j8DPEEu83QPzgZA2vcpAJ9UmbeCzc2uVVvY1fmxcvM7NsgN0jJ740fEc0OjPZhmymOY+
4ZLOmmN5eWfQC9JYhXh9qxLG92V5hO+ZKm2Fr+Py3dTVv/t81oEn3UF7zhJTzOwhTFtpXuWjiRRy
2asHRqjSk4Tp5CApA8sJpkZqZZo/M15LCoq6FdgJOJY9UImEJWx5QPiFdaH9Ob56iH2u4FV28yNB
R2uy64690xgQ1XQ2aLhtX3pJUFA2ZZngZ1D5Pao83N/STJHP1tTbYsXBdpKB9fKHySgOMrIBNdCB
RvGe2zh3SNskQ9tDwEoV5OwpNpHEo9XQ+x5zTcu+vak6Os/f8mOP6zO33ugyMjAspVWorBfpy38+
nLF5T9m701LCKvB0Z0IdAunUGyugfxfUjT+tgaybG5jOUKn6cJltLLhJOeTFiptO/neijCj+YLI9
s3jBmEo3bnejenu/z4ZKRt34K3pl7aeOOzOfXDhO3jCTcpKyCCJo4Ty3z+V/UYI0uBVgUUS455Po
1d1KcrrvXBUPAfXtBIvA68Hgdz4vC4ucRcP5vbqYTLqfTMBxytSzHip4+N2oge01Nxtzqf7kchsq
YM1ztW2+HOHIAaeddmtlvaqrvYD5UAD3AdOYGhz9eQeVVxKxbv8D6C+KwT8yWC3RMi4A1v2AsOui
VqXScQXq5AcAp4qBTwQM/HVwO5fwglqee02Eicahu5HZ1yPP6VTtF/DqtgojEHufAHwn3TKV37/1
CsE1pC93ViOPrCLg7w24/RfLNfDylyMTXWxcsvgGN1pxfe5eqiTfhZ5Hrs3osrmvoMgEg6IrEch5
N0fFI9Xv5GD/6Py8QhkUU/0sKNXrP4QJEvun1zlDBTi4q919UQq3MaXGia86j2mwB/QA26fZrzly
ZSGedkgNqXnSEw3eozVRbZe/xWMc5ty4m+9ziVFyxcZwmu9nUnS/SH3kdHJr3SzUC6cj4nOcQLvI
H/AIdpGANY+HY8QEG7RUrRyiafoYIB6yu6FuH8WnnHqBB/QPlEbxHOJOwjExmytAIDRJHP7p8sv/
tmXwGwzIHVGltEQ3wwIGFNAH57O0ehfUwuxfd4NaoKVTtDLtc/fuIZLPjmezs+vR5ST8DE24lo3r
aFRDwxqbYSXZtMCGkg9owyj/+4aLIbYBt2s10OlwssBM5DM0SQlnmDhdJEgxira+8qreYnQH/YPS
MRYKeLwiYnEzWCNhDmkjyjOjc8tHVrGF8Bbk1307gfphwa4KMxyIDWIHv/zVBOF8Sz5rutQ9TeBU
eYWeAS/u/EcVHINW4qFDDx1KLEZSL4iJ5PQgjBI+XGKUDMJcgfd5ONhtl3CiOrBi3dN61rQulAhM
RSYirARxdt8XsxYAUXzSRES5oQmyXBG1t4q7cylWonItGZCQbk1mT5FH8eBthVI/OZrkBCyWKlmY
fwlOpCmw9U9P1daNWT6EWmuRQhNnGBciYI9JRNydkknXwuDU2zIBel6469HxirYGzszbWGaxnDs7
LFXoi7+5eT1bmMlv7QRw/gbc5uogDctac9kww2L3vcaQ9KcansHL/04mNMvjRBTwiaT3NtoDKr4z
5mL5zPsA+FkMhnjQnu2AsRhibHqu1OOTLLQnuok1+EYocdHoa6PrlSVNDmOhziqriW/1ALYm5lAD
Kn1GbMkHQJDaUVABoGuso+KQvshGebEOMq/getQlpoMT8yFF+4+xtFRnMdhB5mVgdUTCw55RDSfx
75Dk8UHaRPuVVz3Fi2pg8TBYPBF58P6K+r4mRIHml/Bu5ZZNRtyRP3jRj0ebbp9+SK200DwfHEA1
uNcaS202hR9y50+z0dPVIv+Wi4TLTY7BJ+FncskjfPc/asID7aYlR+N/j6Obs+fNFxmQqgpPwPbH
glaQrHWlX2refC5+dkOKfIfIGyVj+vQbrY5qb5HRc/h5pO5bMr6qvBFVaeT7Gc+5txCAL0sRU9Gw
lAtSVahDYz/e2VjAYLirDpoYUFkD60lxrq3uwVxq1KejLdmVukYVn4suWwgPAlaZnq0JPGidmrF1
t5PTVFHdz3ON7aZglDIcnTSWzVlfPsOpe6TV00l5YovNbDEsvjrtz4gFPZvXTaW5kRay/rI37TeI
R2MT9kkILr0J3EwPXelpBO0yS6BbBTjEItuKHhofSl7FampSw80A6k4C/OGLW1emYjw4nIcXXBt7
OtZwtMfh+FwZM3+ovcD2n9b2zInwax6xFnng7WiMsMEiBX789NSBWNxfObexAzOSc+tc7VvUXu2i
i5eUMuQURutEp/TzcDObRFoYZEKri6Wex05/TzCPE8xgy0xCZysCsasyDadDTC7zR8OQ4a5AjWkZ
UmhmTP9sw5NqIygaWOmTkv4VOVnlpd0HrUFW8KC28NO1hNT2ma2STXMiLpLVgMMw5y+p8tpbtca/
32w+07QtYFJShSNX6I8YQDQVlIPApDrjdjd+StH6nzSOQfD4zNyCjB840C4v5qF1pwRD+ugcTOni
GBVnYLXbXZnYmpEM2aaTuVFBdDKcVyPHAneoTsEutsDEZuc681nRMeP3KWFI3fKfinsQMSuG+fyr
zQrXzxsZdzcGIpusFaKxTpfnXFFv+tHsA+pfcdpKTwfikVT4kfhjcxPxC+Eq4W6nnp4f+MsBJR0g
EGi6hh1H0h4MEBwJ8/P2O7r/7aQyP69bWMOPbtjDyzimKzyzkhh435ExVvxwUm8/Z3a6oqjLBII8
E+f25Zo8wNdRgevrau8S62/0zn7q1ZP/DVH2Pg0h1kGHa9ZNIX8mF6bmoDNnE/BUmKGmXBNdJBrF
lHngq1GiwjOhNrlqPQoMub4yifYML0IaaAHFWoPGd3BK/5YQ9hldV+X3cjbbJZQSIpfHK3EHSng3
AFA1ihjP9nQ3LV5sRio4rOp44QoIqSjzMKcqNbPa+69sVu58zmxW4IbK/uJy0t8UUyFB72womMNn
jhOqxKwcVbyjUAdQBv0BZE0kxkBHJE2t+UNHRiSfdthaHAogPVWDKnLYGnaM39auzU79K91XaUyS
Mlv0nXO4Hl1+KEUG9/gFZ1+8c6nu07ysQU0743KgMf3yK9PhZT1kk8VbcG1gxx2xPvpqtUMEzqMz
acW9i6StbQN+OasDiiDbzp6d/HFYwxYWG2GOkHOOI5PpWQ4c2xT1AqA5+/dt5NN2aYqooxNrvh5x
50PH8UcPZk7deW7SQk4aRYOr7GJkZt8BFgbl3IR8v78MjFv+WfS1S6i2R85+RvzRz5qPpZD1b/qF
UgJYtHVFyZzxwkP6HIcte84ALGZ9yxMuANRAkU6bJFye0UfC8tjFSmoUXbnXihDnkp3HENnRnefK
bVEC5/PNDKtJtijpOOxbwS4GyKa92xqLQQrzxCChFF+C3+mqLmg5g+6DpgCjLsxBfxG+Qtmc5z7v
WnlRrzZj/Mx8UF5b+/FoxuTuyxexCPPmo2EBHNj2uYUvnZOzFo6zYuYyGvrluAsf1RMR8+0JrsVh
qVYIReJ6K93SJns1xbWydVfi1rzVavvW2AH7spCzV+8IrmzHt6ru0m8PXdZeym/g4VJ+X/S1b0Ta
UbBjOUsexXl4i0qgr3PacTPhc3/d/BZ+n3IrNNJ/q+27NyKzSlhfLrIDLi02ImvznsFc99uam1k6
U7uIdQhbHQ1CTU9sIHyCc8e7UGB3hv2b9AzFJy6j7sQWMmcFmPgImqj//OnlU4TjSJy1q4mRbIIK
y4pY9+TS9vvjD/YJsdjhgnwqV0+NCFuXF9DloPWKF4y8WBBZwe2+yWX0ONp7Qz986VRlwI952bmn
T6/KyjIkd8Mj3zsfLken4Ry+YuaCVRJYqUxRU3Rcu6eBI1EylRW0EXdPM1busw/N/4MP132Aluhu
q6SpTtAvq2Wci+Kb0pdySfwvE9Pox5gW3Hxg8rJenF6Ul5cdhcPXk8hKKrf01THgFvdZBvEY/G/z
r9GcjUmTVmZ1mhXE3yA+Cw4cTsZeRePnWw4mOfcXFp7QhbekvTnemrfTm1bkVezWb1QAGl7K6nQr
OAs2NFdDiLGo2ganql88vOz1QABgEiMYol1QZGvsIhi5GywBbYuygNyqOlRH0zzDX9QpVh6Qn9dz
0mShN16WqGPgdtQf7SL74O2v2fIVjCTIMXe/CTGhkxQbIAzC913jVE/oKizI3Xfs/2AHLq8yxn+k
yVlnng7rBkXdjCkE0GGsax5077kIR02pfazDZUirRBk8PDWDPe+GYt45AT0+P5nWTLYjUrJCqI7V
6+cn/F+BmoCcgsK+hFTdk1+b6CZhjb8p1WfnC/6DZiNwhEQ/F8dDYYHqjhTs/UCUtzFUb4J3Uw2G
YnyathcDqd7TaM1NW6J/zQUbTwSIASOcaEAwXYnknYLcGdmBflkUbb5GPHbpMzG3P2sYh7Gu2u3D
LlUAKPhScVTrS/onC4y7ixpwpR7iDDLesEyzJ0laE3ukFKlxQiIx6oAxDy/wapLtBQu/GW8wSeX3
iqk/Z9yGT9ZDJ1HGfht+w9jWyvVbEFVw3dlbl+7b3ije9I2GPEZj4SqonNlN8T61qf+8toGW04TP
PjaEEmsHGBRrhHj0glmUcZLHKh3rMDS4zSAV7vjeXhCwgkdtbRxm1HnmqjhPMcoiTwXy1wf1FOvF
XClpNFgN4wvNbRJWOEe8CyROCYs/LQl3Oz9CB+NQn/QYyQaH3NlokGat9Xn0f/C4DoraH2/D2E41
W41jkxiSByhZaM5aU3SszoLWISVNpA2bXlySEeD9BSlkhr8Bok0h/8DUK7YYhW3+9HL+8MPeQ2UU
RNVOyARUfFMmMVKfF1AIe2/SfcI2jF/m4uSlf17l97LZE8Ozrm5U8GNvXMBeEUS+gcgpWcR0CGe/
wGAVvufuHJeZbfdXldmlbiiZhiRfjfEwVM53FAhe+V5fklANmtO5oxE6Fw4IsdQUj5ubyl2FvmW8
zjDXWrjPkyFdQ3SiQtxb3fMi5HaFzP/yu+N61ew0lVzQmUXTuHNS/d3jD2lNNlthC8HZHScXGY1S
mpcsg4vNiY8IrVPSdWHceVedDs3Sasj+GJwFA2tVz4yPvB+5+TqYpDb3FmmHFfGpJkPYnoTbOgaN
z6hsH1l1QxCuwPWrf3dfo+OS3NgAORx46nlf6MrAYqAvOk/Imno+IxO+muwW2J60KdcK2U0YQ8Po
Y5M623M7DCjTt8BsfGR2G3JTygWwoZbwePSxWfIiWvmeOsK+gPOVraPO+wQ9WcxfNki9tVUN+s0+
gC8h9YPETIQ/t9gx+Xu8qVW8j/9LyyPg0XnBDSsQdlZYpGRQVHd/SNRM1pzudIq0kbkPo7mLSbfU
UlqXKe3n4TcyatmOp7MtoCNNNAY2fh+5QNtkNI6AcvX1ImWDaW1uFk0js04jRhhMt9kfzsOdQRqm
WPLZUsFofXtfbgrBlXoT/YRWJEdDav1Mmix4oqwXcswR4CeKHvLVMg/OV8jHYDSjuokaTwluNn09
QHxcxK8tOx+5Pvk4PlZnrLnDGmtjb4d1n8D2kCAa6vXRxYR6s/3i95dd1OQhJKeJk/jDE8I6cGJy
4ydyBKp+NVoN7Hl6+y6aXlqkqjhZcL9MfQSc0riFyzMnfb8pzBSlAvJ2sWB5858emucaAuhSO6wP
6sVXomtmVqgDUijRF5PcGvKN6n/WZyfLTflML9cP2/7K5og+369XDSWaXan46eLGyp8C1s3Vt+ia
wSY1V3DZnDro0QUlmlPfC+whAcjYLxaTbnXfHO+yak6n9l/lD6VKQ4DjyETccZ3J5BUYNImcUdww
ySsZNOEqGjPYwxOiMiwmNWu+04FINmObQcHO4tABstGYTnVGUQcNMMoruFH/nAySyyiyJZF/0ChU
vgru6Go6PAezmPoRpy0Mi5DV3W8lBoxa9erQ9NdWdGbMwXmTxt04YmxlCwPPJ0cGTnQMwztxzUkV
ZPqCLHiG2MBDr6qnQmYQmNK0vwGOgHU9BD37suewf3M9DpbZ6RZV2a5YLeoAZn42mPKu8fReHLLG
HC0pRG+PUlsZpiIa9VuJDlNB0FpC1if2wLs5Exysv/NCmoYEdCXEVD4l64BVnXJg7qhG8pKC4Yya
wiHJZem93pYxt6EQh9eyW9ANiL7kAfRtLaBgOoT2DFUo9QPyO8AZHJf90MSNs25lfpfyXF7ZJKad
CGSdyb1RsO0nhTsV28DQfHuD48JzRypJwFAioY2m+873tUAPx0RFjnUq5sSN9gdH9CCscRBmk5Es
3pUkPqHlwku2OZ5bWrqKi8f6hOnP/tl8kALJlB/aZbx/DyHiQtDVMwXofp+CphCebFEPwD/MY26i
P7pBXGVXO3eEkK2FcPBdLIHwqlbmD2raOFdc13/pr8p0AwawZJhYmT1uV6C/E+x/O2ecet/Jg3+x
81AFE8xoDMKiTX/VR5wOMN6hLke4A/i/uHwxgTVbakWzllz/N2iaWNMxsuVhvTj6cwbDEGr2h31N
D9xF5HuV7EDTUesfVDAc70B9xyOP23ScodKQcrlrf0rgkXDJrH56hZvC7Fl2Chl1j4NBoUA94WN6
tnaK0adU80VzUE6eeL8YpUJQ7FX7xo31Kdc3KUhjDE+VsBmeCKdZKRRxF1tHV1k4+Q0eOGmmY3Ce
lgc5hh3fmRMgCsjn9E3j9uLmoFN27j9wnfNzIRLdU/5DZ2RQDtro97WPWz1QacTba1NEpr9Vcoi1
e2WeIdnfCV+50hsMS9a7rJWMFOF4LaTQPrjrU8J0fo1gmp5yUysLSqkLqtZs8/JJB+0rIVns1e5I
XS8XQYKK1c+aCnnW/XBDQJstm/cB3j8P6g7b/CqiFrJQn3hPnhyKN8McPpr46Ij5gIGXq9/feJ+o
bwQ9kq7ApKbTMtf0nxUV3RRGSjc1pyL/6PHDNEIs2WpYXnRuC0zBPyf9GUnD22jCNF1ugjgnZBdQ
Q0TQoANaQu+pfCBUe/zSjM/P2Eo9Pnjd9tKmQP05uuikIO6AEOWb4ZSJY+X4059b5+QON3B84OxO
fJob7595/5NXCiIh5LbUXy0Zgi8vleiSO+OE4gQB1X9f4LQo8KD8MWEC1yBadNKSlPXLMvGZrtNs
Ptf3dOqw5k0OO84lAtnlDzcbiE+vvqejlcOaUJfjrsfwmsjYIVRDt4nDkZOvGmFwe/ny82jJ86d/
SAb2wJ29mxB1euXtH4xoVsRg1hNpqKBddxLGhzDV5Eqzq4AqYHm8NijrwctDd7WiJ2T1Tdty2w66
zNDAIQVIexZa1KNiWpXHkf2NeCYrhXI8e0UJ3YOiJvM1OedaPuSY6WC09Gg7vAaNrF1YfwrXwgDO
0jDed+x7WQuEbe1tYEz/EgZ+FWZ0xQAHvRPvlqCRe3pgyQlEZSeLi+Jd7Rls5OSb3YMAgLy9WrP7
Q7x7OVvfNR5Om7mrmCXPjsc+PnpPxLuzO02myouRLmT5C67UmYpbpesktauNfROnh7I19rk1sRaE
LAkYG6OEa7JNzw/+ia3qWZ56IOCCNJV+cO1eL9YPKuTNIZIS2cDLkqBbX5/ospGUhY1xg/VvUjgS
NGvd0XZkSK8TeZRiqta+ZatzbJASSB7gQcdg/l1vOKk4g2uA06VYZEn1NeJF1d5Vns7XI6xv9mH2
lU69/hLabJLbPtPCMaoBB6nei9cl/2PG5ehljrtQ9xuXtKHNvyHB/5rXwGZr6uVvSLCyVV8tzJdA
r6z1/onndALXs3EZbLSs4CWLqpXAeJaVMVYj1LebcDtyohdUWUGTD4BrvNWL3tVXKzQ4+Z19NTUT
Aox5D+N6DkqPcUKctPl+9wJ9bnu7/G7SS832c1PesOZ2uuXzGGscRb1PZ9Z/IWsehj/32Dd5dS2V
XEmrG20LAfHgu/MILZGcI+jmeVB6aAzd/MrRoThYBnOewmM1btG9Y6IcaAD5JKpfAMXdVQYs/Ydy
4i8U2SIUUrE3FHP2M5N4kLKZWZKp9rM/pkhcKNec0++SVrWdsqf66LvLi1QlHNJpCEqZCufe/arL
K03iCRnR3jZf5Pvp/zbPr7NRREzuidmdygl6kVMtTH8tJ8MdtMQEinK1D64Dd7raGV4UbsyNa/4D
6NINJ1QDAdUfp/ypV9/AcK7Ljo7c/WsDn47joteXVhseiu5SykPnslNbZXp7OdRze9/K9tziBz8s
KQ4sruX+KeZ6BfNpchuXaAeUMRqL2IWXibcCTYKAnYQU0oUU3Kxxc6ZQqmHHPmx8de0wzQmC7FFT
V3j4cTP38PpTzsRV9RByFJvcLKhhsRObxHbVccy3WE8BjSimsiwuxsLZx60r+uNttlQQhB/k15ps
n6t+Aj7R7sn21y30pRRosdumwEXcY4he9OaoJIW/3F93c/ZmcYvvI1UwKJFwdilEAqA0GxMQH2lP
+cFFf36EorLBZ8Qn//OTYvfQbhGGyKKNecV3GFvUVpUICLf9MuEUCQXHRQ+EDUMbAsY3BiqFD7yo
XlYtDr/hBWJhB4/n7YLC6FeDIlpJfbK76lZyHO4NbGS0cVS2ov29p6hn6WWbRYBToiWLclz7SUUC
PStunkgS0Y2eBcE1NVxCBJGayrApEW1seCrezKc3HO2Rv2gDLsLdfxZ57TSN4OftI8AGV9ghojqS
PQHW92y/6cBXwF/H9kA2ZdWdbtOfzZjpRcL/rEjndTrjLzHLJvrh3LGVXETzWt0Xuh8Zs6DNruA2
mxr/fOODZ9d4TjsPFsgw2OKqyVMJyMCgaXloJFkRa7RcdA3jkzkljEV81gXi87K+sNs8BfoBAvnX
9KQnr8A12m5eyKf9DtHdO3rDou/6S4thfsyUsUG2zO8c3F/TBxzClKPgXRbmv16RrvtnzOj87ZZJ
RxLAfRrAd39S/d4mv3pbVYD+WO8oq8N613ZYalUpDYZRKnxPO+/JCU5zUn7LS7/pEAwzMMNioVm6
79VnSQG2O+BlqjAhe8sCb4tOxCkQ39LwNyXF67GoqAA308pYTheHxSxFMQihq/ATMdh4CkjVDYRj
FnNjtwd4AJl4GZuRbHgVj6B/yxEqGbuQ6Y81Xs2drBzmcNe1BMYlmt64HPVyvcAhkppRCiIWpgO5
I5aV/ytUcdVPNeyv2epb4Yeb4Vu2NECvSAMf41sglZ1UcjrPp7BM2sVTHCZb19N08DVkPNIwQtzb
cgZg8pWYpfy+0EiRgDFkK34PVN95j4vj12OQJpOAzXLQJ5qntTYAMQzYP9v/rI2S/34E/2D14Ixs
3JY35+bMD3a+p94uo/8sOQjJcpmDPINb2xwSM+Io25/NwoubnLAcPBXbNocFg2IFN/vxGLhjOUmL
tHoNyKAYrV48a1P6rMyUE42O5o8O8E1vI2GAv9pn89zpamO/QGHGkypGtvQ5+5kBzGof0ttjtMWw
tktfv/sl41yb2ilsvll8RGKYoA7r8m82ieAb/st+7qljLDKc9G7cyXCiWvoG5TYY1ooiE1WRr/IR
Jl+8bGhXoADlV3T++rPayddngmS++cxm0Gr5hUe817ABjVDErhCF+cZ6wdeKWna44wBIpy7KuCsP
/ySOCpMzWSg2aeCt4yTp1Vycvi7gql3WZ5gukyTbAXsfyG9I2RD6F1w5owJF9uKpXCMHJ8HT/VAa
VGV0URSZmHcumv5LPKZWwS2//IJjCXJFSIzuLhY/30maYzinHQV2VMbf2fV4/pjaDoW4a0vZJZuj
uY0BMQDmOvBbDvPiiYWIFwSSGTfsqZ2oHs6Bwx4IH9qM6NqTMsbWMl74ysxKuH1Thk25Xjd4pm48
CxtGc0o+m6+uJx+1gT/85SFPQPc84EY162/HqDf0TniRh9HxNbAi62p/SrwPZBkkQKA6VKvB9O/B
sX2MYuDEOsLTvTsCjwATZ0E7lnqx1W/UmjQSQH78oa/YHgCil1ds193B1UDNkWLBHkn//+PLAFe9
nXBQjwfkdNprCqbG04KylIlSYmoK6CFBkGVIg/OBRoVcnvaKon6qCKfakQInQUIM+YvckobEoHnu
dRpCRQiZOgEv7mRATMyOOnpCsVyiF3QFLiGA4TpSX3N4aaN+qH45vNdX6HVfs5N+qxc55/i5uoHr
0G46TEHJk/MVsBRipVY6ozn/f8jRpNjOGkICIApLvaBL4QkmIWP0NtHCwKQ8o0lFmCEcEg2/Yw3M
3zyz7hSZe/lIi6WRW6Sgw3LiZe1W1bsGNlNhOP6E9EM85ojF74697gwX9cbnTTtv+9sQWWy9hg8G
6yZ614BNIokcdMfzHn3afm3B5sQYARrnx4wvE/4lDcaol3n3pp5EEN2bXI/0JG//mFrtCc4OLUFS
q7mFhGsfnNV5Hmtv76Dfzjx5mybgLipm1QcGz14nPX4XjBAEbrLX7siutVzi8mktelMUp/57nA8W
07OYbxmvAKp5KsH3c2ZRA0BaEOdzlmPPFFse1dYSwrbf8TfCHyUtrhbRTCbf6q5ZfMKA3UzhI8x+
qDaQo5E820Ypvk9XpQ6Pw0VBuI2UX6N8rzihSC1oCuUJqcV05fPWYnlFowKiP/uLTC94agvDeMZS
7SCvpa8gAL6VgLrByAVjGGHPRfFfajND5jm+YgqCzSmpqlESBuQOLCoQwz/Jq/0P0LbBHGS66jzI
W99Ilu9165fgTxyaOeI92/OGGNFKKE6jOyZkjE5KHwF18Q4+AIbpXhdwMIjuj1iqB6gBTUn9YtkC
T8aALHgm1OGAmX9lT91ipYQlb8o78A8WImMtX4lBC/TxD60KDRs1UKwKj2I28i2dqul8m+oLQfoB
yF4ocBOzPiDh7W9mgXZm9FCK4tJfcpCqJyeizhyIn03CsPxqPhu3P/pLOfFKZuvx2VmIEMWkzo0Q
k6oTYl+UkIR9DRyIUrknuQQqc/Vze/iWig40RCPUAB0dLPpZ+BgkCKYFu9CbZKHqS22XufgNXz2W
wVf0Ln3yQ134Kfn8Kkv48RLRpewBs48LkBzfSzv6GiXg6TLdXV9hyxAqpIHOQqesm1WitaWKR1Gi
TDEdjEZi9tWC5OZeF1HznQNj3JXefrI62C2XbqpG4blz7IStwSWESXtZAe5dcw6KXubfrCesA2kl
5Cc0ULgdLcLfUZ1LofB1AFzvzdM617GNDXGXK5weNNSoeqbsrvAnhzFC9+rzAfRO8aZCtuJkvMbM
p2z7UeNROinJUXNdkZJ6a5lYV4Jpr7kGTl/abHcnaJboRVX028IvX6i4losT5lLfM3QBrkTRpsPQ
W6FCizSK6tpI+fvOh6Iw1CDp3bo842PWFK4v7X/nIY/HgQbLWXe1Ina47KMdJj83WasABnWonS7X
0fz3ZEO7YlH3ICyLgulZqomOrX9hqrbgDIIYQPdfXU/58nhVkuqPUH0nQaCMUwTfSKrtbOaqk7Q5
rRiQ+/CBScJiT0BTY2g1HAHi/QkRmZqLiLW2609zQQHVOIEA+qOYeY45A3KTaC3l3n0QF/WOJg7a
iQMPf7Lh+eFgY04BanojXPcOKjm99NNsos32Dzf2Ye2nJDLwsiHJSzqpfsUTSxaar8mRvkJRG+wq
yD9QetHlMbCBrh9MvIHHelmum+gqZgCNMWqeCjPYNa0FkyDm39i3eDNQDk5eA9OFTm4GqkvhJTpC
29jYlmr1+hzGxa7d2Y1d58RIAhk1wDxaQTtvoGbCNNFOnopUkXmAi8/+9kchQ8nNxhBZ3KqUGH1b
1KUYV8xhZAqNNZzpmhsL1B3yqbXBgtOhr/d5Ej8Nyuhtc0TJH8D2klza/RMkUVo7SJBgPwuCp/0s
S/KW2u4EJTAajK5uZsIqcxhRbDd1gx4Lh4B3YS39Ny432rHY9Am5JM90VJ20RqRQlmfShG6MPgDt
9bdkE5xrNbV/bfvv5XID0WNymKn8C5adBDRQPwpLjcTqpfbvjAxldTLStJlGnM+y4VHdmBI6rcF4
RMrvGbJuTssFMF443xlQEU75+2TUbZjZPL4rx85UAVKG1fYvd2GTejSyBjgU4+L5k5gnBIgPQucq
HWiqv7M4hpTRzyLmJD/5BfyHFWONvU1O6VDO6AndcO6ju3QKV7Av2dJBZYCTB22T6pU6einas+7w
modDnV9DQRvoWDv3ohDrXS9//rSycFP2dD1vPQuIgpyVOJJq2IvXopmLc1QxtXTYyBdeT2N47xkT
qgvk5/baND+Wjz7aNSGhYQ3Ltx0D6X56E6cIoSZL0KCGZ9viIkJJGTaZ4V0ElxeX8hKexzFukPTB
NsyqswdhUY9A9iKXHgCwEtdadhizwY5gIJjpf64g5FrlAQXsRixo+wvdeGypre9wxQPn7dpSQSkN
dg94atmHqwC31xbdjy2cXVXhPRWGuu/Wn0jwCjXjQozZFeT8yH7rXHuHPQTWUvEp+WpJLECo6NdU
8M4M9Jm6BO7LBvZiBIDD0Y+GJhFpwwDn9CBUrkHayWkgfLEA7Wd0/BSUEXLCku/10rpYy74ppdSL
zZdmwGkmSTSkOvP9xRhCm/NNgPx8qjXVQhg8OFPssljYlp4V0DUoNQAeMMvmCLDXJd7vmsDzH3kr
5iKrTefA8QMPgzaXVB8xe+nMPipattVqzi8tksr4MfRXoiD2zxiGCHu6DniPcj2LfbWjeBqiWUjo
GcNONTzGsWSBr8mmY+JW9Amx7Ht4C+pcyH8xO45l8rBwTvdjKAZLB3P8mBVXLqa/S99NKKZXLYRb
3VnRsiESd918ywarbtPGjlvl6KGq5BHGHqEUbqZDB+LFZWt3qZF8OSx08SEgO25MrG1y4mcbq4DS
idLo2kvmFc/adz0TMFe3+bSZj8rdaKbC/o3rrtISxPbXo23ub8i9/Q8nO2mFoi+NuYEsfyrgPeO+
4caii0kq+fbBZ9aGUyjvrbkQh99eQGsE1Peojo1+ChhYgTN3yZJyriObR0olc3E4UltmwjB0cbEI
X199KJm6IrCno3SCxPe+K+17eMTy6L69m0WalvzhrdkeloYHJnSQBNtbO1B6H665bUcuO+rC2tjY
p9k9fqMk05JZ0Mh8BSmgJn5jxZu/jBbIqAvBkuWxW9X8xTSPFQWoYS/PBpTXotzNDHEmDmAJwlaz
loUvaF5j0FY1Hh5o/BSoYRViHY9QauAkGyXwORCFfZhJkBWtO87vuE55UFh3RCk3bO/vg4ZniEtT
TpawWnj0WIv4ym0V7RWqDvfUonBkW0zcT/QgoBW53+R+OqRmu4U8CPErU687nJ9a4yCf8n+ywDzs
SAjS+AvLaehY858EJXf5TjcY/Z57LIOblpDWrI392U6ZRIdlwgPSimj/dAolXWaetG3jko/6H3Xb
9VFWH6EsTyKdhUK4duHX2T3iqyqC60hnwwl4hu65grrTbNuCXk3vNr37gQ7DablnIDsskLw0JHtA
48mu6Ka0c5jX94zdMYvDpJtvKv2zKDvTww0df0FBT1g3ZuT3q5/cEDM7Eo8JuWxYy239V26LhGOm
9tpMALnX9B6scXNqVGPcvGQGODHhep8R0SGW0TnOuLLB1vFutFS4EUEdk8VOALAYjc1hI3N8eoJG
T5gGNgLkfpP4J1ll9GtZKLkEjIcUDidRjgRwkZxmnfK40TByjGi8Gk1Z/ERFAsQJwPo9RhpTi+YO
sR9vUvX1R0+e9qWh2TLBrp4QeVnSwRbQTbeqSXTgsvJCj+IGdmcxi0tcas0AAtlav47mZoONz696
H9eCL3nSQU0dot1IJ+ZNq+dmuyVq0+1796s1XA+b6dRwCjDA58d5iRJB8ssLAolcVtWYt3IR6Aay
M7gF+lSXUKjooVELe8UDa4dRsiSvow5XAz74xZefKbw1UveQkM+bVoSnigDsJPjO5yR+vKe/m8lJ
Co98TATtDKdl9DSPk9/N/Y/KVmA10VmKsKRf3gQfwPDKStNdVxvF7YktOgX2tB7AExcuC74gbqca
rbtUAmc5Yqp14DyiS8cTHv8uED1CotYcoZ4opA/Mr1b1xaIOdEujcCoTvnqVTtpYbIiQLtDQWiBJ
Kx3bamGewB1C9wVnbtuKIl423Fcm6XFBdSH1EO0oW+b0TNlccB1yY7NM5px5hsxyIaiLTB8nSUjR
A5NsUC8UL17YEhOR+7F2UOlNQiw0u6xxKd9ZJtHgjRr5g3F92FPgxa8O6JpRdp11QKjXPxuTtEg6
5tF7Lx5S9jp1KmlNuNzfSy2xHWxJH8aqKRzmZemfEFAzA2mnq+28BatIWpROV42Ie7TjTCi0SGym
63BVEdAukQImXwYTXSbWz/Zd3OFf3ApHdHvDHwH1LHk56glqrXCZ+Mfhf3SE8dTTZi9zMEQbnNW7
9+tW91iZn/nxZF/ETTonzvEUhyDAVFcNTfTlA1JP567KmLGdpGUIn1Fl3KMt8WYoypSW9JIqoq79
BuortKE+awZQJ7hsEXLUrkMQgDHmVV8OfdrtJTQtENHPvE08TteOJ4vrd4Y8BMQ2nCCUu1QuGWi/
eyz9tl7fyETNALcHSPHB5P1iyxK3laa1my2nhbWJVkHDSwwLE11AdtTCyFFUf9B1LLQyoWdmqjZV
cF6EWCp+a96RKmDLDNDR3Ve1XSGuSAA12LNR5NX5L7PNYb5dJxXDjR/Q2wIfIL/faLLKfkQrVlq/
fCBON13F1EY6X9SQSSsy2NVCEduNr4rSXL8CYf+V9sek8OUtU/gkORXJs241IT7A2CvWozVKF7qe
Sua7kQERtxAloimaeuAvD8f5KVVZsYw+6dqisDJcu6aroyXyaXudAk2RUDiB4fkC5XR/kt+2VWW0
SE+9Jg8iUdkwevoeJBIeBCMTJRxamPcnDx58hyHeXuxlgmF6nFUI62ZNqIuuLmXxrb9k1osUHwEG
rrHcPaC4N4WmwyQzTxU3dWg+GYKoJVZq0z7lIN6n9om8N/4GcTFH4+o79mDMKfV4HdvsqrYry1+1
NKnFsNIRwghbBze9R8cNa3MhywyR4oCcOGTDOJG2WWCoLrfxA+RUgRMi4Qyr8RYat6rUgt1Z3USq
iwDp/IKAMO4nvXAtfe90q/NT5F7ZsA7errZ9b2C507fUJXQvOIspxUaRF5MfhdUmtimoXiD4q6nx
lJCJQT8E/dxXUlby4lIRtnGLkZTFHfGnKf4LtotoeSqKbJEmLb1mn9O7zemwuY2R0W3UkSRXQzwB
prwwc3a1m18Wd93nc9Nxt/CY79M8hKQU45q2FTNqKCxUXlFKUdxU3rtPNLY30JcfapLGaZHVnJ6O
+/+jiujyr/SjRuOHMQ0S+hzDL9pbt9/vcpMLHhhfRgQtb4vQdTEzLXo/URiP6C+BjGMa65tN/xF3
adMuUzr5NLVeywTfMJlwMKk6JV7WJM8v3Obhq8v/67EOrmFpJaOp78Ys+sE3X/sp5d5OQ/snSrsa
u3U780srtcNsoxpuDkNbkSq2BSbkf/UOJxAoLl56rKax8zAGxNgybBz4jX9HeYxlSdoEaoL+ljJP
3ajoxq7SFcAkTiepGeXBA7Hac/Uh4FBiPyXVQSDqTrZw19aFSQB+7PwNti9TmsfT/TTfpza/8p2H
qjW/d2yv6YDHWC4h6V0DWLHnEoq0PiNQzZGO88fjZv47miHwhy6TYMJ7M67EByqCF3tUVZ/8micy
DIMIUca1aVAYm1GFYgDBnOk1A4P462PJCMY4R/LLDfX6/Hyr7VnWD6PhvkgmRO0fNysMA2cW5WdE
wVMy3OySkT7TtoQlAIJFeuajF2foTuXUXZTZggdA6sqB0kcgasOT3YCtFBm19oSIusI+rKPn4ASb
4258dPp6xc1y32j7k2uPzKBXdRpb82hGV/aNGcfrXooNE+fcjdgLhFUPBueSwDu8YkfPDLtNecau
KHsZ1xaCd9idlWpxueK+qvsGk0zXtpGTBLSy5QAtIE59NOc0yxhPEwYXiWIGS4L/LIMYTmqEWHLP
OW4IvU6xczKZysyMxlRR1y2yagQvk+4evo/yLZm2JWByobpdziDMg1ybBjIIokmEEbsWz/jwW4hx
k3FbXL+7nI86ZmCx+ccq3JLUYC/is0YT0Mmp7hch/Ytpr/1R4en6MO2YCgt4MBLS263Cg9EgHG8E
2lFILpo+1+Lo3rFOwg7QsT1qvkt8wHYzHyWt0eKg2OG95wcwYwvN1BzOYnFtFQWHzTOe9J5QnLPq
0Qjq30k+dTTW4wsN43oBBc6NowDvU5dLVFmO72Ik17QglGdnrXuN+slctQA82QbXJJRAyvZXAK7y
v7CfBptaCIVNXCilpnmSKommNaIFWXbxCnpMBtG5vgNR7HdjIXWBktTZobXGd7nwmj/xf9gKW2dY
HLOXPvKd0i8PvUYQWYcAWZdZSEiHqtmPfxTZU3vB6tQRNh7vtrNSFtFml/iqzcZRDJ3MjxVVUqcu
5aJSLHFbrRpUvnkqNxkOMh8JHXGZXf+M3CPwHqyRwA6hhb4Sc4wDMYNI/6tonHBJBdvEK9fUUQAd
z0a/ruwbEeK8dBMfK5owqTHTg26OluFdljHoDW0zghDzcgiooSm1EDgvONm18a9rGwhPTAbRwTFm
U3kgcYGFiU2HVmfNoBhPO8+5clzlleeoWDvWpTa3W9IXErd63H4SbFjdfZzZ1MJE/n5UVYjxpk8C
9Y7vq05IpO10SwES+axd+y/Infadd8WxptwT/1UssFC2gNAalNhdRxC7rmk6AxZPWWO/1ilLX5QZ
aC/eMSLThQoAoDAsf3O3pst+OnoZnn5+kdODnM0SsOapwEbbUA4TrzV7SVV62wLbeqgCg/zJAE1l
t7EqkHhLmGIG4vpK2InZ2MwSH0p4ePcy8Ko3gRAM9e5RVb3V55UyoUArkx4CLsNcD+EQfiW5H3E9
J/LwloUALvvu/zkMsbvAuLZYZpzcmGdhgbQjHV8Hq22VLCZUejvkkQpXg3XlQguWm/Kvj5V98aq0
nTCG8hzmFHhDTK78LdxpADTjOi3CWIAuADxHVNkacjrNJruyJmbko4vSPWuWhwUhJZtIzLZ8A0dQ
68AIMF8SxagLSLoKekKuMo59XglMYtt0DNGW5xuNelGEAId8CEBASHvhISgQAe2Ajd4DB3Lcfh6Y
Znji5TcvXsW6PoP9VV1nRmgbr7bFL2wKxHpaYGJG03R70cjxICnDCXHBSOH6J9I6XQvPx5mthdug
+rwOtkTpGrjznuss5mZE0D/y8cpi43enm3fFzkV964R8NYFQMr4BY3hg9pjRYzltDtuiHDAm5MCc
/T6IJqxRX7iZVuG0axazrwM1IAOFnSk2ubERYvYrXDG5yA9UX6lyFtmXAt0iHfV9ZOb+NNt3kGTH
kAityN3AmxvA4wIOw0IpYYPOIdIpTmdyI6+ZAb3YAKUMORxwNoEkD5tXPq0/K//aDIj8TdrP19Ji
GF2kbdaU6MZSpfpBCsa+oWfOGb5Y6l4XCOD8hcXTCxl6qbqRKnPiVZamu4ju/AUhE9WlACSGl8mU
p4ZEiSp3zfkR03imJaZq1HmkSDZ8oFt+oY/R+MNJjd9x76olbOCx+P3+9dGVSeHZcs1kaHcDLZkU
ESUTfNgXtkh1MA2d1lfbT3eCrAOBfIqBvhgUIAF4mQ/nEFSBTXYwC2F9tORfSvi5zS4LureXglqh
WaBkJCgpJjBi0WymvvOH6vh8olV3jYhD7ZefjhCOnTMLiJYBbxM32/hYVIkhryHzLG6cZ7k7nfyo
H8dEBdtEX6eTVVaBxQqiUaHYEgsZi8daHjNod3P+2kr05qv+skISdXoOahM6NztWCANLw+ShF5xk
Q3rd52KEe9uQfs4XpZO6vll3MrBI0vSkg65Hs8AJnga//k2emGg6OLCFpWIhTI2znm1IbkhPFWph
m1oRw/tIAjqu2cnWz/rw3gOped4ynxa2mkavPpNAEAWqhCis611h6+RzOOIPZrtAI5x8WPN5Fh/t
t5eejHeGgT9pLbQn3qpI09V9wr8EzuI+a3OEfH8otQbHPRluWf+rt3B3SclbefyrxX7fogvIvmuj
6kOKz3e2GNr8R14f6B2a9fssFAo7Gf5ML43pzj6S8y2xTr47Yv4YIrR+e3gVh7WKnUqsURK+Xehs
K/COW3qUFe94yKGo7DFnbn3BGmqceLI2nr08OivgennH7LxF5R6ll1021L2yWbcBLb16kedxpQt7
z+RYq0+RREQfT77bLivW3tvAJDGiEl/dQWe4z5ALSjnwvxaJ6LL+W7FbrW0PwJOdb4ulch+ToD3c
FVq2DdJDBX4K+S22zufDo8MieBgX4cBODyq0l2fvX8HsikFbUecU8gV+ALYXkjN99XTzlp0wfYb5
4vFKAijCHjojbQ/3ACrjFljCNeTrJ2I6YWF29vYDhwkew76lndG+qcFXmW4Mkn9yk5O80seltcjB
zlQ4eVS0s26MgfJrJhZD6z/sZfKHSr1kfKrMMNMXiiA/OM3Qwztevf65JMYmVKvi9oSRo+FI+U7y
sVPkrm/0YJd01vqXHkdqyYsxZKYr4l/kIPqf41434DKiRM0trfgo29tcDD6WVkB7VUxDpqy+xlj/
bx6tKHUEqrnkGa7CcAHS2/PdGBrd9G7hyTSmc0Ww8hO0Zc0CjBZ6jpwarcdZLBRw1B2QAY0uR3tK
qRytDcWw4GUduMv6kHHB7btuPQ4VEHvm6P7N3WKHCeJZxnroxdZTlUz18hSuAFTCqWDRCIJErCff
ql38Sjdr5otiCY1IkmrFoo1wxBfsf5zKsVVg8AJHxyfz+PdKdG0ib+OaWwIb+g6aXZ1I+262rn6K
L6AyorpSSM9LWY4YIyfdUaxX5bzYB6CSyjt61Eaekpdmn7zbDyhKj0v8T4Y58h77ReaGGt9vXI8q
oOQktAYwklZscmAVRzmeDtq36+S6sCWuRDBcWQv6X/FxQTsQC71Ko3oOQpX+zREPg/jbzHsCh3/v
/gGP1XtMcFz/18Q0hNpVSKTAnCBwPB/oUxNOaygscXsRmdGtssUlSDqWgy7o5B3RQjh5WvuXgsFk
CSsoKb+1xYuq2iCBUqlRecU49QtddbRKmjpNcBMUPUCZE5vYTEziNs/fZ/z6o0aCLFpXxrMPzauc
8phwdkJwtcf3j1YMQF5OrDvdxxQE9IIMSyZCLl7DbSYC4vqVtwDYAn3WUlU1RzM825eOLs0lpVAh
G7RYBRdLlA1V/ECPQom28QqxzKBq458gsckNtFFJrflOOLW/b+Ye7qZqrdNYR+D1aP8IxYTdoEqI
NqvHKHS9sKeU3eHNRluiylehtkmHChOCK4uac5YgiBtDgP6FV/NTAxSNMHTxj4BZoJjN61u72D74
od0mGEPjtFBhARLd+t6m1u3UvzYnXTas/GF5I4Fbyj7TSkM420rXZcEfU0Gq40yBkIaer/Y36Ncl
gIXJJR7dAxCnSlZRfCpqg3Jg7o2H6qZXyI2JyX1hypirqcx4ZtgeO27cfuU5rcKyiqw+Jc0Xo0wm
n7U3323ai3DDMD2fT30qOBg/7+4z4/fiMVP910iXK7hfIyu+SdW20u5GX98KaNMPs2wE3CTyWPQA
mz+INY5jrssxnUUZKJoDdpiwyDWWslUu5bGQN91ctAHqDqTHvD7cu+Jko+k6xORTM2ZhQ3MjGkFk
ZTIAPhWxT4LrNLtQG0Wc8aFaN772O8o7bJzMBQ5uYkbFOJrRKEBflv1aY+wP2y2y/rfL+XT/PNm5
bJ6vRs16suVEbUjYtS3VLvkPMQKBIn4o7AQiT20xHsmX1vGxp0KSzNoRdUh8F6yKRbnRgJ/YQNgQ
8um8ytVjKLivABGW/LbzxnkRWIqOfbFCGQWM+CVyu21e3cGHwhjV78/IPNx70Op/Mbe65XvyFHzd
TCMIlPWLG2aDvau22T6eualFjM1EBJb1CpX584I7iEJqOSXZw9puX0iJVcHg7WEAaOsw2OahDpDu
Lcup7vFoeBMQ5kQM/fH28b50pHYDPZzJnSsk0u49nJtr6MXEaKQ74QK3HhLTWdNwPOk8W9wBJjfB
j4ZO1ll5AVya+UYfB3kHdUG2muHfNvOQWgBJSjE+XL2JkgN5n/8fRFRoa7lcx4FmFV/4qpcZMInK
xmqzn6Liw08gNS8ols84TatLQbqNjNlUL1qu/EtfUg1ddmvCKkrFpWYcOASPf45EF0bQn9/HJAoN
MoHj+MImbrJjT+7yPEHiPvMmXEtQkYE0rkJ7dZcDHwDS0Hhb907XQNQbv6w7j1WR7g4NCzvI9Omp
ZVKobqRu83kyoNOEaT+QLKPHfRJAi6s0U6PXnZW8HOdxq5GWd1n9OETaiOPYpJHOoAmgcnlBer8x
hXoFqmhS97Lo1H6XHwsA2ref1LwbGOeyfr0=
`pragma protect end_protected


endmodule
