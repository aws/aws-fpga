// Amazon FPGA Hardware Development Kit
//
// Copyright 2016 Amazon.com, Inc. or its affiliates. All Rights Reserved.
//
// Licensed under the Amazon Software License (the "License"). You may not use
// this file except in compliance with the License. A copy of the License is
// located at
//
//    http://aws.amazon.com/asl/
//
// or in the "license" file accompanying this file. This file is distributed on
// an "AS IS" BASIS, WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, express or
// implied. See the License for the specific language governing permissions and
// limitations under the License.

// SHA: f463fc25b8464dd6c1672ff28a603eec67bfcb40
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2016_05", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
tSlSbRy3vdZWR6V9iPruRAfBx++bfwHMPNXyDBiMQXKbxq6RXW84XUgLKuf5Iwlt0o2gF1Dj/gTq
sA3r8Q/yFepRmgx6RtzYrrcpvR8TnBjIArKPLN2DDCmL1R364detzrhgTV0a9l3z9jVw6xgFYqtK
sygSfVpTzke/QPyCbda/4Wl3kK33OzSmKcCzvVNj8YtmypO8EHQZeUr71M/4w08eJIAVBV76JZEz
crBH6zJG+uuT0eGGwIJPOXWwwRM9FDWcATDb7eLazztnAthtHV43ecqSak6npSJ7CbYR23lkcQAw
x/MliqcAJr8SVDasPmAd6nQLpPLX1KRRE9qfdQ==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
k4aggTMZDHk/LG+hZv1wS/bs1zr4SLxpuPgBzXEtCV6cjxRP0C59cOCmS0Oz3WxbzuBpjfA1mNZ0
NodTx749VgDwGwcUMqvQT3kBcQ8z32JQZRRA3jPxo8kmlj1gY+Q2ShfnnW8RZoyDty2ddW8icj1s
5BGuCLqdYmA5CwBTc7M=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
LxQGy5orN3GTIEQAKtu3jis73FwOoQjgp3IGksZFkMiinM0idPwy8hxFuSHizP6pYuoCLz1iMEkC
lOAlCORIuW2jxy3kLzOGr+fNQnqFfAPDm97gG2n0jiTyY3rtgNDUS6UOUVJPWrZRO7b6jgF4/e7T
BtR82lqG9CQ9H+sGmfU=

`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
FFJ15xRAyusP0jNudgYOnTxyyWxOkRJKkxXdoSWgxSjT5EM+rrbJSuJ6VTt01YZjPyZnnf7YqHgI
DmHFcrBzFg==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3056)
`pragma protect data_block
lSXVLdqL8dn78QwozroXZ8sMwDNw90Bc7fGnRILUzuq+FPLDzKMh8set8MStmbqbH+/N5cGnbac9
n2iw+PjHZoM7ka10SJkDZRBUOsDsMkoy+gqyjn0fEMSGoI45LFdTqrH8E3k9f1W8k8vhs9sCIw78
yIXVgBhqx1mjLKq5PuBcnSsOcC0kA7BrIiMwdAW7/kyJzKrX1Bfg5up24yzbcZDdftD8H+nUAin2
1ZsF9p7ygBUwyJNUkF7p0s4PdQt6VzXj+r6dtix2RDTR09kovSwcggk1YJz/JOdUaEOZbeFTS/jl
F+B1RE4Moc3xEGm93G6SmyuNeFTEkz1YEI39C7FNoKTC7Um+KuSRcID1HgRi2ehTwWPod770PEx9
C0PtjT0AJT+e1vAQ7nVWK/7iGGDdydOZV2EakpumGrBxNdQOjd/GVO+YHn9JL4CdPvVXzoVAWaL4
5dXgXCYfHXMUCz03F69iIJu2s1aYzn7AFJEQVQv1DV+NEYHVSVk99A/AA9DeYp2V9rAZ8ynorXNM
SCn8LO4Z25U0otmamV//6b5HzOkkuUi6aufRSrhmUaAzo1/bDpre08p5JRtljGBDvl2lo21vTNFR
XDbsxCTcYiZxssMBIIMTnClp8uw+sJyXk/NaV6wlxh5n6NT5/CVULhj7CpVbum3tq/1kmecp4T6S
xpVWFdEMhgTXz3Qtts5a0e9Wtae8fkZp4Wfyg4LucY2lBGXslrtJFvxsLfz1JTtKgJWrCzXJFqSz
jSQ6SVZeuvbQYCdiXxuCHAs2QlxpJRAzQZU6jOTxQKFyOo+0Ei3JVrn4gqkF1AnhEQoYd7BGnyaP
45xpdbVmfUkmEO9LH2rfyy80GqgXgTouNzZeJJBfqeizs4qvp40kBmI020nwQ1/7/lnSC176ZS8u
mRUkuD/X91mNSZyk0+VWCnzeWfpRs+0WOHWWsb3Vyd+QJzCNlJq90Thp9NxLmBOrPZgIlR/o+7NT
YBh89MHL6UXlf6MlWkzeeqPrXedHmOzuLgjabbDlYt6UJmxga3FmNv8OpGcHxugX24cvGXBwUTN1
0RnPB3A1mIq8drVkBhzzX5kLg4msJFHntOBDmP6azpbVIJCQZ9wFvHMLFUgQ/X1GRm9NCeEFdrk7
maV/tqnK+n+iLe4HhvxLvFC31XMbR9p6ynh/lWFScqBaaeA+luDKggEJS2JQY67GT8WoRLt/la3L
mcS1AdpMXkILQhBG6og3K21/FECPfErk5BP5V76Ah6HuKwCXtAzCnrO+WbhnUjcNZiZHkc6003Nv
ZojnJ7xGfT7VWnjR3qLlrxcFJAmUQMUN+GulzZwKCrqfOQOdu+uw94T98CpQd+EJ3jEtLl+EiF27
ASPp/Eao+fbcwB04buxa3cyXWpSjww/bWdOcTVVRfM4B+8PxZQbpyW7OCp08oo2jj0xHubv4r9pI
8lAzpfTb7j3iwwcOjJqhEEh4CsGAo6D97DVjUWAmhA2cLJJZR3CSZg2U91fftOjZ3PG6D3NTNUHl
z6BDYOnHSWpzmcTJLSBCC9OOMg5puuJ4PLSuZ243cPKqLreokhnVBr3T2kE9fl95sD8iaPaprGMa
UaHXf3LVXFHf76C4dEmMWg9IbR8aA6iuZvx4nE8NXsiSk/S6ThEfNciPs7aPGVK4vbqGMq6hZ1kP
6SSY3PNMK7xQihpY3Xz4fJdVhIKjVVKawo8SgE7j9ckc1vJyzh+M/wOCrEfViixyyVaT90EC0/mD
OHLTg/bJ8pZ657IPgXzUPHpvHO/93l7S2DZV5qVuprMapO9NEirV72fG3i+wqp8z45VhhQkLEmPM
wMZMR45ZR91VJXYjkt/8GvXss0bkLwgHn1HDVgRvbZezcbVhZhXn7kAZtfeqiCmWdGCw/ADz2N+G
OVZ8qQ9qJXV0wF3zAlpJi+jR+Dn5MhDlED6ExjzgV6sCWH0sMwex7WopzxSpwmtRfDC0XYWOx+Bk
FukoM98gdYxPwOouuuOTsOCTDlQou42SbpvGdnLGi7zHcztd2uwxI7q1Gl4IRNPlKmYnUUeBPpHj
nfVm4QAG7pamy8m3MaLEWsJUaQmk7kxY2uSqeGZtuzXBUaX9gODrnzcjoaSCYUxsnjPqnBGYIH1s
3f4eOi52y5B89kuIf8h7nfdeEF2MJOfdcIAEolZ9cuKxsgFtJxnbq6410vw/mhM+fBU98XzJ9+xB
oiW+ORs+QpFI7Hf1PIec1V72ONroIJY7JXhoO8iGxqJyxP37uIKaqKFZE9EEhKXLDfUVwKmS2cKp
Skaf9lotOa6PZL9o8Z9/ANVLkK+jP6g8qXSx50mRQClo5EQ4i2i9yM38rY5+RdgZmeWfPWVTs56o
sTdy3TWw4TPDWgbcTeEjCT5ab9UUhC/W7DwEiSu2T4D1nhDb9aU9k8Zkwqtiu0IlhPzK+8A0UVtQ
8mOgj4sGAFche5Y/5jxKcPdAc8sG1BGE+T+n7wzGuy4mcAz2nLapbiMOlY7D6cYNZJ469uWevZz8
zgeYgZ4lodNd3mB2eNbLpeeR0J2HqmXKmp1+wlzX5S2PJOJP8jWF43kfiEicyrRfCMoM1ZXiejGl
f8DotwqAaDgrWBtfAIwhAJm9q/dNlA6kaEM6pjg/rai3v9mNpdkXlsz8t4VOcR8F0xnP+xFz4FNf
8WACR+zq52ypteVrso0WbnLyt9h9/dohNA3VS75PsTwIN5LEh0asZnE1B5qAF8qs10ERrqc4Uops
x9AHcfW6AhUFx+8FZW6/EVQJRzp75QJtQjOzAgAwZo2QU7IE8Iqny4vqZA3kkCI/7IjviVNqjNQ0
q1NylPBjGfdPJFEFJQbrQjTGYVwD//xnbnHdSn30CmYODmh7UHSpD47lkHBgkjWWynpJYUv2V3HX
VOeDHlYV6F7xAq4NbmAxs+/BgfSGYIZXnD9l478+7izNHjhK5CMsMb2uQBhE0quda9OIuVGwzZqO
0ePvSH1cbTI7WxE1b+jE5lpg2W/RaDFQMatARa2RyudEuAJLESOvwL73xDknJTB959DLancILHcI
UVRuxc8jxzdN0hufCvIeuvjKyMFBrexOsl9viXzI8lBDr15HnnY1zzEabPw3DMc2bv4KfPsAtI9f
MYbYnwdt2MV0tW5HGBrKoYVDl7PHU7heENBszDQgbwDX01WVTehpmqiLKT6JCQ9U9V/wZ7fgCalo
WL7JmbB4h5CzktxN1RVVd1THx0gPD6dG6fQOZ6dlF8AabABCOYFbOI6BbCQhwHxD4j/V5P+aBGDk
tyvPrhkwU/3xbjgvfaUvdJUw2NMAcCYcs9di4F6+IRRHPcC0vjw9AoTK6ZwaCGthhCzXlEqmoZUL
5xbIO/x9zeRbqr0+ISAG+HxWdstilCmRmrC158hgEIIzGGer2m0xiQNEONyulY8ovaCwNZ+FVVnK
DUADXf4ibW7yb6CUswrooCHvbFv1CJXYCG4HUawLzYSnAoxPYA/SBSNVsSAKs5/VOsvo6l6AN4av
l4zmjQN9DcgEwIIVBsr+E/SCIyff2a3Ys7M2uBOuo3ZxWJJaL5Sz75obHxbt6IMI7ZrZi2mDwpFY
JxWFy9zyynyZi5y/QUdzKgOnmFF1cDr9U4eDaE/NKnoXaAKQ0AS4HF0/Od9AtH0o6gqzGz0xZUJ6
q0RXNSnhakXfKLeCZuMthAp3ncTMAXATvjxTMaQnu+e9sh5HDKZOkCh/ZweFwhetkWY6AcXa8NFn
uGuPiPwck8TB6xeRSKz6fsHj2Q3E6O8V/G8JAkU5my2BBYig1dM/zEbL5SxGhtbE+EPxsRz4Iz6o
xuwPdK45oPQ/cy7CkR7LYM+/nFhmKRljulF+HF4Nc1tjElBnnifYD9TkajcorKi9FY2XIPzeC3ko
dXaYJhq0ynWbAgjOSLH72cEwJsbODOw708NuZVE9aP7+PYNwdybHpUo/hPveTapwlueSwwzxKPxt
tQcZ5beK5vHcP/Ca+CR7/TVbZOS3He91YUpsUBsCyBH5fSBB9PUvo8mD5aP8yAZhmhox1rvC1Rok
1Pj4+KmqLo2u9cJ6T8vwOKVdcV5wE5oy3/elT/JtVrP6ITQ=
`pragma protect end_protected
