// =============================================================================
// Copyright 2016 Amazon.com, Inc. or its affiliates.
// All Rights Reserved Worldwide.
// Amazon Confidential information
// Restricted NDA Material
// =============================================================================
//`define CL_NAME cl_simple
`define HL_DESIGN
`define FPGA_LESS_RST

