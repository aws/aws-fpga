// Amazon FPGA Hardware Development Kit
//
// Copyright 2016 Amazon.com, Inc. or its affiliates. All Rights Reserved.
//
// Licensed under the Amazon Software License (the "License"). You may not use
// this file except in compliance with the License. A copy of the License is
// located at
//
//    http://aws.amazon.com/asl/
//
// or in the "license" file accompanying this file. This file is distributed on
// an "AS IS" BASIS, WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, express or
// implied. See the License for the specific language governing permissions and
// limitations under the License.

module sh_ddr #( parameter DDR_A_PRESENT = 1,
                 parameter DDR_B_PRESENT = 1,
                 parameter DDR_D_PRESENT = 1,
                 parameter DDR_A_IO = 1,           //When not Present to include IO buffers
                 parameter DDR_D_IO = 1)           //When not Present to include IO buffers
   (

   //---------------------------
   // Main clock/reset
   //---------------------------
   input clk,
   input rst_n,

   input stat_clk,                           //Stats interface clock
   input stat_rst_n,

   //--------------------------
   // DDR Physical Interface
   //--------------------------

// ------------------- DDR4 x72 RDIMM 2100 Interface A ----------------------------------
    input                CLK_300M_DIMM0_DP,
    input                CLK_300M_DIMM0_DN,
    output logic         M_A_ACT_N,
    output logic[16:0]   M_A_MA,
    output logic[1:0]    M_A_BA,
    output logic[1:0]    M_A_BG,
    output logic[0:0]    M_A_CKE,
    output logic[0:0]    M_A_ODT,
    output logic[0:0]    M_A_CS_N,
    output logic[0:0]    M_A_CLK_DN,
    output logic[0:0]    M_A_CLK_DP,
    output logic         M_A_PAR,
    inout  [63:0]        M_A_DQ,
    inout  [7:0]         M_A_ECC,
    inout  [17:0]        M_A_DQS_DP,
    inout  [17:0]        M_A_DQS_DN,
    output logic cl_RST_DIMM_A_N,

// ------------------- DDR4 x72 RDIMM 2100 Interface B ----------------------------------
    input                CLK_300M_DIMM1_DP,
    input                CLK_300M_DIMM1_DN,
    output logic         M_B_ACT_N,
    output logic[16:0]   M_B_MA,
    output logic[1:0]    M_B_BA,
    output logic[1:0]    M_B_BG,
    output logic[0:0]    M_B_CKE,
    output logic[0:0]    M_B_ODT,
    output logic[0:0]    M_B_CS_N,
    output logic[0:0]    M_B_CLK_DN,
    output logic[0:0]    M_B_CLK_DP,
    output logic         M_B_PAR,
    inout  [63:0]        M_B_DQ,
    inout  [7:0]         M_B_ECC,
    inout  [17:0]        M_B_DQS_DP,
    inout  [17:0]        M_B_DQS_DN,
    output logic cl_RST_DIMM_B_N,

// ------------------- DDR4 x72 RDIMM 2100 Interface D ----------------------------------
    input                CLK_300M_DIMM3_DP,
    input                CLK_300M_DIMM3_DN,
    output logic         M_D_ACT_N,
    output logic[16:0]   M_D_MA,
    output logic[1:0]    M_D_BA,
    output logic[1:0]    M_D_BG,
    output logic[0:0]    M_D_CKE,
    output logic[0:0]    M_D_ODT,
    output logic[0:0]    M_D_CS_N,
    output logic[0:0]    M_D_CLK_DN,
    output logic[0:0]    M_D_CLK_DP,
    output logic         M_D_PAR,
    inout  [63:0]        M_D_DQ,
    inout  [7:0]         M_D_ECC,
    inout  [17:0]        M_D_DQS_DP,
    inout  [17:0]        M_D_DQS_DN,
    output logic cl_RST_DIMM_D_N,


   //------------------------------------------------------
   // DDR-4 Interface from CL (AXI-4)
   //------------------------------------------------------
   input[15:0] cl_sh_ddr_awid[2:0],
   input[63:0] cl_sh_ddr_awaddr[2:0],
   input[7:0] cl_sh_ddr_awlen[2:0],
   input[2:0] cl_sh_ddr_awsize[2:0],
   //input[10:0] cl_sh_ddr_awuser[2:0],
   input cl_sh_ddr_awvalid[2:0],
   output logic[2:0] sh_cl_ddr_awready,

   input[15:0] cl_sh_ddr_wid[2:0],
   input[511:0] cl_sh_ddr_wdata[2:0],
   input[63:0] cl_sh_ddr_wstrb[2:0],
   input[2:0] cl_sh_ddr_wlast,
   input[2:0] cl_sh_ddr_wvalid,
   output logic[2:0] sh_cl_ddr_wready,

   output logic[15:0] sh_cl_ddr_bid[2:0],
   output logic[1:0] sh_cl_ddr_bresp[2:0],
   output logic[2:0] sh_cl_ddr_bvalid,
   input[2:0] cl_sh_ddr_bready,

   input[15:0] cl_sh_ddr_arid[2:0],
   input[63:0] cl_sh_ddr_araddr[2:0],
   input[7:0] cl_sh_ddr_arlen[2:0],
   input[2:0] cl_sh_ddr_arsize[2:0],
   //input[10:0] cl_sh_ddr_aruser[2:0],
   input[2:0] cl_sh_ddr_arvalid,
   output logic[2:0] sh_cl_ddr_arready,

   output logic[15:0] sh_cl_ddr_rid[2:0],
   output logic[511:0] sh_cl_ddr_rdata[2:0],
   output logic[1:0] sh_cl_ddr_rresp[2:0],
   output logic[2:0] sh_cl_ddr_rlast,
   output logic[2:0] sh_cl_ddr_rvalid,
   input[2:0] cl_sh_ddr_rready,

   output logic[2:0] sh_cl_ddr_is_ready,

   input[7:0] sh_ddr_stat_addr0,
   input sh_ddr_stat_wr0,
   input sh_ddr_stat_rd0,
   input[31:0] sh_ddr_stat_wdata0,

   output logic ddr_sh_stat_ack0,
   output logic[31:0] ddr_sh_stat_rdata0,
   output logic[7:0] ddr_sh_stat_int0,

   input[7:0] sh_ddr_stat_addr1,
   input sh_ddr_stat_wr1,
   input sh_ddr_stat_rd1,
   input[31:0] sh_ddr_stat_wdata1,

   output logic ddr_sh_stat_ack1,
   output logic[31:0] ddr_sh_stat_rdata1,
   output logic[7:0] ddr_sh_stat_int1,

   input[7:0] sh_ddr_stat_addr2,
   input sh_ddr_stat_wr2,
   input sh_ddr_stat_rd2,
   input[31:0] sh_ddr_stat_wdata2,

   output logic ddr_sh_stat_ack2,
   output logic[31:0] ddr_sh_stat_rdata2,
   output logic[7:0] ddr_sh_stat_int2



   );


`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
S/IHssS6MP2Ufu5dJBrs0as0Cxk2L2nU05Sppxs2JsR3IjU/VQW8kMuqoEOi3yf7nn3y1/ttd1jm
UiaL3iCNy25zBLcM/4YlIbmVDd2VVdJaa3WAj7MNf8IGRWd3J2FnuZvm0L04mNl8n8rf6MyKpVVO
oDjQ8p5auOsLNTUeWNdEUBm0hKvj/gw9MhE8JAOxdJdaUnyTaorWpDcW+iU2gbxanFv7Ft1vwViY
WwCZYT3j+F66La2rLcG+J9oqH7U34/QS6WzomWee8i/uzmZIm04fVCCQlVjh9xkAbMqI4wQDHRH+
yixOcmgNyRYaHxnM564mrJmgTeN4JYfsx4npIw==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
fIZVQuIz2kMwE7MxSFV6bFIcmtdEYDDxNbkLY1eUcrlH3QSjcF1lLUbpco0ETa/2ftuWg37peXky
egiRGOW6KgLxzjUOIBSSIDWuSyCgfWn3e4qKWbXo3O2pKlqW0rnJMb5hZLYta5soZQSey8AD0Pib
4aGFVnVk+pYYyINeR7w=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
k2aBLMOEBT4UxxJHl+OzgLojFKCLtqewnsZL06srRzsnqvp8Od1eo6Zu29QAq49jX/8SSG7q92df
8enb0TlmEVkqe6U18Y/2Ijtu2K03FzrTuat60v29Bp+cQDsmFWSRB/NrYZH8rrKu1e8iJp9431Id
GjHNdiRa5awt+hb/lbs=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 62304)
`pragma protect data_block
yAFjZ4Kgftnkv9UlYI8pO/rhxHcxLna145K5AgADPYPi1MPZdZiZxDoIQl9nLu4wiKxZwtmfPW49
PF0XRQSdxzZssvyofvgn+Yi5pbIY4K440xauBV7JTBcoBlYGTYKuBhVPVOabI7bmeLqZHYVuLpgG
0mbXxyEv833PURqnTNiF+DaGawNOdybgeZ72Y6w4teeyNL9I3scxEeHtAHYfiTBrPbk7aJtRDp5z
enoyet8oFvTXTrA8VRc+JhJDjDOtjsu3lRxj50pEWm72IjqYnH+aeoVQpT0jEfLdUQvOR0aTkYul
teNRM35Kfk2DXhyQHgg/MBndwyZ6lZlUV5BSxB6HNWCuZCE6rVDAA2ineDbFV4vIJvHxfrYeyVsH
VUxbOGmCOCRcRbItV+gwI9dyqxECMDUOEqpES/WfvTODjyYW4Z6vawXJzmuQesuLRK9sonPknStR
SLE9Gd1fMHDCmsn0VHL3kzXEt6upG2tQ+2cj3Ba2P1tG3YYxApfQ0k3StH3hictYVGaIuPr7z/Dd
gWaesV6VzrjwT50/fQVfPfC0SOw7e8D83D7ZyExKjYNemig3pC3c7kxDpxpl0ikWtAEabHR2V8hq
c/ElJNBybJ6e1dmftqAHsBR3WlHG/lReTQQsx5xYqdm77G/0bAMebqqVLEg43CSzFnoUBP5OpbKS
Q45vQW0QCDuqVMSgv8L3lyZSL6jRge1vqPfkx89ZjDO/MuqvtxjrPMOs4E2h7VWGyQq8wWmXUgG/
5ObQg2vLLTiicT7F4Zd3VY466LmGo2p/yEsCd4PraLxBrjlnVUIhlrUib0OKQbd1FIEXAtt8FX6R
CJIvCgq1a94AN+h8JW78FqzelP4AYCZALrWB5YgRic8T/uh0yiJR1ORT1n6SSkffMfQU62taoNn7
GJgnpkuhunmOejeTr51Ck6osY4SHD88OqGxpG/pjO5bXV41ifsUTAxskISCw7xqpQHyu7Un0KU5M
WEC1h+2B42BAb3fLx2BEdJANYmvUnhhC7IAU7+HphpGmy4LgFOPGcVXE8xImP92Z3IzfhUpTsIgY
2k2x7BkF7vuMg8xAs+VdyCMVFwlVU2VvzOVW8TwK+FwLWJkdJF45N2WRh2982zvkM/1AVoGzl8It
6EC9uiHLh+HzcseIlEHNw6eVQ3M4ymjvR4PzANU0y+RSS2yiUxUiH9t4mGBQ5hD8K7fInlPGQk9y
RcUmYEMDIVpH/+oLoIxPAjBOoueH9GB89gVS2H9DzSQCwIeDMIkMu3LqQlKueNm+T6unztG5Azmq
8AJdkP3h/NoN2Yw6lhbis9dc16tcddsWuwxG3cB/BJE2/QJ41fe0O1+2NE1Rihy+vF5rQiuWw/r/
BewWEPSVccg/jxoBXA2aEXOKVhEbDVgC+Fam3GCbHtH/il8OnQ/sTNNSlHpbgS+HV4/FgGJq5LVS
ByhFfugfpg76MQDkvh8yefHFW4SgM3GxwhZj1fXmo4C6wio5vC1GdAaxaYFEFOWT7xiLPHr48ZpI
T6yCbxWgfAs298qQBBuexOl1WDfVk96WsU/6rULmalkkVO4YkdRQ8q8/PxkrsbkaDYe2k0LfPy8y
O96laJkASJXz73u+ekJ/Wchj+4T6kckqSxtGHI2V6OyQtNwHircGnLOS+Rfm9PFzZYhx/VRmbBp/
hialNBRJ9YXozMNJZ7V2GZKhEqWYDnWRm2rLnmMi16EctmksNgIUo6TUnvFTlot/hQzJYM2HeaXZ
3sMTn/HMvgFEfXtEFrxOObQhnHjnd27Wts6EKdekbNTxqOsR3UZvgo+0K7XyfrBYAItLAHgIpRIV
dpD0RqDVg7hRcZ7VTq8hrRjuV8N+Q8DCt/9F1NCmGrL0uVeej9ZYZYhdSqyroml1dQXTlHLam25j
O1aymuJM62xdSOL96mE2zc+1n9CRXkzRHXG0IMgBPwrrbvnn3+YwdLdOLZyE45WPFZDC7bDm5Vq2
J2cuD23vXLk2NXupzraXuJN4unbEvGRr+ovNycF9RuvT4Uk92WOpdheOlEBwF0HcqGpEo0Bn7h1d
Cy6Zc/ACPgSep+xn79t+P6l81S3hXvrthiMyzSna5XHxkw68da2iXW+7KC+vQRuA5Lxa+srozTzv
Zwnv4dJlB1vK26vomPWeW8Y0EEXeuJU8SGgMAW5+ulQbDWhJR4Yaz1OFl6JUwn1UbDk3s3U0algS
+Awwvzxr7XctBHstUqsJ6fZcrojGj4cR3pUk3dLjQR5ecRSUTU+gnM2m9cwEEURFUjaxZh7Qm+Ps
gAln2zGcHIr7/t4ixyIU79ch/fNOvoQab4hJJgWudhJGva3OTTnCDkBH7MjVAw7DHheBiLxVGQPj
Yg6k3311/nUZYp0DOp/o5f9pFUecJPXFoW1h90p4NibFKKfqfs4dm/Ql+gBXwu0XGtv1+mSoN/13
HbZQxC3821uPXf5opKiuuKEKgix5BTgAbZlvP758NRMlHyXgiFHl0FktW1Y93fz7btPmWye2xe1G
IdV2sgbkKRsHE8WFcrnNLP3uwRCha565KDYP5bJSskyGuSQDc/JzbED2uBefvuU1izUbqxc3N14B
fdXVBRrj2S9DnFFWcWTwsNMhz08EKJMr90/9Yg3MjGwDa0s+RSAKaIbGa38PiZiD0rT/pumEPTUx
/IWjQL6/f8Ey34UvPeSxfQlCEWrHvjgTFwDyDVwWSa+XmICo45imAPWTpewXXkUjvHZNDIJSnJn+
5zpOt+d2AgWaTODkJXxfH5zSNCxQjWzGUtbRnCmkvHr7cIQwnbEfg2YsTcx7Fn5MCXBqZTPORvDb
1swi4bTB2dG85nvaUcwAJm6eggxmxl0mIHULcCgL2whoogPTyNuKk1RbcLQR9F9JigBbqhZlZ+Ma
1GmClrjrhOoAteRvH5eYaBKf3POMosk1uNTNqdkK4w5GWnxWQg/VLhumEnWImP/P6vdtdSR7jERu
SFhISKwd2ir+FVd9i909nYKFaL7xRKQRA4lyOeiTrPYM2u3VHlroM/gwEHpUBg03DqRJVKcdwvTa
JioM7BEryI6UXKn6wfFDhLe6oKCDAxoodQ/enbAr5EuJm4VUzANXXemnTuYvpf8WBYHNZ9rSJ/Kg
HLCfIXJVt23fKI5lUaY+fDKDwzaF/fDjMC78Jnbi93SV0rlxEjPHcQ7IVBhk9/T6Ff2bpo2f0pK+
CT82V9xM4aGkXHFr660uxhb5oagbqjdPXaRnHoE6WaB3rfnTV3VBUQ+VdPzvCohbLRQs3d57l85c
jF8Xh40RsiLD8QVCXmX28j41FSv6GmkpoGyVuDGXTPcfiVs4dXTcFgdhwnF3/16/zOvBcle63F9E
xcATJodEbD0BqkyOaEbkhIRTCNAAeDLbWhxAfzS/Mq81tssAduj9O0KqFu+UoZTzgCkqjS6zxf+M
gaiPWkrKkSxB9jdayCiI3coKa/rVzluYEqLkHDhvgAZr8cqagnZ/RWkm4ItuoPRZMiNNbRIR0YTV
+s9N/IqVWUniGJLizWhAOiuoW0xScRum736dTYW1SORzT8WAav+3SiSqKTQzzH0ET/kXy24GRL+V
xWSwPvzVQzweO/0iiPDd7VzH2EFrRzypxLJa3n/CLa0cMCpVHR6f/a1eQLVRM2iaRQX/lidG4iJA
h0b+T1xRCZdSPxDD3LQ+lpnU6iRj6WfkE+GanlLmGPh+SZuC1oOXgktfBs8J/2J0FK+VNBIjoimU
AC5dlconxPRgOFIxNiMJbnnkskCPLdB2z4TAQA7UGKSqlfIW0lrA9SjkxxR9R4b9PkamKofL30lV
5rYkLRKYoMLIkS1LDrPslizFk8ih1bQucu7ONeQseQRCIWPGR1KarlIDQlYAIebKnUyHZ3iWR6dz
FPpwscIowzqNinGl0BKTuMaTj9kog25cl6XA9PLDkZS+1ZOLJpMGonMWToPE8IZBrS1RcMCV73r4
xzyrVE1BFoUohOrF2k/8uhlMoHiUbc78HX3+eCjCQ6Hw6zwRnlo8jNikPbCtZcixcSrm/A5c760V
ZWWGbHaKyhPdXyUM+/woer5bzuwabLwKIxeniPO8J4IO4dMLLocG9w7vwyDUGd9vAoCkcS0cBhWM
JwoGXSwjuSn3dabJZrHEvHjG7v2660LCqKGJpAmyO7lmIaK5rMUZUGGzYUuKp3Nn7PzETWrIEYQV
Uh2Ay2EXfixGjce6xFwei0TSDm49slaWdTA6dFhjl+STfb7mt3Zlg7+ggXPC9yldkB1WAEiipMBt
GvU1zkxVdo5AcT1InQCeD3MxjarxT3nGV/up+EgW3oQEzLq71VzEq3Q26lQ8rn/+I4D55ZUqIjQO
QOtOM1cVmOOJcuk48DiczRKfUhQkrejXSTtQ+m0+ld9nC0a/UItXmMWohfu9lylmW7vQ1fJQO4Jl
JVJxdvQwO4lcxT9/X5D9o6zSki9HBt1e92+UBKQVvC5UOYp72SyZBTBoG2E52zMBWhUU7WvZR9IZ
+8xtMpbbkYHDo1OElnunx+etM37u9zRT1iXIu38AYJCRcjHRBB5LQMCABRvOxC6r4TmoZQ5hf1sP
i75yZGTMiGtULJZ6c+GzEJIZEXJNS5jrs2aXgkAOB/0Jlz0V2L0kd6oqNwIvbeJw87RzskYGAkqh
ZEfnHEFa0apUUuRS5edaEmmvMCwf1CDU/yIsRVy5xdePoWV11v3/zQ87DjUtFmtiudfyggiTh7uy
jTQbuvg8mQMpecdAR402ziTpaIz/Eo5rahz+iQ0WpnbnL1c4YqyGX/yrHzFzyUjcFZor7X8mMzS1
GnmUhOTnsiL4OnZiReAEg6ouhHAAP/I1TyeqyGofJm8LjqozwFtIoG1Zakig2SoJC4MTMP6IBJ3H
oqBwBuTBCmzPIBu2eGd/+1UaakdgQ1pENxP/XNVuqaG11ecteU/R+4W3td0mensULXg9O25C0ibo
5YeZtRqRQVmMgDY3UhfQQp91SzMomACU0YqDkdOjB5uJdM6LQ94xWU9bWtJ+gFWJuAAh5xsp/U2A
JDtj15Ub9WlBeGq7sFy9PCe3/x0vZBqNIgLKpZvWNKdVojJ22XXYIFh0LRZNj/D81CmC21lsJZZM
wLBgbEAE3QMcRDIM9WykGcEAkjkVr0EHaWegtvKSS2Konn0UHxBjQA7+3e1RKUpybJVcqB7a7Gu5
ehySCdV/tHhJKVxkPAXNHv5eVeeDFf+aflujK7y0PKHZRcdesblJpi9VLjFxARS+JvkgOSosTTEy
xVcFB0jiZBhU+AOpoSmbI2kcOPiwa5lzGAAUPpr1wIETSVHJyksVwj1HkbpK4OOiZjsPWz6CJomg
AYTZMRs+u+CN6MezZ6WrIIcaanu+ELBcX0l5WmYDJCnByCd28h9BeeNrWJycQ8/Sh9y4ublzdfFr
3ou7vd3iF1Ol9pVH5cBJF7OfNCepXrOV1IWNEuwiAZ0SPCObknB0WWALZpGqH392hPjS9yiDjmJ4
T8lHMuuwYBLHCF17kDruXj0pMc3Df7aTyzZK3y8+z2lwBc+9FkWB/ol8FHlIBGCI3DlshAw8EIBt
pNgBKsC8URf2XApKS5r/lLbkUI+mKN4tucBMx3sPKKpyiRijkEJX5RjL5s45p2NMIb7O8aoXpDN1
Ywdw3gFAy5zkpRLfSu+DrKsLKn335YTlqgK7YdxSZAsFmk7mtpThbTlfkLirKDQQ2z7Q1vlS62kh
7FLVdDbHas3RWgEr+TeKvI+m3Ol59sYzhauQFWvCGTnVDX+QZIXRpE1de5WFHv2m+3qf/t6ros98
Xx1AoaBNyu4wXWMgBD6RKhspnLRK83C0pl3c3HRYhcV+F2PNHIyG6SCx/jL0sTXO9f/SuUTA4Z9S
khJZsfumibFWOWYcw3S8kG9D6VJN8jaJI6/ArWDrsr6hn9iVfjAAdIRJ2EwZZ2SuT8tJUpkn7NXf
vdobX5ZhXC7FG/kiU0pVsDsoAsge7/kug5nFcrp11ZakEzhZeDQDLuPykuPLShcbEVFjuskAIe1R
fC4Bhh+K6ocMr+SpfIIiBEACKY/UVIL497ihgDpo0dv7Sf+/Qo8ei1OImA7QvjjGbME0bw89NVL6
ZM8PmE9I4Go3GlTd/6KKSG/OleSAynSeGBTodSFsTyGBW4brjWzcTeIyD8rwZ8cpuOZmj+C235Z+
FHwiu0yh9a7Lef14vwrfdAqmcyMoFDATH6i/dutlUVJZ/5v3evvW1ED/E8UAnF1s5gf4PRyoaG1l
57L1o9NNbOMdQDACxzBTTia/pH2K8t9vbr520dXZfKVG13cDNSarTMnL607FiogG/67ADuUFMssY
UQJGX1iDEx/wy4P35B7w56ev18IPfWJdcLEny9VJR3i2128bzcH88FHlNeyHrL60PPzrIzTPZhDX
+TjfDaug56H6IaPOexRaSuMCA162xHKUdLibuMRyNAAycKx8mESAShtLb3ecOsaE7D5EMC7lB6Jq
jPWU7Bb0/nGXut7pARy2QgZL2H0tM9PWW7RygsrN9VMl3OipZiHFKW3WkIqpi5IoTZuce5SVZI0s
Zy2e1A41U6bYKLzjyDPZvtNR9SYyzgOcSAsa/eAf3vOvGAMkwKU00f2DZxlWIRXG4J1QqbEZ2vi8
NUWPA23c+wNjlKNLbT8YWHUOi5jxXJtrhOJuEyV1M4iuIRNKtPEhTb3L/PwAXG5bxp4/tz1zUasF
LsIsKhwXghAWtTMHrSUlCKyvOSuk3nJzievqsYDFHC5FjHs3+cDK02V52h4QJXqbvvTsChAbUXHl
JAY44Xvuwz7h385uA7tS/8ZpLuz7anKw5PDYx//55S4Uu51AsgDJHqkEC3eQWKHTotZHnqZOM5Fx
sZA55Kghb2wybdogWy4nZo8/m0cVIMRvQxCmJjc2wCKesP5KvjpeIwzCPOsiarWEVt0AKAmnzdO0
HdaPuUJ7lSt0QjXkL8yD5bRy5nVOVoBfZIhGMcT5n11I3q0yCvIPnvqouBRWJpbq1JyV+dNr1RbY
mbXb+QDD5bAjPTt7aQInm2fLADN+v5hmqrvtdshE6v4S2gaEbNHdsrwxkOFgmUNhKgEMiAStF+EP
v7togiHvna4oFbCOrZv6JYggjvRa02+GhWZtKcbWjhAyKbusbWC2av3PGVzsYGuUd7qclRqYYKQS
Y0lELlcc6YCuedJrqrgFJU0thnTTb4yX3TJRvHClt312idBItF235xiYCMHDkpwiGxskKz9fQxFI
cswc38oc48JRH+T0C7Nmh9qczuI8/iceQwxJNHx9yJiSngdQaqTp+SwNLOdScwzjybTe5DKcF9GY
r8c9D+/K2coYC6qMkvTP2fWaSzx03eXZKnILvaNRoK6vTCdQ/15UglbcFyhEuXNfuZzaxmFsaTgP
sXvSXLmrjmNrYCvL9BxcRpxismENbK1W6WM6wP1zPIIwjQk4KVveSMVkf5xUS/UwqNLb4RdNMuzY
avlyAjM2sWwIn2daW6NLfIid8VKMa5dO6UEISeFeJsBh5V31TC52LHMiTbruFFcOgsGjiyf9vWej
CdSAZTRxLE1Z81tpP7NzIsC9Ck4sYxH4Hg2Ne7eE8IdfstoUu4m1zq6P62OuklgUPL3KA2f+8oWr
PVop/T0DppfJjpwPo4tkmTTYjkksexDH7vW1hgO7jEdKgvUv/ePqqlf2FugSF9xXnnS75JqzF8lG
lq5bHYd9UIRUIuZRvG/wOSJ0zr+oGC7FqSOm/33Xr7BuGQBJgB3E6VGFLwZdstE12IsSzTCJQ2Q/
PU4+cQHC6CtW/vM9Uhyr+bNxsXbTtfn/CIALLfGcU6ipK4092/8zwU2VBdypqv6bJ0ouhLoU1rYk
I0rdA/3x1x3sNv3ZfREoitK+YHm3/a4T92HD+6nhZOUVIWI/tq4ff07X1e2jwBotfImlKYbG4YVT
EuEeOTdSxL4YQ+QKi9Z90AgeqmerHa44Iq8yBb3znPF+jmfKQMPirR218pMARxvayVUYrmuZaRvQ
NSI3t3rPvvO1xiQ/ccumO6AY6faWN7wYkXzdX/BpZq2jrNUNmT9v2R+yVC/JHFLB8Uk49jMrwiOi
jLoxdgA53dG2IKmKAoFily0bwH1xqARIct1MFgFv5PkV1lCwbxoJiBIlDab8GIcZoOC8VJyCfYqx
HfitKnzGao6YZuccsLOongg4Q8uobiVUGRA0S/BxgaBMvGYuNubdR2jEy9IV82l8fkhmhwPLFvHx
+HdrP8cdXthomf7IzE+TG2lz/skET236fU/+FiQ0VrqTWAP21EJ6bfLXDSAAZSMDhh1YRBZXW1e8
XXmLQk9XtyQr0ncCNmVOCNW/lvNUpEOvf5S+tpnVdByy4ngV88QUWIF8wnXl+MdIx5C3OPbFebGu
0Qwfo44s0xhRloJMiJN5kxU9tyQUUzDonT6mEIHkraFJ6f9dfx0TiN/VLznJnRhhP5fjapfLV+xv
VPDZzxbHORg0N0BfW0rxC+itJ1rfulqZLuOpFE+pyQTlA+qt9YRyVGGm1oNUHBQ1jOhvXXBj/75E
n0dSYkakO3ekkSRZnyI7KfEl0EFLA/7NneG0nmu0tz/1+rXg5NGHBplqLucX7HE3zUTkx7X311v3
pzawG7pdsKTE0qEGl0iRuqzMwU1O2U/MLCmbrzdXg1/7a/ZX1f6eRD10k9Ppix2oWhF877HIHn+X
k3/qS6IEzlPxgY22A4FXlLaY+MmyqLWqO+6utk0OrNhmSEwBBDRAojvPdz/MD2+T8x+aRl3+ADya
DM0KnRJ+bQKw2PIrpCoOtB7RqBtPxtcqXyiEdLIjEbLRuhZxGRG1VZSqMA6xBGXTvy9epHUgqggE
OAIzxA/de93k6YZ1Cn0maBcmGhhJy/DVvLOiw8cgF9b1lFCnoiXVdEoJ4360W13c8v+uxWcF8/be
FI4N+LWajwbVb35xxolx5S4+khmGL5k5OUzEi6dARminaORh+T7zNkhZn52Q5RiHHJgbzgRBC4Mw
SqXcvA83UUol/wyBwXbzn6JxwVbVdpkrNQ5L1oI10C7iUe/XrsFd6t+mwKyQUP2wwdRRE18teJR4
i5Zn9vNv02APeOi1l8hHLLiInVutmIxvx4JiwByWYA0+SpMgM0RlLfFQC20bSZHYVPCqwT/5vJp3
9awlz1osaNUrlzTirMCOArKwMvMPK9zZcH3M5k9cyxDyvUniuNZy6miXuUIhg/IjvGjp1kbgtFPh
P1j/snljTUdI97oxQta/zYigQddCVe7/po1CgS5UO9W2aJ5kloDHE6xTHFA9BH1uat/edVhVNAsw
KaWx2OP4WXHWzbOwD5SEb1A1g0PZ1vuhz0mTvep84kX4HasKoEhwfiXuCrGw6XTkuq4U3pvUApv5
ffLWP3RR6LmiSeg0jlH15ts7ODwPQcEEnO480igkZmtzLrqs7M8eVSnXu7B4D46cx3aqF4iftmHx
TSgTVU8LRIVIfecJemQhFANhSUH7Z5uBXsvc2cA+tsNKZeIXwfGWio9fvsjGFkZgMsxDyTvqQgKI
KYjeVKtZtWobAZKMKnbtTKVt08SdeGGfR9bAIjAWJOo0iYt+ysP6lL9fOCq2XtWH4++uSkEUpSoa
5h4A4uFgyRfP3AQxJ+MDnaBhOpt/vKaMWTPuta8MfyNXVRdA8fft1cXbWfIi5PJce/Ck5iyVtgQ5
wRD+XLC3N1HIncd8UzrpSYnMLBhDqkcbqu+yJvOKIdhq437hZmT7Y69BL2ga2l11uT30h95NXJqE
neFXqFQ68wbKvp2AeHMLpG1v9+m+QfTVpl6YT1sKDzYc/Sltz4UiG0MlaegAeYvv720KJby7PF02
YsznK66coKdlrrPitb2aIXAMd+NcTXsnY5YRpYlh+KGqWlamJY+9Eb2BHB7W3Cr8IaKc6cKlCR+h
3+sFkShmcIoZzDWhlA8qDbY8X6j0UJ5dPAwziNNaerMiPNWikRGHagdvd0Y2PSXqMTBkX5V1v0lN
qT7HMAfpT8uQndS5vsZWvJNxmu6cqPuZZXfaHFc96JYs11A3iASOL8Obbl+WE5qsMhkDB76odsc1
EkzyvY16kQdJMwH6uffaxW5z1m6FmaxAkZC1554FC+UjapieWnf5by1oAWbWC4Em5I3I9Opi0ZsN
whVb+RVmeKhYUTv2H3HFrCZFJagyAe8iAmt1NPVwbioCk8uVd+Zf12j+rv9us63r6oQvmPTqEsYI
fQ1rAEfGsx2PNFOMsiBZ2xngrByUf+y1xfl6CJzm7RwDooCKSPtpUsD7e74nu7vv0WjsYTpBoMHN
NQvSh/Gmk1zzln78X1zMyW+oGJWuTKfucvd21rhSXccWoadBwCO+DtF5HrS/KsejEYVVU3eow5FK
m0/ddcb4VNOVfGUKrgpwyWnN/rwxV9mB+Bgswmt9PqBHfXgqLQd6EfGqXQpkeacFLTGxmMF/Y3C6
M4Dy1d+QSTBs9Ym10hpXvHwispwJz/ZAyqsHXo1chPAYowF7SmiYVMETe7pEvmyO9rvhq+HtE3g/
2TNppxrIlrH7TJdXF6jVgjQOfChcrCdI1hVzcunTzMKyhS8UjZLwYiXSbUvnix164FVMm+OrbEhS
7CsvXkd2b18YMppWDKVDDEnbFKLP/Hp+f7QzQq+QCjeRge87PXE9aJKZd2MZaRT6eRE1TNeEHj3f
5SoJii5lVivEteEoNf2zJCLvcJIjvywb7+5euWpLtkbUr/Hxv9jIB07nOyoeP/EA739lMRzXAYUF
BUwXMBVUhG+DmUy6skZfqSq/CkPtou10D1Z9EO8J5x84kqIe/SWobli15FT9QGYomKvvlVEu1nQH
cazkcxO+2Di8QKFilSIn0kw4Uj1EoLyGh62AO9VFT6DeU7SF2fEPp+tHs5J6cjPrMP5eexYyezhW
gtlo+51NfEZKdQwrbHwTXqFqhDn/pnMJzScvjm3trdkxNxhZShUadd8VHSfbUo7XntpkKljY6GQj
1plM9lfcg1fuCINuod1yI/U/uRcoHgyTid9g6AQ/E3tgq3b/HXr+c+lWacgXFnAlZIaCrd/dS2Lm
vBaAf6b8l9K4ORga465Lz0P8v0yq16+PfMtgO8i1nS9KRg9b03m+1kHu7bOhSFbM/sLKnzMvKzSo
DVVj8znXXp4lfP2gcoSjtCajkdQgCzlygkFQKc5E2vXPEupkwsJneVBVPtMzt6bxfwK5rxAFG9N3
3DK1xuAAI4ufQu1cuVST0SHKLB+ZLTDF1zbs11FESj47Dd36ycRSDc9QD49V0NOcKMomhvkqubYE
4i6D2BKFj9E/tw5PB3RoHlhCOQADEtdxLssPRyfOB0/v/ZIRDPmI5eUQNiOv5S2oKqZYYNEvVqc5
oF5CcDJdKCDKSELNoGaa0BogMmcmex9xBZHLMj6IXOeEdKqBWnT4xXKj7x9LxvVLhbTpqeoWinNz
pNqKj/7Hf5Gkc/v7b8ycLjtUnzGHxklEglNl66+K+ZAO8/hMdoXSm+0VeI2kZ35Y+M5P6ptCFhPE
WmW+DICfxmqZ/FcjeYQ0qLsWryDZg24rtFtQfwAbNN7Dsk/nZdclw9iOE5FX94dBENb9asYiuRnz
AOt9twg2Sqe8atU0EnkMibdPymMO/J9MuIuWa6LaiI3ri+YmqVv3KbDqv2xhL1/QNWsB0GGhC93f
RhjEnsQqitnVdZJcZP2W+oOFj9vYrjsaID7kI7pDBKjecbfNAMVxvYr82/jdSHMT2RiEa7DizzL3
tJxEupxC2NL43GvU/VC8oDuGcH9m3L/6buvfZftI1HA6nePJfB8Ql2SFU1sLO0O8HZKGC9FrV7nr
k6namytpYC7PZAx1/mAUNHtx1Kg5hTc/d6zwqSM9otlgGMJ2M/WJoLnJZxR2MXUgScn6j1fd85tn
D9QfrV66M5juyTd0ip8FAhJqkNi6RwuwkQ/y+swQgxNIYt49K1GjfFvtxCBPoiymBI/sXXzj5cIi
Kq4uGrYPk2l3T7Sq++0Dlfby1DdSC3Bl0N4RiNI/P6+iJw3ZbZEMWmU92fJ4hcPPqemrk6FC0fC+
ltdqx1xYiSNFgVWVDKSYH8PigFPPjc7b0JH28ndC7XPqBRCO6uzkpqO0i4NIaFMOwNKzWxGdUBgi
II3SmFznrtdhY+0UCm0E0ZaTbC8/hienUZPqoDtHXY8hfvwjojocFAdGAQTyEmnqw7NtXRPzeXyf
r9UOFB6d299LXHnXOyDYs1gMtyLZQHgyR+gCb14vRopPOVJMyJNb5N9lYMKpaOugdbxDrp58YQR0
OULfxc7Gena4ZHpl+EhNF/m9/j6pia7+2VHlGlATj3J9t/3+b0au/TQc5hISvuWzqPYkHSCWPxxW
83/5OIcrUcJ5tVs2AVJ4j97sfJnMeSiFw3U/uloK2rF+6HNeolBOyaFZNxltN3FEf8yJgs8aDkNj
POF8ttOXs2+UtfRp7zBT9xmgzG7ZsMRTp0N+c/DZqdpCJ1Tm6mcgwcMOsS5WRX5qwjE/gDXNsUcO
byiTGFHa1U5qWlUBu3MS/2RjelcAFIj0+2H1n+ysNRqdttqKPiJa7cYv6Iv2yslptioB6+DdmXJl
CywgBz8lhXbD4SUXOXOZXPuAZjWxXl1zk3gcfTjmmYePZYrL5fEq3nrpqMXYSw4SpSMZ+MYO28vl
l13gO1SVljLKywGUTuE8jDpwkcM19uVRI8t8zX49Z+7ZQior3p3Q6CPxZPBsCVWCLFVW9YBKpwkv
hPhBNTEjDtKiPBEXLI3KSkdYT1f+2XRWEfurVe0IwPY7k2a3Y08jVAvKTjnehU8HADQRdAWhecky
5S0VxmBR34ZA4e+Bb76BkVTCljNdLBLTFiiGK7Ma6KLtF1NWoExvPFq7xzbYEWHyPlz9T2d+9YXX
UrcVuxVTRH29uFDq4qegqyoGRI2GNs25NS/n7uAA/gSIHO6v+hHsx+v5EcJ+lPIk8zGp/1NELuQj
upF8ffEKP2/muoWLe6q0OqAPMIk+Ac3s86OvPmYH7aJpnZOa0w4TMaH/ykh6dk21hz531hAeYnKw
4xzl7xJyTmRaQjKhfr1uk8ohBDlc5+QhptoYgRcxyd5Ix6GV0L9kJFrzIZ1HRw74zbeWA3tUFzNe
FEgNLPZo8XLvcIzsvnZOmJjG5kVrzgpkysX20vY/lIYM5lMfNTCk/0tErzYM0tgLdS1kYt+zvQA6
sG7fUGWiUnYyKpHItWpsnQxHwpAFb/Oqc5LDPjsH/Ue7+ITduUJo0WRBhcbu+zYUmpA+KO/Z5+KS
BFu/ptDj3SmGiO2mjpLvOZnBHq8bogkAbO52oJUvaasi9jnUKeWSIhSuOe1mcMAQrSwF/R9nRi/Q
aVIMT//FQnE8vYtCHbm5L9eMefoK8kFSuUGOs1+tNA6UdIW4qfdBeICMeEQoYpfUCkqw5I43PxRu
weKud9jp35Hb1o/KKFIr89WMxBpPFbt0Kaou2Yhdd+410MihUvWyhYkYYPWSL6tnj0YNevbADHwy
J+Rkce2eVEoDed5rWES4JEbRIngGWxcjkKhZEkaNd+7F1PR3SNpkUO6scKAZmVK0YQEmGpxL+fyL
VVy0zJCA2LLzAo1rOmEh1pb3VI41EgGEA5jeJZeE7RF1PiwUlpel2j9gOqDVqDZKIkZc2nxa268d
GtGdhEURk4OZbZUMg9HyQR1yNM9V1s1XouKkSWGYCoUMjMDQOEZ5CtqikFb7NEfN+f38f84Ul44Z
TgBbA1Aa3Sor5FzDgwlmZonljuE2VVzNDoeQXpy+AsiZRSh8JYlRCk2iTBbEIMgEiUoa6V+6ThUp
hcXUdjSURpreaVJ9PRcd7ygptWf3HufFw1K9a2z2C4KDuKsRwW0ygyRQDp87iIgSyQW97l1oCA3P
IqHQRYwqSIiTfCHEp5U3ciTB2TV42Y/Z8sCs8G/G6lPMG0i5es/tMvVWczKDfBoTPDlj/+IaVdW+
2Hi/CIXR1q/vp9hEc3AOGcpTCx6T2WBMpX+UmfP+z8gvqt9oSb8XntzWwUDLI3Y08Zlwng2c5r7u
35Q0q3sszZE6cujpEsuJ7EP9ZLLwX1fImNgRqI0J0AZw/K9d8GbGLgFAhHo7FfFPQQf8RCaol3Q0
P/FeHuRtxUTma+qnXomqTES/o8snF6o8Ir8qmiQWVPJHR9cVgs1MdHz+6WBzArcSnyUrLk7I+v/0
O7M7bbQdTNTlCzciMYSegD2DAnPxNXUKb1ClhnwVG+UJPDFIP7C5gk9BaE1hppnOVssGeAMOmCkZ
ObsMQ4ArlvtC0xFPur7VPSfJRQT8cAXdMtBvzl1Hjx1189FpZixcr4Iatu+1H6a5Jn6Unp1uXBQr
yjFqvKJEaasQFk37jWfLQExfWxEQYDme3cdXOgXZhYOPP40KhA392ptWDVY2rmmgBxNLWBx+63xK
rUjzrtNXqLnZvFEVZ3OfByqGNOGwDlGw8B54oJYRZGSRPpit6F8EY8lrS7ErqAHji8kOGJU3r8UT
yvawt5P4MjAYEOx1Fy14Zvf/ILGpw0Dk32hkWNDckzWzjvngpDp35lQhJ9HwwtTHlQ6l9XYyJz8i
Zj+CNtTcJyKSlYvWtK0mMLq2FJh5VawJ9GpDjlmJv28wlBep9pbGuh2h3+f0snHdBy1fI0jMk6vQ
9KeRxdp6HmEE+1js9hjhphfgUDVcdoqRhLcEywEMHADlJ+tjGsYB6hOVifYiGsCiwtiUiFXx0J9H
M5eAXbsTP5/zmvACkiQO8hkS46O4zxoGga37qz/KMMQkl/1A0GfYZGHtU/R273ah4P9hSBX4fbtC
Su01rOzQvTlf/J7R0G6GHwX8rKhAOyRuMTcKoeHYqbR3hoTcTTJp69oSmM1xod5QGDxcIaidWuVi
/wZMoD/8REYgOUojpqgmu6ZNYG4OXXGFU5KuaMMv4TTnyEoKiCl45y0uZ8uz+zbDQXnwHT9iVvO6
OTv0nOomuOECbP/rfzgKlxTfE7WBILDywv6+6OaJtemKS1XJnhFx8gNhY9fxn5N1/JicxGjyoi0O
KoE+PAhK5tT5a0D/uhRObzSA855l1fxBgNTKbu3XQ94qpAtXDMoPJOYSzC7NuYFUp+ZybQ85FaIb
ac6K1S/he8fMfiGHn7IxE1xyvTtdLk4n7A+fkJJIxwtNLkPSei30uPekkJz6siHVaRLIDi1JHKCu
FFiKQLTusdgl/gPTNtlindUhMXj6LgS2aeME7VJYjL7gxxZHoP1c+39eoiNElwWVme3X2pS9xmFG
MfJTHnT4e+H6KgKzl29q7J0JBDNoWrvMPPRGlVfFY111JeX7DwIv1KF+KggxNSnzIynNgIvndoul
5pxJg54+wNopecCdiTQ+BOd10k/gTac7iQOGG4Sr+KgMTBLUn/H69dvDNkw5qFavs5PxZaWtXE5V
7FWqv3o/cpcV/INXz+TOCCQegD4JhyEKUwtDzeK9AOxzIHbu/a9q+pwbcmLtFJ4YgrwBctxVUkIu
dCNxNLHZBVgDsvP4TGG3xSD7F4jambmtMwV54Cufc10N3P5joCvz2ZvuYKzXrlwm6EQ2fe3GS/Ez
UKJx4ePQ7IVdMiqeMacUonirAbXHjXt60pzmcBhBxVsIA7J18L9oB9bu3mhlsDIkdBjBsAuGjH9U
E59tx2hNRqozlWtYxSHzl7Lf7FsgP2tY877Md4LY/71jqe7HDSe43LErPd0yLyCwUxbUG3HZg/Yd
U7j48ST7TNMEPw3c5EY7woJpfuVg8IUPEqTnBLzp+rHC4Y47m/ZAm+nE5Il9IiY7leT78NFRtqET
2nPH38Po2Iw66VkumQvWbVDJLdZyacObG7v6IPMYhawDKo5/cnh8toRjYyIRgoJez2ztH+abcZrd
X/+o7imId74cIs1FxnZApvr/6VBLRoqH6tfrzKN2j/vZ4kO43PpPZoZ3V5EJKTqVWuZP0g97DkSY
BJtG+l4F1yPIjpeyw2EIzL55YcBuVntoQip1fBorM1MZt8cPBFaXH87G0TPlc09lY7csvXGFIQav
FgjEIDvDgPUwuu9s/u7v+/0E1gpCatqVszh6+z/Je/4NPycUgE/e84FDWx01yxsAlCQfifinyx1w
IKZtPElOlTfjh3Kv6bB5QIweCw50MpY5AfSQzGNZWdClgDjNg8k2D6Zusq+a/y0Do2g0KLmnBKBO
7RIEnvFyMntvkwjlpL8Hn8F0t5VCSWk1hqaM9XZjWSAv0UvC+i+NVzgxxE+DN3AYAyeSbax6BSVs
q4+P5BadaBkE2PCTck1WZclVfXiWl1TgxUbMb2sl8ALhOgISbDCMbiVrD0GTXUP7F3QDNvtc+VD/
wvPT0fRuBYXcVLb3+OCWRzwsihFg+kUUeuJlIaI5bPz4Fewfcr63PahErNnKnzmQpQPUDjfNi6Sz
LXqMGpV4acVZgQ2ky+RkRLAZlLEfXfftnLmMfpZB2M4muaz+cpsN6AMOxEMVZk9oTKzfMmKhcKFS
7KZcnxj7atHMLGAQbMBFMzXbTloC94dO8xa5IEL6LXg1ZTxTNb1/mrpyxWxnII4PhTU113IXsDtJ
dE30Dg7DWW7Lt4tykPI+mVVWh7EdtRjgRobHggODbXebrPn+hG2M/w3WoZjA3Lmd88NvaPH4W+aX
UL0FdTkqhlZ5WZaZWqDkKPkjU18t34/xuF1kNtDXc0pumN178VkdVyKig7GGtqnXCMFVS9mA+E9m
3yrlBrg+u9UVABgmJVKgWl8vh/6QTNopyD16yCQYhnJtlbNo6otB/seVg61tVaQwYQEbbtvyxTWi
pn1NuBKzv5V7k8zXKQv4cdZ2sFnnHZ5KooLrBtmC8w/pXOSaKU8iVWe9bc36TeMbh17ftWzQ8uvD
bRm8S1K3dtf+L1l0vj2AagB8XKC1UB//RzI7d6sl5Up1eIvSUbZdM/Hj18ilQrhsvirYChM5394F
uqHmlHulw3i1gPzIVC0F6qaU+mQcugs7YTAjwpkZozba9C8t/MvhfgelT38x1iH191CGVSGmTHOz
vUcpr1COk8b2J3ZdMpdtv+R0bZQlf+WCXXXyGzYN8k2i+2mH88+EyJL0gjLLiztbjHIAKQQU1zJ+
hp303sP6jCe5OAJnc/XYm7tjKrrnOF4S1VomX4UQlc/dYly904+CYUM97vsjbLKgkVwAe1QZ/AF4
BlMvxoGTsAa7X6KSrtlB50cdhCeKXeTlX8Z7qBKXKqZZfQtEa0KagFOinVg8Rk9JK9vQvP5pfBaW
BzeKWx1/Qq4XdmSax4QK/edtkCqLRVuczQFuKBVWfDgvElsKcdmYJL2vOy5NQbL14gazYM0iX+QE
Ckkqfzl43v3spGFnM0P/hs0HsUNgsTxn5ILyAlEbb9JdtXcb1+dBZboQO1MLkOJzugWNMHOCiILR
gUF28QeWR7E8hSemNngsHtw07mtiLi2nY8m1oadXjBDiif6cg8+XyFhjd9AvlPsouwQddJt3fIH4
HRnx3rDGSktYwIiDid7PKFddsJTA0LhEh+jlKKU14ZVvJ7hXLg2pif8wopyS9ugzJ+hRvRHrmORH
16+PEk30U0kjDyxv0wl3h5GJnuMEbfl5cG7SIAT7osStiSm90rVMyuLYukGwdFtyFV7KDO5dTFgh
323+bKbYaRTDKOZ12+sTHlb2FErMG7ISFudVczz4m2+2yTU19Ak5pDweOeKrhsaRPNc16CNL+H49
rlxHIqIjuVDTLX+MVwM7BOOAevxaaXUEHMsxWdyjtWlQ8QaXCQ0+Crp1gZC5vFRlYOR9m1A+zkez
uxAryuLW98L4B9ZQLslWHiFCWNJwaDTHDkA5lFr53YRdqIC7nARxOyCRLQTK3cno9Ez3f+iEWApH
vz3J2Dukn5Bt3p9VYaZVlgS5Y9qvc8EyyCbI5mqxrrpsbpGaAzx9GjSrUahVfJzoc94RTOMV2Xtl
Ugocq9WrRHeZwGgqjNEnkU6qsMEHbzAFC8656YC+EpKaarWdrVKxeGpKMyVQWhTNesEtCBKO3ax7
TEeZljDVGkjnZIQ8RkWxzOomY7iJT7Tcu3QFm+XQTj+S3iHO0QX17aT21ExuhGwafDddZ5ZHAAXz
Znv0y8hZKs3oN75JWYN37rDBZpYK9PCOoCmz1zOx3xma0OrkYIT/35bDSiaKOd/yYxK1dKP9qQUn
GGNbpKGJGqbpe65I6nLKqhGiI7WTE6DMsHRqQefEj5yHMpA61H3fWvum0jLyHwg/YJhrchmIk3Wa
Psc0fPx3ChaK2Oet5QGilnXXSDR5+Z5uR0MM9ubCSuFHeC2foyllfCS2Ub9xqltsjn7Nj/StdkQY
SMlbL/tbL1oX4bM6rox+nRexxtSENlVAVjTk0jTUqP0fgL61voo8ZF8euAABlioODyXRYKQM+Fsr
C2NFy/5KfXOzB0E4G8xeo3y/kwbcaCxaTBtGdKb/Wf9r5FzVvBaJcDzjxXeMErmLV2FbnpEDyuvX
e4KoiAPFanYG+/ppTQe1v4ymS45QpvaeGXvmaALeWVC6evgu10+dFsn3f+MdWIK6OfaBpZDehxvp
f+xOMPA60rj2f7JL61H5/YXui3ckR82gCVDl4tLL98oFfPXtjUIt3ZzqjQUeDxWpjwSOuCoqHIQL
+nxhwPrP+ybdI+GVtlSajnggS0MFPyeMcfcGfgyhXYonf8BHmDJZZ9lDtY/ybKbdY01W9cXIR0Ba
TrxJmfP5R0jBAi4KlTcZqvqWtp3mn3H3MS4fkIy2upe9BgDTfTYENipqjfE/j7+MLhrUv2hdwPKq
n3jXqN1TRA483WihnVfATs7N7Hzsg5e27iQvfzqOcI18qEf4eO3UPQgCga7sX3frQKensoUq80yb
fYpDEGX88dmOG/594DouzWr+2Nul8VY+hxA7JDIJQZqnV50c7bCSfxtsN9fSLgjf8UZ6Rj/T4iB6
Gz9puTI7xUxxaongnBrBglzVDFWijJlq8UrfjIjRcs94QnGXkEushM5apMQfP+Q4LfwO57vacle1
Q40g3NZFv4sOr5atURhINPlR/0RETsn6oCFcWInikd+coB1JIfyBh78UTdyc2Pw3/AWD/K3hRzAW
eJo+MaPMkQghGUTUqKDzczQqiOfcJlGEgAv7YIqAFFmcrlnAeBa/mpSgYMczuWWeHLHILuo94zpU
39Zyqby1VnfYQlyajRO3E14rBhNhTQps4BsZcpap49NNBvIjGNdIeK8IZ9zZxzPQqlXVfuDUdWst
oVXv6cL8elQ9DHQe43rDt809HAxfKhNZiYrGeHlW2EIYUodcKJPjh9orl4bdiXOgY3Qur5xG58w8
keDqIvA2LbzmX7HOvf6nUNMnby/+ZUcLlza3Gk3+y4zDAZp4Lt3P3mcHTUJ6H3+QJbURTQWTEPzF
GSP/y2OrkrmULtSXrBKfSlEPZfD26b/urctlcEUyxdaQNJ92xZZ6Ekr0RCUHDslGGHfSgPJ36h5r
J6noBOZfHq9EVnluwEAh+9ZH/8mtYTMUyRCO1cyCe9134Dym7WG09TJEx/oMTnsIo+q8vf7tfsC0
HLW9O8cI5CTJ3V0xGGXoqBTtreWf7P1/WImqMqHQm5kfEb0K5hy3qx6+YvBqbA7scDol05UMmZJ3
XHaPax+Yi6hP448tfnHBtqqW9goZxWz487Nuy52fBZmUsHdNkq5GKDCN6BQ+0+WkcW6k3bAseLtN
eOgfNhdKh/LcOg9qATnFRXmP50395dnwIIROwcUgVFUmJQV1Lb+4TtHlIk6LYs6r2oj7iJDonMk4
YpOOpstQW+bB21z6wmJqPQ9sGkPip2TUBdVskvwWelyUudiA3bLvLZBNQAcQcK+/U7hBanVUM4oN
QRipyrgNhcqKqEu1ZK+FPOC4rHRwNBxZF9MBAGn7OdRwXCUES7Ov47JIXOfpxx5YWgKMKp7Ew7S8
fhRHmkgV/dCMfYMV4af8hkFKz8SL+RJiu9VbPOcaW7+kmYlNS/lbjiwng1n0geNO5PFmv7dpUgJO
/zgku1Wg4gUo6vn8xUr9xGhsCaEqzjAt2Vs5+CkgMIDobmaKRYZRZ0ugXfpthQqhuxofzYutTK57
hcZgzTKClNcwLPVlDaYfSEOYucEOIxFZdB1xRvkZBEIItWtIjS/yRqaqVch4Xs+ZgtUoVB4IM/kF
GAm60iWGBQ3CD09hbvyqGvIEm8ZnEBLmhG2xOdyE3gjgA0lzGeZ1XEkph3ULfwTDWRk6D/D8WUfc
ARfLlq8XzCAZkfuM6LQwLnUPnjSISv+srVUrPCG4V41eRldAOr4Zrq/aJpi0hlnJsn230deT/oa3
PLkA3LB5ln+DCu0Df9PJS9BmdhG7w9iESSo51oAqrmgikr7Aq5FCN923f028kNNPfFs9G6wYe1CG
vJy1b9k1A8iI0HBNXa8nL/VAKVeFizngBEVVgtk39uHPEaPDOGS8s9nhK1/PDz8OpB4T+SzJdxUh
AAae/AwrDBB8YW+DFFAZJJuAhBEO7uSLJ2MZt+1HKd628vm8aob1ju1uxpUUie1dZc7fjaTl/4Gs
1g/IlK5DA07GGOtwZGlTBa9JZVnY20oUW9l8IfJm8nswAIfb2LAZvtNnKVYlHXfw0+HSS6Lt/1lx
Y36laiiFISboljtTd5pY8geNr7DaHEf9a8kDmd6MrlzoaGQ23iATlax1BIYyaLbiSMwlbElKmXWr
ylxNFtAUrEgtAUmHopxydPPtc/He7VcyIVmDMx6dcLoU868c33zg340BoFfxjVonM9NClosopgjo
I6Ncx5IQzy5SJEoNqxAVDg07A30wQnFmZEsg+TbX/WjmgY+/9iy3VtKRB5hWej/zqQbQBAuqREVj
2Zcm8+XJyiyf+RfkEqiKHYhlszzYFizOKSlOcyXo3pAxa10ognwj/LxcUVDmHbBmJrR5LGVD7Xdw
IPKNwCK4vbKyz87ONQRQf9f/gnVUFxiG1I7BVw0Sc/sMWLuftkIEZ7QPz3BXzrnKohUryvH4o01b
L67wSJbLvGXY2uHMnITWJVrkowoG3m+D6Y/4qi+tM6NDdLBfPFwzkCZpVuL6jUEfVG21us9xYz5P
MWQB5PNTBUbgPX6Bpy8K3TrWkCMKtpugQKDzGmmv3bYnd99NIxuJHEci1ikJe6bgUdNzxsqiEyX9
BO0KqhWD4iSMY0KPWdZXw4mk4c4JvfmN6DgZC/8m/C56Lv1Vy3VrT6cvxFtdk0BZ84DTHXDo9FnD
bwKV21vvGSCEPaDv9hoWyErk+WABLNyarJYEPVCvqZjGOeAP3c9z5AmjS2wp/E1rpfvCFfBcFGnl
Ugnj0pQwJJ/SC8h4SQ7kSUyOCa56YKdGPEUgFFVxBiXPXGGHKGzAm0zfvnIYBM7ZSxzh3H0om4xV
5ll51xaAOwp7/fUdCmERNxiNaBdmmBnO4KGLz5RNMAAj/wa57kRBXuOuakcK2c14FKspYgMExyyj
pdAuOp3B+voLHX4jZ2K967L2YtplduZYqa0IuqzIqYrvP5X5amGTfd8HQRPhDjlUMD4ZLLFsTLD5
uB5ES0D8/6nlqNvV8TwqnIwSDRbAihW4SPDpeAJz88aaLq0KYPc6t09ajuh1ueFHlbSwntoYwBpL
risdUo7gGH6BETWn/AtCpgZWKIXzh7wFjoB5dTyn6Rzy/3KI48hdtcl5IVN2TS0s2rXGtLEPN+P9
ffCt/GqDRVp5exXRr4xCqYHwX+jpV5F1ykvT2mBC0ik+dTWGfjK7iiv64z9DNnfwBygjLgBHBj6M
rG0FKe1WRAVAwZvVmNtTx+8gmNbpWG/fgnWHBaLnNKEZ3y06L30crr5dnI6THjfJqxYi9LKfvGtj
J2e2ntFjdPxmk+V0/Xq4HLMb2xXsIQhDFRe30o8XeIRPQtJ8Th767U+jy0wTL5CYropnnvt83ay+
LvBNRDCQzrNj7cPmdz4bDQDLOCCj9pvru6Bezgar2FjPzqKtt53crcJjJafQsK4vV5M6Lq6MYks4
oQOIyznu5yQbG5NzbdBOfb1ps9PmtfyPoDzLrLdguc2km3ZQXuIkVetBrBLo5bbL4vBaWtTnJ3zX
OBwWhdxnHMIcm/RwXTNseE9oTTBAjJbp/yP5rjzZLR2rpKE9ZbQu0L5aLAS52FiqhBGUz2a9pJu7
Ma/dK2+/9D/XxYlVsQUdUQ6p77rNziAoi8Dk5hzx9PB0Yn5ZSvpAJz460KaqZFgyVyH8TWDBfA1d
FHK745iYp0maqiTHDtiPfAE1mG5sm35gTEIpiPmaB6qAUlEV4bok1GwNjG1gvrGeNkiLyVyX2O0/
dAm0ayzQN7ixSzA2brCFomgDHW5llfIAVyWx+g8X9KsZOKWXYWCEY3uvWMqdvcSnqtwd4F/TS9zV
Ll/LxBZospefi3pLkjTCqvGlQQ6YAPuxJGIvgETAgYX4TyFjY1z7Wbycca9q1XACTH5YRgNWIUTe
J4uMDtEW3zb4f3FDW158T17vqThnKinHA8ezmQel+y9IXgAwrKRDPugAsFrQ9BEUzKBzq7cSQvDu
rJoR6D6nldLBF9JEYMXGD7LInlnAYqNQFTJtt6vqOl/6GSG5tB1qDCSewcc+6m78Wh2Tz+j5EbaY
a23CEmZRC8qDf9RmkT6SFxiAO9aPqDhsBJCZcIUyAoyjvFtOAly6mO+jFIJij3w1r4M2TbB60rP/
KxhrWGBkUgveSi4RcXU5VDCSkZ3vwk4YZVN6/NUySCRvPGaJUVOCu2tz16WUEFbNPIcRQDfuxf3V
UsGn9F7SncvAdaV+9m98xstMiTt3+9DBRhp/B9QW0Y6jsPR7KqN6PXwTGguHo0Ln0UoTzfRoF3e5
j1EdXV++gwe2glSHfkxLtpP6T6JjL/MNgjeyDsgMxQs4dOB8i15xUN20e/6ldjTSGlGoQ2ONcQGd
pt7jiqoiIooPqmuRRC3pGlrBvmGEF3jrZY2EKprSX+McFZQzTwItcrhYojtMt0GzhqIXl9bvzw06
4k6K3pbMjd0bD1z6/SOAqF0zbnbyaa6FCLXBQ3udQhd6AJnnW8MStYvHnrjvB/r0XVS4lLPKNQDf
DqUgfuh9oIoBkSS7IHyf0mmmNJzny3tkSgxS16VVX32AraDahJspopdto7unyn/6ZIKSYmlRIP/T
qlzIi9B9nsWW3K7RZY1iRmwlnDPo0JvkHlDJkcVVFBwXfzI/XPmXRLwB43UBxwXe49xDqeTm9RRQ
SrRw4HJKwQOrzTyi5cOY4fNnm8M+aXa0S3qaXNytmDEiwSGNblqW96jmNs85EejR9HRuA3LCqj9F
5Ig2qPKXCdxllps3O5gl0r9qwF4ECAxpKM7fMl8Hlx83FqSjaaLzx1BveHbnpXYZ353HU/JS431c
jXsmZRu5pHJzIDbdnyKEraRtnFt5ibtARjtsJaEO9u028bss9CO4+//nTuCyWE88K+VI6uW7Iawl
3nFPwUNt7yHQgYUXC3ZM09+0+xGWj2hpnNVimeHnRE1nT+ut1ECdcihQrSqFMsuI8ylrisp9q3FH
aOqa90KiSxnYekNRW1BRTPbQ4xKtsO49peFJ+8ZiDmUCA5MUivP07zJ4dAvKGHAm3dGSspxSOitW
djPvXxj5sftCDiOOz+fKk94L4FQcqwtyFV6CkXc01l/Krg3ZCIO8nP8Nr8Wd6EZdjz2DFrcyxb+J
EaZ9SyhCni+CPxoAp1KYce4OxxHovAHplhMFETZkd+8MCTuA8/Vkyv49EQRkIp5hsND60HiQq15n
zRWeHFUdMYdNsTKDPTC9UDoQqzaMdyhAEriyWU1eSK1dN2RG9pdw8hs7QZenMGwkGRXj6bUmntxx
uz4UB9K27FNUQMPeE5nahSUBrIzh2PVZv38D+mP/aUgp416Ke49PbIzfMUMnIVo1F/p10/JNGal2
g/7yeWYBv0d6taIaBFRBtTbNwyd1oHuMT7als22R4nl3CK+u8JvFqXpGJRV0dhlg83kEdu3cBTwA
qCd3xDQ72sBl00jDz1DFdn01+flBkFUXhxHQekqygFOrcAVnJjIyTNUumzp/zbk8OGw4qLSvXEXs
gMomRjE28YxSJ9BFuqPpgj+kh8LoyD3d5Er3D6zLySDA3S3yv0GbEiMERTt1lQTWrtXdhIM/HOAt
+Aq4+AqIqHrwhP85a4lStrAHG2GJAh1s/JXNf2/j3E4/DGGu6SgNzxtgO6V2Yx523FgtVa9D9MWb
n1CfoAeGvQp2j+VUSQ9dmL6lxML8cgxA6B1+EKRxd4qPCiqwDLk11wjZgGGMrpvUN3Z3Frmdv7N0
u0Ay8HNr2yPkCfCUDy4bEitLKHAaFY64jwA+E54CVR3xfBJ7rQPb0z8KnrHdPL9dpb5zGIxFGceI
RNBAvCnNNYdt2iCztx1psJ68ibwphQI8LRLnu/ddwg0AlTAPQuNCGHz7/mhvE0V93w7f1TdzUKms
mI4Knfwqv9Nnbs3ehoPvzcxwEM4YoWPwfBDQKLT3veSFYA3c+vMrjwH6fkjC0Sbux0CEtTekzQo3
OH5OekvvykLdGVCsC+LPkY+cMqCe1uWHfp4zemnonDGl0NEnbZt+K93cJO+FTiRIaa+I1hkt92MZ
7H/ALYZXOvSNirBX0kcXmVvy+JRcbh/9r00Fymca7bgYYTMjiGtnUrJx0Ibav/B/s+hMzAr9u4m5
qfFA4CvYeKfiajmVtY1pdf/oOPjJSVu7U5Uffv7GHmvX7g64cjI68uwYRuJ/FCxTzDYbM45DkEbh
kosx5o4l/5UPXSCtWvJuHnbWyLyXbWO8/Oy7aXckzq03V+BGHyNUG669t5c+6Gz07j+CfVZhPrL8
drdi68Jp2/eyrdGpIuj1Re0IKIFSTQhUjJT1PzzQ+MW6SRdHErMfVmQgyLyjvKsDx+LYMcAPojHm
CIsPn4RCzJOwNmiD5gtTXkZx7TwcrbqxzfPbUjTgNPEPCkxw1v7hU8/B2Bv8DDLeDZrPVFmCq/BD
vy9vvDOagm25gFl40T3f7xEo1tSgBl5GyRX57Hj53Hmdk+OAEZECqk2EbJMei1UggTeFFOvYPEQS
Vs8xe9speA8pFRBwWRHFse3JTfPIqVKzo948u+G8r6jvrzzcm0DrAFrRjXayrD46BkoS0HZbJW5r
3pK0YWsSIqYJhQWPvSLtqBPl5iYa4jcyagjcCahUToLC0mN2nEffcctibjTD1YyNsFo9nrD+CJZC
5mnZh0S1bUTwKP4lS+8W7wNEitpqTlzk8Q4t+r4aCw5zEHF7j+aPiMkqsRKo723/YhdCdRhl1/i9
SmEcudFrQ0Zs8zjwbcfuZNVoPqOzr4Eb7lZ4vRhbKsTyL5JTcQlVxmAlqaud3HJBoWBfzAEdswbR
jaXL4CmhvwfhSWTy1Am9qSTDcs2otcDUgoUQf0FxxYFZcKI6c5kDb6H6GmNbwqnTcBNaYX0Uqchf
/9So6Lk3d9PoHKVpY1wcBRdFJ8H9JE28APFaT/GmFklMDIm5qLVk+xtDWoYpsBwJ09crtaN6zy/S
DPdWK9jMgjbUXKMQQ8dEcs5aiy4afvE2VSLLkppphzB6kCcE3fQ00JsmrfIQAmUgEQPerBNLyvMA
0y9/y2JtSq5iLmePg+Yd+Vwp5VDgdJoy6KJMfPPaowqD34ucq60wuXYTNS3sAUEPZjuMbhbHH9EI
rd66/8nk8Tj4xafwIS1bXbzPgqR5FYt5UghlFcEMOYaku4HIjwzUuYsXbupTYP7TYddcCzyNSFej
C9oD6ilYsjyJ9TO3WbyKsNIWp/W+14wKSOFPJh9tvBIE8qZ4oU2QfSkfPgLWRe0Nh5MGo3ZhfcMw
DW0V+7gFbPB+jwAvb/J00m2WNWM5NBzun0uFBSjk9FxNsRiLAx7g8tFZs4pddbVjpDAaHTsKRSGB
OfUZ7/1EkFs/S73sdz7Lj9YGku1RWJkqLQ03N/veSs33N38mmTsoWwUhWw09Vev3OsUmLaNuJb39
5ac2aX3ynpdBMhrM+mnV186YvEkQcK+p+BHH6rlw6VtalqeVaAq2DFb7Pga5xXVyZpR2o6+i66ff
VbcJQIYn8qL//n+npM0SuQRT4xr0dRoazecFVLcbjnLTTbILB/S1zgyMpmsmMTvDUH41qC9pW0h3
boShSQpj9n+SBgSzliVZDMFAT7keWGYqzBCKUPYQsRDAEGSNiCUpBxfNVmOOthix40ZZwZe2MtS2
WVT8kRVNckQwbtj6CctoZt2/pM++LmVb1wcVD4/10chTZfY3rLt0ENtBZqFi96jHlyu2wdr/t7yR
+7XlcmjoykZEQpo+45kVZ+Jusxxb+PJD93K6J2NDIj8qQjuMaF2p843LXwkvtGo+5ydtunEBieng
AdKJI8BaLSMJCynvrnj/AX6Pve7U3656n0LU2UOWrrqCAm73BlG7kG9CjPoaPI1iuJG41tuUuPoi
th/vtAhQ7sMcgnZbleiadN7OmWTBf4978HjusAKTiv5XSJaO4QdIeXW7j3YGJdx8vQA4l25i1xCh
XFGgYUlHuH8cmzz+SP2y17ZIT7wvkV5RBmYoi6ulipGKAKEUJ29pRAUYzCmsWgU9m+ZF3gbUhmPO
0ClaFP1cOj3CT6ntrq4g/aj1eaqDsUQdBCA/hAGs8JqfqCKZBjHztqKKOY5eSbJJPqiDtiw683yC
5m4I7XYo+sQTioISf5/s08sz4OfUMTEcoDIkmbEf7nhYzFYfhLsHmi/daFeE85wXBNuasyXM58Ta
Fxy3NPAVxUK1d3v6+04YeXD71vNbH9Z/ozGz/P5P3A0yEmCjRiRH5kCg5IFlmSXlVoVrtwJ4s+PK
acdcdDCB0lAdy/zUCiq+cqhScjsVCA9IiF96pZdmI04c+rbMA5nVYujcmNDGOZ+mfRM2oY/RKJae
BaKW+oXeWG8WaeHLoxJUXAT+LChzgoiERkKNCD3v59E2PNV84oNnXCfUYxAKjBJ4aQg7JkUaELkI
XB67xTpSK+IH0deTrmRISXX9s0QesyU8BvL1NLIG3Dg1jI2gFYN4Sw7/mB6U/tX/wE6xSMh7V6PZ
8kPJcJNtKKzdBGH81G6jCZ56Bv3FKS+jWydI/lvKFsWDDKHV633kTpCRTsdW74xyN9ywDmOseYVq
g1ScuqF5+rPTv+QYGnHialFMksnuFebb8avrnR/Ftnv9ub56aYLEmD7O1gDoxwT/e9EC+ry+wpp/
Mqx7dnfxm2+h0s71mA1AoBhWR7f5FEGDdKr0NpWyvezT61/cnVgejMMALkDL2TZ1RmFbo9bPRy0i
JacE3zwGe0dKXjlLuIRaozvNpUalzNal4Hi6KcJsTrO9pz4Q9nOvZi6FWlOQm3gjUtgjDmWm/lkZ
W+CSx2l35NgdlzDl0dc6Km58zKThV3gydPT7aizfeWG93tnE3d8at+WjXJU57tyIY7HNOw0pMFA7
6KhDXPfWp6KpsJpO+F+bJLXtqIV7efdlOI0dDXqdzQvlPxde/ELnrJ48Nwmpji3t5ZrXweBN6MM6
7vRxGqqF9g29PGfrobcj5ZeIUpV85eu4ImJJ9rj6Vj1e5R/fpM9fOF8lnF3+naoaA+e6qmZl6lF9
VW3r4fk5vmkt4HJyOYH5LjtgkCJVAxS9e9HCP++8fOD9HVFoWnWT0C52FkBiRmCAqWQBoH0gYUqz
TWVcsWgfHFfeOH+Cb8L4zHmwFRmkQV5wdgt+b+UzcfizeuHZe3MZzJ44ObNJhp0sEqe+GgU+B4vx
kX8RCBPL/AMXlk0o+trMB3jFj2eHbqinHTyErWi5zsJrz1lMONWA7iFqELRjCuXIvRgoC0Luy67w
PYQub5DYP6PGNxFmfh67g1NMS7XVOK3R9r298SIYn6LoFshVUXVQDd2k+MUka4oIW3xinGvIC8Mg
n9RDpNffrLkthZNjhGKKijO7Z9W/ay7CaP+I/ApOtPR6CleJj5V/qQkI18jNXn6qV0IreYLFKgPU
m2LiHzLDuuEP8PtMybIETIBMCliXHImkSP/2mhRdsNzZXsoKTgfwQWqCA1vbdmFV5GpTziFI4s49
P+S8ORH5JfwcMM+JgO6ud3LC2Dsu7A42D/EgkjfyzYJONtUQFYvcYLUAh17Tiqz27CiLOBzCr9gs
deW9Xqv/rZdg93IQu8kKrR6NJTvGC0zeh+FOQcFhwnKfYusETEqDR3F6LsVA16uLBjeF9g64N93G
h0MP/oKROYeJVWWwyWUXqeh42yOmf8s7bPzsOmjCAQP5QNCyPmAP+b8h6m8eanp8XT5J+FGHPTst
U3OAOtzk7UTqYCQ+LPBFwgYFIMD4GzI5AilQIv1QSwctERdGHJzU792epbjvUjFuWwXUvpGPfawx
Ufd+4SG7gpb/37lpfLDBCgVzMyOpSc5LWrla0J7bDBPlMYiJOqTkQZ9inOIWnVIA8AbTE+89+C6n
sqQvxFGyxzH/f4fHtdXaO7yhk1k+QdL4HQQrwiy2fWg3uTQKiBEp7+fBaGMhrL2Rs+sduwsQNU/U
YG3PlVg3T08VCx5PAJbzrb/UViA2T+wgPcB9gWKS7XvGVWtOV9cB6NRrunqZNp0f3S0ik48gPSqc
NYUSlxhx6uFZn2+BoU0xNe5jM5f3M0xkWdhXf02fgdRqRQbgpWwNWJ8M92Vo+LIIgNnrp+A6enja
2NvSvxbnNHNAohngGoR0b6HVAbf3WkqGGlJNlG5uPTrtpmp5Ml2j1RLv4hj01HUmpzTVSqaIiylT
FIww6CDXidZgRF8gfgpxXSvRucu265NqI/ZUUVTcqTKWLGmw97LVc/U/LIa9Bj/loP9grVwr5oIO
EGZkaEURsaq56seKQ91DIp/o+wdptVQQo+21zIs/UYUddETKSFto0SJVXNOs5bnKrJbCLvbhMQRL
F+RmM48vBnpb3Y6uGwVERJqYPx8KlLS6Acm/TIFHtM4UuQVez+kzJVylFdq24weeSWhGUPKHmr7f
oPr0dYXrDY5BQikv6Rao/V/frs1v1IOsJEyHUGNcvXZgDWpcZwnSvy5XrVKQyFnSjqZQSC5fpYHR
qIJwI+fosVTQaEvoDuGyvZWvO7o5m3TOEV2sLuI5a7igtGRpHC+GlOffBQKO4jT086zDGivlytWe
2bFKAanjUjk1H/OGscg+HiBrOf+JQyUSZ+KlrGsEV5Qb6QiOrcAGi2ZKwf+MDoe20tABkEn6rTI6
0ZUi9zdEbqRqcQVneulmz+TTAs5ohfpVvvupVw0CeGCu3raCeoXRN6O17oE/2xsK2sJefaJXYf2r
nypr+J6D4mtVSNIl4DMLWJ2QoN/OzAQ9hxT0hz73CSjgJVuMSyW217womoj5ZTdJfYPM9DgEB+wl
sgzk4UIyPyD9jHpK+Lfzhw5nl0Lm3hpNpvwTSq92z7CD99sjzKgANchiYn3TApYLeESnwDWdf4Vy
GYNQzLNwkjA0UChaNp0prsMactL5bYq1bqq3E/OkzHL9fPOpu9Cy7TOaFGrxuylh6Xvy2QZYBEDy
ktGIC8v2PupA2w31zPSTriCaLJ/QEZgBqWTnxmDVmZKuuomz2ZeaC2ZdFCePi9pEH1JHQmxo7Tzd
eTwwwyQ61i3/GWM55El3CQN3CK2TT1a+RVtK+IQf30/aamtP/Y0IER71lgLhlG218KXxDUEM+RBH
qZl+1aur42F90tXsb1GG7FJlUdW+Wnj3zv6ny20KwaUcwi9t2yVMmqYRFa3+cswCZKmH6xYUsvXP
FoalLYarrx1QSN4DfNRFe53Hr3jbKr0VyMxcrjvtZQ6S5ae3Nsy0odTDAsgAYyCz0Xr0xWODR24S
HmlQOtNanee0FT43eB4g3XZwzfn6x/Tdot8MMI6Yi42NWFHdpQkkTokH3M05NOLtTkL7HvHLsoem
90bG99QX2MLMwG2aGZsuhlBw9mFy0iZLVFkA24UHfF/hH8pKxPjI83GOCNp7XdmOlWNr3mDNdnk4
Jv8kEmLU0ofV41HzfTiNx32EjgurDsuTShujeQbA/OoMvAy0MX4Zv/i8a2VB+j6AautcCYeOWwiF
iyOgcVW0PlhRZRcgkXJycdP4Uf6q24Q7ZRG4yBYKajD/LkcA3aeIyrtlV1Iul1xkNyFnKOjhKf7R
wXDb2oi5RHsflZ6QuOIZj9eBU3EZOLpfxpXjJ8Y2NIvLAU1XQBtkxHyeUEDqhBjFwaSppx6Hzrac
b39xEF2vKhcYR1DLexBXp0GUuZmq6CryhpIeb2vhFGYuKveS5eyPoFUV/YnZ5YNL41T0RlaCLehp
m8n7gP2VPxp8P/Otz7a8WR5czJpnEybKXSAdq/l2RPhqPnb4V0ccvtNjUTF4PaCVzjl50vTxYbwQ
3sUffDNF1hLkyZ+wOOXvsEKtIjxZYEkmHDXUfeO/yqOhhOylQfXOVrfiMIJlKjZaejUmUVepWaaj
G8DzbOWyHx7EOjn/6wAQrsB0Jtd7Yed4yzBcSjo5LbRUiO+eqeAMwOLOaDLNXoGrni2TJWEkvITP
WJZVc1Q8oVuIa87xdfN7n24Wv1h88qnQUs/nMTu7LALSy9DyWEcg9SDlopDQ6WMDRPtwBUTqPoHo
ZTNiYMh82GR9OdldEX48cTDefiUjbDLmXjKh2ijN9DkvhJcTDcNwaA1chj7oOFbUfNO2AUvsgum3
kPJdI44r0az7Ghmx7VYpR5uMjaxqyJ6LC55BlSKv5Lqj/Hvbv6HiQMXCWN8fLQ3We6X/DNPP2iCI
5r0yI5gW16YujuUpE9U7qYnO27WJJlTBnAfErEjly2ksE4OlYCQZobuN5mgSjt1wX9iBsz8spux2
HK5RxMDx/FzQ/x+F92ihv74AF5LY175OF7Zt9YfsxDs+BjrYQZ3vkb+xBFzJEG0ABAeRsSCissHs
1U7VVph5ckSeTw4kqFLqSPjNDuz8jPr6tBXaitmqD0e1Z7hNSRJQl/U1/py8T69zO83h/mmnz/vt
WfCwqj0cM/KA7aHiUFBjUmbcK5LhB42YCQzLIVxS4xQ1tt2xT7EHh7AX/3HoN8nJOUOgeQDiZAao
KbVU1QneQvOY5CsU+2oMxUI0tDhQ7MDNnfiIKO9MYiN2bI8glD5coA86NxO4m2f7HaFgGV9EYpYa
iGHF1Afyg7fmsrQk1CNhAXGCOmzj44tueKsY8UfWydV8l/KJwy7ViTc8D+13iKFwj9y+KdOW0URx
IPQyMnZ5yQC4CrIOnjvzLjMtPtnu4+3AirpoXgEhVKECM6lHrjgRxA4Vu1CUDTtQDS6NqyZZnvhd
vi3X4ktMBMswU6dOOKwgqWILe4RGeKDVALB2PHDTa04kWeBFdnYIVDbiLvNsFTN6n+RnFb+YoEJr
hH+JFCARBGQfw6pZVdc17GcqOzoUS8JFJGssdw+4CCSoYG92mT21RQA1YXAjx5YtCh1gD/aC7VTw
yyBiBQ6NU2qDBeFUxiG57XEBobbbdiiSasR9VFjiDIINPtae55xlrx4KCuNjRkrlLTsFT7rzh8be
qkwBtfQe/p9e032wW9fWhQjGq4ckwcM9BFjz55DVJZby2hruzJ1ewH0cB/XXEEApUmCVDTqss+pb
DKVKtKmYDS4APpZUh6HwuhM14+EHeDcuLSatyaQOqO+eza4oad2tPPZlOtkWmBTuv5KAy/MQMYje
2b6EWhOz/UJ9EcrC9ezDHpeK2wOvgxSkZOfq50DyDC0XrXlwesmAij6AlTDsFwQ3mxxXaH8ovHia
JG1h+2OE8vLOJS3qNokbCDMByLDRgO9gG1tf5Ox/7pHKN7aEVojTtGADXG1Z0IsGjOhn5ian3yJz
QLefphR03axMo7mGw9B0mvqm7O2Ah1B1LK0IiUgOTHPwfX8qb+xUQ9KamPohGCoP264pqkuzatQb
CP6JkF+RoqeZZtFsBxYLLhfjnAi66C+5bA/phSWR31dNwd/cwZr+GwVILvXdKufgLzl3rW3I8t0J
dHgmg7ACmCweIXvrsGIN2cDcKLME9LtCFqDX4N8WQvlBwzOUyZ5fQzRlnzYeHEKR7qLVgUx08G0j
u2Guve8j3XoHA1w1kz1t6wnv1du1sK2l2UER+D0T2/F8lHXLaUpotBXEHJ8Nlghov4g7Qb6T5hd+
Va0f6DV8Xyyjl8pGPhsoH5ExVwgkCdL5eKKVoYNCDuKNVd6dLpQMIoPfO4XcKnHJ2Mjsecbp9O+5
XLGEVHZSCbvNG7DM4cFbp9f52K7lEme25LMbQq8nyn0qKZN3mYr13bhDNQ6NqDP5RbUB4ItndY1r
rqjuewAVXFKuB2MvEx86hvuo2Dp03VPF91g2hwW4oWFP+epunwTEWj3ZvQjnw5MJj6CzI5MSaX/Y
YuG2y28cfnHwfq5f048botNnEMEOKyWIyOuq6a8zOAXssELIRYav+1oWVoJ575jvC+4ZCR4SleBb
LID4osmt1bKQO0PlaA9Bn0rgjRLTKQOtYwtoCbFfqctbbe2q7axAsR5OUWkpAPyZVEEsjNyQ127M
F7EO/8OQ+pD+9I9GSZTtPa4hZrPj3M151sds9qEw22Bs4zKDSDmQbAK2ToblfEzaVjSihsJql0wM
B5BI0DX/AfuK4BQyRurlwwYl9fbicPIWryOoRBCb6CYU1AYArvRoXD/B+7aJu3cqAN9/6Ic8fWkj
yBOUtVOh616BVMC2F3PXhWFZtKNXIVoeur9RidUE/0dJcOv4EyclZ2om8GZ2I2vpMuv539078vSq
2ZJycuUSuc5C1ilD8Gh3QyY2QgWxNIa+tZ4T8atHP3HT9XnNYopCgQScg5Za2C5EoZVJWVIIdKpU
ws1cFJg21/vVga8AjKOZnlyfjZrZUrGwRBqV61NCiM3MpM8MrG7x9nr/3gRcXJTkX1P3ab+A/piR
f84tn22SfPHoOadK6ksRmS/d/4VAMjcftftz/iReEc9G+mm6z04ijC1psXo3H/ICxxqFicB58Aow
q5NBLZT4fg5ozD+aOh3f8FtscxEpNCJGH7ZUqIDo60a16iFRnttSXqmD3wOzCUkmJrNbnPMspbZ/
Isj3UVxvyxael7AIhVdYUu3kOCfJKoodpCqXsV0Rc+8rw7euEcExnq6KEREl/+epn0KAeLwX82TV
d7m7Zd+zqfMwNIxy+nt4ewGrDyRp2Tf7pnysRqqLx67OnB43h2X+hxMJWyRumHScIdiImPqM2BTQ
CWDj4VqviaznJVHH4sq8s4/YhE0Z7ZVjz2RbpehHzQ+43/X833aPPQiQPrcU2bQRUPxPFMAMDCnN
0cAYwSw7Iv8VEtM4EN+WX9V5Ugmv4I4xJk0q8HPFazyPFO0GCpnKKletx0dz1ZrbJJi40m7KF2Mx
pu6N2ZfcdX1PCYrX0dsK276Wahdhi2VOrnP2XRMYpMopMLhLgPGqAuheFR4Qs0eLYaeFpWEorvYz
aJSPsEgjTgLapXqBsoEIA0Vh9GWVpvoiWYHecpf6uNPNxrbmPbZWTUAQSs/gx/HE02Pur9RlK01f
zrKomfLSl91ynVnKi9G7IDRPpg33Io1s99doxq0FY/HQ8Q6ktz71NK4qh9yE/m/6uyK+znDJ8I4+
B6mz1SNo3nJGto76sgCzQlaQESjzL9WhlpJgFwZB+It29X0YCr/i8MTydAA1cEhnfdzzjCWfr4hD
hiwoLpSjPETl9ATkX7kP4+inSS7C8vjCkUfdIwHv0VdYQnllEMVlTP9w+9zNtZTkk5oKVxK0R6al
MVRkXuDRpMTQ/sVHOPhHssxvVx7s35vCPj/OCXYrSQ4Vw+NTTB8oFVMiEl+oTIamqZHcUhoPNG4H
weRx/Tqu278MdwfwsIAxXNf6X8W4g1gjB0hjA925auI+qEjFw5D+IaN3nf1UGQD47oIjOY/hTJsJ
wocK2DeEHaOw8gTRI4449bX2ZcMnAS1hPVs1WGMZ3VVldEdlGvWtIsL9cQLJUiJQPYa8LIiX6OCR
abhBDnDGa9wSfUIza1uZpCmwlCVN8Q/zOEFPhb0Ek9OwvkQWemxTbKnsHrEjksPuf88W7aGtBzf7
vz1KviF/2ZU3ctya/3juGdV8TT+d0CqHVOes7lJ/xUKVOwudB3YOgZsSsjgilyGfbwfWW/1elHT4
iCXZjJwzD7akpARaJEL203dktcG0I/I2dvxPOSlVfwWzVvVlWQXl5rOUspZXiAwzWjfL68xbgyiP
3EDYEQM6KbvMEr9S/fw6pAhLcQfPpztCZc/uA4nKe8IUWg2TTIfWN82SflbU+USguUhAa+lz/ujq
ZjXg2wc/BEGkccn83//S0oi6iW3VemGe6ER08H+5bCmatSRN5/QbVkE2BDlVT2uq4jtTlHYDbeKT
cOtuU2e+OYjUPCzizJiDdKbzzVvuIrWjr7pGnoR0iOLkxFMOMmoiAP3PK0paYrYLIs9oLU1ebUje
eSy2ktEAPRdQ2RNVeUJMzvWkxOwIHXhmh9gxNO6cmVRWFLBdjsKbV+8mwpgVlDNDUy7UzB/mapN3
m8WiUZzYnqtz6QJoLzAvOu4H56T4ufds1DN7X5OY7v7bYF/RXM+7fYGIsxd8gFoulHt0FYgU279Z
AFGhDoEybzPTqUf1hO+tPz4cyjs++5KKd30AAOnR94NUMJhD9uGTbszYCtG3z8+63BMamdoBW4es
x3uOhabfPnGNhs8RWvGjceJpGAYp9+b1UxAYrbClA5v6GKA83xZZS2nEVAKIAajuvlh2R8jiRPCm
5zpbKa9eCDj8NeJ4bBAtk2Y5N3g5n10qgjEpqbytWfyTU67rJfir/mj23tercDWkvz3ErAdR98FT
zuA0+KAbcOHIcqWsy2SIOWcLsS9T9jNGu29/HaM64hiNApMtqRxc+B6yqvnjGPiNJ2kdAr0BSvWV
UhI5ejkincxJ++RqG2e1O16wdN82Jtk24q09Y3vHLvDA7+8WLoxsNDafsnF5v2VGz1Qjjxsove3n
SMibXWDU7BPvQ9NFFAzzdnCmOH9ZXOtJgLnSGqmkw94t5G3fCkKJyRcPT7oMyoxsB6ZDIDCC4+PX
SCX4EQ6hqaReXEY1HUVNdq+DKPMjVaaK45ugSOXUH9rYY5jkZw211Mgs8q1YR3/hKFlbvezaijxS
+d/q2Les2QCj9Nc++SvG8pi5oJqEAFqYXsgQeTgtQjeluTiVLFHY7wrcfL7avNrosklSoctS30e3
efO5vs2HfhntL2cj4kJ/g3mFkvmTzfwFOO3Mj76fR2N+McB0+emd7uJdx0brMGZoCZMBuBDuphn3
Agl1qxHZYCv/uf8QoVVADRG8JfIUUgqDzBoeVjq+0vjIyfmMGOe0M0grbOJCAa2WKak35eJvyK1P
Fw/ohZSKyzfblIFQ6/jvZtXGO248b/C0382D8MtgZkULieN+PZ1rrqcCo93PXbcSd1JqI32N5iKw
1CwNKqWQrD7h9uKfVhHkoIl7ETg1mKDsMS8DL1QPyYxdFavtUf3DwNP0BOeFXtZIGLp8XGgGOCKP
6vZtNB37YrlT2i0vwWTAKaX/LL0+Csj4N9JQGmGitrm5T/nI7Ib95gZRjyGOR7EJ4C9qopPm/PvC
I9q0rDL5D5ZMxpSohqHTrxuBNUEZtxm09gXVHPUV/tkkzJ517Cp0IVbngpsLeNUVbLeEG98PHT7c
BDOjUql5rL4CCLbMVdLPJsrpFEIVYywl/6/MszR140GA9pLCfE3JYZkkXgrVNmiCwHo9LA8jBF+T
lTYWrNE+GhVgMtwLGImubYBHcEpRlurFrOHJ5pK1wq5bg910jWl8Xvzzbje1oPaEgk1AxVVYRNrr
eREJSjRqI3k28pmuwJZqWdDTOpGloEqCrQRly2ASvVl7iTufCMIrA1adGaUSXpzAvKvwFRpQjmdd
5skz9+0YgzzAgJRS8yaYymHiFvkdGeLzj68qyOyFU6e73mT2/qBJ84vDOFLpV3ZOmMok2MrzwNud
6gCbzXsnKr0uaBAktQM5cGyHxqSIWe7rJ/+qGcVZMP7zxrnb8LVQjDg5wlRagLWksFlOEfN1u0VE
LzzDdGo67nhindo+WiKxDI8L9+5YZcoAwT3E+tqegQc7E6dB0rSbG0BOzB0OLgyYqpv1Wr+Vhp7S
nAAGsFYu1PAtt9y/+vsBASAE9PG+GYXvxl2EdTRlAdWxjAO+El6j8S2kQJMgs49FplX3LIRYJQDt
Y6L0x93R17okFUcfeeTi6Om6Mkm3GonGtADHuPgcjVfLGsw1TKdBZBxh8GqrkCIWsBrbaTNK37z7
ilMTaxyKhHprNehbr/ZmsQmcrgI5/vU7MUJYrQUwgXl/o/vM5V1SwFA3favYRM3GXeGDOBmxKaMd
RKGD44DWROVsnG0PAux+RpS6+svVodd2nAhx2TQF/ghQx86hgfs3W710BTYdcptYYp2P2QpVq4PU
hGpzqNYjEWUQXumzHvD92GTQvcHhAfyqZQkICgVIDTk5Sb/SDpwiWSRBCa5gotlj8r7DmVz8mmm+
WcU4YxwhXK07U2ZpIm12jRvGfSREnAqyr/LZ9wVG+vK4/KTFY+jyy4c11kOzjIhrST/syHm5XIG3
VmpBi385NFoj+DeY2qz3DK3Rk088QKxLQT/sjVhJIIL2j79cYlc5gUH5AishiZ6UQZfmzMMx576I
yVjKjz3Wj3txtL7MYm+73r3lKxEWSTcLEQ2c+x00q1dZ3hVceb4Sv2ywtU+ZRKbU07eRlJylCB+O
xQHAZuH0c1QqhRstbKhI70haa4YCiV80EgA8d2Co73YUAzd2XCOEcFI75s/gm2bZA4WhfRez4v+Z
l1R8soHQftBXEHwItWBblvbpxTcRFjRJAUZC85LMT/w9vq68RvvCM0Pv4RLKFAuN7zzGdAKU5gVc
ky2WfoCkFiUO1krgN57XyoeVkV9ZwLXkCug2nxfalS5XThOKI/b5SrP8lamvyXWVzytz15xgufE0
e85z8O/9PFPpu42s8lwQwLM5u0e3vj5tFk3TVuQ1BVAN404kr8aXRaGdJIsVqaqLTmX4SYQMFHNK
sabxz8YuOHKs75SsxyylzAjBC9QBjO0OpFYUsVWozWe/p4h7HAIaXeUqyykaHW39nV/ECBxPKWia
7AgOk+AzNx6pGJOLWZuPuQsD09YCIdw0JIh0Wx98N3ClHis+NSPqzePLcLgDdqUrDPAA3JaIkqF1
McdzIhL4bN4VJsbE9MPzhzNdfMq39DD7sXiij3ljkjb1pZRTfY8rRFQTXCgfaDXwGD3M5aRNs98a
0TjYhXgfK9hcbmLZ9iwIeANMNXhR9iW6EGy/zmV57lnS8f3Lcfd1dzbMz77bxVlkOufFxKdp3UGd
KuhP2h7uVvT6cc2/3ZXwTQI0imXxxpwQtEFJiPh71GDTh+Ri0VvGkKKXuxMrSn2laG3ObhVOj3cA
RSldWJo0AhH4oBWl76yTCIY01LXdQNxVukWRKYE9/yWRe2/7vsqgnDsFwePAPY5Ou19Q+K6w+ht5
ucnNIE85QI1pBZgXv35XjSJ6srYKT2leYBT0oH1iltOjQisHxEg3hgpY41L3u4R7iIdbIWhf4GV/
TQfCH28BcEL81J5XR5abXbjsPcm5rP/L+OsvzGE8wfslmqjc68qYJI9CVDHchJvjZKinYDxEjzXY
SLJv9qw27zmEUFRAcudDgPcJSZMbCBQsfYay5xuw7tN/8QfvWxHScX6Y9Hb9vKS+w5N8mih1WQgT
AOGuV2tgT0J5WbfSMrM27IS5jZLuP/nklwd7sKGjpTZL6K+CV6BhHteM5IpSeRh2EZ6QwtEz8fl8
OHn7K27e0hVnwAkmPXS2HiIeLbftH0/NswmIQmjkpOPzG14yUKqVvUwxBEhFOMX9LCwwFZE62CDf
UXNC5QKWrALYamGL2l/i749ZujXi28i6xXLHgdgUTuoEf+0qGcvsTst5ik4wzRyuM387t+rIMr1Q
vMlRioQ5jlKLRF7dz5AZfM3fTaYnnYobO+aildr90kROOnepIK/5JT7kdCZupGDZ00bqOaFLgNhq
EPGPOuwNhAQEcN7k1vR7YWMl5e+SN+MnM9f5tUO+2W7bm+hsTqSRLFVpN8wA9gYOQVhMggHj1dwK
eKJQzma1ZrnBCZ7o3InlkX9iizwQI5vPuFOERMzj6wRa8gFUCapK+gMWtM68w56vA/x0aMyC2Gh1
uCvEsTm8ifDQObaRtv4KP7XVxEK48N1cB0OML+6pY6Sk80qxnBSrIab9WRxFARsRc6ier9lkryFN
4CTpY2Ef0SDO4CFJ2Y+TDCkbrGhBYxbXKyE6hFlKwz+9lE4vnqKrrSbcqHP4vf8DVYKmiP3B1ks1
wds39fyWiy0kp9wSXbLxi8YQQlXWn2wfcL1H6DQ2I5C6t37nsL8CX+NeAKsZt/wuzVtzg1GOVW26
PFbNkFeddl680zvk31CejxFvbENBgfRD0FjG9vlPM9uFCXpY6QNBqBTtwlk8UzuuGYK3+Qy2xHke
mV+zFRFZZziaME6BkS01eJc+CMABA/EDqQtGy2ISsEhFkdEnWXokbxNj8oihSlo1NepjTiP63c3g
RidmJoAj8sTUWLcQQk0XoCAeYDjIO12YYvUOq3lTlBX3lEmjula6VZHbFx0JkzO1hSnL68tCEIij
vOTjIx0PSNIRoU4kXRL2AYIKBbVjBYZhrZdBKGAbbIruYai9iks065ZGXDYexsPtT+khYDYh+KVw
eRPmzDmgaAeh98Zm/Inhx/LyP4eaNFvBgkgaYt6FBzJsl6kaQu10mkGFnHhC6mTOTuCMn20ffjuZ
DHDKxVkBNEs5KokgFuxYG9OVR2LYN/imPNE5YVfDsN0SeJolYbHYPJlyC/ZVF6ecweeuP2GKIQ23
pep/1bojl3KO/9UnW9xDS7WzDzzZutmg4CsSz5FBfYL9FMd949G3t6/nK+OMkbnBskdI68YH+kKz
eP0TGRcSfXSfg4mc+8SpgtR1jwzYWwSwlLuhbtcDwJ8IAetd5luNQrU5rUfyczNFeZPLjp2R7jdb
CmWAjPvFrGnrpaIVPc0ViU2+SyiQV1QfWI5fPJ6uQJRdTEf4E0Ynmmte51axPwm3CzODJXGZaafN
YIov0J56hniy1zqByr0eN9sWu7b7WOHsIEg4gRfggMsDiogRjSTLZ+G23xHY+44oLKALL3WXSs9e
zvvnyQy2UkOQesEjxs5kXh/5uPmp/0RcRbqbOOWNdjr/TwCDI1PABmZOrdMudn2mt0nG6IpXzvcw
yF3YuXEC6hNE0xDPauxDJZEH5Us/DCWIk+DlgVkiZpuZuXp53PDt458T4GzkhFtILgFlTQ8DJhfD
FzMsv43e/GUSPOzlsbcNeaPHC6AKq0yi+gGcnfODmNPczsQgNnsgYfR2Sbsqgr1kcO2QBrvrXHb+
FfSRs5JAtMKwx2FRDv625QOhmLWF1y+l3U+x80/qXKRc6Zu2E7ZxQemaUBRo5EajSC9wS4JaRao9
smhm7gI13OWW2Yi58mANnf0gkWVLWOWVrMRIAZfLuNeYTOmAdAasZx6IBdcLOpCNkYYYw2X+zNJM
1GcAxdtBUyn+TeQ3bYzUgn7x7NPROShYg9sg1lmDRjAckUq95JVykUKFsaz3SWdE9HBr3UILBL7h
ei7LxCjGzWcsZFGtPqej4f4qDAWTCyDxJsbMTou0FzGTTONcy2iFg/iWYvpX0Ei506wce5h6Kuor
HUQBMpbJLxEBHO3e0uFSW/QM7HCWhhoiDZKYX2SjFG4FMlpGwh87uYEJSrGVOHka4Il5CH2GstZT
uEwkwE/j8KhqMh39NK8lM19yvZTTVdd1HjeHCbXssAz/VwYbJxIgomAXbVKDL7nzAmviPL2JB3cE
xe/Gm7pcnRUNjJOpNgYZaz0tky5ggvO+2E31zk9cyGFaj3AoC6xZ63i7lEcJH/lDhz720VExYj0Q
9YQAQ3k/tLt+YBwDRt7FWdPIB6S2p9vNp6Y4DECwy6afKNYoPHQRfFMrU3RF5sISbsJD6pgp0Jo5
SVoWBr5a3RUIJLOvpPy1pGvS5xPs2x2x38HAWyKHfh2Xp3AAvpbUUQ/nfyzh8QJXbyJMY2bJBEiJ
ZKvNRjH/hnV/r2ma+3uLTkuGrOnB+/YopTKgLRq99eY5PafctC537SY6ZNV9s0IJ9x0V+4xaGuO2
d32bhUcS41GrQAx6O70cySw/Ly2qRFkDzHorgbsJ2XvUs4T/FhyMMurD5DZz9dLa9TNVDRk1EnZ7
KbR8AXVXa+/vlmq/6YIH67bCxhFI9nB816g9hDtodBEPz1AJuQHN6bHPAgM0jzsU3ST+3McbA7lM
6813wa+DEk2Q3EnQ11/wddPEg7pbUxZe+4HQQeP7hPTf4ypkfTcdMSz+jsDeYW8Yv4kDYIxHlt/N
A7kRuGfLRht5A7T2kjJGBr8tfJfLl5YlAjQIYxOAx/5oc5VhKLoqiYxJbL/kB+dedM8wE7b3ncO7
DjdzoFwxGss6lcmeXeMjgCkiOHqvslpNEasoz/gQ6ekYEHg4mx4JfSZokYK/GHYmD/gNDM9CipSE
r020r4wsBDFY4sJRXlpGwfLVRkQX55KGWQb5qZcXC8ni+MgdAGJX4GjlpA96IPKZUWpgnp/ZukLF
FPOn8ZDv4ygfI6fYJDNZHjCnygllGy+AhCOWLs+s4oXl0Ra4HXaNDHlJsM5czglD//oHOHE9s3Cn
a6GB8W1DpG4Ko8Fm8q7Eid7yXQuEsMsb295xIP14x/rXXP5+nCSfGTqO9NEap8u4G0d1SCjodndh
Q6xVVviCnmu43WPFS1647CRhpfgdZT+o9ZcndfI9zknv5OaGTeT+JiGqHeqG3HuoufS9MIL8RdgX
je13KtxSAuRYPE6xXT+he+SWTcMk6QbBJQOx7VGmwgt8qRnnOiHUINaF8M2HAGpVTOKY1Iz5xGMj
W/q5pxIzMswXD8iNOX/sTaosPmIQ2VWHUZhWX8pYCXDecODkc/TVilcXHj63p31XqGRPV20xdhZv
0cGNHOaLJzawh3D4dJf264u9XEzJJgq2ZRy6x9Ni63aGqlNW36pdqbALtQjYghpbVoA0cvjTwuew
4x7KEndsVLQlernxJZ0mVoBStTrP3eyTqdjI2URi/36n8t1/1LlvsY/ODnhQfl9y5NfPnhAa2fFu
abKaXMJvmQ32D9oBAX/v++OqvpKzyUAFp5JS8xxWAY4VOcZeN+tGBZ/b6yeUVJknuohqPG/1M/8t
ASamBGXbYrh5zWoTF6qjq3XBWZzj4SU+Lc7CPAsUh1iL+XSxL38yIFbeBHPdTbsM9sQuRxTGZjps
wxZBKNvfVRs5urSEJL7k0+4+aPS/l9Bmxau1ys2yjXqjExuhjYIK+AsYXfJF5rU8XIdfEkBxiIHd
mkFzG35Bsy4YCcsohK3bW7N6hDaaScNs8uhmGhBX2p5jRuqSIBPJEZD73nFFOpjTuVl5cB6c7L+z
IdmnwB2ogb4m6cRz5S800XrZwm+13s31roQj0P8zxgGLxmbSNldIVchoCp0jO89rnhEx8Kw4t3Tq
/QIfWcjHCAvqOPMWWG1RD4NpK3ehQa3/09hGKjc9oU2iD7C2H4K61IdXDV5H/8VpMoBk3l1zO2W7
Q4VN2o2TXa608izM9ZH8AckByUt+3befWPTPiVEWAHoTYHbkUh14SlNKQ9ON+4hkWYyNHff7H0cQ
IWg3lr/niAOpfZh9eNe9Q73WOZuVCpiLoVenVSVKCAmdIi/YCImkYXQ+6HPtuGDxqYlKjvgGImPL
TC/RTGkRZnmghOZ6V1UR7+BiyG79SE28m/oGTQudcDNJcLkU4EMoiUP0AJVTLPJXGviHed8y6e2z
3cdqCrb4227Zgtd45pSSET/b63rAmqMu0hOzgZRFgkwQIgiZefBIP3pQxuGjl8qIklIeEkgjWmow
62MB1dAm7gwKHhdEpNj5fPDNQbfphSKs8gYCBEm4Hke6P+7eYrZjKXJT5pQbSUNEQgwnQP7qvSwK
zOM1hWwE5OgwkV1YamBOl5Girii150IZBsqbx9++PG5eCInWp05F3DNIhYlX2AWBWBk7NCuZh18e
bOX214JR4BEA90JktLgsDpWPkKYw/AQnR0ok3dEd8sTLtQRmtWhK46TLdfw41/GHqpi1fLegKkfh
QPzPZc+ZgRtr5VnZM9EOrWqNz5NvfHsXTdvIdPKBaFOLajTbLOJtfR2Ja0LEgeG9+2LIT5Wj/4g0
SugUIElcTjf6OiF3fiveWN387eu9O17bQE7173Im64e3EQVIjpkKkjEDqkyUOgAxM3MlYhQqtkcP
jfiVfPxnNiPLisMWq5BoY31mdXoSlzXS+wFJARju61GXjT3rZiIiw6Hw/aNaeEv2WlL11DthhCvT
3DbTSha9K3bydklFnKBgivCS5p91ndtig2dvxf6JtxH59TCe5loywJena1RcR9f3QS+H+ihklPgX
vm4OCBvwkYVqrRJvHVdaouSXDsPuv0M5/ZrnmZTUk6COpUxb7vnKlrtG0KMsN4uU97xPfprIhv7k
hSObhl7rz6jq4q4bDoZqaaQJr14vaxWU/MJio8aRm1iQ79HdgqjuhT4ABYX52i3BfWN2dokuwlr+
MD6JxWZYtxJjEiRgvYeiLoXkcPxdH/AuZhXHe2+ZenH636ma8yI8xd+0hBvrONX0Soi85Zemi5ij
6R1c4IoGFkywSKLn/j7PAOgHVTFZGlZ+h/HQzdP65v8dV+Llioiu/MM1pneV0+qOCrJjSTOJ7YX3
m1z9pCU02R0o8+DgOX7vJj8WuVOyOvdgrwj1V7vhDRQi2B429holk2M5zEKgDeGIXlnNPQmK1NPP
jCQxk2tnPeQKBY26v9E/dvy/3oArWXF36tzwpOsCtVHIMlVVq+bxOWA7MHNdyZoIwKYdDwTtEB8Y
/oG920JJx8ieV61EytCtz/YKOCSDrCbNaEtJ9YM6a1ZP0Ww3J5Xm4MdueFT31LDXzgwdihQX4p8j
PvFc6H1urpZ98ulfp3CWfa45oD3b2emxTRXi9bl8tWbuEkz12jlH50ZGlHjryFjm7MeBdi5Jr8Hj
PQlaDmogV6lUWtIZbV1ovA8iPG5jhGdtZqQ3DWog/RQl/idiqWykWwVimNNoCo3c5gBAp+cLcDra
27DKPX1ekqvzQKLK4RJIVAK+TUK1Z89kdvpZUnYbSdUNda4t5wFzSyxdfRAY9hdzdjl8m3fby5B6
xFB9FOHxGbv4LwhFaaX0rADYa8sqnurq5TnHM4lh8Vqgrv23zVpBxgWUqPB7u6vhalRLKs6k9wnV
/vXEJQb14tycF+bAs3A2H2/RaqWiekUR56v/C7M/t7T9j9zXN3kjEWv+YoifnCeaIviShGuiSxno
wnU/gGxWu7nZ5fH73jg1PTwb4G+A7z7mdx/KSDKNzG58OQN7jxM8hlXugkQXttilDpLYqbMHrWlH
f7IHi2Ks0gn2bDrieAWG65DTvAlOTcrsQoWEtK9MB/R4stonm+3s4n8GxXqQebTuvropn9IvM1q0
yCuMYn8QC0HsAXaE5SqRlx8Fp/qd5+sTKvo6IyNHPhWpXi8xLG6Bc2HtR3nni5tsTKI/EErm43K8
SdFZDec6dqouS/9EHm+aVIjb0p+KC+i1A8sdX4tbkZNvBzpyzJoK5xJRg1647kEeTFE/tRLz1YXD
9E857eq9gZmIz3jcJCjXCKb6MX2p2eWhGtyuZDVnZPzEcb63hd5vE+rebq8NPodqCKrUfxK6Cjl0
avQLJmt7jCS04z4eBDBE7+kloabKcimIQtEyn5EGWu4tu2wZv1CCzn+O18mkxtmHGGQPMQRH+hbB
CdxthVHPZmOWCSCPrJJgomsK9tQKUqM/v/j8rZiG3T5p2j0F0AaVSmF0U6n8l9ZtbMjjbwz+VD8s
4ORo7eJI3ynBdLtXTZ1upkzkhNMlgLhXjKeR6r+acFXExdUNrcZRt09aJv1T6rAjviuJQLK+u3yJ
OhNL5j+Wt4RxOm11SrkTiRfCx+qgpTroOisEl4bAaJQjXD282plXctsPUFrY+9c65dt4FUbzOHQ6
UvfCRm3cdQS6lBy55/9/ihfH6u7///sBemv6I6dhS1tZlCOO8vlzra9yrghGi9cOmQpG/IjYCKhM
i9HBRh/1DY3gy22kpjk73n99p35m+QHT52AUuj+qk5K1yVjGHjxqSne0GpVL2ZLulSaYJN+qqsJ8
xOPIG9HE2ajYwOrpQLc5IhhJ+bc9tzvjrdtAnEAIdUnvcnKQhmhMx1KQuffVjS2/e07K6+Y2SL+k
RkXJEGHNor08FALV5K7+wOhuInuGUyJQrIpgfQ4elGIBXI2eTyTbxgG/IdfD9UV/X4rqA42Un0II
YluS4PadlLlMKMO7S+e314uIlmIwl5LQ5xKCjEls2nP9I96HQBJTr92fydIGVC7VVYMaAEmlnKhy
wjediIsRzRlzGFEnEAR8MQ+UYKjpZFg7/tqtbGf9eq+BbRIitdiwUkooddwYHV24M/gk2Z5QrKN8
bgcuo534D5MP/mOv9lcDhDVHwq+e1MMDRwrGYs2ouw3hkjy4AYQMIBLpzQ7b3s0tFDQgq4wJw+WH
2UHvUfPsTGxdf/+61NQ1sRGQou/F3KLIbeQEl9k9jeF/NKg4YszGgiM2RnZftH/HIhlDY2dcc7rt
jJW0Y9wsNRiDs+yiajfL77sArbxKR20TSnBS2QEFwTFv1iETwt1BEMqa+1co7H1o5Gikonhoxrje
VaQvs3n/p6jc1zDRdzVrBD0Rq8zmSH6ZK8BTBAxNrGft6WQuHACHm5B79BIVAATAtWX2Bg2GnxUd
QCBE/zMM32Xgs0l7BBA/FszjvCoPtU6Dd5J2dvcp0Va0+wVA6cVbHIz9f5lstAH1f5+bFUiBdON8
I4F0Dit1OHA1a16B/hiETXYo61uYebVUPaHmowE0tvLlJ93URGxq3CC6A2xnBuLHClSSeQYc+wQs
Ay0p0rtpBX8kyB7zpg8LYVPxT/MrdRHgthQbifUNSkcAh6kX2kuJ2WfTLt0gawEMEfcuKhw1Vk2Z
RM14q3lYZzT04aS6+duf4UVnq7Mr/AgdN1A5UUFF7l5vngCVzCj9jKVRmwxh4y2+mK+vo4B6P+ny
Zibt+jWvLC6dYABIU4+7cF//F0X9z9iw40QW59wwOlZFihSv52egw4H8fWvEl9r6Ln5y03fDI4fY
xsmoFmY9qOk9ANwJDiZiPJ0S7G4GKuivguTY4MhKbpKBH7mYVdkkJYwIc4EZmdPlXzFN74QNgVfK
xygKQEfTw9ls0wqItbksXkAzAXjyawjU40WfBWTaH92P5pRYaEkfNaOHKOARamHC7DSsaqsgLfAF
Jz9g5TYc0QU4bqitO4Xjy029RykvF0bDoZb0Kc94hlswwsOJ5MMIKne7gg9ZiR3IvTy7nxMlRFq+
T9nsoxzp0q9u9bzLY/RnO7K2+i/z9TMtr55jtBFIIg2ZGAj2J0F9BF9qTq6DJwBAe4em7daXLHIg
1FjDbr+ejuIU/lQQd3q2AdCZWS6s/s3bP2CwSX6V4ItLndTa5o8I1IMKUcO25vclQf6GXWe76DiG
tNf6Zhp1eL3EwmlIDIkJDHXDGbYRc7R9hpMWrn10VtvkdmO6I2DLGxaZV6vlfUfBcbMcyGFvtiCR
l84A5gCR38mflWZ7UL4V8PCm/VrywQXJBfWFK6+vMLImvNy5wxEfgyazO4U2SWQOO/H9GwiTmUui
lBewHEYzc60J357IRyT8LJMMAQdzPcitHo1W4D/1IPPsoM23u4OHk4/rvXQ+8f/A38yrVb0+qiKC
tseSQaoWnjIYdo/Fxpv527e1GCgeEASv0ecPE4bRV1rCR8wXOKmp79RmG6/UdQFqT5NCu2AnvQHk
/6KR6z0htOv1m8PgcZ/F9KNE6f6smDLxPZqNg6x726sdPEGcyJE4pWJ71sGS9St7PXIYsnkaLwE2
3xH8MAGo3kQbHJ1l2llmrwEmboZS7kXXqwyGTERwe/9yv+F4x3tG/JZzf1o2uA5TqVAQDoSnVTSC
Y6SCyb0GFufaRnBTaYVkqFfiA/zpMAeGZjnem3q1s6b2pkGU2uF4ilcP7ucZ8xEa9sLP8YcRlHsK
DAYUpxvK3MKDNLZuodJD9BnPuku8mR8nCDPfSWddgG6OSv5jgzJOoo6GnaFUhBdNhyuF7QIEnVwy
uGw8fmhO1p2TbW68C6Rxx/WA9WmnNIflFmYVeBq4paTR/O/IrGTt5vVDDpBA7vMT33NmUcVA85Cb
Lc1id8Rruwoa4sXY4Q4ii99Ji4grJJNRYib+d8NHROmiRusdLC7GewQAQxk8ZQx94Qbc++lX6JSE
DljgBHsf+/slV3jx8edo7Vl4eODpyobV1EmDnSeH+Zu92xz7h0j2E2LGn5iJKTbxpWCL0qjn0OK/
ULMGZdoGoZax6xpb81/iIhWqwQkVSjMc4QEmB0/IKf+I/esxR10PnY3E/iTWnnrkWqN4lwmSoEK3
YUZyeDoccIjIm3AlmOudsNiUq3Ot22N7YQDgo0WPC6BP3wNXrc+ImUI0kFNL3NxlRojFxMCG2ftM
EWgHhDHaaDduINN4gxjoux/Sj1WGjlFRJt+4eqSGfSB/vsTp64FqkNoG67Y/7AITRA9VNoBxHZez
V/riPaMtsSPKvHMIuCGqNJrSOjhbVC/F7msAj+iA5es73ef4ucfTGbET5Q26tEtmdCSGngaqRpyw
cSGg8FDApVmgk2MBDBZyND3LtSGO0vmaKqy5XdHNWU28ofCmWjHSJMm6huCpnXOFuorOKbp5erhg
5IPUX/XE1l8a7FwRbJr2aW8B5sC5nLroOq/caZaAwLNLB9hQwFcTsZc+S0/FhtlyaaRbNKQePMdu
+y0YjMqWwDXv7GZbjG1+OSaJm3jD81fHxOKmwj4RyZryDFGv65UTmp1Bkd2E7GnSPW+zWY5cWqbb
1Ywu3AXnmKr0z04rWj7TOWbvNLJ8icGOvLzoWuceuVmwDlQ7u44q7R+t6bQuiX83lfZDrRb7iGKx
2XkbYTS880fKBhDS2z65Pn5YbUl+j5THqHKvGPga3HZCMdQfvSeUOuSnXOEisWp7wRSpvrg17ktS
RF21vk329mMYEQAZVKGUDFAz9ABuyun/I0j0OiB39PKtfTPqjuRuT8W9VYzGZLZuTAQaZ+CUm0XK
zvritJKB0UYVxx72Bc0FB3EXEqEi2cPaXpcHjFQUo/izPFX1q2mykyTkmoTNi8EjdxG1/J/Na34d
dN0DIk/iI13Ar8phvONW2NFxFMDtyJeL4lP1pI5uYQawPwndd91KNuDUjR9IR8DRcuz+BgVB/N08
H/K+hgY7rxAswhzWt5q8ujSomEbkDUGRgpN82t52a4qn48jIKuDbrrmnbsxQtVzrRKGD8aJ/6N1P
GIg8Nlm5jEhhaIdrHwGQSJz5iNBTnOBBhkCWkcZ2AlElLU/zrkVKPxbDGzOIST+pYawFC2bH3tmb
uEY/ODC9/iFCDzr7u47y1sewRbP9d1hA+yCFZpJfMXZnzfqzrLiMIJuGrMNMdL7xCwLXSbxmmK5U
CgGIklMysbX6vB0j86JAz9Kleceyo/1q+DfxI+qYngrQd2Jmrd8RySLoLqOK5qQhRZGhuBjNF0e9
fRAlVfEWiP3SxNxFhjrnj4Jfi/nxGKNmBShfFvBJpYPw5refSWPCeGEiBZHBit7+FyYSuJWlU2Wg
AGy55wh9PCfJQhWNL8tE+/IvOJanQ4YninKxGLR5eEEp/qljBt704YXAl0c/OEkeKc8Yk/0pixaH
I2uL3i14aZpBHS0IALJSFPlGamKvOcjF91L/ZrDdSTGMa/PuoyJguLv16lo2G5uThlY4/lOub6Mp
Z1g+1+pNGFc/07rbZI39c9BOfUPZEl5CJswB2ZzvWCmpVD33XVVMB1pW6AfcMrDLC8qVQpcp7hNj
Rn1qV3B53SwvM91doyV3FDJaziMCwpjyd0E288Z5N3mymg0svNBqY+GC/uZ63Eh9F4T/3Rtewrrj
lpBSuewFTxE+7a/cA7NAX3s/pNmQ4ENS8MacErE4P00Bkx35a1p8kiDPqHStQroH22HjscdvKnia
z7kGszG7iAaRbEtOSqdqzDgje+yek91EHAaJRI9AWBDiSM9lamF3XSLeUBxB3hP9ht5jNWzggj1L
nMoILqM7iqCtQEggf2S5f7Xb5IqcNKDsTwkUcwiMtKuM/Vt6lzdLKWXYOZQPyTrxPKpXUqkL2Tnz
QRfvF+BuUfc3LCkCgqMxdeC29CwnNS99Qy5KoWUJfVLpn1rpLoo+Vh53tD1bUvZw/DjmjTQou99b
X3y2/UTVmIqyvneB8HPN7FiLTSWe/4RWjuB6Ue4UJ5+q0W4hwjddGey5g9cRvNvmOQ0weET+nbVT
693DfN627qovVxx79n0hK2VXJAAp1oEiIhV4iQnvAbItus+ZlPLBZAZLhPJXFsIesME2GY32KM9A
t5Wsj4P85Ya4Dv8o4gzZPlieeoa2JWP5dryBegtmD0XB5G3Jm5A6/WirSi6NuHMl2NBhM3VfbZ4J
s+2X4/ZgZXyvW8TZOGoj0BtnOIpauZUexMLiBn3miYSctR3CuN4Cvn8QmJvgWsPmNPop6Wzq12KA
oRIL6p+4c7bNgjgT8qZbRtkver+bcOVZz4f1dQwYFLUN+q2qyUm0ADB0ebJ7jISOinTRDALYaWFB
fukeht4uW7vYStwTjVVlv6hzava1FhkewPpzhP/lJtr6FRq41waCRXQYev1/hdQ4fqKoJyJmp7QM
FzAk3mMHCvlx4zf3VjfT1x7508n+bKOodu8SgY/AbG5IxGNu0rWN1gm9xLagKgfJuvq+AUVpBa4j
8WqBrxdA+wcYyuDjVjBYHVQi0hlGK7nZYoOJSIDDBlyYcqn7L/uVj2OST6OCSyDw8diE4S+R6lGY
NuITxbpWnt7H7D7SzquTvcT9MGMJUv3jQNsu2mK2Zz1RWiH2mihQIU3eQSTillOfb4y5gncCgjjZ
DFFLgiYzbFGPHyUmaUSwEatAit//GWAsKqQkVSJgiTRk00Be4uzEjuYrBPl5EQ78t5jZ9a9Hd6DT
IHQFQEr9lvcV8NqAmhr7J9Swz//V2IqD7qDm6Sxim7QbjPczhVw22kaHSQaPL4slB1GgUmFRnrVT
ZVrvaKjVgLKbbXzDAtI7I/C1byA4BtrwxXC75B4zoPZ23FEeC9x1bZ9q+OurtTrM33y8BJv/jZ6S
nSipNICmpHRshsY5LYhFg+rl8UoESlWyZE9U5QFwWmKmofC1tGIHxwXW8SIKu8gnXU/SVp8T5x9A
zbHZMQAWjjIiZZQLIXJ/dTQ5JhuvV+gHdD8TECisXIj50Wfb3Eii+XlGoPJq7Va1dOxHq3eLY+mC
Ge3RaTl5/IbZ/wYDaFrYt2vpu3X9xz3G6SWWiidf4X0wuBSJWoJSciDRqCxrcBZpdmRXY98j07R4
nIZh91fysUir4ZcxcYjWKH+sr0r/VZNPZhscZzUEMxqQxt3zkzjbMXorFB1UAfH6siPkup7VbzCJ
wwPxmhN+/lmuDEDK1Cr+5O8ok0rDOHBJy0YE8m8yGNtzMFU4qQ9ga56zSUR1gf+9c3UvZfLrgvNQ
IGTEXqcOQP6LyZdhyZXZcUnhj3w9BYDTU4TMao0RzhAWinHKaBwzxfbxW9utlbXI9ChnIAalSobN
Lv0S+bQp0JV05A1V44X/04ZXpG/sNK2vLxrBERbJwndnGQXoDQPHmXnNRedzH37fEFDMBDWjjSNo
XzDao36haL7YYFKL1wMHHNnRpRW52gvD1soKpUmHyJH1MOssvyJAf36TL7SRDsszXL2n0c/oX1aN
Yf79n4qtD0FxPhL21sz/fN5Y4v8IiiQ8LNsOJoYqC+6tURfoALhyagejcxvWTMHJ+qHhfolZ1jWq
6Q1AKfDQHgVRSYqg91tee5GDPkQnV3vMX9ZIOQ1qhtYmDFuRboitLUb05nL9HPoO3w6pb5X3pCgG
cnjHNy4zd4cqreIp2Lq9KgZX3DgrUEOeuJoHDhABlimJU0QFPj59XLd1gn9jE5j5dZZPbi/Tu5Uc
KsJAH14fxxHU8+oJ+TDfIZVtcoTG4iJ9SAVRxL7c1atcZHeb+D/xrRu7YjSg/HQaN3lNqfVRp04a
ByV2KvfOpkreZEJ65Eq7jU95uPU5Ai/djUid1LjySa0ArGBsQqCNLgDeU/9F/mFVnrfIpxzkfBwy
1RsrUFxWIj3DD1d/ddOfUwJAe0S5RXCLrf7P9jtO3Au6dS3K4ZsPMOESuxTmXneA1dznyL0aVuf4
54SoEmT4NSuzqLBwRXqOJW/avnFwynzHxks0mTnAakObpEMP2FNah89Aj/J4+8YwiYDSMQ6m76qi
fzG5v1LGSrrHwNaxIHNToaHWGathiaCF9qjdTo3ruvB3OTO2kF+uSUsckmjYD3lFOcGVY3qZ9iTY
LKJsAz9jsA35JalrnycJE+fwhKsSQ56v7ZPgG6Vqu2pRNvdfrufSRiXVfDK8AZnreJa1geNbAKWZ
iEXsB4/XiwUiILZ++b6P61KY48XQsZ/RZF8S+QP9p5zQVFwDoNbLMi1qzJjKhz9/jbMAABWztzQS
UKZidSHEML2tqSRG1BUpQ5I3LYO7tQl6hgkI/5hYV5SEdmmWTje3iWUFFauU8A06H7GFtGn2/Hbv
HyqGR1Dfy38nIkO1GkE9JWa4O4fJSet8D1wGxyp4XmMRoDpniVdIRFNuwzBGSd7bd1KP6n2k9qi4
mxiwf6GCVEXNf/VRXcXyHEJ1raX+2Qcz9IZz8wJjlLYKnVBZG0B97wC0ITLcibk8wDNSwY96mHQi
MGJJs3ohNK4yhitY0O6iGckG9d+mkshtmUSASaMHT6hlQnQgT56M013Kaf72MgZKycV3Cs3kqGt/
epRrfd6A0MgyMZvk+dMd16ls05Im4e1CxnF6enJbJHIIxfX8h6H3Rw2vKdG5W78SnGs8qSNCqXBD
I/amMxYlH515K8FHstesxruNXL+9NmmFYBQNVnX3nkhxc67Akj5NMGbwDTeME8jB+LtAL7NoPUwx
klQ5qDvC4aQ4XT7JQZFKk7PodpBs+s/785nUXeLonfYptBjbV7omuKV+Cjsasuwz81M4qu9J0Bl+
7/az5SYnQ/tm6i6ZsPvG/fdPGP9bIeLW8QuH7okVwzCslBptUZprZZAyEVd3Cz2W+78wLrKnxGxc
FEuGE0HasPP0mcMxEReEtIS1cqReJ70/YAtUqQCf43vYuuE0bbayTnmB/rFYQ6IPsECU3Y0HgB6M
NpGGAe4K4bZSYqiwLxxE0SLW5EbZr7uup8OeDZJkIqjWB6a8aRQ/w0xo42hkUNYS/0F/GCOYmJq8
n2KmXNy6nNSk8ZFV3g/fgeNqt6dBGgwhaic69/pxzKJT13uScuWrbkIAUQw9kLqHjh4WXUYxDudx
SIHVel+u/0QQxY3lkXaXiUAB4lJXb6/Ah1ePI8peBlOGcy89RBXU+YtlP0TLG5rTXADxhopBiQEQ
u3pSqIs2GJXqRN/jFsgd9l6lsBaORHOu0kDKQYWKHk3/pH+ms3dsgxrOUmW7vMA9aPZlMJSsrKn5
KxqKPA+gPA3mVQm2gXodshiVaundzFF+gaUlOFDQlon0lBEVzcrzrKZXA6uhbK1tWoXRKPJ5hrv6
i/+oX8m0vov3aHd2tw0dXKTugkC0o2rq1ZVaJhMVTkPM5PRSMgaK4VcNEMEsRzCtED2fw2KuyTcw
uAakUZA/E+DJcVjGHZgXMRAebj4e8mkJNsYe98Qil6xxdZo1XJqSp/BsVvUpLci1NoriHjehox+W
47G9+8730eOZioQnpyATpz8Qd1KiYIST8i7s4iRgz7l2n46GMIC0hH40FUhqXOYGHbp/NesBYws+
t3XiRvvtgKSYGChLXYi0cSznByg7naHBio4tPj7FlZMcUpT0CzvLisPpNkCOgl+kr9sjVNrKdZPY
GeV6Bp/LhlGe5jX7dYbCCrP3q1pNAs1lOoWZWHGJSHD9Z9bnU+G6Axu8uHEBhoFxi+odfEcBfFOu
LMV+bExfuGfrTdWXTVaNoPcoer7YfdFEL59cNLSoXAbRxNSRQ69rUkkMIOiuclt62WXjfxOuXEJJ
lK1e6ZCbeUc57QDI8FnqxcHnjH2VpUVPbwU2TaV6R0+7uzLnWq9eSr3G+wxsdKONnIc6KNzfiI3p
kBkTIpvwekwHWzLVOFyIn9jG3IYSOVTjVHfB4Tt78CONUog5XSAbe+gCxn42RVgUlGRe8R8BMV3W
KHokNynM+8wBctfbupFXmwCpWij6vPeBYnJwp6t8390hr5T7Fc00C20RlpU0WW+WXoHyKZcjqYQb
oZtemliM6x3jxyH3diAtKv7C6FaX4MtLIa2kohHU8wLwQxqyGtbrwrE28Qg+L4RHwRZDOYBjC3Cv
xGXw5VWCfFV1S21iF4hMicirlVawer0DdUq7/ps6AFd4BQ+qF9ulwhAznV+huD22WCEbhPfgAGjM
ShwSs8Vs838gIIUUkdV+bH5mjgDf2nWF4t+g4pBPkzH8+p2+rLj/5qzCClr8oeHNxLPL4383RWhD
OYkZf1vXO0ux3fSix/uz+j4BppX6K5/sOLk7EWX06Z2QN89Mg/czr43/RHMwq+jd3NcVcb6KTF5C
iGwYa8R1YokicTAaYx+HskJht821iDjJ6xG+VHHihvWPJHhESUeUnSUmd/WKg4s7BCCDYpJKa+K8
/uqNvTdGymMaUIAtYomJOTob76UjS1X0tQI1bCFvA1euHueVgK9pdWCa6pnSZ8g6A8+Fsp4QLoDU
wVV6eamOGqvqu9EIIwVzszehoqS5PXr+61W1ByvCQrPw5u+bdxXHJs5yFwWXeKa0k/63QDlwT9WL
mVDBAs7D3Rl56c6vmpvvhJBc+AtXSVU/m3bKQBPtG1LLVU4YCCOAQAFTx10LL+kE6SPtIAqtYGU8
9/4u5wu6sW93nbESrdTgBzUPcNz7tnDCbFhAhFwjtSB7Fz7bstbwQ2UwUqQNDZgLscdeTlOfIaEX
93imE2YlRq9YHiROz9XmpZRoPl3lRGkV7ZGC6DWN2sM+gbM6n4yMVPYLdz64gekoiSUowSfZBK23
LyH3lYSoP6pz5XUeh6SydK9PGJJLI1WJ0qzeTJZkN8iDfZ+eZIgy9RR3tVhwPJ+bBmQEVAbYLLUy
hHL4/nhNwJI+8Z1yaNZzdtJAWNk95+gK/NiYl7Xen4qPrAhp3+J7NLmcGLI988bkKbaTClmfLYoH
XOWsIac7m6/xUpuO8koLTJXdsT6YQKs52jZ9Q3el6zt0WRCmIwWWebTEPpUMhqKb1ceprPK2xges
B22CjR45bW3hD6hihxWxEjryogT0cNajvrJADOFI3gG/OnPP77LuGfbpoM03XcDpjdFQ++ebHbni
pAOeaAVlkWyphcrD0zVmBVwbTxEenOEOqJUX0cQPsWk+n2AQ3RSnWsbK+HZ2zJScr85jSPK/oboe
GowDi+7a/k6FLet+/KNu36SNXlNvNvQONSwQjEDT7X0v2x6EmZv4szJjj25+wWoyzRsw9qUUhGAT
4NpzZv4jG1xWzm5u6TxDoOkmpFnOttOLRqViPGbzfqfsR76jmRv4jQzf9IcbGnMMQFZQJJQPiYNU
agMtx72dNDWslxDzk8WdToq9RybMrzT80s8dgVhFcHGEEE5OoFcHbo94rjyRRVUhRs7Cohvza7sh
snZr8h+yfUxwAhKTEE7LYOYYwr3qRaekJPjnwIg2ULqD208NHO1A9Xrbehv2IBWNC1JpBtE60ZLr
V+PVW1dnucTZOEjU3CmnaCWUr7SUxvR/hbP/69mSH1PYabFvIThRrFyptQNEXvnNnQcBUnKJuiNd
T1lqSDco5uniQR/aAfYpyqZ5koA2vUE3FAty+Ws3g2x5cN8ljnKN0qx3zWLVUnGpR/U5QK4wO2IR
LUY238I103O51vghoOe6T7/Hr46cLUY+9F8kxJfQOyvJBjyiCAiXRDUL8l8sGDDZcHrPUfgnh8v9
7wSCyDA7pNU3zAlEB+RV+KAXjA5aIIkT9Q2c3c1i4QwP4uaf4FyGHuJo13uv8IrW0PgiZ+gU3f9j
4RXynELWXpXUx0d8GCpV069kToUjDXAw+L/VFi9Z4+jCUuP76WlaHC8UBA2xvaXxsJU1qn5/lU9k
DPVaDocKNTgnWYHkICQqeO+pLP2sU+thtjsefgddvJh073GUPEIAQr5U3j7JQobFFxW1nZ67RvMy
OEZrt1xq9LqH2Sx5N/2ZYIoFWAcyrhRm29ECGd6mWiAYok+B0IGDC5fpt3rKiGGslCYfZfb/KR4t
e1u5BBcMg4GFi4TOkUJOsQcTp7ZsQeCiEwjxyO4lf054y0QzRfRCghedcCFCzX/vaVXvmtnJc2CA
Ur36iYUocva/0auBripGSLIoSYugeaF217BqBOGj/6RwPVGV3/U9l++uDkxrphta+UEluXm68Qvw
+05SXZ3zWZG3EOtVCwfrG9AsiWjpouteou8j+fxARuo6hM/HuttDQwDuHDnPKXZ+qp0rbVxOQsUo
ikwXCdBbpiKdeQrGx1AA+dAciWMvrC76aPTfAPOcqsTPr8Ly7ZmphOY1CE09Yjavx7UVT9TCM67P
IthJSVcEwIiw6vgtxzfkQhxx56PWNMuoU7lp9zNm/ECPn6705t5sizZUaHj9S2XdNcm9RuluG9DA
1qK/c7XpRgK4PJdLkqT43ExD1JGpRpvlz45yXnbxHFfiN75UOYDB+mXfiuaxQQgAl8oc7vnkNUo/
yZH0pwj8iIft3txhDvVW+XtYxCc9aUzR2W0nr7OJ61X/Nd4dd5+pWrGzRTIsenFSQsxe2EgRPyrL
dSoTQuBOWecDOfotwN1EaO0pCwXHDffNSkJtMteRVgleFmAp9JIPPb7sOPoCBTjg0U1J402a4Nqk
+AD+jvTZ3SPkhehfohzFIM5N0qi192QhEUxNfmKV8eVGw6Q6Jxyky95ZnJpOOhfsV/yd1UE+3z9o
JLJVFV4y1nt4M9KdMSDNRizCosDb4hMo1PHpT2gZ3NjPBCNCv3qofYvWW4B0YFbbZm3uS6H39DCq
U11Y5RZ3EKeprC4pL/8ENmRS4jhDYxzVvKawLPuhEVDzwIejZlYnIXTclyq1Hrvy5yw+zBMhjxxs
+NmmlyqJ+QqCJ507h3RgfY76YzRePmGEj3IsYnXHZIc2VokWupISn+isrOGbPNB3YV93VS2Ig+7J
FiQJvgTBeks1m7aECc2OUR80/yZmhW5sgsRtI70DQq3W6NczZ4sDU8AJUbSj31X8ln3a6Y3+iVqz
kNZFon2ilxX871/RB85KH0Q0yUuNyU2LprGhOQCxrAapRJ9sLhYjd4qiKBSXtDfd8b0wSku4Wda6
vvatQhSinlMi9PAlJ6pvxBXegh7Jh1gjzhYrEL+5PBZsRt0qmXfnMc6m3xTenreJPuMR5pDae8EX
JEo7l1kHbwNpJ+wGfbiprs1LXU4BfWHrMdcWkBVmxEnABiX6xSLZ93YRlbvvSo8hAmh7urPs8oPs
Tyfz0sYZSofBmB2ft4DEmflK8+WjWAEdnPH5C0PS2nQht7RQSL6F9MxMhRWlwbXDXn5r3Rkgt1mq
seoKTQlqF3e7QOI6cv/RVo79OzwtTiRGJQRiYXVSy0JrXMdSisJyeh/EBpjU3N/jIL1tbfYRo3LJ
CEJMysy9wkJDfg/3lFMpSzi3jZxccP9msLlThJuISdo+pagX+Wm+MQkymG07rMQThU4w3K9Rf2Ah
kpaFDlgaswG6d4x88wBcDgjedK5ozxSdC/ZKmLHVW5t+iDQykq3digkw3RUyPAVTRNcgM+8J/k7x
zlkRVZ5sbxcFAehsLhdrohebu9A7FRmDPd7nQJF6+93M1RRkY3cxEv3hSD7MmCIxTNIowfslCQvv
3i7ccnYZUk5VQCccQyBSe9m03S+y8jsKkXPZBcAcHiDRztzhtFVI6TCIycO+R2mUWHELp27OUbuS
+/k3GP1T/8sInvblzxbyTh9jVFE2lxbiBEV83Mf/LM0FN5cJIxnSU2gw21GhgOdvEKd4adx4vq+R
OVYU/6ZlsyvwVZQm4joj1duVjCbNaoguqu+bcbOubWlbcbFvifDrFsiZ1us9ZxwTfbGbJn653o5q
cYf4P6hJMbkxEbTvRAUa4hfKKvI2kmcW0/Bx2uTw+CuqVPDLtq/r1ZF4l1Fn9/Bvxedb0pHlJJtb
Sk58HQHCpaiWU/94THzf3wUe0BsrZ5otdSXXrqcstSIMclBQrbh263u1ndoq9CDoTez57B5c8kk9
wUbHkztK4426waMB/NxAZZfIyqtgijndZE0Zku6yx+cSWILRs9XAck+UvkxcthYT9T4VFptP6kVn
YI8XCbVp4AZwsq5Bwh81ppvpWEglIdsgA4b3C2l396M6YnwARsGpLhK4qjLbj+pCQvB7g1igk3M4
Y3+ZDoUkFttozmmqnwhyajEMlKEw5M9ZjnwSLmWsE63rApIv8S//59CXiz1MrZR3aRtI2bOeVshh
hBDfQ0ZW9C8lYAVo2fQ+J8AE/CM6L/K66WnskvQZZUVjrLuJkQrBcyY1L2xwMMOI6UIcikDnqT5w
ItJPhc5dQLHdwYhSFOBGGxjusD+D5CFtrdpRdKE7c654/pzBON2/GJrm4fKzpKRqC4C79TWCsoH/
tHGoRZmWLk9zldADysuKv9Vyn73JpWzFRcOHIAYiikgL4YaDGobquRVLSKbrfgx5P8YpgyAvNvJ2
YX8kmFyFreVRNfLNsk2n7GKC2Kwce29tKoNNY5xZzLB4XXWgsSuNRSFwpkwTph73LX2J+C+wXfJe
Z7qEocxHGHxzPK/U58WCilhwaBtBjWcshLRFjaxUvWuOO8KdxP1VKj0Yk1cNXP2SD9E2VLNutkVA
3sLXuESR/leVj3Li4T2tJw6RdmhN2UIQxGQfYfBFM5z1BCBaaZt3Bsc2o7imL5ya1SWWiJ0FrUBo
Q39Zoiz4+gE6pZRgr2wSUUv7dpBAlumdPMp6ijl1YNJ6+SXw+VY930DRWH/6jQbnr3fmvlcGdZIO
zbqDtsZ8fpNGmRWepD6QQj29nyipBhwQClebzqsNyS2OG0IzHm7A44dcsR78AuGxB+EE61TDyfTr
ARIob4zGfiIia7u0dfDIY0gFe2ZEKDBJ+LTVQpInFzk1W7edyfDxiBoJZxNgs7AksuSrjrW8lxzk
doUYQPJ86/7oNOvHdydhoaxxrZc9aRCnwAbtXWiY0/f+ZKL3Ky8LOW9lH6YrwQNIJZEztIFYxQsF
LXstLeEb1EwRln6qYbABmjgMhcd+JTjlBC3kF4c4nCD6CeUUf/5dnFZ+d/Ttx1YJIOzhU2uwZOGw
A7qpw14kj82iktKyFc5tJ+L/6YaD5Um1JNa+ZDyN3UHMyDSYxTEOZMpDqxV2bJ3cnA5qIe9QWaU6
H8VqEKy4y3MGRw76O8Q+P7dWuo/WiGMun8yUNsmlRf9esiCsepo1B/wXpj5/INenH3EKmOneHuTR
+692xWCzH1PxU6E1lR+pbBd45C0Z5dxFe1h8mfmYW1AHpIEOJozAmHJuPPqkNlBWhU+4Mz24JcWi
VLBVrAmC6p4y7gOlcXbpkrZpg3wYSEu996FS9Yvl6gC3bcSqFM1icjofvcI9Xhp1jDhebv/bmwno
iSV/rrJTmBZWGjcnYt7wSEDB5xYOlWx+TZ8rtNoVxYPzMckVruaBU8iRzWxfDmxleZrYC6qTQrBQ
GA+hNA2YMwp5SdanBiQcwzu5PRRIquJEjuqgfWNzwxc9yMyj1pOcgS+kG6Fc+P58V4E9v5WaMWlF
ucx0QrndNd95E+BJCl+ofb84OCpW6vXeQ6CVlUnrypoocJ7p4IPsYCokD555EHVkODL07iuEYBxx
FLcy4VQPU0l40DuVhirEBVtxkRZET+Ny399i7WkvArA3lIHqCJoxb+7wAoYjBtWTapDg4u4WUwIB
LAylP2s0j5kD29bHzBvob5YLDHMrIy2B30sg56M7xFxdx67SVzeG4yegr2oxh2B4nm1W/ANsE3/O
vh9auN0CuZT+u+Hw4n2EGFy5jrobosNwoTaSXAezzanlImnoXbwdA0G3ZpKZ2NJs6jYk8vrAdm7H
ttr8w4l+dXp9mcBiUCOzgCW/aeYmqr7caQAtcnxdKSUYHPecH2YlUBTnnab8FiOtxC4OR3NNcdc+
EaKL/6MvYJiJ1M+XynzbGttZUk8OlYx7BkCCqTKQHL+0K7UdiuubdxMtwaRlKz37/VpI/mrhdOJg
sLQlWl/bx9VQ64MxtozMptIJ+SNwU4cEhnkYMrfXeJAwG+vqgdixUeZ+EIHQtBwgJ+WTZR1cidyS
ebBwp087I9yapNX6SmoylWXsRg9MIcv0M7SfKBCd+IxicaqedAjqibss4iwdmapNHOfurjJAuOHt
vGs8eC0eRBNd6ExHmWhNPxFGoT1GTFs8F8jN42oP0kMHhl1NPuSd8O+UeH6EeiY2+hj3OKg3fqv0
lU0qmaeiX00QCnYazWlpLjWURYYjugEmaDrB5ft4Wnyk3c+sOmCOaW6XpKj9+DwDhs6xBQUHRcX6
HVlPaRk8x1pgdI/YrMNR+gjwAcsPs63E9uq2k8hvoFpRqrcQiCQnd4IPbJ5IYbVDo1kqLrhbHnEB
tZYvVNbE2IJ69uG9ZRp5vGOY+z3ZBz4jxnpmx6xmPFSWTWbM+H1pW1JmNDOF0KJ8DDLN6NwI37lY
FM+GOOgv2rHFx8bsYUFvLa8jcfjuUfF+FJ9SAdouhBP8BWfhGW0UKc9zVRc3HbVjYH+96lAShBPn
PiCHg6pgm2OoDZK/HG5gxfSTHEGLC0F7a1KuYAsnNAJoGXI4iTW1p4Do22z5u8BSFbbSidh4rlR5
MP93SWONDfTz5t8fHKWo73PFmpJljPKbFDbLn2N6JafiUkJEq6koP540haooOANMQ/C1MqrzBtDC
RuRpZak+PBPUETmHtNXGd2PvGckttyptFyQdP0mvLHNFI5tndvqPuNLCiked3fhZsfzvCbA44Cns
F7YFu/KmH3ArKpPsiT8u/aP9yZCiDWdYp0tVCqLEBzXZNjdvf1icJbi7f4VF374RpNjXw/4VvNSQ
a9SpaesJ9cxj4OYTXqkzl7ZpccxAdoNPw6IYUSdBMDW5wQkFGA/AIMLz8Ivmd5MufEJhZyLTwzYC
inrvxzLxbJltsmUWqEPvQpddEg8wBnIzHWStUHLzyFIh+Ep2zTGMHML+oCvtoHILoCzxWH1GdhYw
xqRuK29u3l4taOS9USA8hSZfK166iTwUe3gXz3OBIWGl8XZWCgyC7z3VrNNqJhKznal76ijRnBed
cjpzsBp1h1gXk4vw1hkJ4vKiWvOun0S8FjvuwxIcAUbe+perETNb7NTNABVw2n6teh1Rs3LwMTMa
zGOUywSyTTadSUug9npieQzGclLN6EOf3y7y2f7vIndS4iqCki5I2gVvi6hNIOXNGdbnmFkKCSQE
WebqzFvuT85DFrT+OUeRSxJ+LEKuHUW3y7whrSWIpfcta++/UAJrpcF0VkJHqKSBMG/yK02YEfSS
uomX7rCguZHG7AJOETIwiQN+KLN0uxV7fgg0WtIRtC2YlbZpfvkJpaASNom+H3AfjrKyDlVehp/S
aBa7KiV/1t8k68gG8I+oqUcsc4OYGNqQFpXCijgQxFn3cMbIe3q3xFqQM7XJVU4uOuLyqdbCTcwZ
HI0myNVz1GutzHRjtdySWAckKgjil6jRq3M1lW3xm5OpQyOCYYz9jkS2bxc+sB0yoODIWlQHS882
vfESOUhcE5YZyreS4X8q8hKAAFF9KIE++ieqzqaoyaX66QvdRc8cyRbVJ/+IEzNbPuzs7p6/TLcm
RwdS9AxIknhiUr+xBprSgoZ2VBB17dbMhan7FbqWzpADlbA9RqOOWns1AsEG9aIh+JInRVc50CWL
7Y6snFE4ZPbNX96FHKPK0W4Kg9Yl7woFjuBDzna1w9Qu6VWmctx1phRO3X/rrmCUPagm5+V7PhnI
3o6jI5tDYp61j71qCVyTnD7EJOPuFg0slVD2rmd2pSIN2+xj06EI4+Z1DoJ4635orZJzNit9qeBA
3hh5rkM6CoS816KgN8/DoEDcl6r1eFVOoN7AAabPbJRjJnC5zP6mIyZgfHJ3LNfFVw3K051So3lM
sMQI3ISy9Hgsvf2VyDrNGaRmzI0FwRXyKZCO9gGYxHKMNb2zen5i+sMQC85sTqIG74TeBclNXRXl
7CduC2uTGT2uqzumpO+JnvrE6bVHkMAVlYiIqCmBYfmzP0nAFtSSGCKMRuP/spDwu93NcXgkdIB3
ywL7Gu5cAipZdVeNzO5tcEN+ZejkxWA8/17Fh/hc4f8dQ/cOOD0ISVeB4pkIRlJDhpF847fziA5J
iF86z8dn2rwtM7slRQcdA3QyPMlmeh74ZOpiZIg2eooe7Wy2Jf1xo/EcLZGyCoxG41Be6eS8zGGj
rs8IYLXH3hzYFaUDRF+U/5Nil7lUgq12LaTMQYlRPx7J1srUQvRo+C2K3vteoURlF+XHUztnAoAl
Fpfh3QHRUpiv2b/GE7jwW5RPeI+O1UJCxGcGNC0u0AqzPO5Rz5d0gBEO1vbObQdcFM13Lf2LafXJ
CQNYiNExI8Ph2nCEuR8I6WEk+RdqRwpUg33jCLfG6rk4K0T5A0EIJhSAVRneaZC2UgDPnR6aQeY1
yZPNJoDyKar8xpUmRwX0dNdEKgwPSPHYwVUYiB/pnAn04xIwC3LNGpFNfZpCbZfkWb4HpTPkpWZe
iBeSsfQnVOMseUMp4KDYXnb88umIH8HcJXaNlhujwDgVAWYISyK/XYrbpivkSQ2brIhl5OgwK3CF
NMBdjWxqKpQXElujI5rQqxjHc0aH7lKfaXjcCTwWtkW7j87WKDGD37rgi/vT1ncKTn9UqyAuEvtV
P5Ssq4V0Tx5okvDFrArupluT8Ozmu2awunbnfAbR5qJ/aLBSuzz0pSL9cnP28WvzPh3tOGwXVSRQ
ddVm45qUDVYA4lF/7J/AAF46omJcqyruJYcrSUDlJjPfFUaI3tO5L7OZ9ICWKbPEv3mX+xFvHDvz
V2MWB/yZQX63uGUwbRj2rFBAzuy2fyXMHpNJaEm7IYZEco+88lvN612YAhq1F6TJNEQ9sMeWGRGU
IrSLrgINur823xAeTqLpPs4zj3aW+yJi9raZdqVPIYXeB9TA8eB/ZICPQbwdAC6ELyFjfqq1goEp
mkCYjK+1GSQXF6vd5biADhZ8rptySANpKTw4c7nuJ0Wy0BKOKzvENkolO1T01mwVFiMyhwojMS5G
BHwRW3rD5yRpAfzBhB9/MCBnk++aynhdtNXFW7iz+lulLsE0o77AkHm4pdB5LR0LGp04oIrxzOXD
rZLS/tNBpfp9DUlchgbYx3yoSJqrwwX4OKHkkBXRbkwON+YsTGgAwKySm79jfqYwDBWjgaHQbqaZ
WbWoehFwDyteT6+975BuHyOxRLczGlQIJASB0hxZl/ZiD3aSzpSO7GAZJ3KjLd+Tj0M/OOTFTg0X
uQKRewyzAmR4Dv81zxbQWMni0gxHqQwbXJ1MNC+WMCYfomii4tpYe7fif6RSXhrCpiyUrq8/eYVL
RCzdqR2eOVl+vIN5OKxKpMxbCjc/jXrmyH9bxJ6+tnJqIX2w1NNi2CINqohYe283YEd9LmLV6O9A
rPB+gqcf9LxBxCXL5iRsyHdk7JMa4i1owBeLpkwJIREWWjWsGh58Qhf/5l8IuPslHhHZ1ac0S71s
LKnyIUNSTusFAFG68ExiEJiOCG3JqLchwjVwdvMMk+QkRMXywO0LQUHHTIYu63PdmPBq6KPy8wsk
0JfrmpI4cunJYkXnbRFUk09n7+ogwX6KlTBGOCADyhFpIe8NBg4g8T8sGepuZ8uxioaeCPP31YLH
XHw3Y0cDA3RJk6YUnGGPhfafz7CmDDe6iMbwoLUyIIRkwYK5kmvz3s+d3uqekRP11N1RecqDLsn2
Bwb4m/AA5SdQaDRFuHhM/8tgSZy/R0Xf7+RhaguaJmyIzI5UZuSIrxDPl6n5mUttfmgBGoag/Oht
rOHUPxW1Gy4ZO50ApuvD7S98bN4srpfOpsRGPIJbr2ri4HqXX3vCnxNiVLlD0WKxGXPOVEyVoahQ
wN4KPjfIf5dwzpIxNzzhJK3itwET2kFupH7pVanoTwfS+mE9y6cGSAg6TpGT3Da2aoGnrpHOdMvS
bUUxKWVTGRKphmX+uXs12Xx5QkzN8bgAaV+MFlXUCF5AAzFOUwok9DKbHvK3ZCf4h499DojviPSs
Ldic1y4gePkhJmrYa/nCAoLMEpKk0/PqMReNJxgujUzvcH1ymriVT5Y6WviU23RFlDXKbWSO16Qc
aPO4QbNZJHf/wFV6FgdLBTScJXJ1t+8Bg5dMWD+VhygZfYEmbW4IsGaJO4/g2a07deVrmo9WRV0i
+prn24sVmhnxEGyWHjSWl/cURh+ipRiLLGg48aI+P8wuFlZGcWogYtxnX7SgjUYAloi3Jw8S9zEW
7C86gOt+pAK92/3NhtOATsQe/lHkrde6fi2EcMWKkBZNfHFJ+GU5DiXqKij38oNk+PS5ueLJG04w
+S8sH5QI/C9Dmm+2RazrvbFRJWswP5A0HFDzq2tjfRweEPRYpoBOgS9cGVy76WpsBxMZD2tw0QTN
PrRSzw/Iw/rT4IY0fe/+K7RGn11o6cZR7E9b5G2p5Elt3WTWXM0JA7Qce8B8g03fPbSJuCH/eLyW
VOtB9d4mim4KlsS8pXbXOSuvLGmBTKh47ZQod/C7P7AKrKKMWondQ8J4eGtcMRql/YwrNBC1Y9WP
WhRiWnlWATrdJujxxPBPPS+QS8iSUOkNOxXE/vfRRHGybvE7jk5y0f6CtR4ZgOpnbAmeE4zaQ4yV
wpW3g3MuLRb85nXDs71kQS7IkGHGZrxIj/VE8CkkuARdRDp347z7fhYuN+in/ELB2CCbUOLdCJ3W
2PGRGLo+dcMvmts8XTErHN44feSHZYK2eFBteN+AASBX2qW6u7G199hYY7aRrB8mLuS/Sbl9Nx8c
pnL0sXOqo9Unb2tyRv6C53dvVZ4Ykgs58P7pC4dC47U49o6oUo0px6nzhWyBeqKukGCQHRZBVWZ5
P49uUNQcibr69tHmPthaYJMbM2dEwDg0M30LrSOMnhK+7jS0D46elAiG+DJtkfD0RpoejnIGs5q9
20YKBUNrWdMOS+mcM2CpLf4gP9jG0D4n0ZBDf71Ezdo0k2zn45vcZafvaihJCeap2tAuuRUGrbq0
wBODZDqIAZanoOSbjkMuK2XLNoZg9bIVVunF0aoAL08uJmxLQwm4s54+bTZ3uwrSp+FcWjM6bcVv
SWMSYbXaZbHTxJLw7eT8HHnQlJYoleQCzm6lp55Fhy0lsM+RwnRZFmgsAyng0fsYm/BZM+t2rcNI
L41coz/lqDq93nfaY+LWo0izpOnykzBaDEqiEga40dLzoxpV0KKdTIqlodOu84Ii+tr6mIA1MfBS
I1HecC8c8lTeEcEG6lClA6uo7bU8s4VzHEayjcEac7Zn9ZevqrzZ+f0FXvekwTQudPyGM6af9DGy
dpmN9B8YNMzat5FQiHH6RlQ/81N/LykL/x656j4bLdthyG2+BpYtnFmZZmKVezHE3TdRL6iX5XkQ
Qj/VDiITQ0Os5w4WY2csp3oozMOB5gI/Ta+klapxsEBKvV9jhoiDUgDgOouVzOJl/GyLJic3Oxrf
MOVcVJGfzOwfllDumQQ4SVKCr7virL5tmDonVjnbO72A9DGn0rXllqqyXPvDW5Lsrnw6PZou0+4v
tGm7VevrFI+U8FmaH/Y4mtjVN5ahQuaQLYfQjoPPU1+3wr2UuCKPS1no0XSaWSO9hYyIDBSDzd3Y
FMrksxOb3G4IYStz33Qp+ANVam2qSBqA5afnLI06brnGL9mSB8vHfISRdo/Q5f243aa/JJ5Qm907
lK5dFx7EFQ4wBHEIvBw9rHv6/CSWgDMtJu8dcDoTV+9L/cE5ytfWtoHkQfQJAIuVWMDKS14BfkPh
niSqMTDKnTkUUBdRdvAEizm56IPj66RqcEMpBm4ZvDjMpVb3eKbzSczo9hE5Q32KU0FE3ZKGcJox
E34OJV77HYsATu+l5wGq2vSIu0YhuVr6POvRgUKLix+2RgfwrSwJWzXj4OaampuPYqWvuOl9rxrc
Z1/99c7PLTsOgTCYadb3+WYw0R8ZeAzOC6vPHvrVmXGl5vuUqJmQaas4lXe6M+BqiG9L+mBQZsAX
z/Y0U7d/K20ixyHoQVq72ZCSlHDKMSAV/Nbi99vfhoM06Yy3juMwqV+70Evat1MzXaZazFZuP1U+
ZMsLPMgKH1c+cihLqpMZ62tKR0FTzoP0g84dfOb7HhSRcYAmRASzZQD+mRMGsZtSG6jxCjCkrCoh
knMLhEqhGG7AlyV+NiNvfKSsekSpycu5IMZvNV/6VEsv3VwAVn2iv8CfCH6+oGfgjy1dXUC9f37D
UP7OtBIAzkD69Vqu6Wt5KZQX0BgQrbPpXxR2M2xoZmVh3jhJJ97nmxqCa+x7moOzBW21+uB55H48
THpgmyrTQLbqZNDzKBXhOal1VVt2ljwwtcathDDJXjWrDZWkYrs9vZlLRXgmxxhluqzMc5lbvn8B
B2GDMBGcwei6GLNxFKL0CpeOIJbOcnW9KI3KF0ElYRsPqhPWK1f11osqRfLa652+JZm/wzRQhW+W
b0j8HBeCnPexFLRwKmX63Kkg02eT9U7FAUEXU2MlGfoOs6OcN6ghlJujdbEcVQ4tXa+GtMa7vBbZ
FCIpZdCLOW6tORYy/Q60LG/NDBTOW79yKkCSDpQyHylYTjZkXqpko9gxw43lOTq3oZ/xQkvoQxpi
JzsYY4PRWd1ROz1Z0sZIDJO7wBXQoYScsMHkAaTug5JJqyBPFiRQ14Mx10rr/4oY8EdtCvh4VSjr
RRjIBsY+eJpdK0eEIHElgzYmmNcndDIz2SpNmAmEKp9nlAkoYkmAhut/Uz+GdffouUA2yVTM+Hg7
0akvnk2sptxEpTc88bhLMMcrYYr0YW6nWYfqNkgbR473m6ynual5UY8ozC3RtuuBMBFAKopMgdU7
ZU8Q/7n2hWVzFe/adtTJVWZeyUSY574+om0F1GmdebpIRItHCSSLUxSZEAtzGoIOATS6xR5QK9OO
Gd9WlrReW5YtyI5PkBqoDTWGZyDSr/1Bn7DNP1ROBclcCiaM9Qi0Nd402AwLKyQu7F0iOc+tVGdn
hxxbKkiLWlcFaNYVaHrfInfZZxFZpu6vhsU3VysmhziPKSMffCufZdgJJOecbvmvBGSF7V7uM0/z
ud3izzyfR5hVmLQN3TXjwprT/GG5QwMbc9uB2E3Zh8FCuxFlgq+tIt/XZU2tFN+7rVKDghywpZYK
MMB2MY3jK0WKymxxHySTA0B8Obf3Kk8n/aUmZhO+PzBsnlqooGFtpYxRaAQVQj3H+Hyfon3JDcNH
/7gB3QyDD2v3wje94nfZQP79OJwWndfzpO7Wv+wJ+QQTCPAeXSylIG+5WVPGZEJIi9ZbzD/kHZsx
pqyqLCPKOVg17khxuaOphtpm01U37mV1sf4NamDG2S6pxLjoFDhC8jabGcNioNVI37mqdsSbxipK
QUbnnzqTbmNbIFDOYZEgBMycuP9wLLI2zMcJcL2jtf7MQoxlL7ezdk+BDBdpbOFVNp3Nf8FaJd9T
Y9+goyHndkRl5eQZkdmWkQbUIQRC7P5hGgPw5draYhoZeEx1oXmeMVV6EGkvRDb4WXGiRd3rbxFH
RVhwSXmUJbYZVaGwvpFCKfTW5TId1E8pJ84wbFUPfwk8H24N4CPKDSnYLeh4RKTSTDm4QTtbWa8c
QSNhNiO6qlnlTDK5TN4IagoNu7RsGwCNsYK1WLIeK0kS1BL4v3kSZgxhDE+SDOmH0Q5GJzobYT5S
0Vguqn9jTst0om52pIRgfxn8W9LmgDzY0mZlJNkPMjnOEzpMucpIocuesepyEZqYny9sEKjk/ex0
CoXROMG/jMso56JaT31PTbCs3LIM0iINuoe4aTmFS8+OSc1UohGZ0aGQ/R3YLFEbaxred8b6H65y
Tg0iWRLWzQuv5+uepyBJJkYHom5nUP+8uusImznGPT5fsZQAlhl6nC0Fv0F5A9Rbf52k0yOKsYGa
uCVZPNKLSCVqKP0iE5tblAo1svZ5FIcXqWmrGtfW21G8lzWZPemN5MaK6wnPSTMIoZrp+13wiZif
xk94z6cr9V4/qHfH80cdpfqqPEYIGM7c2R+qvUwl+M6VlqGUxjNPG6sCclPD+yU7RZib/nxRsFlA
/DbLxlkHvHtjpLnqfav5Jldgo6P9uTwEFMCOHf8K85omZih9XphI8FuiE6OAO6spbo1nAj/8iEwM
/KDvnBQIHyj40CqW+k43DKyZM3aL/IJzRtGcosqntQzDRkxxQMp0veXzdB7SqPooeum6nSvjvAVy
VBLNVFvh1gwKze3mEkTdlQ5Y8nhOPfXUl5mIDGZtIHwLEPPWza/z4Tt2GGpF2RL5guAU04Bgl00I
M+Ftrg/FnEzsPuwkWGAUXOMQfdXWqxwdUt133wFCCFKkSqzezVkBIvHWPwHfLPgRoXtGPKqGFXq+
EKllY62n+WEIcxXRY7I69cnoXx6AuWhXkfb3Ec5Wvn+PdTs6Dmv8acd9GfWqMNiQH8YzEpmk7RQj
T6Zkpfdqtv2KzoWUq+7bcJcJleV79KnNmf4a1wtuAEJYFNie32k4I8T4tFfUkbQ2UNRPck8blEch
aN81jRKB1f2xZS3uRD3LYo+0UhmFSqFSpE75zBmY6YgBRw3YX+UAfskYgsvJvNJorR1WVBnvzAyl
2ObhiFMskbj/Aj7pGNgC3lrI2p8nILTE9GDuhK/lIugTXqI+jAm4ofhH2pVuA/l4BzdwlOR4eudN
/SrPVgUdB0wYLY/gISam4UBEzCmhIPD+IxduVTPp2tooZfGThCmSyMl43jgo7c/BAFAM1bsCvoZj
Gelc3K1DOpnFlSBIiEv1Q84mq+3/7Zi2hhikx9189jJgyPu5ms1kZ/L/diX0am94MixVtM98BaOL
Vkf2lbH0xc6K51BW59vinyzpD2GAFpd5WV8XwfchzcPzjdlyHJjunCHdHIoDaLppogXUKr8c++p8
ZmrUII8Ne5ou9qvyHcNpUCdGONYlLFcYzIvyiEs3P2dcdcQ73F6PBkXOc3USr8rOomkKhjC4uCc9
8Bp0q8tA7dX8P1nD95vcIMrglqGfJNiopIUu/7TLlI8qhSZVWS9XIJa8BiyOHx5xl/1PEesPgsi5
q+rN/CxnMyMQWStALauSp4j23pHXGEn1DWR+iNxklx1SCcvUG6Age7yFHeipaiqv9iMbk8VmaDyP
Y3h9M6+kzOmPtUbD0SPUb1tL+nRNYr38kv4Pxb66rXKFkeYRS3cXAm3CaF/JcY9ZdS8mhT7hh+rO
fYHfAN4ci+21YTxRt6AargH7KjpNNIjXKuOR7OKg6rLxfC4ti/nSBP32Tt9gDX1r+TpeiAEPiTEm
FTqxh+kGRaGZZdso4LsEhjIoa8zK8dJDATbd/lYEThE9KUAvKfc2EPPRq++MG94jgcHpjG3HEPIW
DN5q5DL84sUacJbOxhjz5dcZrn07H8pnI0H/P6Km1cb0DuX30i+KU+mtSLtFpqYVVMBY/ekDchsW
rBqODDW864oXiII8T7NW646UpVTCLStx5T0sTHDlvUZSd+/AGaOhSmVqlZKB+b302leNwiAeL4FY
c5VhUVEwwl5upi+SRS6efkKUNQyKGtsYHoLdEYxu6WUVa43SCLaFFCuPGfvnTl7PnrDp9lnSt3VE
QjOuG4SWRcPHu7TLgKbbs80RdbgSI4iQl7dX9CMY81lBR7+LLQG6qLItdjt46y7WUwRpUoRYc1Xo
SFf9y5Wzex0M1wXkHuxjIDGS/xXf/yjVdgvyFggGWFLJRjyiVlwqjmBYC8G2NUt8NzjruQpWrJPK
l8vYio3MZqUQuMoJI6tSmeVqVuvgrJFGSB1U+hVfmB72nTPdp/Hdc810PntPwWxE0RkDz2Yr4XE1
dcFKMtB5lKCOq+dnALbPPt4wEamFYtmlaCxcvkCue0RocU3rm/NnMPcOdk8EoiLSYh1rNqRXfKC4
WTo35CD+bEEFp/hZSXNzOrtColv84oy46AcLQatd1S3+Vt7s01JDFtfR18LtObew9S7KhRkTkG+j
Lkh5JSV7BzpFuUdvf3+9AU6T13OtFtmeeYY8o6tZqaAstpuudx3sW7r3LUnr+ECnTRz+vDdU8KjO
RKPNwcmemVNcoMM3+e73NszdMd2ELpUJpG5qhzGYfZfwV38IvZKdbVZYmDYuR9BvmaVI55y4ePX7
7MTzBlY20DgI+/DU+zI+X7CwjbF4bYfvJADKNbtMhFyiz7ybLSjoZrteHOCmQaumI4BSZbSd6b6Y
Ezdn+SSscYK7pvyGNzHmanQhHuJeo1Kg1xjI95jYgl+dmjw/Iq1b2zICj7PQJjYd/+0eeJ5dNlyq
5LHpKuHuTa+RzRxGJ1s3uO74J+tf8HH8cWiv5Hwz9Lm9ZNHKWtxrxZU/6pgRpymieH92jBXO8Iyw
Kc4tdnsMEqsFoqPUfjJo0h/PO0Gq/Ccpjhl4GQtr/cLI/IQMi7FQnritMsWEBB2qEaflAchR9t2l
BLFRp6BZq8QfW0Bk11cIO3mXL3YgUgc8tTU+SiDeaaTGZ/iLPq4WNhRYTmKiWmuj0wyUqy2DqCK8
tjuS1qCjncDyf0nzdag5KaZPJt5PwbjdPrRI2419jKdSchgaoPwHq2Jlr+Y2V7GryYAjuuVNAFRP
ZaahQAlAipEBy+swUwkGfkEIlvkahuspxSigo2iJqjmRSdcPrNMGRxTMNES6GXLygVPV25dGzrVK
KKLL76dhkoo73Ak6XOwLqyIP5hF2e7UdF9+Wvbi1WDKvo9Q4r3IvbW123VFPvtmDEEML2ZNlcE0m
a7s94rbsyUyaCK7Bc3NmtsuKxKnZuBX+jyT3jSZm2oc1ahooX8bWn4nBYELi3KEcdNixSEhEUplq
lgRmEl+grwYAJv5KbLw7lcorCGgluLHd6w6MtV6m4gb/g8Yw3NbqwSJsIyqGiVMVYx/LJglSIK6v
4+VHZwV4Qhb1eFjmD33fVu+1YUjqf87CHBJ42OTgNWYhHvz3d/vrRZfL+fAkiMlslkag5H+GuXc9
ANBHAxbBCUMUU5EiQcW5l7wQ7UMx+xwijVTd+koJ3pBcJWKMuyBwIM7fM7EpL3xnuOXLSsAF9RQr
Lb+8DLJmCnk4fGZMBmWthX/VVjkeDD+Z+G/gMcTRMGhy6QBdDIMn3U8UnFwnTTGjtk0DUYuO/wBL
54YM2TOuilbaIYqJ/J77ZYFXheQHprKJYdPUN3QfZWxtGT0kpX8zCqf9GRpHL9aDArA5UIiUItue
paU+6bZebr67LYO7UkQFIUQWyCJWXN2ILkYHjXtnMWglwX2wwqggDTjPZnV5im3pq62pIbPfGDzD
hMYF6wUQCFGzwDbcrzu3g11S60mI/rIMsd7QdoiS2XgBt3kyoa4pIluKb/MH7UaPQSzaGN2IJPy1
+1kF+aM/LE7u4kTcxCuyzTlg7EKkVpBKLBUpWaAlHYMMJ3VEtSbP/kPj2ccikDtoziDcUFe7Jp8C
4FbNMb6bBrkH5gWMNAsXNDKNi8cMHFnRb9Q0I3eoBm9nIoq9O4dr+7Ltz7DneAGu788kCbBK8pHX
cvtm+GxlrnnekPiETe8IT3HKFvPSLUmwBWOWl7dL8UEDgwqGpXZmdDt7n4ARvRmcHBAwZl8CJObe
qfcb9jgb9SnKgpumNARfbaujFCgdbBBJQ5zCmLOHjR2nTf1i6KKInLhAqv7t01GC5ZyiVha9HqoJ
OhSDdplrPkzH4fq0pomT7fOERx8HCoQTHL6l1J1B7EUOIaS3xwBpdrB8dWgoS8pi8pagTsdYbiwe
nOmY3RSLT30Pzum83fJPZpFSG7okyiw7mdb5dAEaSLCzb11zQxf0uHvPXqXo7nvY9mpgg+60GAXh
QxwXK/12LmKt2hLjRrGutd6FvD404QtJZdqf8s6nHIYLK/UrbbHQlZ5ll9foATePoSXKLw9/QT11
kOE2qKYYQjVEB9Env/lJrDCDuO5KncgZVHoCMFl2SW3AP8Ce7X3SxFIexM2un7yTdQ/5KK34iKGA
Jg32JM5jsQtfzWA636RLDu0B6Hug++jUnuib3IyWN9xztQisiXt0p6L/NvRYpIiX6Hlwpd67HuDq
kfmtPIiO72XVdqViOA9NJZgxD4UI7FQkCUhm8kOAoRwZsIU1KySQqZR/NyIu2CxMtlhp74QgO49+
mBIDB2OVkYIxrVpzlWzEFHo4AYMyzkmdruCVJeXyjhx7iLbu26bvjYvjDvmhOx10AJZjU4LuJDLL
Kfz056GacbOOnYwR3I0eOmuqks3vrEOyJm9w9jLAFej89NonaT5Kqm/boewbgjoOEzKuSdhhQibP
uRJjSpB4SB7zObA9Ea1rfVw1n+RaplRjGOZAmyMT12Wx4UoBGaAGNvBnL08C/46htsxGNItR/aW4
zMuixQHL7GJdj+zUCyS9C7wumfratgY4oM3JEEaAP/S4hFG7SCuXGygyRGUV1m1X7iNKclsWGbEU
+8QQyHev0gLsjiDAPxyCAImo0au35I3VRBNxFR6vzjTNLrHfe6148v1n5vhG7e4JdvanuEgPiQAB
bSwTgUOARAAs9a71YRs2Ffa5MvbtO+7mKc1u+AOkKrieOAShHX89sMIeGnANh74khMpVhLYD3xi+
m0NEajnuN9oRDC7VDV/rx2wmAvpmdh3pTFSk1KclJD7CebzdD1w0ePAzWRY3v6cYDOnBZ0WksMxP
rx13RFu4XEoMByFrcIA6ZXmcijDFvQhiNF4+QZpefUnzFx0KeM1Pr8T8D3p+RhytKDtJQsNkYn4J
wHle/+5wKxAv344a7DeVnn4drQZHJeGQi+y2+xSwlv66FmV4SShpMcuSraYKt/GHXt51f/v3Bps+
yrOycl4UWiFtGHm02PaXrDlk36xBrO8qBnIWd/HFy3ibl9m2YW7sy2+8zA+0GPpww3Rmz/k0wqD0
zZMcJeLKFggUFOZtG4IRwxy1lSF+wuoXlwVwz5maBTE+M/E+8KczLIeBt1g0gBW6eAx6O+2+dZdG
VMvx2JKIv9qVHmk7gM7v0ODLcfxOauoQs0nQGNxWwgKmYAMnS1Dv8GhCnzzulvNotUFDOI34vWIc
W9yD9MzSDpnw2BYB+7yiWSvIsIqi2Tn1BZ9DgPtGwhCa8H4EbLIpwoH1aR5NgAvpJNBvPmBDaV5g
P1UnPb4vjkoi5g0KssZN2y55HWH0e5xfDMrUrgDOvoI1CrVfBYa9spd4GDN4yQy1t1vSP8Yk0mxt
vZEQG5Q2ykJmEi0gOp5J/FgL0d07F4ePO8SLOI1sH0DURKFO+cOzE9AlwWNm5so2ulIuZ1dCmE0c
bYFfSxRxrKW98EEjG7Xp7tWeyExSumUYQgRzb2Ikhge4LMQMCUOswmLdKhw7OygkdPkLG7x+ge+F
hPcqTCRKGAEhJsZ7692PagxftDRZ/P/sy2SbaHE2MRSOVa/QZnWy4DkpZMLl0RJB/ftWXC7o3aKu
0sP6+D0VviEe17XEa83zZoNaWwYDOtrPREpo/lX8t391Ql+Nc5N/U08kCZpNsgw5Jhp5z+J4lHIK
RDKJJEHuASdHFtYccoZvdjlRv5M3ueby8Ew1yRoGprIUmH+djPURITEMGSStl3E5uxCKMYKBFJWi
hlYDpdExIVveBK8qw2P6JvEqBLb8DI5JDz08LUQM2oygjYsAB3AP+mvAlbqkY+0rem/wOjJOiQCp
Tu54kz/HM5yMYSWeVkgKB5RYKxvyUaB+xZEdoUlmMzQPOFmuYe6hxpI7rNQZ31peMnjhWfDf0c89
4YwSkde7YGk4fsWu1TmYkaDgwEI96/2SLN5aoFq10N81YFJzcsx7e6a36gXBP47IGOfO6+XibzRB
woWbmXFmV4Eh0Zy5SzjyPOyVHetN1qEC4Cjxsv41+XO68cnFMHE+8L8nkHq1J8MmDg+pb2DCZYBq
O9LeWli4QSrlFf/GhllamQX7hEXvaXE1072J0J9KIGYHDjGHDq7aR5kAxTMUa4/MfH3cOe+G8oaJ
lZcYr+N3YSjCrtxp1TffEG+5jBfCBPIiooz90Yb3KDG3PsExiJme/0ATXbNKaM+SFliOIllkp9YA
s5Mv4zDkauGCOH0sZN3WrzIAGsmWZ3MCqBE2iZfnMFkqUJrSpZQD6U0IDZiGaKRWReLSuUnNXMo1
3bvuDB/mqtd0EBd4SFWx7Gux0Woc7CV54SekXMxZGA66sCsHmUuaHp22I/aIvLbfkZQ/j97aH1DL
g1OKj8o2E9jeMessh1E3Po9xdFor2NbKYe8+e863t3ljY3J3+MuFWOwuM1xBq5/DHrwlFtML87wn
Y1aC13Brf8cTuYoe/iYHXtabvmSDB99DN5p5rSmrFevsufTABfAvTAtrkXuXU8VbHwuuGj0Jn8RK
fkogMY7qmfIs2K7+U5xAb8X0+9hW0d1LLqVn4FT21VWwnHYqv3IsTdQoG5bQNSHAsvck7E7hFtvv
gXT7RZw3S0ijo2M2/UMppVWz9XVErPgCUMUSQiS/0r34sKuKIYRcjBhxTjJQvEeA0VzOSrkufvmv
dEbD1EvNt0aihbGl6j6aPvuQUPjC/z5qJ5vNqaftviT5MFLpo/3ShxGY/CFTXdnzIlVlvldSy1Sf
pDH1+m0y2vzz0Y+MdLLPXN/bVS1uD4hB1sBFWG8BltTa6bhl+ptagFgpgHLkRaoSrXaq0yq2vFpi
lZAJb4CNNnigQic92v9uPDXMEivjxgXpbbt9ruLOwqJU44RP9Wt6g/h45ZFMXH2RNkiWVpTh7mW2
WjyjDHULzpKiJzU/iz8broxj7FwIo/n19/Y6OtcABTNxDwL4hW8aXQH+bNyUtiwx2UQmO14XwcKa
oJ5q2BLBVhhIJSCzy3dLYAS0IqbXqy4e0DTVvU4JQ/zXfl9C7iOs3ygTPY3KHr4tN3M8Gjhh/Igg
bEfOcnJRhZ/8E5CCCKOnp82LX78gv612S2lhRI1sfgh+TTnyI2MHFJJgFmGhaBs/vJ2CZZ3ZzOJK
rvrf5sWUR/kS2rD7KKFdqRMWQpuzOkjmezwLItrUj/9Q5xcAKmkgYzUKIfjDPrBTAabLhNdcC3I7
HN7goH8Szj83y4YY1CLEyeoOXXErGcdm/ErlK4ZzNjVK50Nbf/Gfpra+ZuU/jlxBJ3AKMRU+0MsG
BSkH8VAMS2TPATrXWf8DCfK+JrErH3wQakkJm7HuVCFpr5QRuPaXNvIWGFtyhRZwjWKQvg67k1Uu
Lp6STgP2V0NI2DsrOa+xg0p1JQ+GN+JM/Akn5ydr07TF3A8T9LKQ5hldsF67kqJVAg0U8KBiw15v
5KDOR4GjRvQPaJ+Hv7EWmCHZMXJwfqMwYVcvZ2El4kq1pB1U8AtQ7Z3xoBawmKQhj48pEq++xOZb
oW4jlPYDxO0YfRFW1P4IeWcA25udqS/oWQTW6enuUwyScSt7nRd3tw2MhwkSefU4+92CFer9izsy
Y/yebIX9DKD2FtqEiRqFIzta5sTSh4Kju8rnsHIlwitGYG4YytE7xRXbaZg+sLOvaEoAkqlW4dSk
hjjFPB7wL5c69PxAtJIOx1XgMV1o9u6bGInZObuz28mlhg/h6cqMNFerZveUD4RHxdhOpmFFWVGT
atO61p/wsLOX4iXkyhe2ZsIk0IkrafbjWLxPl9HFokRM4wM4PR3A+Dbp34CQHUR7UUQHRfDOsI+J
YdA46Bl9bSc86skP8JeE4fka6nfy0x4WREcbxUbWZAsdyTBpxJchXz5/ku3O38ZEFy148RxjEYP1
t2LRXyePyiW09Ibs8A4qnmVNIK6+GMKY4/kp4qw3FXY2dlbF8XuBxfIBMxxGwqyuHXCrlOv4DPa8
UmKlxzJVDIsZqBFpaHMtIMcOE+2ypav6CqgPl2ITGiqcgOcsmcKpsUJp6hbPDfC4MmKiTakeEGtD
bzXhj+JjaJRCll7JCMNbWf0vU2FlqxBiTw96QvVsenreXiuiv3n0EJgyzcXyNQfBn66NKKuhBW+X
7Hmb9qs/cic2h4oX9eB9SFr84d9OBDnAo3uRYdRiVrMNCplyb1ioKuT/4rZkV2C+jwww7G29leFz
Aw04d3gZczbTvZMwzd9MvwTw4ox7wrXZ92DCiImttbD+L3zXcxtVcBhsOnWhydPs8mgMSnw9XrGb
rqvLLY+pfIjZ3abr0RnOyda7Zd6FHSvyfR8Ii/xClKKBz3F+y6h7TYOLw6fgGEHefu2xPAYuPsQm
bJoKr+VbjyxzGtcGuTECuIDcmEumXCXmmhz7gCiREoAHpq9kQltCNJZNn0L31sdyTD1Q+NeQsnOb
/wyGmktVDpFXKiij7p38mphLOtZsoY5OMkMSGFNaWAmBZ5aQYCeX9+1qE6D5DV8xmasWEpvdSvVy
1aiMS2b9OkJNYRu0MlfWWi70+h8jLCcWexVTwBORUPSogZZl7uQSY+ZqT806o2COcJpMcPAhz1NK
Sw8kSf7gHndMxgx1wo1TjLnEfJxmauenwod8r0MQRcem91GnrnBix61DFTJyE8hrMaMHX8Tfd/GS
PBSaObP7ez49AcSvEPLSm98S1nB9hUnHsDvUyIfoKghpj3cOAjRCE7SIYlM4djfBo3kJYCLB3dQU
hasDq1jpZD9qgWRaPKHqVVJxg4dVxaSUhyimjdclPB2vOkxfq6mITOKh3ID+8Bp4/REFBEoF2Hsp
BOO32ipCgpxQBKYW5endf8uJv4xWlfC+/OiTUsBuKk5qzP2qlVY5MdO+9XMI610VaSJwGG3WrhxL
mONx/ySskodUludAL3GeU5OtECBs22qLKxJ4KQ9HfdjdFsU2GlTxBlNDjVMUqFMN3kr+9JPelDOt
ASHZyQcfH1oGIa3E/+w+3WeCPvFNnvCLDFUfn9oEr+niF2bttXU6eIOjkC9jMUo4tNS3wFp3eTqB
5AP6nk/GFSew9boIQO91u6FjSNVujaVDopf1xy6qUfx8VM1FcnpsS6VwnxCPe+NfznA2i4fXSWtO
oWR+/S6o3r6//1QJUaXALCzEqzSglg4X+CwBlzNES0lzpQq49YSoKLT3dh0FQktdsFBnHuiCSSQZ
BY0X5/gMOSfphefglFGSuRfiMZ1yy0rM11eGdFIDt4uU33ucwPWjpveMlH56xiGaEMdfY3VNNRZR
iSI/AUqvgLiU4n3MjlznpfH2/BwBFmFyocccO+A/bhkY3+vkfSDZB4WTH0VdhaqdV3p/Yoi3bABN
nF5GhnoLlKGv5FDlzxPA9UZld4LV7sJmBJWSMu5inohqNOVa8XTSQwX2/AlcWfCyj0T7YiNrMtup
isKBP5IC2pvhUeDjfejOC16pjZ7Fwrxp0tRRGJEqIG8klstwYkrIVhdeL+Z6riqcEFa335hL/eZd
XU+0t3/NPJQD1u50dZy+FFZf1cYUuSeLLh2ES3BnRQNgZsLor+KFai8oPEUvO0IaudfE4ChF/Z4F
i4ItRcSnBIHOt78DvHZIh2mTvhJhCMw0u8WCVeFSBtyOOib9BmaAI/R+FibfLpFWNW9bKi8v2nnU
kE7sYl/7rYp5t6uj6flGdFNG1G8kOkhMRZehXOyXayM2f/nNsZfX1NfWWqN+F/g+Uq+ZDx0c3r8/
TcWv2s9KAffsWcPZ+VX/6rHjw43z7OoUluDAg1LE5VCWBBaVW95gvKzLnvxzgyomCphGZh6nCOp4
sccJG0Zq95yTvLuEskpIu+R6n7FdRDUs8dO7RZeF7XnRB44kaIEAMM6TjMXKn7mEaw2NkFlVugYY
+hWlrShNoafUPCJ5+1fnu5iWm3in5W9bmdmLiO+PGdhmK7RYR2M0EdoJoYyNHm10mcimifQ3a4lJ
1OnvkbSbl/CHZ7O+BiH1D0pOKzF38iUW52sBDdQ6BtwzlsTdc4FFErB2VJ940F6c1lTNYag8pR6H
m+5J4vdbbH3usQb7QNCmsoQbIQG9agrohTnmfS2ZXbLsWLYyNiDTu8YwydiI4JTYT95O4yt93Y+9
RecPVXVE9cBOSockh3XqjQcx+PI33NIu2XB65VGryJJLbipfEdhJrE/kau5m8yi8g8xPvNxrFLLW
X7dexna4uuxoENVS/BDfk+V6o9GWuznrdVMuUbu2eUGpVTthITkXEz/ptUAXwODGlzeUnjQRIGAG
M0CFM0AmgdWj8aS2h8C+IBP9hzgGpR6FpRAamZINRlGJhglLaEV78xkXGeq5MgR3/jn/EOAVAY7J
FcG/jhPPiQdwlnYNekrs2BjWPifFAskUfEirG15iSinbHfntqcDTEq99LmwcKWyOMhwhudjjVzm4
3PaR8WRWebqb7LPJnAbObuPAZNIq2Ksdl9vxS/wI4em8vKrXNe8rWZywJ+4CPo1s+cdEkWW4MDog
pw0E7daev9wq+Zmu7HS94IfFhwJqgtyiWxlCuOIxDMZsrHYRLllFPNDNPjxxcW9eUJzjauzTETd2
o4SWWstt0xrX8GZE4z+LiAV2KY7JqY5K7RZBnNhkUXs79eiUoVcjTKRRDwXujqt2w4ztgl0k/w5k
rBkDRXrX+2EwSvcahHLVTeKTK0P9f3TzrRI3J5WkfBrP7S8EJ6QCl9GG3JOv+kUNDYynZ2x1buGX
Y69CeZ4s7rbHuOLRPa1REYfwfbDM50LnGyCm/FryyDGQxpasep0Ed/TI2wjWaHC3tdKe5mIKgWYN
FjdBs7ZBeQgB9u8dR79Uio3Sv7qXzhhUptDqccW+qNnP9IlfIpJ8Ga93uzCYKgLmLwbPP0g5maiU
fkl0ot9hq0vnVzkGpI6x5qJQ/Lti17EniHyEdyhDQXrOt/S6Iy6XGJkY5GqP+FuPqKxyX9UjCA/V
MFbBmyB/qR9j2OTBzNuuWRxyocea3U07IXs0rHfWHlaJn8SYw9dsUf3NZBENrIKKoUYsreyknkdI
TC1fXqjezQHreiqbBfB5km7X11c2vYsAgWPPDfapciuMaIKCXb9YvYUvV09SUhCLy9mMt+ogpe4e
NtNNfS37qqjcbjh7/GPg++oTJjOmJWujoh8lYQbTdYIYmy6tnxw3CX3/Yr2kiLwquco11UhoqTq4
1GYIHcTbVzQDd5ZH9Od6tv3nS8hlABBCK/pe/4pXiBJ3Q6Qs5pJ6X7eJnneUlHU0mu9Rvmns1ed9
vS+a3JorBO0YNdHgI/j0g6ZWE7bedAWGS/3pi6VbBZIx30fLC9FDcYavcSB8XYAzXP//a6i6p+th
AV0zpu9WCPi064rORtV7sy1bEAhTzg2I/FwfsYQwmj/63dRA9Jh2Gtm/Z0C9JNskeSzqwR4itQuk
JJmt0wCk8VuJxnIPxDxGwnRUWH7SGp54G7WNJ2/TCSeKGBBFUGJbPhDcStma23KNaIVvBSPQIdkM
MUtmbZhHOmKLK5YeFBQgIhn5wlhzQlZArLSQdtIpTrg8Dx5/ki6QlVpoCvV3Pu45/d5c9D9/4DV0
p8Em2Zl2RZuneXpwp9XZ0MTUqZt0PDM7eqpdlkoWR3f90HT8BLOvPChX7NdJgUSAZf82INGYZ4o9
MvmQiDFPA/dlM9nMkj1O7nR5iduYaJwU4v73SsmQ91D57dOVBBv5E+0+mc9PTe8b/Kb0hTE5n6JW
h7ILlK+RcDsipbCyIk0ghz/nKeuI76V3bGKiO1Nr5LZRJhpQZSAg1I5ocynWtoPCAr9ZqaHkogE/
J5M7EU871wfozhxLggGJHEoGRASWO6vUKpR/G1eI0h3c2pcmXRHtQedJsViqjuFpxr21YDTRd/I9
FtYsqhsOT7CNDpbOn2wo5lXIIijqPkCSrPS9qkP2rWi6r5yh824FsIR24UOEPcZu0tfJhx6ZATKh
Y1fYedEQbFmKdmBjg8R8KzfS7drp+yCaEHNnZQmDNvsp4dXIVe9vRcFOeifzVytg0nB3WjKu9yYt
C47DVytZL8NFzBTez+qCjWTR0/+bfSPaSGLHBHs6Rh/0XuYjfQ9IQPn2Bhtg1NvSM50L4LB8K9iL
aC5Eq9pEhUOxhrqyXWuAVw5/XGMrLy5/8m28yPQ90X3O7tWicPBL96BW8ovEhH3xCDww2pET60rj
OoqJqOnzGE5dnDBzB4dLVqH/Q4E/PgGDEVMv3UzFFZ3kEAFUTHWgQhvr0CnxUPK0VNul0CtWJAdh
FTW85YFI/DTch9uAArPQfx0XrQ7fVr26bGBOXb+MZ9nPRIzfBc5Psp47oA5p5IawTpSMdoc5bgYK
xi1gKZSbL4+/2cy9gRs8uR2S79HCwKAr1WwJ2Dh4ISSf1I25k5njsFTdeADwlLKdc4w/e3Y3Jg8y
KsjGoWl+YmnXdZXrAnFk54fAdD2nAWll5u2gEW/SFKeg/MZv9+SSfQnMxTSkk8BAs5QPsThF1KM5
RVd1ZNAgHDwjzv8MfxWLE94ciPv2hjhdTFe3zuyGo4MHiiYT17EjrP4y5nDQlCDU3PfpYHRDosmy
rSTePvzw/u0JT7XNp1ynLinvuljbx7OJZ4Nf+u6SLGfuw33IFiyJL4hP3zFDa+zG4xsXZCo3pln/
v8wyatLy45hjsSumSYxgrVA/YuP00090rul7BRMBtUA5omeqBHSltLD7Wo/trFxhkwokGct67lh7
3F8ZYQPP1DHTfziR8wqAzYbaEqoYG9Yq754OhiGsA5hRYZolJuwXZpVIMSWK3e57YNnjkWfwMG1d
XB7ccQ0YXLyU/sCeIxwHRvoJ/E6BfeUstUgUUsE+y7rf0KMS/steevXUuRJVNu4QsW/QH6q72qg4
JRjTJaAbs5p+7OMdvblXt83qYv7aPGgSjrXF7mPIFXxPkzdlsc5AF5jiPjoPqvYXAlQafKlZ++d9
M3kplxuL8Mo3+grl9Li8T9DSBBjB8SQ41htyM4cHfJrh/4JkPjdYP7x0iAYsaSAIDovzGitUysCD
hTGk5aWs55XrqfQJpdwZvu10hSV9/W9Zh/KQqSeCl6WZsyb84pooE0A7aFWbNFBC42B5/lOS2ITv
Pfn++8oiWjXD5xRJlv+CWQS8Mf6fPaa4VgNzxqJJolEICzY0oaxMEX1LUV3Fs3bJHtvL7+9Z9yIf
Zh/2AF4c1a5Z7+PrlEH9I/OpUazFXt0A6SJU27rZwHu1/RXuXxToWuz/AhmYmV9eyARKIb3CRZn/
3xIjrWc29zVbH80TVUCv/OXR8VxErwBL4DnGKswzSkR6oZ8q+igZi/eVcS5GA+c8zzJ8kKnfvv2i
JxiD5OdbG+HHb9IxEyUz8SbeYn9daD8Ja3oV9BD12/5sAYIYrj+WnA8YdL2T3ZCx2Pqq4R7BCrEP
mBV2VG8BNhggAQASWs2jGftw19VUi3rUvFtylR7nHHvfqjT5M1Yeqa/aMOT47I3f/t7vz/gWJ0wQ
Iwu/XrNhl8ujw2IGqJM8EnkpwxtOOtAhCzmywLzdK0o26EgosD9xVOP5bQtIplQDMElp+rvxiQas
7wg3WeCXJmIeMaQ2Y2JfCklx+eZX2Y+99g4GelN/+UBnUkysfi3NjWDfMptz79F9o7xb10o3ZW4U
r6g9NrhjROtF14hpls3xU2r5IrKjUCF+ItS19pk3FSpZLRWAPrxnvUBQf7keVk/JQkyQtteQt+54
Nkl1I4cqECrfjnQjhyZQNnXGJb1Cm7EhNddLv+c29xVui7RUZwf2xulQJ5FSmYSOQOgFSA99DNBK
q0zJz5jhVEWap3MzLMBjiuvwbawHUTv4+OCkmnrKtLJZEU6US9sk4hb+GDYCtF5kBoonbCVN0Wan
v2m4DRsaLGJnyTtxWmu3AbGhhv6YAR9OHR6HzOuoKZYLIjJrgNqTF10OXn0pSjhl4IYyibrzm7LI
4bsPliHIu/RPi9C8qPw8t72rsZ+agvaNopIL00Z4Zyr/1j/V3GFPVIDPzo1Hrfz+3J5kcZXfjejT
R/qvcV1T7+XhR4XYiHM7PKpAvj11L+ucvTew57TUjoYiA4PBLEcpacMyPidR/TcLZXMbnjsxGqMu
sKvA1DP/6aTieRK2CKMdb2qbZ13yKnQcQZ41HHsmDBIiT39TJ2idtKDutxQYr6EnL/8AvXO2otfZ
3dwUm/eQchf7SUuQH/Yv0MQkiyUAnCPr/QyiOM4NsaSh+0dQ4Ww5pE5QtqwASmj1rwHdGthrcusu
BQyOaVobgfxl4d5vr7kh6wJhcSFCmYLoluABT4obAZbz3pGoFmDLz218D0keTKTM9YemwpAxpDiW
6K944zDNp1d2RGedPBF4cyx4UX1Y6PANpkSaGc2ZAARwXTOUlDaw6BQOcKndVLcL2smHv9zr2PwY
JHGlvlpV6kR4vUaCygJyODWEBxsBzyq5siG396IdXBt+loe5KmCAc2eooJs36WLrcZC3mV5rPGZT
Gy4pRwKHnVjkXUfC3GTz8N+yE5OXsvQ6yLG4EAzbgfuCwfD49jVfyH0p9VdE8EOKscUxDyCj9aHA
s3IE6Dg5v+Dd+JqgVP138x3E0HQuguzVGsvmMK/edCwbAuxmYZ/iBVyTSLipR601GMYqHK8WfzUc
6wwyixjSUD8sM7HhOAXXSOzVeoy11vfPMDlOOErfRPNtJs1uiq8BKqmuwrrkZLHv0ki9NtGsroe8
ObzW1fzGWEnK1AlSJFhbDVYrv3KCl4jj1Be+ZGsKO9a1UfLfAqHY7B8fdBCB4BCBnjnQa8c+HRR0
Dott1UJJfr7QvjqUZKMyTn6uQpjlcSiAiTgdrwHrJDQUkVUiEUJeCvNKQPIaPu10eRVbCEBbQt/V
7XH5b9x1RPY8sUiWD4faGMc4ouXNCBJueLU6XAr/6aEGjPcmkT1Phbu5bCHvX9QA/Zx9Z+HGoWDC
TqlpfVcjMdko8T8sHLksrRkgiQbv+QtCpcqrTj9FiycYKwNXrgzCZ8Ph29ByOYUwyru0wjUPhZdz
ouhYVvpWNiOiN1kobMtEKFrcRYev7d2kd/zyxQDasZXs8Pps/P9d3EvOBpWcz8slmqTQnOVjfWGE
1Vx4/9rUoeyEfSgnm5RGGCCDAbG2aRC4Vg8BvDWFJK66YLB79UDiByOOksgtwDroTG30btmi3JP4
6QWJo/xSu6yNKpJyLZ4yNeB8j6lQJrvhwNX4gBjrQx5KfAcfRtDW68XgdvBSJ8XAiP+TEnKTwesN
ZJGTsSpQ0fnn+zvwpsi5f2WsARY53X+Z8TcBOljjdPLPdaGBqGwfAmFkCjhCut99g6S1+9hZiInK
HmWWpgfhBeo6hFeeoXgcqtsV2o91bt7obYnhxk2TagWJ6/e5CWBkoB71BB3mXx6wshnIM1w1Z+ym
6C7zw5tpB31gZqolahFntASud9XV7P88G/2yY2ve5OQ7GCMire17atJYZFoNuLp4z2+ygm7cdu60
u3t+j44ZnJAgefdDW5wtPFgAuAPlOyTQOQizCJcbQVdmy4/8WTXEPIDrNjsGmFUkMuAp4NNk5mJo
FI8br4IqIVsi1rwmNbYkmr+sMGwUAOLPasGXp6gkUo4SY1T2tYZcnxu1zepFZwGPHcfhmGJZEvv7
aoCQEuqk2RVKvIAQ5D64XkNhO8rNg/RNZ9EB0ofzzbILXiN/6qiKaIaiu6G7xrULw1LKJ/ha4rmu
TcQNCvOnXBeXmRTbzChqS2Go+CIbX0pe9gCSQerBJNaS0xEILzLuFr7PpqmMGlpVlAKEnW4hKb+y
sV/7pNkRTPjggkkZaN5YqelHHCkdX6CnZ5PN4UDqdJHtqzSIUvbfKAZghYtHP6inJwMr1L8OrLR3
ugbcDOy3XM/8+we1BUYh3xj4RlBE6IhSwJ8YhKN+qAnzqtqQr1OnQf/kE3FbIBB2Ft5O8Pp2AtP+
xVI1sfazXOypEG0D9KCu0JAvSGTkhVmVnsRnOvv6oL6Bs7ZIe+UQ9nHj1N8pSIEaGRScX9QrZN+j
fEnjISk5kHdyJ7yj6PuXHvGM4Fy7c5+SJqYiPb72QrC04mX2sXEXRaJn4063RArhC4f2E+6x79F4
Jb7W+ziPUHYBxONLgsIzkkCdzJ8udbl1Wa1+fUesOL8rb0dAnGsiCSRrG/Ti5QW2Vn/ndL/i8CKU
C0k0tE51qL/5vOyjcY80lhWY8VpTI/pDwcuH0yXCxSdoCg4+v5wQWHBiyMug0vF0iPZQhKmx3Z3v
TQ6Uo3ad0lFaecA40gUtcLfhpOhTqwcZZSSjVmlq+KenvDOvgt90eBqPswtp/ePZACfgVY9zvduv
W6560GICqU0HppzEVPZgeHQ70DgZUu5Q+NBpFzidFFrY7SzuMSz++LX5GvPUyAz3xCoskspzP0cR
yVC/xvhHNqlA6HHyXFKfgQJ92HOzeUnOrTchRkO4OkY1eEf1pecsSl8wOve2jQ3Kv80EE7WRBdJm
dQlDxW+DWiJi3Xmsq3UQzI5NRkGAyM0HIhQei6yw7peb1uiCzpYkYCrfpGXKuokFtSsrm42/MRtU
NC4hdpx7w6iZozh947cuCsrysqONvlqoNU1/zdeAjNewoZVmcrtGu+n0ZNB21Q8GygczOaeLeQZ/
xN/I4ImToQFS01wBxPVJHuVkQM2wDQp7Jb+eZ35YmaV/QqQjA0N1uKun1fCjFD3i1JNjhFYbmB1z
hbG0sYouJF4oOJXXjH14Nm9ZdxT/4EQUt7bbvvSunSpBhjGjjf9xr/FsavlxabSVv8AVOl6adV1R
TmGxW8ce7Nt/jRajVxpKIYAHPRtvbchjFxWvZSfA8mljrLKac+cDVfniFKJKgB9Vb4WOGD9UqBLY
lJZ8Zl9vCnmvYZJhayeiu7l8YijjI1xE8EhYCPkyw+kF6ILCuDapGI8yO9E70L6eVaJBHLDHLw9Y
XmWeQF2sCA1A27rbZ4f6WI/rd20OKSVeeVcsbTx6MPvbuRfqo+yYTRD5Pyylj8h8DRtddD4P3gHy
buZAL5Bq+5DAq5id5h//Eq7kLLTHaBp85c1xcGkax2sZ7bWYjES9PCQACEzD0ujfqIYubar5znHZ
x+KbKYVMkOrXhJdzqceilW7EyoHjPPsjHXuaIHF2thMD3jJnTKahzIUBNIYfqZJI2pOISmf4kKc+
GNhPsdJqPDOEmQWd6+GMgmi2Yh29aQ7qrrtKa+T2+0LtijrrQPm1KW96Ak499v8EKrtiPGjSWF8X
9L3TeQOfUN9J9QQxWx3SGti09lsiNJajfZdXskyaQ3myzdV3erDmgGE3t6yONyXfYPNSOv80eg9s
ncI+Qes2v2cMTY5Sap6lyOBS5oM7NkLpLCu9OeoVKsN7adPJX5/UD67KwgmDQHYp7ysuCcxifLvY
kRsC
`pragma protect end_protected


endmodule
