`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
KbG6GtNx8ZMbhcs7r//bzOcFPRqkQ4r1WKwIgstsKlNcNI9ieZhxWs9/UJBfGYRBaKwwqa3tt9by
TPl1sNnoOM8/hekE0LLpDnRCJizhCcZDYpWIaH/+/gERVzkFIcI9YfBtuCXS3goupzaBBQd1WIZm
/a99iaxBiarbaI06VjoInansT6oBHilq/DGcuBwNlk+jSi+BzgGxRUvGC5wgCc9pFFmjH4j/o/eN
e1wgH7Hp9tarlv1zq/pSyZQby1KlwRxiYo1vvzd45tQAOr/kvyEz2MWxVBUVzylMi8VQ9ho3dH9g
M2ET1SaEPWcVbWtfZM20M1rQvIhcD1KOFrlbGQ==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
ING/jFwNlEmr5xZiAomvAKs2mqDZJlwrIK2Zm0rcPFghL2bYUBHcl6BmiJGR2swsUH7/EqGP3OUB
IOBEaIJBqx/kwv836E2f4gMy6dbMl/tqjQG8ofc6qm7AuqKJmlsKIXNB1vIwnGhYxGL4SfIeWDyX
04ERy1MBMVSRzhO7uss=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
N7NvQ1hrUFYl3FgwfTpNQK/VSS5AaIerYD1saXdPDvVjF9Afbiljw/kVZrz/s60EeB6JU9ZDok7N
dD3C5BBCONacniph8kRMp6qUIbD0fUuyP6FL7CQvipiuYAF3GT0XYNmcixnojcA/v/vZR4TkdoZn
pMi4coWGMayk6tl3QNc=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 12016)
`pragma protect data_block
op6kLjtrKpfGtRpK/dYfPVFDi+7q36mbz9VjITd3zrCbXjnbJIEeMwjj4ghmHskYKeRFmUrVkwdo
bmeXLLmkgW9PupLn50Oo2Y6ABXUwHOqHFXwOh55DbwbygM51s4chAksLI04MaBWvH82hXYUdBtPb
j0brQro8HvNcA1slJ6jyyWrHJXSJZgAT3tQ1yN8+oN+NDbUBQX0pjNfD7FWVUTC/W6nTTfzYpodm
u+9SBHcwqzNgCctegUNG6U5uTdEq+F1ph8UdOgjHhVZ0/f3mkdy2J6kuw/sHPymKcGihVXL3LHO3
Q0gqGKR/e4xxTdr42gUCtXC5SZrobqBzroi4NIkYZsxhaH25J3rZKzPBqJ12Fssqn+gsJOJNUTHS
A0BW7WfNWHyM973upllTdeCYGOHLs3E4LL07tUP88NA7xfO04YpFMlbzZf7rJpVtQidrHrWERL00
tBQ5j8esJ/w5oGeBgSbYkBLNTBU7MuxVcT2+6C9GXMbLPWkacOEmzURjEWazycD273mDPqx3K3sU
ChghyWJjBY/wRb2dZJBb2rxWTiLN66KW+H7BnT22LWXj3SniJJj2MNVbAzZT0al2sKbogsm5T6dL
NJ2UPCPtcODlVxHlF3PQDkyYoMGqxNMLUwaZdi2cA28cPmpoY7KV/9rEruEjnunQ6Cx7h7ScCK7G
C6spGx6SV0OR9IxgJ2+SPxehjFNDs19rc7RdY9H8+eo1uywugg2Y4c432FiZc+DMDLJPtlshggnS
Rd85c/7KmqxMbItsYJt2zWdBjD+CoEkKIZxwuyWFiEUVExSj4gEJX2O6zR2yxZx2Vd5iY0MHOeth
118v5R5EVW0WMNVs6n2OLcZ25x8CLUwGom1a/CuWDUWag/sxkOXy+tISHQc5IkLblW3CSMv6+3vp
ZxnlDFR/X/wDjjoc6dWz113O2n2mYB+yswfpYPMCE87BIJCPmdooSRTMv+p29Mii1CUItEnxfkQY
H19dfBSGQHimvawa2VFMfUJfeFMfqpuLIclFiV/lFk0sceQ/NzSNParG0AwT/dhNxjIaSfW4DuSt
G0ntWFEA0cjh8Q2mH7Mr84gFm2T28NJrigZXQnJh02L694aF2IbC6jugcyD6KXvSBAf1e2Ksx8Ge
SjZ0xmlU9BKXVv0CU/VtO3P4tytUNKYwiRH7Zq2XqCMhY/4dcRhpqJjl/Bwo8ygADH6SycCoIaN1
QfIFDeyvXSUeggBgeXG5wDb2ZJMRsv9fsc7X1ZuqI+a2o7Jsj6VkpFpAmFcOfEFLbRqZmdH41Rlh
uNCU2nBRNXHCV7WvGVl6BZipdd9aEtYOQ1PIDO4oZSnDtn9FUsRSvMRsL79DY1jWX3ePKNDVbm6p
E89E7qCpXkrHwme9pEHUNgclya2lagqt1cjMy4kl/SRxn3PdTH62bA1Nc0bnWpqYtF5uEf2LDUuO
HQtYanD7MtXJ/ddkSM5Qz8VD71SeY1dA+tS8zXWHJQt5/0PNm6h14C73YcAtgoYH0GYO7OPu1shV
eCCF3VSoCa+295ivAruPzbikEBtBJf1GZcODLnUcywKsFusVsy5s6ZyNx9GMHvOmIpjPo3QhQNdI
lZZGEheCjAHO7wliIJZ5HiF36MwFE7N8SmSG6prM0TRoYRqdRRqhLqiJJFpQj+CGRxa3fuwQ4w0M
074PmmVLxHZV9lS9UF6gcjsAaBCBWbW9RwjEJlrr0XQLq/WAxeGZcWHtFfEv26Yg8hO3J5sZlRwL
r1a0Qg2HaXgZxL46svqAhkBgKOjybce+b9Duqqclb3tiGUHtOKDwUsKokzJclaIGifH7qhKIX+B2
s9whplGnLuAUBWiNBsPZv0DRseTk4xuGoAcEcXxI2mx+FYqLqIX65cgtKcZ+zO9a2WacKerDSwRO
/qp8XXcwkn8EKxwZHoflbS0FnX2upNn6XqDmOfU4rR+GuSNhZJD7p/LhVc/JoX8XxmiBQowov/gm
MSBZMbtq4CSdSzwxTIETxTGCNizkI3/Ax6snDToK6uNcJQS2xhyTuSBLy8d6vnMpJmAXd7gV9Ixr
+3K4QC2iX6Hif4XMYfN4JL2UlBp4cazvQa7nxs7nCOI/nGS1LWIbDzTGaNlL16Dg+PeqsNdJViNq
9eGZ3RHyPrQF3/aOaGlNXWdWxi1yXUJux8nzL0G4g060hDL+dmopXw+RXaiQK9L+RGdxs1DhxG0A
C9VOQTvzHqmXZjEFLTJ2c3+fW3k2zybUt5Uv1GeZh4fR/cSDAxJH++IX6gNuavHBKos4OWvGFq+Z
2sLg42e+8KCyviwsbC6uNr/g5/iMqsHhJa54PscGhJABHkgv7GYKbtwEDUOaqyZ3YJqA62Js0eso
u/xLLOsiaTa48qbv3W5rNBYEf9I4uIzsnj8g53TFfqaeNI1Yo/OXBTTET7iP/KzO+R2DYe4gqgv8
m44OAi4V239CrIGmPBeG06TWCmNv7Yd/6Yq6Ul3Zl6fYRAopg3ikxb5CI5v+DEAqnuaxYgIh7knn
ZyYOaP7FnTFB4h+7zv5ORa3UWNVlKoIFCQEZG/+wqUFWaKio2U5GHHAiuApWOqF4gAft4o8WkNSS
iAzj43LZjOWtXxpU+36g6+dFtkNQHF9asacH+3fKEYDyR5+O1Mn2zuRRIXRhwUjGrhfvENRqdWxi
nkzjQ22rDaF2h5+MbBM13aRNxPlgFPkE2Xr75WieDiTzd7Np3kO0r3DnGJhS4SkfMwi1ZbJXJdfv
JT8pwiw8MLRis6eLDJv4hJCg5D/8I6Hr0z/UG498eKce80ATZKHTHl+dHkCOG5MK3HCk1q2+IIn0
pjkuV+j/8yWRecO12Hjy6zgkY174XtEe7J6u7quFTv0GJTqqarSRDzOBNun65BUTK2iZYBz8f4jE
Ezecml/tkkfHDRzTw96XJegKYo7GLr36k4b9szbUhBYn8L4le198Si4Fu+f6pfjn9ms7C8W1kqLP
n88nQcRh8byJNwzNxx/2OU97GKUJ3Xzg4maFDUMbS0Udla6lfOihNUu2Y9DBrjoqsAN4n/eYlt+T
27EwiBKCxvbNBKnbfTcszjQBNXoCheHK9sxDiNQwR0E/KbS5wKQNQqqbGI0+OCQdqtKD6dQHDya0
4oHxN5j3CkLIGNQ+M01IPsSli+DHinP78mp9+RFf/lkOqcYgQRBqQdbBIdLnJ63Epb/d9Nbwmn94
3E/r0jkCl54+0d2raGkI8Nt1R/g6KwPC3R55ZDONypIJ8t7k5Sq5wVQ+NbSxQcfJbqMVp30990sp
peeGvbsMJ4UW+yw1YaIFNU5aw3amNBKhMuxKhBEN7H4pwJG15vt5dR2ORITa78hrx7mrd1g9+dxI
9JGtgxhOjB19OfjmjcyIYYUuFHkpnwNHg07DqMCKSa4TzO3UMEJoO/sa3DDP2LXe4HCDedAMDoAA
a+c0V0aw2J1M503PnTYzx0zrUdXfuCmtGKbN2o/JIphsmXwtm++l/o5IrTe+2wEwB2pZDdkKj4hU
kUqhVrG3pezlY4Qg5yeSzvYxjVa0sQzmvmOGRfCrIVeLEA9ju+JtzFfvqLcD5nfw2mEje364XMAM
AJdRmIIdt373VF3ezvGNTIEVmm7+PHGz9d6a8F6smqFaocgj6wMrBffreG9wegAuPyqULHxH2HYG
f+ygxPcndBA3/7m7z+0dvWWzRPoABCWNPDb6/teLllH7qG+pRrfiUpejAzylJ/aHxd0dFhhPiE2z
z0gG2fEUMXLRgOajYTUAEFizKp8gSjzdci7pqSnRrAXu22nf9j4FXuhuu+X2tHKeU/TkNSMCWnuY
NRZGgGsNbGgAFqQg+rcZ9oY81LS+6N0dV0Sk1CRnYVWX7lCBW7MsbDKecdi2SPRDEgNs0N4NktDe
Xoj2KYeA9vTeqZAgsOKdlMy8NFlR2IDapZzQlieofFO+q5mwGBxzz7fEimcfNVXq75ohnHRvJfGi
aDvmDQ+TF0aFuFwmXlhq9GNe/zJRnhZnglsR9zq77VvIu+uGl7Djg07bi6AYyMhkUwZ6aJeNwo4c
i0I/8z1QRgid/cM6u02F1bg/BMpnDRWycr4HFkuOoNI6GoEMSmZV3XAw4+MmXb2mpBBm2kwJ1isf
gePo/Wy965BKroNBKnbKOOB8qDjUs59bDC6fT0If2eV711H0jY0vklX/+ZJMEuaknt+JHLwFmSTS
dUWxtxcxzjacRG1CObF89WYy/2yDLXvuIZtbGyiB2Rs8jjAiMoldqM63MweVVnM4Crl4TuoTz8g/
oj+cGL4cI16oRTP6BZeDrhHITMWny4eZSZB4KcyINhoOYJWo2PnS+cW7knrT6yNlHtrqeV+D6lFq
Za8nGFbH6Ix0NoTUSxAK4aobD3CtFswRakgaL+zBzGXSxYqzVmJlszcNmmoDxX8Crnx16uOxKrBV
qop5kkf53O/Pi8qRfwyZyk76ilGtQRtQAkUAb2rypZBe5jjue1ormkCaJrWfWZTC5Pzi+MVBtt50
RA3dQN5dHK1vthp/Mj6/Inc9K2j7BjMDt2ydPZRRKNd1tfflUMbYk1torFuZVKQnDLTGiMWW5vEq
2rjnSb3Fsk5TvGb10Zky2q9B0TinmE59luWxPb7M7X2fHU+vSNcqKcuPwKMSvhsmU/JL/9vmWWg7
v6869CXDJhYlOFW61APtw71LsA2JyO1SUzW/pQUvNl+tkgkAOyUrf3fEzKomuyuHRnrpkCs3p1xd
MIYgPJR9m//llQx2869utfRnTtymaVZZif8CNvYLk0fbnjnQtmUWFHmAvMH5+WVPXRSACFio2tX8
ygeobPwnDa3XJtnhuQxjKFL52e028XXZuJY9QIAs02y1U3Xxu7LVNEXQwD9kBmuuMc8cqNAsF+3E
y+ylPUOGVLIjZVEbdcOnEjXgtbLevYLtjlmYnngCFWZQQY8XhLcbeieyOUm7dJ+Y9HVWDyGllpvB
IIl1FzxGd9nOzClcUSsKZ6PHOz7ecnFYp/sgOMq+68/hPSg4oecxTVkiQqsOrkA4CNvXOuUsG3cs
M4hoZg4Duqgwfb0jJZQCxzCYjYPR+4rz1n6Bwgn76LSy8o7SphaR59f0eGBErLOG/eJR6HKJuYN/
qKKMfXCZtKe3NN7cFxtYd5lGiGGcZbzgOUkC3StR0G8HkfpG8nyXYWyFMcIQVyiiUCfYaifjpA8h
o3uRNhjrqhTB5ivIPglv8+JR0kokYp/DPfB1dZ69P9iiHJRz752lhAj1YJLEsWQUfYZh9kumCP3F
0gEm+T40hA/Mdmd1krYKfX/nGPmdyYwJEGZxsnMgJD5he6nWuBwfwb1zue4IP9+Riggnk4HDzWcl
JoB4Y24gL8K2Bb785Hy86eVpn6q5IY1bJ1o4u3tRb7ScE9nDvE/h3fxV2+jwbCnSkLu/dK+LkKgI
egjRC9yudMucy6blPKGgx+dPL21ZQmBaxIjaaK6cCmi0NPudi+vwh9Bx7RWH1/hDMtobUA8xpddg
PVoyrncDdosLidg0DbTOJR2xaGOAXTJGlefQuwwaVQZtnBnKwaicb8Nug/UEyGjP0o8lSDhe2oKY
MB1ivys0G6a3zu7DLn23HSs/gGCRbN3azqY+eZLb8BqZdjX5lg0PNZ/xs0aws3k4cdEweNVeXM/U
c2Eqn1M4hoMr46kgdD38Wznl143WGvNQxIoVECaP6qJPLUSLdFau/qysA/tBmZOvo91Qrhm00YEQ
CGOVQ6P26lKTjavrACf6eTAjaEZePuNtzzMYCqD5k6Nx+CAga0bKkGvobrFCjMMFcXG4f+BgyNl/
qTIVHrQh/ufHG5edp+x0i2f6YYWTe+D0TqX187od0aVnT18fXqGceKClDg4GI4d7T+tPur3qNJJt
JoaHKY2FTJBClUekRNKiVFHP5BUy2x54AeHciQhkz/D0/7cDV/N6HUp8hhYsP6ptN2xtSQ8VQwwy
1uTC4SN86wmozkz6Zrvf8ogVMDIOoGpq1Heq9f9Pxz9OkgQjQaG9Wph7/tNnZS1M1gbTMbT5sL9t
3FmFHytHbY3Kh83eM94dqAWuhhZzbg1PFAlSB/zS5BlB08FBL3Jqbfn49JcNPTUVP7c+6m0YJaQF
TB1/5s+neHf+XZvsotRn1fjMYho6hj/ZUdsfRgAcyq6ZcxC6FjpAdk/P+z6w7X26dD885Y72H4Cn
fTDrfFMvM7c168LwAY1es4bZAtkkjRNt+y6O9c/X26/fB4QpEutBr9kbiMz2sy6aR7fEZriA6UkO
wTc6M7XXN87OBLM1QaJfBNiHCrn+H2B3gyu96s7VNTlrMb4q59Rz8M0qQi213EO0j5WyUYssShYR
d4qs+1PPPX2vPuz4Na1Nz845usWA+dWR6LBq4PVM9WXXvdlhBlIZCRuRb5pN0HGA9zbbyyHqSjBU
xqmk2kK6jsuELzhyjVkbnrmZby9iet4gHQyTbd09pRN3lnKY20SCw/Ob/HpSd7j8+wAEJLTlutQF
/ov0iGYOk3+/4nJ+vc/A4La4W/FpqLlXnpFg/Jq+9dyINTtjczbGCIC62hNPDocGqaA0iW4K/2t3
3N7fU/mMH02eUS05/8wc6uc4R1r1eCsQ2GLDExyIpZ1igC0BXXpiKVHVrv8PFpjA0LqPhL1k65BQ
G5c9fQiHsM1SB4+OJFS3zgy2ipEug4/yicc6TqHVpI92r9PiNezpgwegUfBdWtVwI7uoI/+WjRSc
qjyglGI4Ya+1cwTmzeXwWb6sVKeEbttxKeDN7nvRIH1/kAes6ZJU7420gYV8N74rRWLn4A4dSrPI
6GKMstJQaIukatLP93tpI4BANLkfwA5uaUa4XuOHxXBm0tI/FwCYS0x2LNWMN5FUcp3pJxkGeNk8
1/FxNhpVXT2SuOgATk+R+wKJ37i5QdCEcZ7rHvP3mHUWn0bOijsBYtkuFsHr5BTIclnputQIcYiL
Zz2sBAjSQK/NjzsZNfZDdtkjJKRFbVZAgt7v9xeSRSwOTeN479BYTP1I20cgC7Ju+r9B/Q9lQC2z
c713pdCizSwHYq85HkSSdsAxkcH1JiOKJuk/RLaf+D76quP1yebO2k+RZTnLiaTl53QUB3HVL3LD
+NPVekhVj3dxSSsxKJxBUYslhBXA0UFbfBoCbuC6L2y+2RaH/njmND2HBzM1G6i1qETHgBG39680
j3g61iFd/pikyK9jkEc0svhivgcLXin5IEURj5RdqaxG7qQb50eR6r9Z57sqbKyezbNATmxl+g/y
/9hla26FptUKkXq+NAAWXP20AmYoXp8jF+g1Dh2yfcIiMkS4o5GUFhpTWGGv/vHEGZrDGCbO0bLD
U4S6pXZFW2+8qL5FnC8+iMbWBoKSB9xP2v2LnfjAr+NJnJzu0Dw87n2PuCw7gYL9SehacdFc7vNa
XneH9HXu6YnPbSgeas9jCisgEZ0T1JxSbftBLnUCwaKOVHSr1ZpSaABRhnbbyvJrNeNaubMDYnTG
AcAgQCQlyeiDeENnt+8BzuKXq5sGoAzy7P8vWojjrVLO/tnwgYfZsdLrSn7HmO8vrYgvmGkR76Gx
hOUTfE8Qz+j1kdeo89GWnRwSLPK9DgWoOQutV91yCn9XunYls+bybIBxCyrgvqb2UFqYnBcM6NlT
8kZd4pUE5ClJ28NQEUM+b0sbyubvYde+ccg+123JYHF05idvm5Qv9lTp8e6o1o5F0Q1O/r11FJOc
YlYh2E7dfvHkUcU+6NdLvlD6UWsLY6UBkRZ0CX6CdXBWc46kkfV3OVDXxmMl6yTpnwpmlQIjMw7x
oecJQSyLDdVfbAXnkdHC88Zyvvj2G0xeb3rZM+YXb3BrOcpBCtTCSpl8ym674PLynXxy6KtG4j2O
7QZvKDViQaHzkgOaOlMYeNimP3pZ6jCQ3OFb722/pMiG3W1ABpVscHiqhRFhLZOuWYbjvzNtTfjB
GyCLXthzn2pHzYxwI3m5MbHuLH+ffUQ/UPEMtUl6wxu8FlLxeMfRd3o0n8k/TufG9MVUzn71OKZb
eW0oCXcQDdIyUuuiu1LsKSsDP59sdEafuAveW5ABhvKRAzuLu2kS/uk7KBtx9XNEEnScarwz85iG
yEQyyuaOc4l4ZZSiSW8pCYgwDMjCEOaFFGEYNKlIY/mVCrgdWGQd8d1NOp+X6kFYidl3h7fkq2TD
My5PsLpZXlAqRwUYHx1NHmRilymAKk3AVVzYJvkxJRdWqIg+I+u9jsHn5En01G9uu42+E5QeOIKK
/sPefyvB8rIQ8g7YWOgiPP4b8d4hpyVDGGGJ45upcEkfuaoL+5+kZxCEmpm9SrnjRgfNg74QWViw
LRgdzD++0dCdpnG15aQoJkGRcgHv6ZxZ+5yZ3uKvkTB4OPyZTSiar932Wpz8STR24IMPobVjhyy3
eihhxOdvDEYsjCnWf4xwBarfjzhwulT7alCxKrHhAJiCqNxv5qA4azNjhEVJAl3IvFLSGCh1xPw2
hFwvmIBB7Cwm3PGMsg5CkeEE02Gm87kTGb+mOV0xtvzWmoTogDhR12SZnXglQgVBV2uC+T8wDpt5
ZkVV8eK1El6AfXxLqf9as5uJ+gJGHB2nuMrsnt+DKLo4D5DO+k8URZzjzlqd0Qx7i1249xDW3XuC
2njwvWcTwTlwgONXnMlbc2bGd8uWwTejcP85WHbzzRoCB6QR0eYQpkBcy6GxH2YZjcmDY/n3p3X9
6SaPtT0llu/u5TeYu7NHz7NMbO2PxPwWy3yvwr7h2kkPyOhAjmd71prtRXxiSy7zS3gvUlbGrNfm
hoDqitLNVd0GmwxUQDjtjqyhR76zNDXP761F4HyJe2mBA4mC3xEvhNTTeQJccO8+9EJ5IH7IGdNk
mztqhbKTbLrVH/dBi3wmoZF8alFqgtt8RpX2Mw5oI8qal8sKhAWH3kTn/sd5bKSkT01XCngEbJjD
Z7UUF7q7tyJjiHdSMFzsy1Le6astM9USqd7MhbAG+L54/Y1BvxGIqEyrVNMldub85I/VOi8EZ/1d
vp02gLZJe+k3qpc7m65MLnM1ndCjnzh3ZCtvbD+SvEHqfMwBKN9UCFEshZ0d9L4RR/49S+pYDI1k
eCENG6g0bvzNe3cOKhk3WXPii2tzh96Wvg6KyaPzjZ+skWh+AmZeDCHpoVFunTn0rNOk10mWp8yA
XKXrHwBgetKhYVENdbvRV4xwh3mOb8bQslqUIUBo6QlSXtV7yHQa03+363cBS5MEBZ11ddmy2w7j
mrQ6jxXXfOeTyq+f6LkVOrM9SmLLei8ZeydRsLaP9Nusz4Hu6+Co9/BDjWliL4od7iLv71oMhbOe
jQ9xCPuYRZRk5Yy+f6/XEI7sO4jr/YkF36fiC+ILua9IqEMBosWGHdbNWJ9godP9B791HiHI6Ulv
xxvtkkcZQicQYRfbCCOWFD8EV9aBzvGtNDTCmzXkbCJAgvSFJPjnYLGXmnyKC57B2zZjYBwAQX2b
S/mdCT2hs2S4ty9U3mJin/GXKV5h9pnnR4RrKHaqNU659d/m1Z2fOwqw4431sHpiK9Q/3jAcOc1I
/8PY8wgDCl7Dq78BfuUJPZsUOxcMq5KU+kgTHX/K1qT/pSyx7bTGqAXW7GnwnO/BY6iA7b49pgIC
3h/0X31BpX02EEQgr+kHhwrct8SEpS5HMg3FkoAQIIFQvPoo8aFfFNIXAgmtrrcRyk/+WSA7Hj/h
wF3Ox7bkspkkWeZvyX88kzwzn8XZOyK5QjEfrZSnA2ZXhB8WfmgzbDG1gTeg5BIM4Ssu/ba7us1y
s6K8HINKxP0+SD/Z7RlJxdZ/9hS2Ffdea/1IzDqGJv/opilskM04CnPeuVo3uKNpKkrrtt8ArZ+i
Dx1yCtoN8vJJubHAVb/CkPKHDYs7Ad7y9T/JLyrNZb/EyGQ4zDOEyJn1hevCTMZC70972NMMZUdk
PbvWHBzTTklRI2dS/hq8S8cOxXGeDOTGeJpcvO4UAFkDeW81Ot70BDJD+tx87YGI1r+1QixRaC5p
r27tVwVzUgPDaPX7Ssrx3HKlXK3WlD7SgHCXWbf0xA6viy4wYAfqv72nqeqR1xtSyYBHa+Eb5fd8
khCwgw5u7LzgaZGyOGmy6phhdW0mAlHmBoPoz2xSQ9qFOKU76jzXXqCh8Ey2kGMeqyxsA55lGE2n
yrYR0sclFUSvpVZQocuZYtAHO+bQHg7o5oKRXpNJIul+qsMlLt81BfqPg7ayH5VIMNfVrEtfU8gT
XKK66cmXPFFxIe0MvJPMEZGw0KMi+dwB+B1q+tlNT0LwGlnKs5UcM2pNZynYsmKjSZY3YqcoXvfY
OIYymwszy566bon+uiyZqGiYdVXkYRResEYpng1uXGOm+sk/e9bsc0gReSxGgpFG4N5CQ8bDlsUb
b0tWtfp+xxbs0DJPAVaO21aHrsbaUDaPJeTEysFSXC69SLQQit+PzNLUYwzIyJoe/5nh0l2dTV4B
fsofBtfrRSkCQwQuEJCjHwXIEGJW88GujmBCpxFVeOExlI8NVJRqnI0gEOKV0FUDsUp/xBF1tl13
n9F3Esh6o42GJrmdz02PDL+f+yNQNkSGCFwOnf2xUCLJv7SDrknlj0xLWd3Fn0LpxYM30X/7GmKR
BnAufRQGGll2y7LoM0ajFyYMwq+YiO8WEW99ayCotCkqZjSk+uFaPhMr8fJ6vWU7BrjlMjH/frHc
q8mL03Of6gH7qifdRSho7UdGvpTytvQV2XOtb6QrMchtWbPThQW1YUE0jWPjQyYtWon6p/Y0Zcah
SeAuju8oI2TpgyMGDgVkj7NSwl7NA1wzWhJJma0zxc+YEspinRDswK8JnA47VXyaYTB5kATgwj8j
anBRDxp1JjZSNqACavK2K6cOtUqCogTWEu++VtXflq7986BDDQWsLHt/4yWuMMlmcWGiVDxTkjRO
LlqvzhMGStffCEXQJWblc8aSPQFPqrTF6PP4xTn4Fh0QnopmxeW6ZjRybLQAf8u83PYY94IlAen1
8c5JhZWoihIf/YWsDJXT2FAbyy+9HmhyEyuTKTkIaT64GNeA0SOQzuZdjKHYWcn+9z5yT6uGZlHH
L1BNqjFMtKvCLRyxW/+IeMRWxI6poU2SYN7CO2Igz9d2t8awSvht6e6a91+Rkq0c3JrSN0tQZCeH
/oQKi0+tOKy0XVQ4NLcMmjUryJ6ck+CW2Ocjk7SdAyATK6zxC5SJCfHtC8vC9hl0+6b92FiWLMDs
6U6I0rBG9gfzbSeq3WpF7xMQmtXIxi9fWPbBAXVecmRRuXBKU/O0bspLTpLjYkr8QO5sBpMnAmIG
MxuCoKYQ5Rr/09TBPBc9/IUlI0zdtoCCdF/cz6Pz6OddypCTpQ2ffio+tDc1w/4avZzlKgZaJ4ZX
hYqXwr04ZMlI1KCJ3+9v65lOPY1QmJRftouEGb1p1Ke8+UoJ2k3rigaugQEPPSRzVrG9NAKVcG3X
Ad0uMi3RkzzKqT6ttN8w2JJcA55aKMwcvK8FAd6Sma3rKNL55ezIXVzLi8Xtn1BzIqxmYSHau7mU
Jnq6o4ONV1G4rGweMcz5j3cHJQnrdxEdtM5LLnJeUiTn2K622RLmHFN2EHWdgGVVb7QLcKMk3Bni
T0tSSFriieyJVS/TIUFmppMFyobgSGgN/a3lM7/9VUaJuZWCHQRX9nX0Wiesnnm04N30GqLg2sI8
4FF++7KvuwtY+fNDOrGd31/9XmTfWcDDjSM0oTv+APycB0ipxyfocctDgR0ux1chQ7JyLaSbKp6i
36wocTv9Wzb7VlZ918+FbFdx0FMucNKW8IpMWNlqUhvYSCwuwdiIGzyUoO6e6A0/YGAzx25bZGzB
CuIUmiuOZ5N+DxoJdFrUZWCD9LiZV9528hRyTFz8ysqjy9zxC5eYe6ElQrVk6zIw4Q+FH400SeCA
hhNfdVJu0Cs3LWYQ1z7AoY85LO3OFMqCAdsqjuygqUtDoILex0dhZ/1PWlwtTy3KJNi8WEb/VTc1
qQcjxOJopPOdCFkhQPgUmiR0RZI9rIcC81oIrPUlVpLBw1UX7HIrkVk5A58hvp4/i7OEDepaNI0g
hXTpfCznS0SNaZHg/dUeyPwq2Cbz4jKKzxWSARbn6N4RrLBHiJgGabF7gwQhsw4mF0A168Sxm6xY
VyWma5xBZUg5p/p/bBIkJQaibLlDFjUnYB69gxyWkVQBwLypVBGGdKP8aWGzxqdbWN4DjNKAPRoq
N3tDWBgc3PdbJ6+1Lmlc8Vf0m6FswrjqeG0tixK0AIz60QIlWejU9B3F6pJecH3TYM2zebwVeyRT
QO0mFvZSKUtGlbTLjKwEI/Js8c9HM3eNg3gsKH+8duABWT4cHG9z3cHQoQNEAPt1uTs0M3H9jFSR
BHW/I6LdiAI1g57OleD4DrXUJgaI7EagXyE18/XLxWymws8g4Qi62mTL0YuHOtNlxwKkmMP8cn4K
iogDjQqYTHR+kz4euCYa1/H9+5mjbaJPsI107FKZMnn9ld4etqkbe0NY+/AXQk7ioixy+u+5lLCY
4iOCneRuqjBbgiYc42TlphChr2aWD+bqD1TlFxRj3bR0uQVMuSmsViz+SYGed6shEEpBj74lVPsY
g0N7gjBdveF65DIsxWuSSma0ilq1vENL3ac7BRmLlsVbsgWobqQHr3qkyyrQ91pOdY6/HrG2fH0Z
alnrc8VE0amUpfPbL4KUi054Bpo3jBSARrdkTInMwkVEhGOR8ygMg6Y54dooyXkDViY7Dl7mgBvQ
zL14l1J4rmwwI5zJOlGIeirn1GzsxyOlLwTDkQOe2X3yeu27vTudzyQtYR+vVp5O2mgCzvq+5O0v
ewHNdtjyUQ+JV2r9mE4ye+q8luSIKdP1DXmTgfo3Tby0g008mFPS3IBTPc48oz0EaN+Dm05DDqgQ
aYc7KZoUUkcf5EEmX22kWUw7mh0zb/QbQVcdHPDybNFsRYKJZxdPcTfOQSzr1okICHPonU7P/eE0
hgGHzEfAuBkAQ5DXTBzLpdk7PsteDHokXPsjbKbP/jKh9NMJJVjflBq62WJeHrNtWivMNfHWUfpi
oN9+NkvzyAS9CUnb/5+TJQ9g4cUavM3GB6oqMTCk92YzliS+QAaMNir58ysWa0yqJEh2wWusj3Gr
oVsi5CH3THl+VgGNcORJXO7710vov99Yd9v9/wBnK9zuLcM5SmBpNNNHhX5N1Nt9Cn7VZ3qwadvC
1YNIUgQbvXCkICZW/KKf4970l1+XEp1h47oq67rNJ1WromsnBxZLFcVuVGbY50AGqsnP1fXCLrcr
D3Cpvjh9oHGEgM8FfH3Sevu31MEgF5SgQkllMNdd109sPVmAKE9IC0YrYLxsl2zivkovzHx3vAtF
FTryx07eumpQX7wQvKP34s+ZUCSi7nbEk6wtiLMLf+Nm1gnamRZZhdzMh0tF60vOI0RasL92slWy
Kdrjm9hZhvYWbrE3H0QLaehlvJ+mBA8XxzV+1ErZ3+kitGZEFINsOBGqBC1B2kd8fksrHj1OG4Vb
X8Qek0X/QHswzInBU/k7QujumSFJhxTRlM2DvLIjcdJeLlyBZ/4jGc6Sn8UowUR3Q0LkNkm3S3Ga
19P40q3xxzLFsajYwoGBFjX+DCJKHsIWzBajBmTQeKPHnHa3ttp2DEQCLSH7RPuJkc62hm4NZagB
53mbNTAH+tX6cZRLqoEzBPPo0T0IDT3P7vY9vMkR1WeubU85MEXXi5+mr6ywM7gtTEmqyyIq6zon
GpfH3o9BO+WxNMd/K7hyQkuGQOwqk8VrC+yvcatawjDaz0P6L0wH4HDfjQpcWlmsAG5rgU+x/+zQ
xfFI5IrSw2Yl3m7OFVMiFbI9ucAnoHONw9cKD6IANzkkEGXSG9+iQfB81yptcEnpk5nWJhBm+7BA
7Co5A71d5ZFOrfOkyiS9JYDmx0aKgAi+/uFcB9RXINyXH3qBmh1k1NhPO83hfCC5xNlS+LVugzeh
8Cof07OF9GvzMg98vQ65ymO9L4JEUiLnnD9+C+HQlxsp0sL5FhX63zeCEqfo2RznCEBnWxb42POs
cCgrY7OHoCSN/C1dBb/4umnrUnp99HuSMprZ38gayiuCs0pSdJ94sqQOsoE2e/M28x2eI/FbgZEP
zTSRTDAKjp9zEXsDI/Wnl+ZF+MlEqT3BrM05I0KQZsNn5xTUNC8HJSNt8Uh2Luv6meZSEAtiBUQt
pZRFdBaFqRAZ24ZFgSd29OYgg672lONwUk4bOXFaokJGAoByIbg9TDJpVTzpa9QZiwJiOSW0gmQ6
P6VOvNAjeYDBAULSP+xe1eo2OslsvfduKDUjXP0WZ6coscUbdKtZaiYBhsIw/KHP6p2b2F3tX1IB
6FMGSziDaJz+Y+f2CRervUxcTzjS2JCRNHo7orNRZCsl8Sus9aA7odYJw8NvQLLulmLbYSUb5tmc
RRnQXavl1osy86O4il7hscV8eT8IBPu0OjY44uegyQL6unOXAEjMldEyaGL0sCtp5cwKt/gbcpcp
C4o1yLMIlpONtf8jmKAIQQgLGL92q+NHa1svxi0BQETJLwKn5CLsb1yfYcFBfOHH/+mqHoBNXUl3
IfiDA8qhf3zUXlSnC5u1ISmFRr8vIvljub+8B2WrkNN9AKH7Lv28RUc4xBVLuO5fy3gWKVBdrHr/
DWRUMj9vXCfWemG3WmiT3MqFl3sFtUcCq4vlK3RPn5psbiBYRG7GZmmGOP7Fkq8fbJ0h6yy305/j
z4bpsqKIDtfJyGx0IQVz+ZYnDOgIZHIUU/y9Ou7HS2XeAcbNC5xr52OQDQZLaeOlw/KQMKAFZLwz
Oe9R7l6b+Q3hLZ0SUTaWFXDskiq1rdSGlN7gnKh4Pjpt+DkFwBuQh4/BGw8ZxYG5bt1frfUl4m+z
K2m0DcFp/KYlIv2lOcX/SVnIvca1tXdqAW5hL6OpeWqlQFE5X7En1twxMYVyPblZzRe7up9/wEJx
/ZcG2U2CsBLB9dTWjPFkkZL0WjtWch6KY4EPNkoJa62qZYD4sLR/+KZCf0NFxm8wl3RkGcZ+3sJe
RL1lZsEQxlKvfs0aNvYFSmAqG7aSoBw+yDgyiH6/G+bzY+rLJoKWOTGqA4d7fPUDdi7Gef9/PZ3J
UjRd23QHPGYG1jyuv/vAwC9GW2HRWI6dsUWcrt8Rafk6JP81tYrSntNTRpT+rUAyer/C+EHn0HzN
8IqDGgY3q334+9euv6RsMUtGWULPg4rzjmRVU/9Ev66y4hwNHKhFSxuFbrf4fb94gift5UX/t8nY
rgiJ5tukdrrITKUrWg7/lyKhZFrcUGrIBI7AYaScKjuw2vptIY6j2a1XwEdNJ3mjBaSU5cIWjjY5
1nDkkNGg8Mk+qkrJ3biEWxl1DX0ARzU1Tlt9fiO3PC1A+KzbLmwyuGMJqdRs1lpTh7/fzLLEHwqv
RSJOB0QYMgnsE1gz47V31bXNG7iGwvtZmyAqdyYizxrxxTqtvEo+seWT3xZRrJJtWs2sU7wxuFT/
tpb0JHtqNJpQBr0EOh3hNnwQD2ySWetQTNXmM0Mwwaps9GJtgPebvpO3lXFmbsmpS2fmrqu3xhJg
R/CKo99RGsnTDStTr/wMRA98ggKNwOmieU9IZcg1mvz+ic0Oq82CW3w6GBBdKilfK1UkRzb8tECJ
W+nPfmATWn4NmsOXNrL3dQjAbKxDJJ6l1ZmnxQLs6t/BR7mtUWAkMN656w/fwrh6jEWciMCaKDay
R3XU1tWj2MLGwuu0sgCoHCq3Y/uKFoGIyeUhufR238Jd14Fwyk50wOWp5yF1C6TeDP/vqvQVRbKh
7ofk0JWSInsI0ORGqNVSGUjWZosfQnHX8wCXgvnvNecqd7IYtP0psWeXBphJ5NtYOOQo1GlUZjWF
3pSepn4vtTkB9CbeEG9dLXiZVwzywrrUt1FIFb1Ji5HaaJOXfV9fZLCvllUjwPVMiEQIiUcKaBlo
1/anpfX6kwChy7m5RAcY4Uad5Y1XhEOCrNwVp31JN1vZEKmokpycOWaA4HSGfEe/MfzrNDzjSIpT
Gx5kLmo6dvJzy6MYXMN8gOK8DGXNPLYbO+hDBI+aI9Q7k/k1XwYHW/QHOndvzw==
`pragma protect end_protected
