`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
BRntypleKsiOOGcMPN/Hazs4kR7KzQkISbGh4WySGNnASVrRpimj3vNQw/xc/v3xRYqfQXbfTRqV
s9fMSiIyqt4NQSSHeYDVzlNH45BfVSelRO/SOc7W73CP8Zx+VENHInxNydYs6A2TwHTnD3l6ew1e
rhRIpiqU7eqgG3sizqi+VUZem0GfNs5v1NEImyix3fwSJ7Xh4AcpsRZwhziALjJvEjU+CXjgWNie
q6YTG2k23kyW1PwhcHIm+UoWfGCx/9Ae/hMup+b9VJZhTj6I6BntumyGVsuzKi5Z/XrDb+uNLJze
AqE0/oWcPk4Bt1STYL1wmLwknIliXu+ZH2gN2A==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
AXcQK7AjMsPi9vewhTS0Iu5rJ7WJ1oLmLPufC8HdcOD9S44t5xg6R4ke75slM5pxnfagTRTxcrLD
eM9yil6qXQZk/1ljf4BOvxxStFPDo+lmkESICUYQteHvnscT7gWP/KBZYaVD7fYCY4eghe1S7dyI
5nKpheo8ytPcwhmqG3c=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
FrjyNUbE3Kjf/BecrIfrXblSuqtti7hklmxQCUFdEm+toW+DhVEM2SPB2arjflm9NFj5DYKQgx/A
pn/6Ofz+JuqW3pcJBsqL2KgjHaaaAabpxAIxfLKrN7xRnfiA0dWZacDf5C6IXACsA6QdPwxhxLAc
5nWYOQLl0rqhCjW+wtU=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 16752)
`pragma protect data_block
8/afaz9JiUmUlk5EV/+ztxD2edmUs0Yy23fwW99t+wh1YuzCqSWhuPQ12tYv1Xds+oKevYawtbkd
gkl0j7B5QvRzUsuk9Mq/a8KaRGIqRBTUPXvA+7LXSeQvxHbTjztR08fGpaYfqE5z1pggZKIQFFjP
gCZP9Lrun3Pi7K1pi+Tkg92YVJJFpdc0iCtApCoLnq+5xprMnpLkT/cJILk0R8pG7bGCibuzj+xw
q5BlhPMZmEIMrzEMModd7Xiak9ho9vZ2ODAgh+q/ddsQlRyOYKvm6Kk7khyVRSIDdrLMG45FqqAE
K/hbmiLmQEYiev75dFjI+NLNNzCBXS7O60Le+F13yrRY2Vz2mUumxH7NDc7TiHgZIU3bwLgFEOMv
ITH0WXxFf4CG88wtMwUEdgr4M05Bj+NldLjm7Q4hPgSQp8wbmXfFAxry3Pmrud4AGbYhffpP7CpE
cIbwjCgqY451Y6Z8dMPJXU6l+ncwJtpRMeLh80YDYSCds4MBc1Kuvj1rjt1YekKADKDJ+Ug+5fpN
pA+IRUH6ZFqGrjk/kCrsHX+C7c2XXwvI+GEQqwdzvf+s0Tz5/RxHisLJVHle+gmy/lH/rlnBTaTY
JbGhV/T3jWUNRqJSQQPQirPJlXEYcZHeXt/g/FkSALE5JJWG1D+Z7i96TipyldrVakBMy1Qsrj0h
Ie+23od66Luaxvz20TKlePsr5Z6BdiaSdaGKKYog6uraibGXKqCsDf7j9hMHTCCz6qNWpbyor35S
GKwWBZn4zVj5qxy5rOHoeNbjfMGTGZOfY0UmY2RQAS0pAbg77PqCjxqD/PPplx2e6OxCZINYSU/T
dOJuunQBkNs78EWNZH3bFrC5rujbSZiVikhtcIa/D4h1WJA2bTCX7cdCI7olcK7RqUlCGCNT9FBc
66RiHJvEjrXr8vqfF9njOq0uy0Ww/jHUp2TDxVrCrTfwShafJJjTFnwG90R2aqMtPQV8jpI+i6EJ
j1HQWK1Pc+cufDATpMngafUDX+PJ1cuuPkuiNQlr2ngFgzp+gE7Biue6NFrnEcSN5mF+WZqkRzwE
pa1tUPMwu2b5gsYWMXJpngfQA5CiCZWo0VWxF88fTK1GDui7q3RreHHEzrYUlJ3iizTp/bxIDSwv
IyvCXQRdSMLz2kAsKRBxrs/1ESqKWswbVKg9yBEOHhEYylbMDZo7gPpQVljaYq+GvJiXGqBTq5p6
YZySDXnAdRqjYdqJafKTKZx+mERDP9/A6CPHUEJoQDCi9tH8G5aY4YJrbBX4nBvpY+2ZUV8LiU7g
a6wC3flUPE3185AOUfIPPeKWkH5dXCNt5tBimqZtLFJ0RaX5fh3GNcMrGjyj9PbVehMOv6BlyLk9
YdZAuEIoI6lYDfudq+odcJ/+TSvkl8MvqW4uWbUPBBBNaKKbqudsGrG19pSbSC/K/c74vbfuxFq/
gxNwtMg4AnAOG2U+Y89BKHMRTRcxN9aurLF5v/OWBSr308ssidY0ujshYngRtSe98ayZAo12tPok
pck+z5obPFNFMsetVYXpdchK5lAjcY2J8ZN0cUqAJM8JD56648oTvxsrh5/Ew63S7NMZju0ajwLw
b8vKL35l47+emD4kvBk/sQci3gfgJK65u+xgBDEKJWjv18HvRnkdGE0q+Fal0X9moToZwXCV6KKg
HCQCSu9LMC9gXcqbzVi/VUhK+rtx8zZByoXnWPB9LL4D71QAVOgjdx0OwkU6rL2cUcgxyu9b+rQH
HXcdnrfgi6wdaFRg4uQZif3//eVIq+SMndc3WE0r8W4miXmuJOjQ+6Z6NnV4rUEG4IQTuOdc2DuW
gvHbDMpdwIKfM0K5FPHUMR1DwKfN6zXocwk/gK/uxSi8ozukOT7l1VhoSFv5HLYe1kMYKNVdaxbH
E1VpDT/19QFXRcJY//tf+gYrHmmHEFJ/bEP9N2CAI4TIJCUdiJs0vIFqGTP0a201D3icbTTKdt86
r90hsXiVq2MaSEWez0y2bkOgo6C9YPTn6VxvRRTRcSTCfOZtNbVCvyARSl5amFfFu/bEUGfLOjG3
TLv7Bd20F92CZFkgHRirI8KPXiU9QeY9p5f6L2tyfaHscbRSNT540R9U7KOPhc39dXdQ1Uvjn4rC
pxOjDNg5pPKcFsZ8WJf+SeKbj7QhgFiMMbL3ji+ysRstERjno3eZ2A+FmsDBuvp6LXQod7T1bxWf
qxwYLaCrmH/T5VGOdbeJqXzY7AI+GdfEDX1+ujH+KRVJwUnHqMf4GWfwpuBK0Wn4YFGXvA5uFkGT
MjvOGxznjhHPpXAAUqSZ1P3m2MY0ejJLsGYfqG/OBx0Z/D2orgqUcoBeej2bt09i3rKe8ekajAdw
OC3S1rLzSE8Edxk5fcFI9f0+31ETdHTLmmAimo+xqURjysrLvymUVRWfLmGx4y2XDibUuXxlIasR
o4/IV0hjE71JGNNN337WYL4P27nGe6OGbaD7EEjNhTLb6iHTjb3NgS5UvhTiuv4Gs2mPIcoks0Gm
6UwXbTV5i5kJMbSsd5OG10HbbSIlRsi8etSfR1Vr4ICJ4pHqgSs8b9ZFq9IMwvMaHsGGCJzeHmvS
FnqCDhZyuLyB4Ob/L/Khz62kw5EiqRewCoR1o5V8hRIEM0p6sFU5cF9UiQkR7IcTC1z415pNgUHA
mofQUWgvFP1fU5+zbLZGhZa7qwlUiHvKKibjTqzdvJsrSLGEvujrAmZ8Pq/m+fNiioX38eQcdWrO
vpYXMgfzo8NBQNzteDcBMeOvOgRWUWR6fHco8IIjwBWQGVcBoFNnaZ6oF2RIYROXAAxCoxWGhW4O
OLNW4Z4FpOJ/C8mrEFYYTz+hjfmVNQoklEzHYDI4ivLnGpIuaCQQmYggUDvm3Ii+o4V6qjOlR0Wr
NIfv9KYdU+xF04vo72GFew+FsKAhFT2HNBvaBDAaScew4QvrMjkyNjMDi3353wbAoAS2cOkm3Z2g
e095L2OHuZg6oK2lXVlNPIzoReDcbVRjbHvq4/F/D2Lxw6NHlZYv8irjUn+JhfU4qpZ3J98zI8Ir
8GDhhTaXjGYn4JD9710GvfYoL2caaeaTBTVakP5gtoBkQPDRH+E1KEdQAjs7FysARJFtBaepKijw
SDpP1FZ8NJ2skT0+K4VA/X1N44xcO+yMLCAOYRuapqqCBznyICv1CNJVIlxdyHetJ4gDQlZJjvpF
U4DbYdk7MWe385e9IvH/U74Ps0U4ztNAxq9DH5m8iCM8E8m3bgMoYO9aayObxvloOx6+uGrvm4ig
1fKdylFBERmSsGyCVcyI2bGh85PCDmNLLFl0WjqN2+05/M6mRRXiYo7OyfVwK4CqdQkbc3A7f2nL
v7wvfzGpTZgxFIuq7Wgs/sN9wpnXMNco9PQH+jQTN4rKeJjby8cvFfKZ/2JaXBwnMtBuGCohpp+I
eY/uTTtkELFH2GkcTU9CkmVW0H/bIEMTCUQQL6M9Uv2WV7Tf27eLZ/6QEpHXzIfJItWxOaJnHelq
Vyp8AXhq7426SSAmddKBY3en0oOpQJOJe4rMVh9gEFfywoTarENKS3NcSFEtIGDIXEKD/7EOnu1e
T5A6o3dg0B6vxG4JubbxJQr3lX6Y4l1jIHmw0cKx8hp0LfgGaoCbrm9tsEeczffM77eUpQrlcgWw
HX/i5neueGDLp22ca2LueqFr5t/vhNg16Q4JeJV1UDbrHWI1S4WqbQ2bvGMmgXDDF/p8m9WYM5Rp
3HUU50RQSKibgMy2F5biA5w6HVCFFaT+tRledkJR7E08OvabufmU6Tbkbpov+3Uf58F1dbKBbSEL
J+Qg8en991QUrQQtMHy+3DHuDptFiURZaDXDpB6tynbPRIF0D3wVidY2gCcw5f5ndY7/rdGmmSdk
thql0yLu7gE47zt9AIcE9KWfYRoo6dhkZfkvDiSYVHrrTrcZryvUynWK224a/cx3kkJScXTSuUu1
fO4vSt/C2EhRAkn86xb5CQ0yjGR4cxQC8X650zjJvvkGH+8Q/BXVyOs3YUzc8fv6pM6++lT+jEj0
un7lwHsbwHxgY9aHW2sq6C1gih4olGW+peuEvarSUBLfnIoj8BZsV6aJ2r5l0G9a/19MX+EHfa0J
ft//SUnm+rz2xRwifyubTQ6P/K87YItVInZPVe5h+6J77Y0Fy6d5pFdDS0fWnnz7D54rZMjIPl7P
OaH5Aq7y5HZV+uaiURt58d7PyNGHXZ/F76dIKW1nhZ+QP6oSGOtXEYZ2KmKkb3/gmzV7+0jMDDNm
CeNuPfDdFdOFKiUPSHbhs1gBpoVzWKdduwxop6qif2xsl6nuvlMSU12wrMeLTpZvJVsV+xqtbIbd
ZYGM1KtUhCSaTM7jvPcA7RU8YJysN6285DyuRr2NTCngjJ6zdGLWALLpGpbmKyLn0jxQQ4v2qzVX
4eCfaAPTO8bhXBIExwkCoO8rCFlBmzALo3d4AUpYS2ydY8wxKp49VFGFwC7PtKAcO+P0GXwbEpGE
AHxwbYjzvXxMijVa9gnzNO1h5VvCUnKM50yz13ddrI24ayPooqEF1llrPZlHLw346iXiiFLo3pQ2
MEbILkHmyEesiT3ta8mh/xxNsy/ogOQTljK3JzAetuV8nMtcysrm5kNTNyTO38RasB7cz7m6VQlI
h4v38A0wy1JMAHgE8OU53esvLZ0Rd8BU4W76qW2Lij/ot9JYyBEx+RocKDJ28FTKsWQ0rIBGZaPb
xjCSyhT4n3qCR8ZmjDjUGj9ScZH+R/YujFzAljtnd4IraIsF2ygqFAjSYom0si010hNzEsOh8DZ4
ru99kXaBugsfK1iHowkGb8PYF4X3DAaPkokUcrzK3yp7A6rlpIG4P/w8gGP+T8NaItF1vQ0FWY26
MRQe8bsIb/I9yo9p6rWxLZ/RlWLqUt841b4jH2nyW3wbgTjFJNWeIgoIKxhsbEn/yKxgFr/sLS4Z
dlqLcJVJmhc4MK4gVz2miPqan/mEVmNqOdIeZ+xCLzOVcsGaXvI5w4ecF8+Uw/6iDalN+vXk3ePI
WfqO5A4E1wr8mcmdlkxKcdmW9ZeRDQ8Ph0z7lnpgzsBQPQfr0dkLJkMPGevwUKU0fKkK0//5o7OT
NpC9Fta0IM/TOyCmf/2riKufLD04CENqmCPZE0+BkXVwGSiZwVmAGoowaP5bGMy2xxdVgBYhkXns
lIBDwiLdzS5IRcc3ISWZBLj99aopWlLG7vpNY/Lo/wFTfcqdum8jjKhNwTewdr88JXobj0Dl0tcj
qAWSzpjI1XLBkz70owjj9HGCVBgVP1qP5KGhWxjpsJIDm2zodvRUSN7JgPVvVxLG6twZWAuo8mGo
m+Rah6Sh/dACwORuOFlVOZowsuysRLwPspMpABafh79gkoY34AFjThkh6uc6woIst5uPHKX3Efi5
wLqkwxGSDERS6oXaSJYfKNAAea2iXKFhCjXOh5QuVuRJBMxcXqh+Vi3cCcjTNZdp9Zl503yRKjk5
/L4NSNeTRZtKkxSEpHwSCcshlwr1UgvY0sIWr5pEpYP9giF+EVEkD4QtVku9Y2M6e5ebu4UlZCXm
nA/0vio16R+9aPWf51YyNTJYEMe748vmEH6Z0PLTHHZ+stvjhXc4AFXr48hNxIRwkWfGBfy73kPP
mwyRyxjeh0ohb1gi8gjGLkHZmmDpg+RgO8STnUelE9GeWxfNwBxktjOO/trDMQy9+JPAvfMJH/2Q
VFFXfdV8tAs42ifYlzYObZznmzqubXqWxf3Xp5Z9FUq739/wWp9tuN0MuSVPd2ugBn/HX08OZPyq
sTpqQpr8dqLDaieImYSh4akSp/JAYWQeRXsTKsdHlMmMxGI6upkAk9erocTRtsCR0LZMQTfAfmtt
1vi9kdEW6f/qd5iJxurqkNlFW9PFKE6A48ESAmwqjPNZKd1+UicWI9bZjSV69pgaRPQIIpbys57I
swBqPC6GIVVUBw9JhJdWrjWFP4HOTzOhN1FxdAwuSdLoFGtKScq+oDagYHwsUIQEqa25NtUmoCuE
R6wfmp6r9HU5J0zrZih3R3d0huAa911jFVzWeCbz7tBoKz6kiGOhDjjbQb+Lc/IUu20oiXDSD2gx
UuOO+srWJF3sqzWj/tiqlHeeTsdIphuUhZVgJsukofXb6V1aSLZmyQ/JOeph97+Vu3np17z2Mgh6
w28HWKBPc1aGGHubrloIACmI/qo8+O8h9smy1osVXxhG2skZO9KXXXHQZAxyhgLgbFUMjsMltPQe
RV1NCSFjCjyNNBAsWWhgrzU0NY9CWi40UB0R25TgCivA3+7NB51tBzW3BOD7/u2Ag9yjY8TgGtlP
uW9lhltQrMWp6MLobyYUYAAFLFCu3ZuxPwL7lF8YDhIuqk0+s0IIMnEqTZgZgF/uK/B+S+SAHUVD
so7McQFwqw+rua+4qqx/E0pjej3Ba7lRnDQX6ktcN1DKRZR+pmNusz7t603kSzddQUDtikgvxDSq
NnFlQcvWEt691jTKScAzJr5HwEUx5SLLvcmORaJXettQaLsd3ltyVn9tDb6QSmEBQ1ffUAT0Xxoo
NCVgs7G1JGx98WebZ059/KfsCe4l4ZyldNMTbmKLvUfza3WkFw7kAH4xrrbnDZPrBe+RX8kT/hJ8
lekgGU/p9F4OoyFqjfl8Mk6+9EcD3k6yL9V6jCChGN3wsP32PTTSAtmF8ZHHjOjIHiolSrFfjoXR
KqGjDX1aVSMlCly8RtSBlWL43eBaedSVEeiLtNIR9qnwarOLwHkS2LMDmOwj9mlKJqD4DUi3JLVp
8ekXZsmuedwuJ0WkIfGbmNkCXenAy2uRNwKI2PIg7EZE+u1yQYxa2KLRtCmI6LABLGN/Lub9K6WI
x/D6KO/s0DIDqDfx+KVb2PJAOd58WlbRFiE7jWaXPD84bQnen5VOL2Y7s1KlFCp48ewaljFGIcJ7
JKHLI9ZL4Qm/f1dvDZDJwUplG/3NItDPvUg6hRer/tq7ABdXWZGW4u68vnrnZDt/8Urio1NG8RmB
kjfzN+SXSsBXaBtSXspdvqA6am3DmRInlzyRLkXmzcCKDedgWIzQ+iXwKUhOOag4brndmCeYkmwT
XqYoz1D60jb7vs5NLgvjSXGK1OSVkhzCiwXrF41guwNwy3fzz78ksFbpds1f63vcdwKQm57AT1Ui
3c9IYC9eHR9BpeIDG5X1FzA+HPfobnq2faclA1yMJHIsrMykhteeq/9dKueo0CfJjxwsOViLZ+7K
Go8RoiYlAPtBLO0fwpq7Nk35pG6CMRainJQtgbxpL8MgEY9FwvU5zI+heBshOLFFzYkzuJ3iCRKk
lCRXeJ12cnDEqfvTsP7PixnOHqezycKEtbnWw/ZXfZQOk3Qc+zsgqAAIIYoNlVdmcxDOb74ttDAO
9fpodsMInaiP4VTSSuM9p3+3pA62r1hON9UkswTtYvextLakuvffMuisbVA25CjmgApCf6cwiMp0
vCHGFC8KqgbKsI9t6xXPh7NdDef2mJjHQSU3AnK6hLoTjgBE1DKNo5KDo8ZEMtv8T68VTaYglEGP
gSn1irtBqfZkRbxPUAWBw+YMWwhmZiqqM02gU0Za3EAbwP7McSSgls0Ug6hKFKfpW0VfI5KThl8n
KExPNSOKOTqN3e0mPkbo44yTdGQpNohwwNeSsG6O6jJvaalgrY7SYrsPDcnBfXq51HNHhJNVXxzX
Ed4eXiQIqogHQi85coTeEoY1w/zYFFW3T1SvFdTWu+uG+sQ2L9zZGYd1QsArlrajXaiV8aPGP0kF
Yh/oUEWB50/vEWNB1xgSy9m7w7hluNV1R9QmHlxYYWCVuKXHur778gGf8EKiooFmUh1IRVACRpaG
pevuOhx707qK4Ns1vmljEa2jorqhK4IjrSxnAWyKtsSKAoY6aOt/LRseUFJ2JdwIL5MtM8cYliVQ
0yCucDcQSQtUBRpq6zBas44vK55p2koFjUnFABsiTR2HDuF8AIlhTjr6/z/h/Am2mnyffl7tUvyY
5lt+j98+qUBBFG2omD/CcCa6CXkR6zh61zZRPtLBzWKDE9nq904AFtNStD27jmmHZkThrxJbIGjC
EnAPQaaJxnhpLC3JYiuQXwV1KdHy307QNomZCX6MX1qTzBg6vTFkECS4zN2royDnacBXswADLzFB
/Wd2eFDbGfF4tg4XrIaGtQ0efpYJIxVpzplTVOoU4MvKZrbqFJQFtGZHZHeoV+gZA17kpjFMeCAK
AZ4XoYiaT7dBjOZDu4pn4mfx53gI9WgAe9GLOFzJmQQJwiKn22Q86zXeWiGtXcBY7iljJCRpD3dK
W4YHhF8HmyTtZ4vxLRGIcNWA9ChbmnH85Hhs6N/IOVHYriBIYYNhnwxSFK6Au3WhsK8/j7ejJV14
fuBz0tG25itXBYylX/T2lbMIn/ZDpdmppfZb9La2iH1IOj724EG2BRhg0DVKYJUdAVJafP+Ax7cH
eL5ybgi/zwOsal90FncDZ8/Ewk3Sl3Li7+w1R9zThj5YOnZ7jN6TQDxsf3ru21vb3SLlD6g5FIzz
GVYESbiQzOYh0lBAhWVRLuZH30Upvtrv4yXYU2VnJEv9257i9L3P3RtDYhUfoJ7h0cjdHd8BMO5P
z4r5dJONygumshtOt85XC41FCHFgptsLQB7sjPbAgtJvo0i97HE6KjDAGPRtC/OzeSYq1mwWVRA3
d91rL/beicVkSpjkwWFmw/qzXj0iCqYHaHFnQ6oFWKz+poG9LPwJV1THTIMGSFu3vFMo3B/GVtSF
OlKCsBF5ZwanZT1i/TIi7hsLhVOD6tfjFxqbwpOKlkkhLl043TkNJWSQW3/W/xeqw4aW8FNr6b6J
Hth5+xN8DHCx+bGZQx1UJ0pz6NEEYUYmkNyM6PikWbQx9pPsph4tv5QRMspOmeZhFKJ9fCSKruk7
i7FjyNOaeBPBeo/o9P+9XzjgusII1pOfAu8u3QWls9iEsWmEt83boYEVOOEcWqelkVSVewuO3mJG
9ggrHHb+zztxFoWa8fepzCU/B56tEUbahscVJllt346Z1aANwSHszavwRi3bv2uk59W1mGUsCFY0
kUOqCz/LtvCxPOZ4gXIkg7fHu2tQIBaeY0bxMurQqzfs5+IAUVPfor3Rsp5NSkjzELvlyA94ZhWF
wswcFgt98ITKi6awpWcqcyJ0gB+4GD4GsxfL75wqn/Uoh2R7CdlfWPflHKKk0BSqJwbpe7/pkSVB
zeuWIb/8irll9zZ+UdvJrl5L+hRn12a6p3ESRgueWOaz8j0JpY313Unb9g47l30YuqDuQKNDuDJc
Mqdo4Phf0v1+lgzjP4//LfMXIh/7lIDZVb+EhIbn73DRFcmLEo7gE+Zgugsc5oNX7wrVg2iCd54e
+8EtT11hfdUhoMGzSqxsenAjmG7+/CsuEkk9j1N1mSPvOoI70iHmoqdcMH+6QSJkrPqy9/3iJERk
gh4Fpvi6xTUpwSFg4FYCIDdKVjqOeJ9Thaksp8dLpa2iUyl5hREMmWvRONcYzaD4+xi1OkDjDpBO
tzZY5SjiMgDuMmNQMO/72MUiPV24wVJhMnVGiUuC/Gywf4h0p9dQEe2UX4l3DMsdD4/jcxzvfLVA
tpd8lsfOLT+eWQdR+7ZjcmP8uVQv5fOZFljQWr7L5suaQmX2n7gDF2zj+J1xV+08wYyhGUxTSbgP
0L4tLFK8WYfo2hSERaB5FRHs6nkYeaz+9VJ0cL7/dBbwQu/2PVcvv8oFjMrISpgv2rV8aXkUK8JK
RUxCGVseITWbqXE+J84bhRPWjbmpEsEBclWYytKUknNyt2+N7mj2UvTndBcJl2dAYVYkkGJ7JDbW
DjYSi/ERGuQhwe0aubqzFF1owtrCpBd7qvesV6BfNEwLhFJt1uX9wwaBqfn1GLCpnottyYUEKJVL
D5iy+0EplbxxYFwBw/OJWz+Le7c9MCbbmQs9xAif2+RTlhn8wFdwQO93kSuSXR96UwOBCWvyyt79
vv69sfmktnJklRsQiz63Qs8LS/EhnpAtsu6MgWr6cIA4IHINlmpPKQSVGZPqRJh888f/OtnYc5T3
h1D2pXwbxQEsuMr+QVCSo/fzsmcJ/FjDB5cKPNAce74JcuDHHQi7N/9hBNsymOW41KVkX1I/CeAy
SUbP8C20m+y/+cNou3+mIjpko8fcqSE3dM1sBHKZsx7cKB6p8OeTh1W1YdN1/+D179+qSTUgtyWh
5G2ilt6VBgr1PoKKBxnt+Qw3DmPC47OWv7px62Y70nknmsz0Xx2f1jtYdvggdVGgnLW0l5mihgZP
hT0UCoWlPKz1efDCcg8p1kjKDKGJCqjv0Bki55t2P0pCrL+kmLhHzAwWRMS06V6ftgBrP7tC8bEQ
Kvp4uNJi8KTCnvANVapqh8kLJJLU6t2atOOrMyk0WBWCEjqc08c3VxAOP25CHIM7L+1AQoodgA2b
hqe9MErQH/BlVOWRU/IKu4SldiX2repNrs190vHtMJ591IuAJo9c0C9hrqLMt13EoDLG/7ojNIYs
q0OzOPDD/qErC71JsUZDpo9DJqdiK4jgEcbav8q5b8Iwy4SE9gqguQZs7gajxTjs83T9bpxD3qRx
Po3gJM07WL/nD1D1QYjLl9w2/kSFQVQecZJANKfLWeWixBW81mNO2K34glgj79EmyVMfkQibP9nk
px40ZCAgV8rxyycKv5uC2ZStu9gnxz2kA3SB0ko18AN0FGiEAnqW5w8lLRWdce1di5IEyKhN5Qs2
sXjkg2ox1Hv1VtDVlqV7KS0xD9i3vfCAFP230hVSdu8EH2vCq9u6wb9OgL5017FNPoNzDVqdx1bs
J34fIQe1dagAlxr/WRdbjR6TTsCg1EU+f1WlbZFkv9jn/lukdh3OMhzm/IWib47sphsP4lI6HfRr
psC9aT+Rk+ahn8r/NsacJ7pfHpXOQOP/4bYZrKWVNOPAxMqsYLoQshnzHSoxmxx25/GAgFQnR0dl
U49lnGlWQJCpq2DJSxNNna14vltRmwD6fabSqTTMtCwspfW7VXUYgpWG3pYQJ120SpgtKUMDvvna
wEeupSZumX7ElVT5ZzxLJvLWE7EnxpCSojHovu9soStEB8sr1noU8mthdikIsg28gyXg8yL2f6m7
fXzqyk47a8zfS+BsrfnKOtBUhLIcTo4Vw1XwP9xU/Rux85+d/1Jy6zfohHszmb6xh/pKQNmhk/tz
VkEVQKBJnS+g7UilMPqV05oVBCWsQnO+/8bsVBGqYAGkSWtFVLqY0YA85mhXLu9Z9rCriIrZyxmJ
X5e+vf/AxyvTvygjavjVh561qRL1NPEHu/XEGn2vMd5z2iEuOk0OVj7QcPeL7+P4Ea0upNK9V+HF
MBanM09wxQoc6ssHZnI4m4xgddrbMk1mwEsQM9IOLoe6oR2eIyzIqNtrE+M/qpZXyurynsmMlAg9
7wvByA/hX/z+gD3MO6N7Q1Mswc2slXG5zXS9UIZLasqw3Bjc3dn4CfP/16kpYuaHAc4AxHSSurtM
L3bGIsslaZabaT1P01PF337YFVGxbdzhYI5KajOreGQM1BoKYW2aSM+BOy6kr2cJwZRAsgZj8z0G
tPf9gp5OyliiOQ9he/JLZt+C92qZJgGI+hejCsjjgQOoMrWK32jzo6QOkrbwoEFKE/LUFGwP/bPz
e/o4BCckif4bk2sXjIXaOurPwxJrtQvtVkRcwA6/Rl8Np4UQ0uxp81jVqfEXPxbG3Q6tYofPIeaY
rnfRTOVx1B/RBS9xFqgVDbahR2I5KjUZnW2pYQExzJo9UxZfB0vBfRB//G1qGBffhwqVP2Du5/OZ
FIDf8ba/H/m2eeytJNbmlKvuvZIUOGT9x7xCLLZwtEtC6U3K9xeukAZ9n2aSDdeUd4LBIkEX+bDU
PhDc/CzIDpCzf5Cq1gQGgmUUbsSkosvtSTDAOF0qxs4ht+7Vc4ZXuP+bnOOqcw+fpMNE/YvTBN/s
ZGFwuq+9uMTrjAT63meIMDqM5ts8kvyZ9TTH6HOYrj7SHKCVs0fb0NcLs46OIpZW6H5pAAxs02uP
5msgl8QqpK7Rz495elA7kwkYI+YXZcqh8UWyv72N6iPrzRxUKLqNJ/bsjK/VL2JbiuDHJ3j9gJWk
ce2Xt89QPk6Wnw4i1VGOk/gJh+4j1/XnzBUWUYMpDaWp1sAhoQem8eZP5D5+y7cZms0Wbekj/B1H
CLYtmwX/G1//Up7bago9RG60Jd41aYly3m/buECXDY2zC4pmQDByD1Wptlqg6lHzgFTn9Xd8M7FO
1zhi8pALGzvMevmD5eDxWOxmIB3NLTS9n5Ri+GS2sj/UUMfu7McflPbb7hmqUwAHyqYLqVzjAFXH
NsmpOH+Im6SJvprzh/TzGcF5ertzvzQEE1S6iJdORbp+xD1u/Xv7YbIg1bN7One7eNvxVo7lNgba
WTbQTo+dSKipdwCk0iQ7Q1B7Po2bTeN6CkUhfVnxZP19tkNPJ1XwO2NylBwro3twop3vke2q31TI
6RHZcIe6nfY3ZXkKP1GO0TF6BpiTkradwrYvbh8tKqKzx1RPy0AUk1B6fjhyFaIXNzOY/In3Ej4q
E96+qNNQiHSETdSXIsygDAEG9ui0tdxuuULyMS0HEWBqDh/oFbKxDPByVvkwHrJm/1XemibtDaJX
gIRZWXudcNk69pRfAoXw1HN3gxmow9Wj/gOdStL0l8VCIcRIY+rZ7RAJbej4R6Se7MfhbZTa+Hgo
lYRotuOxkfWXfTW6thlyV0BH0gLufteaMFTuNoHBy2rSM6+PJBQs+eULOpX6Y8I6sLuSTfBZZJVY
1HDVYN4jJLkxi0f3g2Xd8kBTDjGnnElqB5MGZ8T47BOxSk4FtN4xcdezWF4TYOYJm9umVOa09c7e
0aIwQRqjjwhNF2BYqj3J7+vfmV2kpGMyRfIJL8lFX7796uCSNAA1ylZrWVMZyt+Oixq1rSAu5J8V
ZVMLPiZGg+lnvjBuj3WvJxGhTZMeXyJXZ7Kw0FUF8ETVQL0hNT6c2L8ChAdGYzRXtqsDhlRrJ94A
GOck5jNYLCgEp0rMLy4EDmIniApkmok9k6zM+euDXayfMxRioZj/1fxbWPywBhK7rHX7K2gmJ6p0
DqToWrC2mAf49hlPb5q+Wr2pagpTq0VaERMqGPcHcOcij9Ibh/HhPWcUkL8s1Bt9VdX7mgsJfFOo
WEY8H3dJUJnHYWASfcZXFoIFfYyrJnnq9S4aFhDSeyaGobkGaHsNTxW14p5tad4uYwTIcu2Dmf7q
rX7biRkYMl1fgkKV2h/js0pkRva6zKPk5moaKFsvobCsDw7IPOYZ61ASz0CtJQbZV1dI92YFSZHE
j+h1UE4FqfBnqAnC9sRmmeqIWWR8fFkPkmZXZBJr/Ntf1ciob53eYWedu0IbMP8nz6wJA/4qi0EP
z4xuj/6sP8387Z0xcWpsnffZhIkxmOd7wLcd0dpemPlgJr7EcLQQ0X/6TqlQoNGD+yIn0ILj6M16
6719g+XELvdtZxzf4ayWDk7aNw6H4wflmvXab1VHm+wgPYbDhy+0IvDxRJerSuAxra3wcHCJqcRg
2duqwEKjX51dO2AcLTClZNoXco+s56EwUiVJFIlY5NwqGXIsIc6Wasgb2gc5+nGPQeNngsqMXQ/8
aanIEgSnFPOcjGoKGNpz0wj5JOSWICKco80s8KSTruM4elri4GO0dA+lqvjJJD7l2H3btwoqyoCB
II7HFwpMFK1N9gmOqXuIfnH/ahX7CP6wAdjzksly8DePQ89+cvWwiXJepeRxoTcRs4/x+n0la3PX
VdMBIztbELnvxy7/2/bW+N9G+9dD5LK4Fr4/M8Uh3MLno4av6X0A4FO0X4iOv0px0AZcoDHr6LxF
gf/FH34V1/6z2BiWPeA6eV3FYAe+KPA36aarykfXmgVy/o87Hay1IUV4+yGhtNng9tuCLlpY1zay
HTAlI4XoSFKjV+yMdvLacRF1b0caXLbEeZTVF7xenlh6vzcUrU19azaqI4bGbBTqW+V9ThaK5Vw4
pXSTcRfRP3KthsHKpQduPpl8+NHwqblnDeeQVv2yWidp3M8bzNPySpaQ4fTK4KMN2wq5r9qkoIbo
krkWUVDqXUmZlNSVkEFJBc34ZgWgJfw5EGdiTJR0P6UdJ53YIKcRbzJVwEmPT974I3tKDdddpHLG
4DcbWP3NDwyZjrw9TxOaHcTP28jOylr3RuDxdkEhNQOU59M981knZyaue+qTlN4fLpF+faE4xuhA
fdo7A+w1e8ebWiR70/GsawpR5zh0RGBcDMgsQ/Z4s3renOE6UNyMvKd7GktzrYJfUNQRGnVjLB8x
ICAZgVQ3JY3c536aVT0r7GeNcHY8Q75G4oJ05H5OIk1jljqS3YBuIahnBKPVe1nMcUbRfHCPi7FT
RuRzn5kzDh/W0YWQo6YxgBi3SXLyCUNBoD2f5gX5qbsT0Q172eiG7IlVK3+Jt/lGvCQ+jKKD8QBZ
SCa6y7BYs4a0b0CZqkG5Gi6Bk5NkQsvdve9aEMo9gIY5nGn8XbwTpea7Xze9FsYG8dX5lQMIvpCx
Jro9u0XuL6Nn99Gk08YpPnrT4htMi9Gpm+EPjluJ5LlDGwe8SOuFrai3jQfOjfzwu4YBzUMi7s/w
SyqDgYxi8bHYGAIQomd9TOajNvH1kj+4XHXeYbQVO9Hva6EpEvRrMlt0bMEfrSxzLwyFDtaZi8Oi
mSZqJ1GfyfdoJK1kt7npljoJ3myFEDL6RaKNLvSFnGY02S6JuTOznkk2ku7Y4Ll1kZhirX/9c+XV
dfqcMqWUvL9gdZNyUO0HDa39losYqqRABR9IgytDzxvNeoB/aLFCIszruLxPYRctQvv+9A6M7s4N
DoYYnscDlX8Fxf9ai9ETggcH/zUWTSupRPMZ177PXoc2ltTxzbDMxp3jS1tZnlxL/8/+Ptyax1bm
f29MA+TGGXum+lvUFjUmboyI69kZkK7MkXmgrL5m/gNz8V2XtprQiA+FRAb3bUxcaV9V+2Et1lyC
CCIKzrIu7V0Ptml+l5KT2cLd2/Io4wAbFxTpHYi77ixnmVDDg1W2CHm5KNBAIryhQp7ObhMEoauu
HXHnZPypRGS+uF3D0ivsFiekfxvrWFgJuZ1MRfqJSGHYpWuaf8Pd7XtUupVSxVIyRljSqsw3wnGx
KjJ6W5/0UtFvjc5R38umCOLH+pjd3CgOw+MP7UBYOgdS8UIO5r/brROj9wKZCG7lgZIFCJERGHil
AVLtZSLuFV8O0L/9WhI25XOxCLhcPVcSV8syY66TdpghbUSLjZugIDadcLyPludiJCxz1aRAg3H4
FD6iJVV8K8xVXFuSmaLI8qxYdgyxz9dXRsUhr786TNF1mJyvy+SC5pr1QUQkCdMLFIeUxnYas54b
K4bRD9FW/DHKJdnBGiq1NqmohcED8/0M+xsxVGEgGY9aGE+jj3bFX9WRQ7cN0Rfx+ZycossFmcKb
NmwhZBBqGMo06ppo3g6pHvv0+1byaQj19N9IYR1+N9raj6LZamln/od19HazGMSF5D29T6M+ymBp
w7prAs7pm8bhkeAqgXlTWT2bGLemokd6SU6Lx0Q2AWslAxRW+JkNbsE3mnIjiAhPPhe6uzi9BA4w
hmtr6un3J0KNpv9NnBPkuR4tlmsWa807dsoRgXeof2xax3feKe9pNGvy1wHJt2jUXSd/v2mQXB/v
kXj2rH1Ils/vPGgb/Rd5Paz1YMZEJtot6Zc6lZItt/rMgHnK2l9FfmVnnJt2/SkiFwsZ/GjjmMyr
nmmG221qIdL52548Koav6WUXDN++jPWyqN2yD1ZhfVn679c6uQO3++14Gq1LYL/kfhzKV82iMDRP
KJcvTftaXl0dcpBCpO49qZC8lXeSkIMbHTtwUxA8e4akiq2td3/oN/EyTaCuTfUkWdfI+dVF1+Ix
RCM7EEaXgaEyIb9Tho0kLpCajE+jAkMS/j6nEbBpcaAawe2UkkGcWpNZpzzFkokRHSEdC2Q5YgvC
N2fVbj38GhaXTaX9G6quwlhbCtS/E5+X0aiZsw2sNDPbhmzHT/uA9d7YIi8qbWgHShShiFStpH3q
VgREVBwOFi17vCSSoxfZRz6QPX1otCumd+/6ERfm5K0zMvzCF9/KB5iOANmT40iI1KpuvEXvsqes
sSLnIHV5RcM8iPJGIpvPW0hgWlFtYRJJ3V0DeWiNTFScglkVuErXC1Wzttrepeym+zG1v5pQubBs
T0eLxhm3R/hmf3PJgzllZuq1Kf4BvWjDOjqtFHrYxZAr/kL+Ro9yOwbXKGpBtkXaBKI6sE1S5zHh
HIvjPa4uf6zx5MdZLq5p4MdbJwHQMeQBg+AojxDzzShASQry+6cVPERe/cY3WG09h6KYnqAHx904
la7FdlSk1udV09dfLOjzL0Qw/3IHEvjB4ts9CRsKA3c33USXcENaBW9tF6yhfJtBKeqw/pLfkh33
Wtou5XPt12B7gDtCEQ886fMCjfEe/BX2zjkw9SHXIJhjiQ0uaCRyZnftF+yV+9A7jnAjirr45gpT
+YdI/ZJ78y7OS+2969AkV/L9j27YjtBKf/p9PDVaVTyFXDx601lAyaBKER+x2JirFV1okrH3Nmzb
utG16TKo7d+1R/mZEOtJm28FirK10iaybHQuaB1krMiaOUET3+9yP7iYYa/rkbA+nqGE64c+NOih
/hqWSFvZmrXNyjTPMqj0GfrbHSMJiMtrJsneeA0N8VSDkpIIhGb7QFSGZ1oGuCSBxicsz81/Y424
/hD2a1xt1t2IY5KcXUD3PbQKHX/6AnQbKcvJ4um6Bvvej8Bl3dB3cxnntaM5My/z3qm6nZvdktIC
EUwMVjq6F1c6VpA8SrPCL4Rry7V6gT8GmMgZGsF8CQ35Z/CxFQzsOgNQcW4fyva9TzSNXrU7J9Fx
Zo5HfsucnMtREkq8MnrD5tV0Pwt6mdZT0ehDBvyF7Zu9rkyQFAeVJoifyb8tXQkCab9X1NVeKUCs
ki4dBuBcgP+AnJqQmcNoGXDQuUrtLG63pPJtHWL1c5ctqmHcAYmUTBjN28kRnSeAoUTpWvpoQoGB
gtYyqM60hbJCDjKO4wUn6nyPVSgL79N2Ciya68jHf0DXPGxVZJ5I05a2SaCu7j6wliud/Y59KabG
eHEN9So8dRAj7BNMZ5lZL+B6+0SBFv9wiJUfL9eT+npMkIbxez0KUfOUNbf8zc3swwcgo+MYdIeA
8wWwAkwPWn0TumFx9cUMkMAqWfkIOBeS3/LqofA2GuPzHucQKh8LSnt/4LzZGPM9h52PlRqirPWR
mvjSLs1RC68ssxmsJ/C1Hr8IeJFTGqVN/uFgb2yLbXOs7YESYEH3BmbpF1Qf/oKJdO7uMPGC9psc
2qbENeyDW7xopSa8mWriqN11Lkf2xKhj0mEaZ5SkhPiMWLskksjznupjg72qNBaZLyNLFCHsNar0
E/4XB61Cr/QA4zMQ2E/d4V72weC/EoZBl3uKpjeSJYrcNWBzho5IV3Z3WtaM7KiFBp2i/roguLgP
IdhnhlHVLATvzoJ7ESuc2R8MDbCYoCUt+2TIROqF4Wgo/sEeLjxAESTnmZfvoGXotEkw4IFhJ5pj
Ev4yVuIhjJkJEgxR5Z/y3nOTE4UxuysdUaPOzRMVORWh4l/BDH+f2X72zMCgLDJ1GSPAXYW9+lsQ
xXKxndFydTfTW/6N8j81WfDfQoGX9seArPY8HK8yiYMEuxUOtqXCO1Twa0mn9mvesdyTYlRhhhN5
gLIv80we339w1hrB2vb5Yl4+9VL2xNbZ4LDKSaZjHW5wu6Zki6ozulMBw670HHNVSId1uEFeF6wP
gEkg4oGI04hT3ZL1G3NKN6TYtDN145yqc52GTRY485FgiMvxmIEGYCYvks0LQA1ARc1mXPlhbNW+
OeydXvJFmsjEOko8c1OhgHU6ORWTfrSYUHfYzx6MEBL747YVihfk0fKFqeqPRXY2Lbftu10utLNy
Y6OeNsX02Mz4hS/Z6pck5KsVbXFoTJLaPetLr41FpQBk3iFbMlGVthVioj8zdWJV23urXsdN0ks6
fxPsGTDksdrVorCb09aqs3ADipWPjUEO+nDA1R2pbzSktJnqRVfSBjYEroar8fPZ5hAUkA+h2Da7
Eq72yNJ79F0eOEnNl0CdmaDREm/vnv8wyUx7NLfE6C/PNtp8y81bB2oPKjDQMBn3M2cIytw6YHER
/XHC11zxDWAE6pcf4W87wFPXTnDwt/3F+ly7kvDrx3MYM+UgdEzuhwAPCRdMDgpp9vk9knFHzfOv
uTV8IIkOMxUaOYzf+MqETZMPCokkuZuvn0r3YZHwNSZa0nNwDzwWc4WwUOGcaMiZlrAnruiuoPCA
xCvzd9p0cnEsvUp6GGElHUtPfqS0J9LKDExlLdy48UnpJl05pdkZuu9iWNdC6FvC1rjNnk+NF0ht
Ct9iKK29yQ9pGMnLZBkqidUQtrSpcvFKjHvxx/Vtq0WaM3o7AIRKGkqAcJbLt8Woym+tVWZHO5AR
krYsn9CAkbxVtP/w/SsHmxYml4OOQLvLX2JzZozmJNWtqrhezeJPb/mfqHK6pGMlVDzDTzOn3YnS
RCfSZObvsN4XQiY+0CNpgzf+si2RIwdCLNr3J0pHLTfIJwigv0012ThspgRy2Tr40YemRPCgDOdS
HLNMS1sVmuow/whSJhyGLdJ4nbihPxMuSo/8lpk3WsBAumzerz/TBtOUXwkz1xEh7ui6cddbB2Gb
neHSq0lsNZ7l9ra8FcCZOCDTtgKRq0ru+XGHR3tTg5Qv9+ClgH3yzDwTl2MFBYxIM0LUuThcFA3a
X+h6DuexQW5Y9f48Rj/0xEhawfPIxFP/n7w/VyVYP3WqjC5clXjYfnDsVPvIy/Asanw60VnDAQbe
R1KTVn795fer3AsLu/dF192cJQeQKot67CMky5pfaHUnhSg4Q3mn3c2QmVb/tjYLPj3o4ON9Lh2C
ytMm1q/50e9qGXX80M1HZCT6jcWxreG320PbZqh3OS5IqYu3Haep7IRv42MuB7sgwsGyoBV/DykV
MYoPQEGl5nQJB2GhHm4NJq6/8M7VdkCFykBaOk5gciQAqrji8T3sP5JdVA0yiKzqntvitqoBkKT2
1opxgmiZJIE9q/wuxWhkq238WuJXnbowh7hiOSSRTWQXcIM0g+eJt2eCNlZOAxpQZNFhxBZodKPo
9mQkVxqE7I9mph7fy4igVxFPWlZgJ/Pz54LbAHO0Ts2xSVOaGzSE90PWl0RrR9z93PcPzuoLLjPu
g0+6SpzXOwZvPj3JHiSFAr37vTfFdFEedauZmZwHFHbQrvRWwOcZrksMA0IPP8XdQr3RBh4fCCYB
QfvGcabLMUCmV0T8CIJB+YdOvQ5NRgSet2PijJ4D6ZHVangvgFL8Vm4Umd5v1U0lxc/HejeERdjn
ViKD22UqrPVi1C0DwR+SV5tiEt4Hj4YqCd3dTEe9daCYemmf3K1vRbmoAmJrB2YIFwXqKYXUqR5P
C45BQPOuR1bez71qmQ9YEgjkiYX+nUFrFY6f18MIdeHK14j2E5WAnnCcud7S3mabpl7RgneeVlF3
Uw+jRu8ondFFFB282ksEtupnO+o01OOenUjjBexJAThB2wTO52YMEiRIv8jpGVkPkADEZJxbHACn
Fwy7Pel21V9V5Ce/7ZIKHQRpVMPcnuLU+f5zLcCZAB3thtjN6qDlTCv8JuR8HrkNAK5RNy9yJBmc
Gn5fNJa+okJbXD3fx8n/Vs8NHqBCiCsY2mwEZUGFLD6MMgMy2w3kbRH2HLbuqjm7jkgFeM5WCT3p
pRjr8uRqxn23DYR4gsLAr3E9EhpBGZ3zHl1FIMpRvZTdDaQ4d5pJVz3vT6WOQ0LNF0ptoPZXUxF1
h1H8o1DeZB+lNqB3LLmYCjnegc6c1ZgSblE1kXK8lrzJtO9hbSZolRAXT3FBdgFl4Cbm1KYWMR0d
xCD3YbBw2D1YlXRlEEcMF1AWa5dZk0JwO/SG0Ze20ICI9/6A+0RkA9OU4bG9noz+XigIfNY7M55T
HU7dVgBCUt+bRkG3BhlN6XkanOt6N0mVqYV58l68gAqoOS2IRjzBWtrOHoj8NgO5DfvJdAtbpx8Q
PvLlrnrbsM6k6M+s2e8kolZUiRIMRZj5z27AmVunqGyj+w5JdrWQEX7PO2fKcrr54C2eENt03RuH
3F+U1iIXogKjuDAfumywVW2UjhltMrEUpJ9ZbhzHBqlNuXr/c88yb/12aG72tC0rO1BEULgEmbYy
iS6+JQY0JP8BN1TyadsXDg4rl5ucWUheRSmL+fNK8p7RPHkNadsY0I8s8p4BBFJHfIrkt0BoalHw
0hMou1Q7JtafCGYYZUwoLjF+rMXPurUkWYPMn87irTpmyFxWDCWo5vhNGHsorP19dykOjNMzXbvH
5aIzYXuys0YttYxQ2lr5QdU4WsQNKT3B8/qmsnqOjwx+yeIl4033EnAMUciXVfkmdWESuKWO6KNi
paTUNNIMH/mo4w3rToXnlFL/9japWjVW2OZn6yJs1tZmftUA7MdmkaUQJ24ktuXduGekdjFmZwY2
xqR+q974UlfHOJpeLOMqZm28k6QyyGXiynVNswVppGjP01jiyCb30txsvy9jhH6RT+Gu7VyJWq6c
GscUJxJ6nB8tirdBDzlC9hDerhnhx8iRjjaP+KIfX45mVz/Qy18yzBdUhqS7sGzEJdjUOEtncw6o
e4E8qZMAWYcKsE7NwsKuhX3f8FjUPqIGx7+eSG/d/MKruI4hGWr64CcIePV+HJcN3+rA1dEmTJNk
ldGfxx3ot5bAWjWo0c/zx8H7RAjVie2xHHBCimrw1SGFhv7PknxochTNVasPsmq5FJ3mPA2pmErQ
1QsLb3XOzyMwK8ikE+Hlv4XynFiyweYsT06eP9kIXU7qJOPnjTOkp6cHeqmXrrrBoowGEUKJeijR
j+QwlMhx3mxyPMUOcDoNGzkq5Ff45s3ox6mt+q8xuU/M6/ElvNmhogqOvl8yv72MFWxYGGZeyGzR
pTPPCQPvcgTSi2zgIg+zXtOYhUmMCvAcfkrI0DWJ6CoTipalmQgXqjQW63RrRBP0oN5cSq+Qq1c6
3BuwQK26RlSG8z24ga5v/B/yY+2BSsnlVbGzueSXvt3rf0m0j2kOa7HoftQeM63NK081Vf1aIJpj
KCv1MbPWsia22qv7lZRGuJ0IwNCEOwWClLhPYtwLOPKm68B7J3FKQjRxG3LJnsdm/JQRyEgUYIbT
GoTsdm7TAHntWCOo+PaalAvgji2BOu/vmep8PiY9SgQhBzORKVpmsVGLfN/uoaVvxAgqPWl3+HVQ
gonUR5iI/q8H+ZVOGMkVvlQURkaMt2/rafaMCiJz3UKEqvJJsk37MQrmjyd85gee/LlN/P4H7+4X
sDf4PAu7vB4g486TBq1/AJzhAv6xuHrk5c/72s9QRmdHT9kdNv9p64QjCrgTBj1VjNYp2kuHn219
F81spSvSRVCAparQFBWcSWnxQNHN3m5jF5PObH73pLpa1Mh0FdSAeOwOv4Z/Bd9DAD6RTjMk5ti3
aYBf9x9feBlWzy+vXYxnP8do7E+Eyr6cttRJRVb/GXEfMEWtRC/4YTJcrCXVZNu8gOUt1HzOGbFC
dmfS4d5dkiI8u424CRZ0yre+CQ3qcjM4qaWjx4CEAg/fOFUFT3SwyMxQqRNufy4o9v8/sy/W7fHC
Y3VsOa8P/dF5ZgXsgjk3wwqdkmOD0jZBBImGHUBxNgKobRAYrp7NUpcZVNScxyhmeVrFt2XWanjW
58tjStwDQ18fP3KlUmZE/voyhYkzWQqdqlAABT9kGK75Tp7XAxYAozwtdk7MnGLWtL0ZvE5Dubu3
GAbc8lFUoS+nlaQR5I+8izoePyGyB7fptfscEYFGAljK1I69yHj1u2yfQGqVlVBstALjSyEhH5tr
uvoeyiyC8oWdV4KZmmNhcn/2ZvWTjRYPhGa3W4NXou9dqgKzChe/1TMu1FGYrIw2d5VmLtXSS7c4
35whEG+u7DDYRtNDMLRLgXHffgLs3yfXgryMwUNntsF5cYZcxSaa5LBI9aEhhr0bRg7Tbr9FYDkb
9J93UAmvELd8Dar35bxeEMJc/3iasX4A1vjSj2Pg/e3KGAzMYuv9/vxThYvtKV8SilKcsBj30ECJ
RUb+WxfXN/NGkxpxb0KxE1+kCPa7EyYY5eZjdQ2+OoklzGaEQCsjStGGFUV6WzoUcByW+le7k1LB
hdZKX1+D+t/H0SiEKIg2Qkc4IUkWhsM0Fd/4MT+dIgwRiebqkTlKs/7o44B/RkGpfg1ZX4Wax0D7
h6AVSWa2XBOnONz0BEeUIMz4aMdDA/1J7Dg5m6v31ts3FjiI+umgLqYfM5wpUOuN+7uk
`pragma protect end_protected
