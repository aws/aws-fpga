// ============================================================================
// Amazon FPGA Hardware Development Kit
//
// Copyright 2024 Amazon.com, Inc. or its affiliates. All Rights Reserved.
//
// Licensed under the Amazon Software License (the "License"). You may not use
// this file except in compliance with the License. A copy of the License is
// located at
//
//    http://aws.amazon.com/asl/
//
// or in the "license" file accompanying this file. This file is distributed on
// an "AS IS" BASIS, WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, express or
// implied. See the License for the specific language governing permissions and
// limitations under the License.
// ============================================================================


typedef struct {
   logic [63:0] addr;
   logic [7:0]  len;
   logic [2:0]  size;
   logic [15:0]  id;
   logic [1:0]  resp;
   logic        last;
} AXI_Command;

typedef struct {
   logic [511:0] data;
   logic [63:0]  strb;
   logic [15:0]   id;
   logic         last;
} AXI_Data;
