./../../../cl_dram_hbm_dma/verif/tests/test_dram_dma_4k_crossing.sv