`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2024.1"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2023_11", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
qJxYIPQ4ox2OXrpSKN28t5hgVHi4rlIxxv7eFQ8D1YNZZl2ns/aDLQYiuxYsm2FOpAO2IPzQbuqg
M5xPjRX3noQBg/sd1mn4VbgOVxG+6cL3vX3W9ah4FWTgoVidlJabJfBXWiuuKK1kdt+PC7lBWZev
q35pNcczQyTIEVkBGqSL3tyZHKuGVKTJ9XP7KL3ap04RRVoPERP6WCicjxRHQD18yDms/zX8fXP9
btORaaaOrvfswuqz9tRmO/+Kbmnj5+8eTz/1r9sFzkqQIfusTd8S5vcBqSCaWy1+Io4IrVEfRffG
YNXap7UNDjuINPaewooIOl/wxAihgY33zt5zSg==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
Qe4Zd4d2oFwg8VnIbboSdF/ffMXPg/L79jPgUmsKx4F6Ljggo2DVPoZFQiEv4974b2jU7bsY8Ii5
clJDMNmcsZv3kx8u5ytMVwB/8Wy4bfoDU5oJecfVOvpPeJS6c3Vy2GD4vdfF1g5ToBydhx83ogI2
tRlOGkvJgr53vj6l6X0=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
X90YZGMXtkIqvdGpzSZe8kaLUZ3xaH1HJrIAQiK503h0FtdvaQCJdwhHEg61C1qJwGtOigzlMhm5
Y/AdueNl4rr38zP8KHkug+p4A3vPDdF+7mTp8xVEM7911AAYmNzTf8k2+jG6M4pxG4uZOU/B7+yo
pJzR7sunWim8mWqRr/c=

`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
IQYEBD/SwWlkNTTZGtA3YTMCfzSNC/OcHUQbkPCk8uU+WkxsMflJGEbMwNYaPHDx46RJ/8/k5yRN
Lp4Wz+9MdA==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3504)
`pragma protect data_block
csVDCIthbNPm1RdSjM83ih9sFDdg4bjfYdwDV+/CeDRJmmFMt+oUlqnnO8i9JeYlOxVGaTfqtEtw
IrBFCe70rF+sjOviKxgdFibasA12bGf4553kQs6/u5IfSxHM33wr6JPT5R6yCNdSdSdcR9dJla8i
DnCP6WF+XhIM2KNwACymn4WV/fo5gwVtZa05Roeuu39hbYO5T8wIUUhmUxQanYViANWwEImufTF0
Ikqi5x6cBKZ5tBIi3tmMxfAFbjXyxChG7xwLAKEAAEJ3Y4bQKu6zulgQlNTXBw9eUuerriWPw2Y5
qU88/rWa8sxnnIV7f+yhU2f0M+UdE6lDtuhtPt64jO4SriSL9ou7Fb/YUyorfTVp3tT/A1B14gtX
LQeshChdhEYLxb7ruZuk5SFwoeSlL0xsi5jWhGIK9Ci87to5YcdVGhkZyhiV6KLSdcwLGArZxb9v
u/7XdQYKZCGjH1kUfcXv7wKThGKwYq695YDX7o3pYEndcjm7GdEqRFwEavJ4SAHgQRRxVrHOm4r2
Td9ExA3t1+u491KaleNwfBt/Ej8qnDpRLoMH6c1xHUaIh0hDAeXiLOE0gHaJB7+7yr9ELDMfEGPU
hjFC3nPbJ2hOfRkX/qphPauJETuRtoPldRngPPPHoaUVjs98yWqUhGegxgd7eYZSYsJGI/fKL2wL
TzNQC2fC0Hi3tIS8JL5vp3v6IOPTbb+VajRucSlp7UdV5M5eonmJ9tyk8l8IXHGROuO22q13AxuZ
KG5AeS01wbM/Lw87S4wiYTx1FJGmRPbc+2ppvTY9ruQOKG5Rr/KZeiY59YpJL80zG7cFokxdg2xg
hBtNPvIIjFlqIYPfCDOznRMiS6XUDvwg/zmIFvwBTk6dRHm6iDJ0T56v5cRKB1y2aSNOj9lt8UWr
PMqvIaahSi5QIHBkAkTFG6R3HoSOgDuNnmJfY35acwCaMOTdbjdNo2lZTj3ouZl0U7tb7yd0Htwd
ph+HdVDzJWekK/rNzVWoTzNoBfLS0GZ3ChwQln4eN4hdbnBWNUctLJKtw0b/JOGzNputNmhFc9x7
YUZ5XJaToyTOEs/sszJnvDBWfwanfaqutJsGGPQPRjIX3SloHg9Gc/9P08RghVOp+Z2DIg7RK4cm
uIZmuK6BtkE3HFrUj93WMyL4hl3bBjVFuV5qCDnAMOQte+oIuoQdHNn4ey8TlyBY1E69/mbebG4E
pOW9X77nYQ+ddobiulNxbWI9RP4FDqEf4+wvtmbO0B/KgKhymxwMUcX2Hm7HTcA0SU3eth8nisbj
ESyZTMZUU0i1ZeAxOmAu2LNkGE0dksKW3agKuio/CP7dW07ASLVC4dCxlGN+byl0yDvkt0qeeO/F
EvE8+NqqKNkoLGShSvp5am11ghRgklQwUD+9/TfCgY66vt5QdPYdfqfUTrMqTuqsT7TgTPjMZX6d
Ps2ozVDatXdl8eLd6QGp3WrnIIg6DI4aUUJ5yQs3x5VELAdjP0id2mi97pMx+iZtwake6PKsRCW1
tCpkk8t91Xzd7WlXRHV+MOYwWe1Egt1O36W6pzRNuISRHi3mVXPON3KPSr/UaeLn2g0GYbPIk4SR
hKa4kC2NebKdFlo1FRJTvpJcmCM9tDdrDW33LvEw048zG8OQjo4zzVXOOwmKqk6tYMVQQ/YxaKrd
XEivMw9i+wOvkOGAD50sygY3trXdW56K0pFabHhchJuchfggqWfuCxfvC1n3Mlv2nCSxs3rUGWYq
w2o+FAtkY/vex8TmJUeU+Fj5IWLQxVK1BkB+/qAVlM8jj5kaZ57wd8/oqZHPvahIU+pJ+jI8S8vv
ROmMIXIQCx8lFroDQMW3iF4sf3p6+Viaoyk9qG7F/bmoJuROGJ4j/3ckFy8tdNI3R9HiLmXv14+o
aI0/Gmf6H8FLyx1qC7Qga4e8zXmDJ7Gf8MqUFc+SXRlVW2R/oj6S69SxNowinD6ebcf658QPtM86
ExB0zLU2XunElz4cgjxXDfr89LDaIc1WmoNwDsM+aCFq2y4NIO0RwE6fv8a+BJjq7q2NzxU/Obt3
bDn1WWN1m/5G8ndnzdwzVbSvpRevy/dDVLIGJmfc7FcVwcxJJ74JlSpcNka3b9KAk3xxVMbI7nyE
q6DMHbxXqHo7x3zJta29APTzM+Jlo8fsTuNFsgTNebUEqQY9ojTcmfZplFl4+DEMkxSAFNJBNtgA
+bDeLpiHlDtR88AsSbWSb0lBgpBI8xJwIkkTzeq3s0+pu0HtuIycU9t7yden+u4iVadJ+TK6Z2vN
qvQ1MliJ3XPRVDiayGjHxjDCUM+SQ7V5YtqB+5XS0fMk9RyJFsQG2Gv/KJj/ehHJwMSgT6o3XgYb
t6r5YSqsC29L7dBE1KRZt32z0+QUrlYpJNP1/+RN5MDLB3DPi7OC/fUj77vDfZxgcd5KDrR9Wzcg
wi+Vnc7i3E9MPduUw99yz9fZIEpvqVIeEAnCyVGVMn3g0XiNOKC4eJ3atVTiNeR71+BIisM1SEO/
A22Q0JVTzmkgoTm10UTsqIxOapihDGlZv8ALCEp0mkH0JwI02Qx03C44EKain/5zBxC4LtYnoczV
KkVBsZPe81x1cNXW9eu9WcK8+M5fPFJ0tz+tf9KUdSeiWcD6BywlqbopUasAcEd0MkOR7wb9aZ+x
SyH1Y2bgZTTFe3pykOeNW8WL2dismbqynHAtqT9evxsuCA4y2By4dF0X2RSf+YTmQMJN/KrJgdBU
irnuetYa6BvvBZZD1OiIKzjBthQmM/ZJkcOW8zYu/L+Vz3TRbjWlV2Hu/kg8OmuYZZDWsE4F2GV5
UnkY3hvJdGvPiP8B3WpDMTdY7jZoAkTLqSq9GMiJ7RYsgg6T+nZXk/4BBHxwYgsU596VcG70Ewm9
QHt3VCGt0/OIdogqLLIBLyDBKZXmDf4NddqLKYjdHlEH/8hpl/X3G6h5900mTOt+/DQ0v8PzgJNN
ugLeZpDQ0hWqAhbTqqCLp6ynPk+v0agwUCiulOepb1b3I1QCTlt6EOvvaJQy49/7lbc8TKGBrLzX
eBI4BBNJCoC6WUAcgSu4kr/GvUK6oDS+vMyP03mnu6928x3wJidwMiFGzSmOVzGA0P3A87+XJSGP
6eKIOAZI2zcJol39ithkhe6+RImdjdYdvDXMLEbg4kJMIxcLO4X/uO/LRq14M1HNxxvTJjwQABgn
17+ESbEPS517w4z+0uCTO77+m9SOVSIYiOJd8WmuD4gH5zmqNU/B+w++TLIorHW1BLMvgNJPMXDt
k/cuHVGr8I2+uvmY149i2YQ+sTqKJ34pWoKZQd0Rr4rC+rOc/mQFCqeZvCLXwGgf/DKU/wSxlK0U
SuXBRPUuVNMY2Mw0QswVnq1GUpD1z1/j6ql1t3GiAb+hL61hTz5mi/Y2p4GDF8o8TbMWQHMvCSB7
TjFe7PdOzu53FmzXcvfwm3nKfHnNdEZ8x3TO26PIY31xKz1Ni1B7Bb7mjRVXuRaOqFTRVp0EVJol
A3Vqz1QcStULGkqYvk9HvPBE6nwi7l+WePoirBnw8fqxVdrpXWSCF0XQkTTnrLIKd1nvJP6Du+eO
CwHX+jbFrWG979v5tGEY7Wi+PLef+oKhATFhdZ5h7NmFbYnXtRb/XTB7+vfme4qaJOJVEKG7wKGL
UH2e0ucOEU2uDXuU+s6DdafAF4tVI+8nVqISLafP3kEnKx+7s9fRmth+NmmVCmfsvcTXBN4juvqK
+m2Cm4y/ZAuaI8tSw1vafiqQQQ7lkgNxHOb0u1tezwwqBZKdMuxr383/LeOIqdLslIt6uMXCom6G
c/ttLK1+Li6vGtbSc82DMWwDSzVGMDlwQ9UWbHkWlksBGq5a47mPQAiUF0Mbi5lEUqJT/ibKkdM3
e0YAHq+XTvN168GcvoU0e6vVVxyueZcmxFt03Zr42JPLFpBJ3WtoXz2bkjLBs7OpmxDgRD/A7s9b
gQo7OMFHJADJpRI2LQpo2CDhs9l7Ee86xVhzCZAkSIKiqdrhWqelfGV68R1UYhMFbg/A9uB0V5ta
JJtlw/R5u4fk9LNzRZ65QPJpUxVXherdH1jRptrI8RZLpG66QGznou8Co5szx1HYExrGpy8gkx31
YnvMHzFrg2UgKzJ1BAOmqiR2QL4OLXgmAIzrYYfHkEEcgl4BLT6MmbGLHT5iNK2sBr0CEPx1Fc/c
pU5lQL3wu0g+/3/GIGyLLYo4fIZCW+m26C+AJQ07EUntGmnJ7wVQCzsu8glRlu+QZtH0nZkx9wMI
iGH3KKJ8l0T3NUiznW4r1vyb+8haOauwqLZ6o/kpV2ERVrZwYcYRknHtAYtUoKv7P5hjO+tsRQsE
cRWlDkefAr0IEPz5g/riWTyrlSH9a8y4j/d2X7BjF26M24PHebZETcLoUrDeWBqCrx26vNslCic2
hFrfpeXYtrWgE/OBvH/jLmirnDDgAJUn52+f3dt5p8WNgtxDabOQiUfUv2f8ZGaWq1nxInQWfmwk
769oTSGHaE6ry//dgG1W8Y1n3rjVVAL/IpVF73++q6tgilzt4T9c565l9zxTFnUV7ERTkhE4RTnK
tvZap0cdcqZjOFW+r9tvN2NCWZXPie/GDsV2MZvKvq1N0xM4BEFC7otnnNrvzryLdNWP6SsGHOpu
Lr2Dv0Ti1P9xSFTBxcOHY3KQ0pjKUBqYqEuF
`pragma protect end_protected
