`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
BaTnm68ZB0A1b7RI6fOLcJfKQKYjp4seNvYc/BNpvXZc2L40KjW6tr9HT6+GT5ekoZisMQQeAR4B
dOaxLO7BGHpsv9LlJB0lv+JPiZKClEa6VszZ6L4u1o5obkHVxp0vYpdaL5ku+ShWy6sgMj3UPm7B
HS6TeapplDKv8W/u/bNSRgYz7L11hlx5BBS169zt32EysZu6W0/3JsEp+y7gqtMDBXgBryrrtW2g
UyIgMZjLQ4IyQesgGY2dp/N+E9rB/z65pxsmrPHkmZCiTJxrgi/Lv3346SryXQ2O5qWfRlmgurcP
2jS2Nn2SyQMh+goMBeFRuSrh6GqztQAXuqGM6w==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
24hASjzmZye06p1W5AOXZkCgkZKVZKVJgRZgVccfI456WPKIsDWf4jtnXAxZjSyOSu+HKz7Yfrpf
CjBSiNqEacds7IV1XIff1UNyCQyHpOWwS9c2NLzSzDD2+iicAe89zFwrJ61CSQhDmj53g478wixW
N11BWOiZXyW/h40evdo=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
e9w1UMVJqGnxOS7yWDR7FSSl6RHkf4OVu05ltfZb8d0sI9e5GFwjsc/ig0SmEBLFV9mqDxuX5jN6
eCeBGXNM4LgpVsxa1aNPri7i0VD+DOzo0OetoVSJtTOD6yIUltsPbpeds4KOh7so05bJ/c6lQy1q
xy7MtVovdvRJGCC6Bf0=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3504)
`pragma protect data_block
yks7hFWqzLHlYSshhYKdJlcZh2gyzobTQj2UbGBvmlTwdGz+puEBkSFvnk1iCC2/8NQtKw760zkL
P/rveCNjMWYLtQpjLBCQQ2tG9HNw+DV4L9sdX5dkdaGGkOxfOMtUS9C9MchsguXiXgbR6VBBDAEM
upBxoUAiMhtE5fwqWvrEmpJcFhK0dDKWi7YLBHRf7LYO0q8aEKSkseOQfpJdQnwoWPFlEcmz8wGz
ck1rkFUvr9/qbd6c2GKupySg23hx3cZePqdE6bSAy9Z5zBYdTLCWL2CdM9IVootHQf1+46XWyv9C
baYq9LyL4D6roj1kfAkGI7O5VgXKnGSyRtAPK7QC2uz/iCkpFDAWfDxItQ+FUZMpkMBH78fOvFEY
nvYmm0ojEyo06X7k7+VIrj3JNzlljObtn2LCzDkjHE8LXet46S2BqY5In9U+5TaIi+O9nLfMLWiA
QtjIHVi4x1OTL3fjwJnWYMb/EarKTX73YCmhfqIL2wRYa8ukp91Px+FslfFLnxSIBLD4n3JrjoiG
PcbCw5WzZcFjC22GQuIr5r1WyeSoPm694gUdNKJ91UbFyeGHiCFsdWuQXokCKzJ1WyDYCYAkifls
eIhP6QhejRS/4C7OTyyv/mvJHMCNDXqxxGLsZXwIFLgwdMVEv/rB82zCLoncoimbG54NAGxdZ8bT
/qTADAQX1cr1W4GHH26pKqeEfeie8kzmyRtzOR84lnYIroSm1j/Y3KtNwCFJ00Ep3FENeHhZfMjJ
5tnCouNgomYZpb+IH7PdzpGhlYoS+kgHisQeJgXaeocC+JhJTuJAVXrmmRYBou4slfvUlqn8YT/X
9iyBFjnC00+oS2tnIcEhHGWOGeJGI1KrNknZ5rPwUGUhM14Xwg8O2eZcaKFo+1VWnIPikacD3IMw
8Can1sFmsv9D1vS1ujoEwJJYaxFKs8YEWX/MZyk2/DlH2xPIECy/GwlBhY5jzTbfpHLt+E6QHIaj
KXgXhSuPU4xTUqvCbayBVcEEm8v22Gx5Bke1tU6LEy/TbiQ9mg+UZwuP+cYgOWV55Qw14FGfVmQD
PYJy8jW/FRlriR+pm1U1NpH/5KpifoocrtGYPwUJty3tYks7L1vWlEyDMg6Ah+1iT7zTbx4+aTkX
bMlj0mR9q3Tg0QOlblokW5AcGrx/3gaK7/03CZXAO/E9jV3zc5q4IpcVSOYzdULxt2JT2cxWjC3/
Nig+PBi2nehRVvVaWIboK/aa9g5AuljcONcCd0Tl+sU1zQhTBqO2VtX6vMDg5EMwaVIPY9RIZyUS
1fzsLFRJXpEWfxFieQJpOVy9td/S1y7noS4ScPWepiR+V2ZqXR7JZBDYNtR8Ia/urHVeXNeG4ed/
x9X/3rE9YBu8BcY+dBTlv+YBig8k6un7UCwpQOACxe7UZFbvgAsq02dSazxmEOPfTGOllVqIhQNL
XrsZ/j9BZe8CDSmaFa65OtX62U8AbCHkwa+9kU0UxTtvZGc0Fo5z3ziibOltpuA2z5vdJVnR3p+7
jHVlhcUcr1GHkWN+gE7K08/SPX7LKTSVheNi/SNcPPBV3ho57Oq8sk+q/BIq5NI1Cz5X1bbTxjvI
1OzreOxgc+6BxB/xXY4nT5PN7jsAAIwjYB4VBeggALwab5/3GYkT8eWb1Z2v4cgl1/PUxvgkn2iQ
0BVy3Z8CvotuoUzB9b7psQpprnTELswJp7FcGYKediNE/gSvs9NevPjWijII9lqW4s+jFctjqH/Z
hRKbFZD9W+fwaWTBQP5i9IiOqJCE5TZdxjXZl5H+hVff2GjIjgCOcJUBrqCmzRPVaTjXuq23Xf1s
x5CXByeCGQPvZgewTtJbVjYozCn0NYwfmKgOU1W0pkhNPARTR4DUvyGIGnoWj81gPgtRqOcvIIxL
K39MJAl09HyeDdR1LoFzNeoKCBdZwWHuLdh+p2DRlLF5SIXoobIYICh1rdPOkOGbz+Go7EDdl4xA
rRa52L7nu+PgsDBfAMD/Cg8BqPqmkcRpbcNyEk2BW2QroqyZSVEQTA3/DCDi6enxjCsUmMuVdcPF
sSV4D072lAg5q1fA+f/JS3tf15DD18x4fZXSCwwhtQU1aJpmuy501zzro5si5bCtPXuuEWPUENgd
IBPIqIruKrXkdjC+69rMQd3d8msbw8Q49LFIwmdYUh/fFBVcBGwYQkHjnxGDMgc9IT0tRCm5Nxhs
47vmRKunGyG08wa+i9EdPK9lV3XIJLo7KgCQQryDys6hEFTd4lhKcvJp4B4noIHLJXacmKZbyy0D
7qpmJOpRWYft4gCfEVxGaiuKkiOMigyZhnGOpHCyppOulTIR3XY02TVPRIQc0ZtxlRFyrOj29/ir
Z9QeEKZYd3bAAg1R4D35yq4U4UaKjWw0Y1Xpcm5j9iWF+GUT+GfAovXUWkzdh+O3Erzgj98yTHwG
D7UxkZFFQ2MLSAiGZ18hvZXT9002G5KDNtaXU7G0C2JhduaiiwW1KxMiv8UHRct0bQdAHSPMw7u6
m//I3Ul85IDJpBMAks7tVQsPEiC98DFXAPFTITJR83ncQsg239CA6iXZhkKcOIy4uIngXVBOM5M5
qD4ba1kySoKK52rfQATpcAgUXZTd+xUEy9LNGtmat/1dSCML5GdWyLbKZ4k6ZHJVkLfhiUbuJxIl
sNnq+0B9vJs8P/tr8Y9+0D5tALqqQBB+be13RN3xy+X57Sh7fv+IzcE6nILiDCcAfU44h3uJt9x1
yXOuEEG7zcYiuA9uYwHCMJW8F4KszS2wMfoYxcM+8dhSDC9zH37sx9jrCbqb8Z7PyDZu2Qwa4RJ3
SuMtYtzTq/XSSFQYAJXLbF/q7iXVzaUAsylVH40QtQnMRAJ6k9f0khA0SmZUKySmzXf2+NcUQyYX
dXaLDCFSOhawT/1ZDjBZ++txRz0C/OzWTVqh2R3/QH/0BbkFuTcyyc2P+7KLiRSdR63pa0avT5Jw
C9kkjtrpfDCZTFQtDS9nu/jj6QbfGHYls85puEPmwN30YONJfcq51A9ab/m997IOZpqccN/zAcl/
YAE0HdGSbG5WMaN5rl1DyaJES55nFocNnSAhDzIPfFR0XGFf/Q8F99piCaVd93U7K69TelSUJ6Qi
tUObShxT7300M6v9th0NJkvxkeEoecdeMLrJOM1HCxqgtwVZzGuBF898RMFwqonkELakk7Wctn/T
4cIYtAoK03e0+zqaeC2pwrn3hvQ9oNSPQDOE8eNap6VZwcGN1UbKAL9qwmNcr4TTp60gQhjj72yd
zgDuTTdC08VieizRcqkzfiEoQ0Cd0gSamRg4biRH+rJE7L+aR4ecoZhE+08xU+rPhqPLk14SkCnQ
2+Fc7a10uvSFEMBAEiVTt/mgA472B511I1iWKGa+LW7pSZVS/KCQyU0OTnxN5MXsWySUwA79t0gg
37Q+i6tWekM3BXEtNGMIjk+QFEfHUol7Qe4UlDwttUKEpLE4K9AaQsHMN29A/valtTGbkpPiZfvG
FLyy1IJ+ADtBjxqlN0ugQkFt8BNUbIzI3UdBVPI0151aC8lNthdrlsHH88TXtQ3iHnCoGlKohItr
vRmLK360+tj81eFayWkRw2A11Uabc1vKe9NmfRZyd3yJc9yOnjsICgobTNbu/vH73JG+CztM3bQF
XrJ1cMy6injLoT20mCG1xHUgNrPTehlmf9VIr1msJBbRjMgHEkE4ZNULvSBlCAIx163H6vKjbTIs
I6y6MkeRlSzdVj+ZSP3Vze00nDN6lLXdVfa+eWruhWsx1w2q66+Un2YQrHP7o2cuDGSs7wdOmT0E
exjoG96i4o19mJUkWgh5U64Qzt6+oXHgahtiKS2EL08s0YdxGZsUEEXaBoIT19j4Z2VQU8jRFjE6
1ygdNH+btrLN1jaW8FV7EkTiq1WLGkuBgq/yem/BOatLTo01wqNwG3hS55NUPEUYB9SWb0pO3Gf/
jLUDEWeCIEWp8DoX/ePSdFXwr0aa1ahCJnccvZfmnpqDEIxZHF0oL64jc/IC4gt/cLoQq3aOa82t
FiLMYoSkuaVplDxKt0I1XIAs8WB1eMf/b2c5wNYh1xlPz3GXu7e7rm1R0Pejhu843K8CzPTzq9lV
s77M4+FkDKOA6QVoZWiesoESwUryFmrW5j3eKLgdOtDNwHvpHzuu6nMMHK00E+bVdnd76xvnw/dy
K4lPWkBrJG80qpZgw3LkN57furAk7e84kAXx9kICBjd4P4DD/IRw9EElLzLbEFapRHdohcumTc81
vTgT4EqJmEc54YiRphiDe9X6uzxnCOXIQ2kC+PI516ELwu/Za+YGYwtpYJGLPw1L6aSmQE/QHH3u
W0LuO6Llgr5sfQJMMRaP296Y9o30HAGNKJp3W++Xxaw0rfbTyuW/P6TsTVtexfyTMU7qZhtQP+0m
7tp5FsLL9uJSCYYVaqS+eyeHJuBL2cUNbGb69P7BMgQ61ht0mrGL7xs8UQRFx5W6P+EZNmMPQsuW
LIpgJaPq41FpEPhzoAmyGqW7QZgZIPoy28VSxZNL5mzAuExxK0/IOD0/TZD3y0g2UIGwmAHq634r
WaaKvV/Vh3nWt87oFXnneZDOQ8MGrle35Ddf387Zy6NIUg3RYy8/8RnAta6+w3Fu+ToFYUQd4It6
FPRALcmECRdrysYHF41FyjbgYREIaj6EmiPZ
`pragma protect end_protected
