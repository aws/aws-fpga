`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
c85OCTvJ3UPanTdBRuspRDm8D1U6LAdFT7WH57+xIfWlJNrnMIqMFw0u4Gs0TJRCNGtxdvITTNuD
wdaGdhJVsQzsBrNm+phRA39xky+C4FgZE+N2aDBiEMUieHenzBWOY73A/PMQuiAER/8Cyh8C1Rzp
UJljL147eC7hbML47cyxuqS/eEljAnjU+KuEHxiFL2v9Dfdurcv4VmQ8zpWNkmR+/p+ovhxFjrSg
tb17k3Oxt80gCJ+4w0mM9ruDRXvyAoJ0U+o/vF2K5rHBgRi/+zZACP+ho7Ybyi9zMJSf6cF9Xu1m
6AZPhGFURoz+8Q4spLdnMO/rvu01WvrfbNxxow==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
JpU0LfKUCnG3jiXHssT9LwKG6s1Ss7oIuUdGAD8LSXQWxw7mQhJ1fnj3/KJ7OQWvQBW3tCWS8BN3
+MqW7NRZuUTWhSoHSlJhqXPojE2R3bz81XRCKFu8uGcN1qjMeFJex0bJ34Io1FsHfTureH6iP+Db
RJMdoUA5Joo8f0dtG5I=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
LtNL/0hL5yQHcFK5DswaMVmdlWgxFh936rTNa2Mt408HC05PGea7CUY3csnyD0PmEqJKELSHOgyj
SlxplLWByyhE8omahuukl4gLLi9sWVzFonKfBrmerbuDLwEXWW0wLX9xt3xMLX9FfZ0xGJE/3KUR
Drzp72YxtTbFVMD10oY=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3376)
`pragma protect data_block
Nez3rlOb+yt4cj763Oa8G1sub/LzH9TmdOpNACrjiYf4b63oIXQebWZxbooccbmFCphF4w1DZ+z6
TEdrhbZ8TPAYQggQ4UmC1R8pTY3r50Edffkh3c6cH0IvCDnMuNpeJNMjPCmSp4GQG3x1+MLw8ruE
OQbSgi3JOTM2GFAORCXo9xjtIDRt7D/RtHYbTpTgV7eRH795ArW6YnPLRnHijZVzpQI4BpSG0M0n
2h99oCmWz8q8d8K2TooJaUcOya8qzmZi6ouZyM1a3tSTuQUk5V2FV9yEPNE70p1jEeGRxs8r1Pyq
bUUY9IwTiiJeYDoEU/CsrkFN0+fgQeMEPccLFQQv10dVCYT/lQ54a9i3gZNRIqtTJff6u8EFYPRv
IoF3z6j+4W73AxrQIYcNqtv1+1Ad23OlLqTdOQrVUfXzM0RCaYXHzuF46GFsWxQUi6Yv0QFUynZo
hlroWISQSNQNp+JFY0CBN0fOJdTC9zZHQQMrssIIeU243238oQQiHPZJRTBZWTHJO1ZsD1mTpH4X
alcWn25MFti2i1Yb7olRksXb1aec9pYLpAHQ+C8s2F8R+qDUqcLHfNaxXDI98cvXMFGOJBlXd5e1
Cwgaz+vnDPaEkmflYJyxW3XbfvOIapwHjcsJ8mdNfYXYslPntS+X3WiZHd1ov9qsyTaYzsLoST6q
oPZHHlcOzDNBeu24Ny/K0lGqzFgtxd9BUZrPzl3Dz0Gq7Vv1R9U/dUW636FTeAOhYVAn/UA2xZCK
rT5r45yjn58IryuLgwkdORw/YH+7xomwxSomGiwEgClQmoQcYpiTG81LOEYPOdE3NBbuCGkYT2V1
wWVDjdo8TcvHeSid5j9Z2zTdbRm5+JYiCbR9YeND/kwInpv3VWhytYzU0jF474FN7YJzw6En+Qke
w3PEavFCi+vFir0LVILtlB4YwUuPQhFTDNOqUBE1FHenumQxMnFn95llbQ4PqyPl/YFD8qMKYSeh
ne75mV3b12e2qqeAdg5qVl/pUdgsT7TUuzc4CI3liMMupOICruSO3ybTbhPYUeujzSW05EctEeBB
Lgt/CkppQhwghcBrMCO7zRKXVjkvYqxPJZP9axOhoWvAZliPJLNjGZUDfPi+73xD2wyeRIeBRake
aME9q17lsc/Ui29jJLa2eXpth8xKtGq5s1Ys7yR1PpXYdYFcjZTOaJYBdv9kQZ1+uektg058hhaY
n++mF/jBRuYiYeVyInLaHqNdxljjI/jQzSZdvbjED+fMbfD2iGLF7zcGibGT8jM8RtqYejynq45A
hSCwPA4fgq9mGWeP9iOGjG0x95nRohvYhyJMVVbfxXRfiHx5BJe01ZkMCOoMm+tCljPPLALSsW6C
ttwD7gX5Qu/iz3InEhc7AjJ01K9SXadWisI3KTvAE7tPt9iwbE+aLvMQE9JU0IR6x//xdk8TMFJa
P9B1ZEyqROwx5uGLlUA2wZXEgCkpr5HkE1iNzePFx+BuonLMfn7ZoZnUb3m1f6QW92hLXD7Nu4Zd
KIdxAnoZKLfUlW41eicFioNTomZHwNhtv3axydVrrUs8sEDY/cER9ZMHXUbwDeNltGNu2wdybxRo
CLB+6kdjNCxLOWDSVG/3zjdpix5eHLCQM0mDKkI5O0cGw/I8xdCar0bpTM+yjXSWa37L+lwZSo3a
fhf4JJWilEoBLSEtBhI+CSKQlLLgI8eTPUvxi8VaMd6+SpfUHU11K0xB5ZnHvn6O77iYm12AMH/K
lxQDoad6lYjjQBcziF2k2D7NRM06vYA5jJSLwyl7J9YhVQlQTfGDInxyw1VgC6f6GFc8BZsezhnr
EzwafmQxXKk3lLjnRkv9m17Lytdsb8VYmc13i/LRNVPmh+cUkOTZKcbmNEp6Pr6VZM3S4DqpbuGY
t/3Fv1NyL4A14cWY/9zudOs5qZhKzMXwQYVVCh2zViRJR1z4RvftWn+R/ANWgT3y3w/ifV8tcrIU
aJz37nY39BuzgiBLaPV4hZZ+XC6RrsNKSu6plNk6dNuEV3fWtIkVTZIFZo/ueyHLWneUpjGOdM63
jB/4nsN5nwhdeliQ8gZQ9C1XALHxuNJIgT8kanC+9t7piyp5Dqb1FxaiRSY2fPIrofDrQc8361ZM
0zRfzbNH6HJEwk6QrmHjxyfDO9wzXM9D2A1b3waQZ9BsD6zjYJDzXwbGkaO6nSbizBI5oazstQ6m
UdMLpdXGQ37gfSuHfvToMVkLGHkJ8/eknIgyPP54ALRk5zCGrvSyFzGI2LBisvxsCaNGART2DxY1
V5orVDfWyqKPATG3mD7fvCvKUTYK7REuqrRkzlgN9YQD/yyEly1Qe+GJV/zjBTV4uEa9fDPeF7to
eXnhjlmfQHRlZS8E5DnHimFFGGD653CcaeEEcMFxYi2VdfJJ2FN9yU3YPPFRkwm0GgYfa/cPTNbv
+mFkfiLGtXvk0aqeOaEtmrCbjVEXZabrOkiOeVzAIGzDciIvQVXoXMqAvwpwZfLJ4zrjkyGZRCCv
/mv3xhoEoGr08oopkyrFGYZgOGNXhzdcCRTJHLa8X+4phzPwONYhq69iLaz6I3oWQzf961Cn/kQr
46yJbEphwLR94xvzA0nGtTny9LQtcA22HqKgEwENEw8YFLkWLShyBtSBKI8K3+vIUm2xHifYaQ3i
1ep3BTbdAmBGbKQTzD+/NGFuXvAXL1kslZAg1gQ3yDHD/+26CrioykUSyoDYXc6GQANN1I9WJ4D6
DGIjPqXG7g23m+Ezm9sfq/cmhc2gzcStYx0xmCrBKFhD+5WJx4zOYcHC9OmNnvnb7UPlIGkKFKOn
W/CdQY/di6x1X6BuHtENmyjqcdh9s+mwZhS9HXOxVgP8Lr7IsvdV/UiwFprmzVBB2kiAMiuk12Jz
fqa1sq8nSwGLIf1z+pjO2sNcHFKFK9gsSH7eIRmih+K0L3HbJ1XKl5QV7XqSI7cVi82sNdgsxlZ9
35GFWSKFaPLpkQ5dgas9RSuKY/GWnqz/A2IZtoSSnfn2rHUsk+uujzU2ttgX/x6kyR6TSr6HWgkX
LzkeWdlM8LshSenw5GzWlbH8WxOaaZ3Ky/H3VJ94gSms4ODE3lO00cu41IiNjGtZ1q6aefJFXn7Y
9Lxb7/5G0RCvT80VADVML18SOG7icJRfCBlNR8GrCtYY7jo6pg8QkcLBHac2/EP489shgDVRlwyB
qxp31avkTMOWswD/OZVnfFhwZlguML4ry6m+F7ANYpGV3e44sLGkEvFEXBRCTthLajlgfRQVhgv6
fC7NrWNXQ7x0Udangj6APyvxFGqCBJcMRDIujuf7PyiTyWHqYpXoFZnezrWxXWbj61CVocQzbAKc
+PCRt0uW0dsskOitNKv/aHqfCFpQcS83zZT6Lmfs17Sk4hbwuNvFEtCdE6wBcBZHSCZmsRt6XwPR
25BHHB21S1otJ9tc1aidSS9lKnjCuUKAQgsfRy7km3R6wtVKr5SnKKkPE/LMad0JlyFoGqm/S8QX
bAf0pE4cZBlIn88t8tK2m025142SuJxDOI3pDo753Gu4Hbcohn5bKjKvZMrj0Yxt0nhu16Q/2WM4
mNnHePceXPmVYUeZR+g5C0TL5e88i/DEJHDfPKWq21mMTF0Yx02dJqI26CcxJ7ccmbDjhW8NloL5
JAVqemMibCFX0/xVMSTnKjTWDtWxQwwGi4Is/A0JUtPrS8z8jGgWXsG7AqRlTOSfDZKYWiRMaa1O
5WsWCOLT0PjT+77D38kYw2UbDMsXVWOY0OgQ2Nd3A1OilX9VdN3R0vMkpfJp162m4biXSCbRkIjf
WM07OD9aG4rz4LSbHagJK9fzq9Ipg9iV2AASGriHtevPiGpgE8OI6Onp6Gj/SRyM+SfY7Ge91c4T
VKUvIDS31F4xb34fe2ABkOpzfIxlmWoslK91dxjHMwTiU+N4NaLRvvadA6nLpyxncWmNFYtyFXqH
Z6chb1lryjReuXsUXyul5GPeyz1HsjRqXGlnzj/9yX5ISXL3eSeTTFvjsbrYUp2GotwZPI4LCFFz
cNHcpO8AA+Yt6ht7cxtrcmJM9DlZkVC6Zb59d4lbsSQZtdwP29MmFdhZGS24/XcStwGNLC8sumda
3/vmO14WS+gRMQ2WNaGpl6c1C/4YMmncO87zoHYg7Lumd5RXE1KrTx+urDVHnw4GYmBPWx4IjLYb
DLyr4XKS5TCzw3KK1n0YMhHp/I6+8f+6mpw4mCbOIY25pg83AIcv210tysqt53WZL0af86RxvbqS
31NynTgAnQVUmxcouoodIY2x70NBeu0LS8BN8THORmlrhoVNRb1tmkBV4JuLNOgDR8TKFhGO+T7S
UiwWBkhxtyhNzSGZa9o5TFFLxs40tKUi5aNQ05L7G9WqWhwn09b+t/m+4d6lfF/z0EyoRAcCVZZU
3eveCDGULY/BtEDVJxVgOWxsnb7Yd8/1sEL1UylOJ0HakxcDq4hLAcJJMpSFc65y3WO7r4svGsA5
Gro7oZVLa2IOdNMh4A==
`pragma protect end_protected
