// =============================================================================
// Copyright 2016 Amazon.com, Inc. or its affiliates.
// All Rights Reserved Worldwide.
// Amazon Confidential information
// Restricted NDA Material
// =============================================================================

module sh_ddr #( parameter DDR_A_PRESENT = 1,
                 parameter DDR_B_PRESENT = 1,
                 parameter DDR_D_PRESENT = 1,
                 parameter DDR_A_IO = 1,           //When not Present to include IO buffers
                 parameter DDR_D_IO = 1)           //When not Present to include IO buffers
   (

   //---------------------------
   // Main clock/reset
   //---------------------------
   input clk,
   input rst_n,

   input stat_clk,                           //Stats interface clock
   input stat_rst_n,

   //--------------------------
   // DDR Physical Interface
   //--------------------------

// ------------------- DDR4 x72 RDIMM 2100 Interface A ----------------------------------
    input                CLK_300M_DIMM0_DP,
    input                CLK_300M_DIMM0_DN,
    output logic         M_A_ACT_N,
    output logic[16:0]   M_A_MA,
    output logic[1:0]    M_A_BA,
    output logic[1:0]    M_A_BG,
    output logic[0:0]    M_A_CKE,
    output logic[0:0]    M_A_ODT,
    output logic[0:0]    M_A_CS_N,
    output logic[0:0]    M_A_CLK_DN,
    output logic[0:0]    M_A_CLK_DP,
    output logic         M_A_PAR,
    inout  [63:0]        M_A_DQ,
    inout  [7:0]         M_A_ECC,
    inout  [17:0]        M_A_DQS_DP,
    inout  [17:0]        M_A_DQS_DN,
    output logic cl_RST_DIMM_A_N,

// ------------------- DDR4 x72 RDIMM 2100 Interface B ----------------------------------
    input                CLK_300M_DIMM1_DP,
    input                CLK_300M_DIMM1_DN,
    output logic         M_B_ACT_N,
    output logic[16:0]   M_B_MA,
    output logic[1:0]    M_B_BA,
    output logic[1:0]    M_B_BG,
    output logic[0:0]    M_B_CKE,
    output logic[0:0]    M_B_ODT,
    output logic[0:0]    M_B_CS_N,
    output logic[0:0]    M_B_CLK_DN,
    output logic[0:0]    M_B_CLK_DP,
    output logic         M_B_PAR,
    inout  [63:0]        M_B_DQ,
    inout  [7:0]         M_B_ECC,
    inout  [17:0]        M_B_DQS_DP,
    inout  [17:0]        M_B_DQS_DN,
    output logic cl_RST_DIMM_B_N,

// ------------------- DDR4 x72 RDIMM 2100 Interface D ----------------------------------
    input                CLK_300M_DIMM3_DP,
    input                CLK_300M_DIMM3_DN,
    output logic         M_D_ACT_N,
    output logic[16:0]   M_D_MA,
    output logic[1:0]    M_D_BA,
    output logic[1:0]    M_D_BG,
    output logic[0:0]    M_D_CKE,
    output logic[0:0]    M_D_ODT,
    output logic[0:0]    M_D_CS_N,
    output logic[0:0]    M_D_CLK_DN,
    output logic[0:0]    M_D_CLK_DP,
    output logic         M_D_PAR,
    inout  [63:0]        M_D_DQ,
    inout  [7:0]         M_D_ECC,
    inout  [17:0]        M_D_DQS_DP,
    inout  [17:0]        M_D_DQS_DN,
    output logic cl_RST_DIMM_D_N,


   //------------------------------------------------------
   // DDR-4 Interface from CL (AXI-4)
   //------------------------------------------------------
   input[15:0] cl_sh_ddr_awid[2:0],
   input[63:0] cl_sh_ddr_awaddr[2:0],
   input[7:0] cl_sh_ddr_awlen[2:0],
   input[2:0] cl_sh_ddr_awsize[2:0],
   //input[10:0] cl_sh_ddr_awuser[2:0],
   input cl_sh_ddr_awvalid[2:0],
   output logic[2:0] sh_cl_ddr_awready,

   input[15:0] cl_sh_ddr_wid[2:0],
   input[511:0] cl_sh_ddr_wdata[2:0],
   input[63:0] cl_sh_ddr_wstrb[2:0],
   input[2:0] cl_sh_ddr_wlast,
   input[2:0] cl_sh_ddr_wvalid,
   output logic[2:0] sh_cl_ddr_wready,

   output logic[15:0] sh_cl_ddr_bid[2:0],
   output logic[1:0] sh_cl_ddr_bresp[2:0],
   output logic[2:0] sh_cl_ddr_bvalid,
   input[2:0] cl_sh_ddr_bready,

   input[15:0] cl_sh_ddr_arid[2:0],
   input[63:0] cl_sh_ddr_araddr[2:0],
   input[7:0] cl_sh_ddr_arlen[2:0],
   input[2:0] cl_sh_ddr_arsize[2:0],
   //input[10:0] cl_sh_ddr_aruser[2:0],
   input[2:0] cl_sh_ddr_arvalid,
   output logic[2:0] sh_cl_ddr_arready,

   output logic[15:0] sh_cl_ddr_rid[2:0],
   output logic[511:0] sh_cl_ddr_rdata[2:0],
   output logic[1:0] sh_cl_ddr_rresp[2:0],
   output logic[2:0] sh_cl_ddr_rlast,
   output logic[2:0] sh_cl_ddr_rvalid,
   input[2:0] cl_sh_ddr_rready,

   output logic[2:0] sh_cl_ddr_is_ready,

   input[7:0] sh_ddr_stat_addr0,
   input sh_ddr_stat_wr0,
   input sh_ddr_stat_rd0,
   input[31:0] sh_ddr_stat_wdata0,

   output logic ddr_sh_stat_ack0,
   output logic[31:0] ddr_sh_stat_rdata0,
   output logic[7:0] ddr_sh_stat_int0,

   input[7:0] sh_ddr_stat_addr1,
   input sh_ddr_stat_wr1,
   input sh_ddr_stat_rd1,
   input[31:0] sh_ddr_stat_wdata1,

   output logic ddr_sh_stat_ack1,
   output logic[31:0] ddr_sh_stat_rdata1,
   output logic[7:0] ddr_sh_stat_int1,

   input[7:0] sh_ddr_stat_addr2,
   input sh_ddr_stat_wr2,
   input sh_ddr_stat_rd2,
   input[31:0] sh_ddr_stat_wdata2,

   output logic ddr_sh_stat_ack2,
   output logic[31:0] ddr_sh_stat_rdata2,
   output logic[7:0] ddr_sh_stat_int2



   );


`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2016_05", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
pgt5peCBHI5V5Eh416/Hj5oNL1WXvbW4Zm5IOVUAxYXSGx8rDHRq24M7XfupEMGkfgHpl7jEj7U+
fMp8gGTA+/Xzh55fObQ9/NdBeeWH3jremz2jJdvAIk0BfwYZnsvES15i2EtP5QtIDTUKqUjxeG/s
Tgaj+HscsTCV+aGP8by0a7nNQqYD91Bt9sJh4Jh8zitI+G2kjWiJRtYv8Y7QhShTjmlTYro7W2l8
2Fnsa1SnQDLV4VJzW3B1M3aJBreGi3p9nguGmTUXsZ6ug77m7bmEkPzZwdIhP0KJYhUubkGCJLl4
UncKlWC43+SWB+JsABD1bzeCfiktilYA2RbVvQ==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
uDQMgkAdk/qAyf5Luj1QYDm2wNnQvEiqA0hgfCWRq3vThKZEL7p1Tmx1c0qvOAsZYuoZQU/ZMH+u
NWzc7oCw/G2YLp91LcJxoRKWlODgRNGqqFY77RR+BKjBEmWRO0YzUowPSZ3luXT6Aqeyafxfx2XT
0k69/Vjc4jI1AkVyH0E=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
SsLQaEXu4ljnypIg+lHgIhIqZ1XHedE2DV4dZpxdpjVkcbWTzMaIstnXg2xactKfvi4wqGfM1rVq
Uv20x+v8NwpuohYKgGdAJpXFC3MQfHTwclRfUAgy/yMtI8VtEBT75+HT5iJsCYY67swchDmdB6Up
dYH9lXYDdCEYdqDGips=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 63632)
`pragma protect data_block
SG/X1784aq7c8v0ClRHJieFI+/K9om8jRUEKGRfVpMGWP/Hjj4cIChrlGAJUWguZMJTDktU3iOpA
MnEnJZBdoqPfTr821g/P49dxFMHDlVTMI5suW/CSZnb6JoOqR1RlKan2mtFLvxsLwkpqB5ErhQm9
ALD67ztXErlwtaM/qq1kRsdv+X+mdlbxLsms6ipbHhgL3zNhh77ma0v2LZeLOwCbOS9fJxHCjhs5
iGiaPYiwRJdw0e64kM9ASm/6YD1HgffPNnH+DCS9BCJzj655YuXj25M8cXps4sTxC92zxFs+NmB8
AqZp5Ak5GUd+bGTKcPqxna+XCOOD90QY+IpQEA9SLKwSW0erc+0sMaHqh8R1U010DAn9PI+7JmP8
eoijfoipyPSkcNNEiOPT9mp6u7pw4VegptRRLo8GRXKEqWpyvs4LnlmjIEyhzyUogLmGkxjXU9Yw
c3xi64Zo8rtXmAlz/W5CAVp8p20ndkrcZnokuaTfZAtEFKvfCZpvktJXj8LS7kqG6bCyDxmP210B
InhJ66RLAYgcAd0HHeoqBSIpudPYs9x3+1Zajgp4qfdeyn8tAR10PY5fXme6E7sJyUH2T5S8lzjh
IeURuz6YY0xEfRlWzyqqKiEwuWJOpG4roizrTLDeJOZmx//U0H4hYklJtYB1owzzsPvQTgRV9o8t
RJ35mSoxFV/1QOBdXocRfXpYVPZWSRF5qSYae9A/T1yYKEZ4mTn/i4IB5RMsy1VVIRiEKhn0uiI3
b3jrpKXlHn3DEizzA0590JsNFqGfVXcXdztDt9mqGTPISUwN83XIqg4/MD1/EeoYW9AUDcgEGS2u
irQtAvQpOz9qAe6rFmaR+v/SQEmNu99j1M0O0UzCn/KAwyZEwJygiC/rKQySwOUtVp+l0NisQfO+
z2ZwQGiWM1rJPtLXKrP4A6IH8bSSbsLFQdg2BWB4cbQzmpYY4ss9sQH5secm6L+VzVXQ50Xtbu7s
D6uuQj56td6OK4NNiBrKn/nkkOF+lnAxRtyr1vUkErD6wtADRkUcG36LN8yHeaMSFFyBoS+5BcYl
o5sNVxMq1sCHjk1Ib8edIpWaQmnYNBX/rZngXo89JsbINnTZc68zyJB3xAKwwV5PF9l+0HEaXWhS
alWnFLWPD5wvVZEerJJvnQPu1vp+gMvNu7wQJ8d/3SAihxFwpNFtlXtxx7AWnFYa7XxvK4HTO+ke
9ijzVnsGW2MHjiVyItHzcZuEzz/PN3qRWwc+Qt69CoVode780O5pLi29gIFT61MCqdhUmIe1VnUI
+fajmL5oobuvoKu3Q7u2hRL7sg/ilN2KR2AMzvrfBws4iPgmOEpsrw7+rhky8Iq2C1Po4zTfD8Y3
rsxBUaI0YopnVZPnqz2Y1jJDHtR6fTYTsVmKstvWyLESL6W6H/lpaWrmbfo9nqvdpsbdcpMNb8RF
+kvdqb9mwG1y4gWgQ7f+2paEJHaKIh9IhjqLDjJxu/MFGxzDUXypdt87uKMionrwK3hk0xehFd/C
iaE9ovNfmVoKO7psplDLk7DME4hu9KQlhHq1zfb8AvqVSMFszuNJKrdY3JM806XdnK31dt3idDav
AUYnmkGYVoVHdGe6ZuSCPZP2FIcDIrO5jCBdhFwIJXO7OjZbFxqN6fDtwOazlvbl9XzH3kiS7wmr
R2g6FDVRUmy2qNDhqiuIWQk8y7zZZTC5huf+kUQ0+baKNv3azaq4UNojy0NFz7z4hso3R28n3rFI
BXJzmMc/LVc0ShBoLd1yh6ZrZlYjgcKN4zu90nmBuSqGkeCiVJBkbmfOTW28hYPf6qOGQFIkVsb0
IDHVJ18bCxr+2oD3QSZ1sfZSrJHAfmGbSuF4EdXCFo4MlQwixlMVZ2RwFJ2zK+R5RIyVU1Keoiu5
lucuPChiSGLShlEZHhovUp1uq8CmzuhV9diF2Eg2oShZohLPAoh2Nmlbz+Mb1vJseG0DtM+ammVp
nE1/XM1p+OMF2FYIuArJC+aIX9EyAAYYxYeQWuzBJtIdtyjiugy7g0pvYZI01dRv0Z1UvArgyRYo
7CskdXNJCH0Na4aQniQDyG7TfhsQW4UMQD+3RUbsdC0DGQTJ0yJRvjYp7CfvzwHIQqme+MinIcnM
kI8br2NaPVBHdRChnwcTwDFQSBTv8VLAAt9wWM47N5sAzxP+H5BPzT1nxQ9Xbz8a5yUo2MynzVbY
z3Qz+XsmubCsk7k9fJz+30sz40tR1C4osY9b1MSmsA8M8Sa/aADZHoJbRzo8lmUmRGzP0LGARQIt
5HOeeohZL8vCD2m8CyDBSkJ4Z6aLV21fesuiWg+VDWsVlOawIWrV2O7acB7W/rgdLNP1LiLzH0+c
E9HRxLKQjkgmuePsLaeSOpNrmjDsQQA2DRDpPTnp/PUR98pyCh/RNmKs1NMp3ThjNccWGLPUIWhM
nYAxhbweiIrkYcQBQLFAYmYLU952IqpckzcPkQuWEGfN5cTNj6SCySSpBUydRKO/jEnlI/DXJmgf
GKOVlI0/jVFd2Y2jlAzgbBNL3cBwU86ne0U7S37BbzDtEAyUFn0xRJBEKgHs1UtcfvJsi5kagmLS
mJpuObbNCluk8nbe3ce0sRUq9qcIGy+VCPjpLh7E13uCBo8gcvqn1vGZWCf51WY9hW6RDJD+oThA
ArNA64KLhDG0qDXrkLP2GA6NAphUKslM91c8oDVZ8/p4mZ68oyWvsrxWUDG8lsQ/lJmJjasJrl3L
CtayWl3o8i5CQAbmaZjjzoIAbQhWOAWbx8SBamBR/oPC173hcKUp9ju1B5xwGNLh0cNVx23Ycl+M
1i1Bi09ru3DI0te2K1Z59B9TZXk9pLWzo5SsYsx5i4GUVjupd7r0HNwUX4W/HI6JfB6bfI2sllM9
FI5x4t1GIdElHNgZnsjc/7QQXREnDACv79nmL91PrAltkWXq+bs1cW+yvW+UCAUaSkbZnAA2HXKE
0crmnHHSiRV421QyNQPjUpq1Yqksi/SQQDyxpzm2gS9oM5l5gB3qWQTCOwQ7eDKdE/B38F7k2hjU
UdSnDnnDeQ9Lo4U9TSPtVeZPHbQCrdXo8fV9XGwz1cTI8LERLOHHHRevVbEeOWgfLlfSZnwRXsUJ
2fJb5kjI+1ixw9eVe0vnsOG5XQYmW68XcG10ipqhXCCNYTeytwPtoqFMfKBQk/u/5jcOskwZhlBm
e6hodJztHJxYcgSRGYekxaCITut0m2ewQHKCtJ5vWVj3Pv+HV7XzofeH2lvd+lKYVMf5McZ+2CkS
pQf7Q9TNIAbYFvKJDJ1bTZQciAsvPf/1UX3ooHuBt9M7mK8lIEF3dRG3NzwpbHaQDBSLP/WvoXlI
lOV205Bt1TSvZxTuCkX8kB/Wf3HOqDtmqg+wpRnRxUmaXXQ3VLfhVGtk47MraZg9xBOyWkzHk+CA
ixIuwPDV9XckH9KkkyrtRLkbtUoCIwp2dYj++uHA1/iSnWG0McHiXz9okx3cLr9K1beicqSPxn6o
1q6koNYkwNdjcFfRBin2wQ9rWnRJyEjulAQBQFCM84p0hez7SJNnQTu5bDRAly6BBMddj4RxoptU
kZq/k91EskaztzvqEWG82TEmJZheiKIjuUYwTiojBridzeaoriTbukqJlmML77WXYhDP5frCAkHr
JVJFRXqSVxfyECKBLxezv2YCY+83tmJva8DuT62aCUoWxCU1bk0rYKuPpDZFUoeAfyMe0j4836E0
JcVelPvjE5MIxW8SJrwpEoLxPnEoNoFubgWecyiiXNrOYomVwgmaO2GdMO9UJ7juTqItTZJmsPTW
DQoOoirMxG9MpNnt5Sj4wZ0YYaNJnjLuYL3xmc+RhRHM8hjdY+JGM3se7h9PE+XU50pzwQ1wTLkD
VrS2tFRiYKvs0vJuz04uhW6mczSJTqK9H5QnqPMtENBApAk3U/+HqZVgZ6D3RsD+WS/so4VqGBTy
n3J9UAQzyaLrH2xSMEgGWGUPUK01se0XKpdOlOzez2MGy6WFXNqPzo+yFIhwRKSPWTEoduEmSdwQ
Uezc4+w9q4lGXmdNHZREOosxtNC7j50fS5/mNi7yrdVLPjyv8VC8EPoJYTGb1OjG0/F+WuAyg7dp
GuNQTLDALbM+Y7PbqX0ba2BmWJLnValfoeaL+QoW4cvly5ZEMA4tOyAG9SqTx/NSWCrwn4UJAOSS
4x/CrxY3P/mBx0n4Cb59X0teqNoWtN1Y6JjnMRfKTTf2VxVBrRAm6D+Shq9zq3z+QzI2/JSSIRGz
ROp65CI6RiQO4DOwCSbB1YKRlxvUgthBXgqlHD3lnJXC6dxUglon7WmsHPwSTPu1srdtMhlHOmrF
rS5/8TZpjftuJ96HPH/BSOe+RlmICV0pYijnxK2CyhtYPCIU6ET1t+S/W/EloXfHRNZj7VVVasmF
BwyVNs26LmcUvdI8w2UlmJklovPhaXUj1JfoUZv1bpuv31/eTiZ963yzYXaVUeiiHCY8zgC9rrAA
nKFQ29yeUQnwR6V03Yk6ghhXiK2JPNdq6Dm8qX54gikRidJBSJRcBhMVcv9ZDIXRaieApRfqzmWQ
DUPU2wrIgXnQCLr8T195QkqEiCECI6YShifrb1Ei9EjVtfrrktwMPe8UhsSD8XSD0evihJ1AIHW9
KqCmCouWqVbswwZxKiEyChhuaN2qAmmeK58kZ8zhMkAc2MQALoEZpJEipzq+vqkGDl+mYxPOe7PF
qkf6Ttexw/p9FVk0vsF6bHC0rY3AkehBxhHmgm2spZ+5KTz9sEyGDoO6DHNYlipBHZT+tWzDjfib
YZMEz4zf58DeyUuoOD4Ug3xmUhDS3zNGptVAx7MDVFsHRxLtKGbUtMBcMOejc4P1ywmeS29oXsK0
n/DkJM1UATRBGL/OaLf78zjBUM9H7STwcarQawKCr898QpnY09tKYP3Z+yMu93WBdCEiHyKYe45G
+C3Q2GLGLFVEJfu88hFVzcUPyQHuO40CNPqj9WE7EiV53btKYIwa7xujFTtWbEomJeRWIoMp3SC6
p7dXf97XazFY+Bd5Q8yB5hJD2EgH0bjfHnen6Ky2/GpET0jcwYyEKUczGxVzgB1NAkFI/DtHss31
KL7mo88KXlMpiA0EDiUGmcKeWm6aIfghiTyzxNLJAo+pTt3Ky4meN3k8fm4ndQMKWqnQN1SFx0sJ
gAimFd2nU/ErzJKFf/ETuQUkhCZx5/qjzjg4c2ieGYsr/9+IJg6XmYxPQJgkPl3P3O6c+J0b7ark
ibjLiH9cZ3jUW0vKuQif/33bznZ4sMDITgmlPEqU+xTSy7+Yg6+e/XzntKJ2kCpdpGextqH3bdLD
AvNie6CWJM/B28VpQiXtRR4NKjAFV4OdeX42SHcZE1NgSsfjzQ8vtxL+5td2jjUnCV2wsV2GjQV/
adjPsOMAtwlfGHjauakqPN6kaGIh5jZRYLelZNRVjNANM8OWrkwI5jMlFACnDLYeOxF5ZV50WdO1
xWTdabpXJ/z02RQj01lxA7xnyDJFDPwsiUN8Fny5Dxfl4UrKQnGiuJcaLeITnX+PEiwN3Y4Q538o
KhDbZns+04b4aLXRNILBU5H9QiIh4cKPUg1pfHJJUiH7OEe2JOcwqVAqP6c1Ztm2rNCl4dKlCR3y
W6NgapF4zX1o45pKYs560P+zLdtZUHNDMq9SBfnBIpL4IPp2UP90FXMKseSJw30gLvGi2UNic/62
y9qIzOpNoPvrKXEfjHCE2xLvU4N4Ve3MplvMhNd3MbHZduVSvZgXu/5QaD7z2E8JtkqbbmS4g1tA
UNGo8KuljqIljhqjX+NkXeLmwMe8UDF6yXTAMEFzO5eP06saFVE5dy2GXo0BjR0Hq4NzTEzynzz+
EjS6/fWOml6vTGcdeGkJC+w5Hko6DbbOPWzzqXEqtJfbRgQNHE2SQWTCk2dm+jY2k53Db0Tm3ait
5j/SPtsAaPiaMprADN8OuNmbIXS8Fqs7MgAjgZgR5FLqMmhIyKheAAEtPmeOzfr6/kLn8TFG4pai
2LSxboz+RvzYlwcJ5ATTb1EFVgC+PBhWGgcGQSu1Y44hrxATj5DYF/g8r3t653Jqp2oNu0O+BBkd
3BsFi60v1oWbbornIEYErkfXytdFW95rREyh14VGfJzJGaFhK60jOxsrPVC6Gh0uY8htWmN2b5Q1
KceJ8K0GONnQUT/1CIUN0YKYAsM6pYJCByW0LJmvGLYDHqaYY7TTaS35nuiXdwb3iPpndOZdAKEF
9nO/in5AvVsLUB3fKyEQ+AaReXEujAIxHD4bCuvLEXWjhjCwHheACClLPRYIli+7Sgw1mGa7RIFZ
0Uy3n8qylOKDmgF1Ru+8YNS7+vmVSpEIjKCmv6uikCDeNsXw+Ii2prQn3/I6LBizRR2RQ5OYZAXt
8HWb01xnszHX5MC7R2pwUC+72wMwmKuc9pYXXMhmTbsBGhBdRcwnyyeHj/HW3/0FQmm29eWoao9G
W/Ge+cq/wdjWd/SXpAuFcbQtvbZi5P6zy3Yy/aijA00hQfNm3ubm2XCxklW72mmChztG9rITLa0x
8Xnuohds7XrV9C7eCzwGpmng7P1G4gH7mBzeXC+LAor8N9Rb04GNqN06HJHZlZyxzjhEVDt3w5lF
4zFFxg+57C2/lFpCyplj2lRnrYGmyg8PT1UyF5L/lcfHVcO/Z0MJg9Mw2T+jbWrsYGo3XBIVFQHG
rNrPsyY3r2hhWHMHChkAPt+0P4o5XzmjJl9aLrXSXGvw4mNg0UE/amZNkgPGC/cUiy4JFlwJPfeL
vpLOKJDya1d0VSQ1L2WvPNa/c3jQwjzsRU3d3oPQm5Q3Sk2ii3RDIu6wkkXnZQd4YRbhZULMr++d
hZjODkVSZM3QfrsRrebDzjZa2JtDwUkQ1E2ypNHOSPfK0wb/Zvngcl4sSFaNq9KgxkhYKRYHmqRp
wJ3Wz7+VgVxO6UKKDNDMGXWX/UCwmAyNAtfdPCpRkIu5G2wbORqSwj4Se6PZbo+RUoV2B3uWy6Dr
KLo6MdPOBXJ7xPEdRk0wWd1waZ9zdDhttM0Yb3Zde0fA6fvUMO89sdkzDr8+fiyF5dvz7Mbpuyjm
n6gl5zyS9npvomAJF0rgCvteO0CEiwJTzA9+Mgo7xr9xNgU0grl+zboGwUqI7gaj1JyYxA2RAL6Y
Sl9oTM2pRPfgT4zVrB4pnAuzxC7GMvXJ4lgGe5hxoxkLWA1zk1wE0dlxFDcJ5efRz4p8Q0IOL63X
deq9JdxsNbRK60CvQuC3kOWz2oe81D/o0dctK5URudlMFKCJHX8uxw2tEtMoxmOP9uNwSP6bDTRC
N5f146ngQmjqxr8P7c8AWnRxPM+gmxXNl5wA1xC+6H3cCM39W9NIiXGG3f9GAQqm5MNJrcZpp28V
FK98vyf7s3BPQ06CeJOLZGySVUx/6ZuOe67m8vbgv982lOoooIPGcpLNTXGZS24CmrtfCcvIhyBY
w6v5R0jh76NcIS6m80zkvKlM8Woi5/JGa/VEECaheAwXOnEe4RYcbS+y/nTiKaNDpSSJseL8/Gug
reTFRpp8ajf+Y5TbSC/ltmIwChdNCut5/Jxe44XbYJgM84ZVI4N9e9lMht+VqvIayEhpa1Su8JSf
KB4m7T12R0zGEt/0mG5R/Jyaxclje+ltyZjWi/QsWjNNiQ1RHdipn0smqlH0bwvKiNSlJ5A4/bei
jWgLh7k9BPL8q456+/eZJYp+4B9NeftEDtOaGRINaC7mu1aabc5i02pYXfbXwiknzfEanrdoWZ+G
e5AGnjVemXn9beN2xbPGdaOKSsmGp97uPg4bmc2+eoPy9slq3HudXE/wUEc41H8cZhNJ48oVppx3
EVcPX85Gxm4Z2KOb8gB8zC5p3gG93DzLbXOqXkgCjWBd8W289A9IiwQGjYy8B0E8FlCPpaF/pGfB
U4XFuhP+Ayj5IC5PzY+np5K+SGC8LqWV0Skq6oCSgKeKZAVxOW0d5Lr6/lCuW3ssFdBZ3CVJ0cxJ
hKT80TbRnlI/CclLcZFPtMau1xep6CAsuVX/v7e9ulPSOOBBFnsQRGETNQs9UobI2x2OLDMIZQEv
MPQ0wVJjiTJV7ODH3fbaTS7zLfSNByUI1R3fJg5poPyfhqKvjYPVqbHcMKJroqTXLtYPeO0f/Mkp
AEKCuW5ce9ToHFbp1pBKnl2D9OTJYO+LEfsIIYDCrXTpUcqep7bESEd4hWG5SFa8bYmqKvh9t3LH
93+fsH5nvLgM7stuhsns9/AsZrUYMFVU+tog9hg1t9oXzlrMXMk67tTRl4z1B86AWIBZw5qFhJIf
+q1zD5LaFUElDzHM8ILBP6GgIvFjLSS+w+IJGdAcsd+cqV6Ks2QUjPp2hqzvwkvDX+eeVBXo3NAT
tLxhQfUTRRYdRE7oV79W0qP9M+yT+NNKQFfKshWk6OOC6JB+j7zfjMqjEi2kCzGYBe5TxOiofqLs
ompbX0biAx2MdwWYU01NSTkT7+l82i55MuYsfn8tR/Rd2JRky3FfnHClI45CxE6PLBeqV+XbYPG0
KuyuCjKU/if4TU5MLFXI3vZoNdWI33UII6cU8s9YyaurskOFOKIJow1npBt2+FmMAWcyuOXj04Ir
uf8tralHuXa5GoE1NDgzdzFkGNqebQy6uAt5g9eel+VufB7unfymICwj7PBhHEnsg+eMIbP0eu2d
zMzb58IB+YcvGT8j32TjxG+gkQYy16pYSr26DaUoWs0NJ6HlyQWvHucex9uFS+z6vms1RWb9jQM5
T0u3KfSHy1IbyboevR0NAt+S/KT6VyrZpX5XpmglRjnaVLq96LP0yrV+53smObU2It27xYXz52yr
ikg6xMCrsSicYvewh+eTJ820RjTldH9tA5iZQt62Rs/KWK9+pJqC80JZxq9bDaNsIT5s+MJFI66S
h0NGdKwLnjN7RmYSEhff6454yhydpHPzShxx3yqAnt/t/H0yrfR66G92x2JxFlltUQNoWofUcyAN
acYNzoc9IhfY+cyoVZ3UozcGOrEVGsdUz75yDlToZZlIrcYyLhRiNq9a39/Uq1qnmS0dXVNHAXHi
yWon5CBMXJHgKvzFlYFxtrol74k9XSxWnbx7qtxWCxmhPe/EOv5oLAv9EC36Z3UfxnXMiLvn4suV
TLjC/CKn3Ug0eM3q69RqiFzIJ/l3xUjhnHN+wq9eRdZDJxD8ZjNmCPCRoIisXDkWZaYMs8ViYVJO
ektJQCobfxwQFbHMZ0rn9LotGBe4v9upUAfo3EBQkRnWz6HrJxA7PmNrTrxa1v8TtZqGW7K0uNW+
7lT5IB2ArN5GS2+Nbkt8XE5PPFxThsP4gDYMy8hkAjtixrttYWWt9sl8ly3ts+TJPBfmYSf4Iz8K
cs3+48tItl7LFDUjHAwUdhEmIW51aXWu/5+SVBy6Sg8zEkIqYp1XiJv2siHNI8AB5p/Uh5gjhR4Y
uXBxHeNEeJKyioHDof+dSE60Bfg7SIQ4iUUINRdiYFJ0XfxqL+w9VBRZeuhGRsTvHSmSM0Ov7rKs
BwNUd7PHTqCAlcey4JZquMny8jNU3KGxajxeNPdP4JY9P9Olx2GWMMtWNFnnO/TfQYQw/ENV8lCu
h2f6+0kbHf8PKEzWHFRC6p/FLRTA17FvRJ5yRw/FCB3mBUKan6e8VttOxzSof95+Uj3OhJB2P6OU
uKtOlab/7IXMSQ9rWSLrDg6pR0vg3kv0yBzz8HQ6X2HWwShZFai6tAeXnPKtDxIZiXaYFt+oJkKI
2dKlMK30yX+5obc3rq75/BvMbLYgDO01hzs5QD2E08gYf/K9VYRRt/vXzjGzlj7kGmBqdGMo+Muw
M4SVDdKbVBlWbThnO0hJFSVauUe3xG/uTKcvdBIDkQEpw/cu+CVDnshMHYKsNz5NKD1od8lk+LL9
L2gF+xEv9hltX57YaFsZJTQMwuTTjeNStxQP0jd18vezfCfZBg6jbUVUEKJMVYnEPUaEV0CEWN77
kVZkEa+bas4I3yvSiatkIGOUczbz7EhpUGWyuH7ZYsVzJ89Iuf9YFjXJGwv1b7T2foczWmY79XR2
UD1A25cZkRxNaWSeiu6g1rBlbnATEHI58WuRads8iHQ7WH2E16lwIA6rC2DJ/dedO+76bkuRR9VZ
OjSbPhOuEbn6V+PhAFF0NFDJtInJEntPre5kTW1PPiE+bVgMt44ehTIABMVTyEtvUf8xC0t2M0aH
HqYZW1ZkBEw5qOohSmnd2ZiPZn2B5YfJB0lGh0/+ndlohnbeSCTH/8CyqxG264spbvL24tKidkVn
2qd3XhwX+FIC2zFmMUuMqtrP5SifZuQqF21xQ1+Df/zQmzS61zw1gnALqtlnnwiUmJsOb7fLTf3a
Kkk4ypUcYc6fbgpDgtP3Ba0Hc5FyDHI86tZwHB90WBvzY3GTGI+PcLLJhQp81OOkPTYYmXA7svy+
xuX/vo4X5+n2jTVqCSccNBQbAiyV5RgcKzmG3qSCRLu2jAGHzldLn1bndy17Nh/e8/AAF5A5MFuI
+vuFw0Fd4uDtGEXuJ2CJ+8kwxAZfumLkx9eTVgLMIyu7DTD+ByL9LxGYxVaPGmDMnoGZhybLwTuG
wfNAnirRVV+2ydUhMnfIgttu7IO5zFukcJCJ/iqvIZmLs+i43K8ujIj6/oCPCMSKabb/pW547qVo
ZhMOL05bJd6goAR+dxlahFLuYDWPLcCotR7+c++ew3rILC1ohWZfOw3Q00nVvE0ZZKykC8lpb2RB
r9hIzqSnkv1XYziREM2AwEOFPyf3SbLynXwB0zE/ZLncw72Hnc7SXaN3oiKw4R160tDEkD4xANHv
0DAPs/hBhenH+6xTj5bfuPGM/DFF/OknoFUniqrgNGvxoqpnjvDFIckw746ELjVVJR/8kOD/Aj4R
AcxLpYwtaM8iL9HcP96jC0AFH7DLtmfnZMBLjbVZArOI25SP4WsHs/aLd/+FCzTGvkju2gV/OBFD
ajfm1JO7hb+S679S6q0eb0QP49LKiBcHrYGwi5IFpjOZXvgFs4qhwbAp7/0pqi8ZS4Dbj40NQdk/
E1n+xeDdygS0P01WuQOTw84Q8GhvODYfzmx8ep+78walJS/4sZGK8XQFejIG6FlTQyQoWcQTOo4u
DMG1qhqyzVwndBrOOgPw2aDN6JslGh+DpzLgAuMqlya+IuCRjVNjs/yzkMhAdFUqmQNRBTOX/gdU
0RVny6EIlkJ5uqoqHRk9ddl2Nf7Au2/cL739hN5MOpPyteTBv8gsGfgJCgzkMzAMr1umOctArjoO
dzEZTIsmeQUHNVTzHPp80COHgaPwTOB0JsWT354AmuAkedehBVJm+EwUNtCuxhWevMOU0v80Z5hi
2jImG/aRSklDZE+9zju3CjUvOAcRpFYuFxss/Uq9wgstai2bkspW07zAY8nPP4rm2tQ0Wc9UvTh7
XuzjwPkJhzs6RAdSiA04SLf79ymY8BjIgZYCKYSV6sBtHipnQY0lhUDsZdRQwscAjfrtXEsnJ884
OxYU2TEsrE5UOS5039XOW10vepg62GsZcEND4xPbzQrjpoApqOUZK6zfgJd4xsm6T+hmSia1Q2ZU
KEkjEoHIRwz0q1bamv5l2QTOQGc8aictZEqhqz8c+YuE2fBthcJVgKjEK05MKUQnJeQ/MW3q7Ybx
QE0UAH+TEsJQpqzL7QMb86CpY4xYCuWzR0/H1x/cGpSQ2v0nD1356+LAa0Ib/exra3X9WrYxFl+N
B8tmRYVb4p27RMwyi8PpxWPhNwZmgGbGTi5jRTfEopPQje+rywfXG9Gdc3xohQApebE2ilw1wCTp
wCSqM9YhCdvmkcnEFcESzrSHViKun5MDwKvJ1Jll9upfR6La628rC8g+G6H77ikVAs36gp7NuHV+
adx8oNDddGv/jqGqsRiEcIstcFZies0xvX++t26c6Mo6daMjsVliIC2vWuGbCoqArnAooCk5zkjs
SqMto+anp5AewIwQEl7+od8JwhDb6+t3TlIU7yHOAEzaFAwHgvXiGpgKUU4ur1UmcyEpcOGXA0I+
CDoY57AxaM7ecQpECf8U4htK4iJA3iNtPo24VOGqCLb/wTmLvSp39wSz2XpHXq7BbvINYwLvLplU
Po1HXt3WXraIotIGr7yUpIyVjX3wH3QIFsJRl4PRyeLULcSlKwKIlZbNmZjwgb7VZOizbkV60kgG
VJYuXjCMio1mxq1FbW5QepplZ6Tl0O4coIWmUBfLxhkjYHSJywDrUMtk7Nk8ozUl7nvWVsuZJLVo
Fy1DSzh2rMj9ngm956ph1CXX1Lm20v1RtSZAXDGAwzhTHveaobKlIMYLs8Fzf8OsVKgGfYnbVWgM
ioLmCIDb2B208heVkUS1jed65kf0iHV53Nl5OErLcQNmpAyugqWJXMGuaLqonzTtNwYskJi4Coa8
RIkus1kuPE9TWMf66xfBmZtjcz5MmY2l6I+ZxUTYwavvNN0ubY6Fnq1IudnxQyWDwavT1OhmWSRy
/XA+Le41rMiJ0LlVJDAMg3rZxgi6mfMwDeT5fX/njw71W2iaciZIybaj/+hc45lj9zAKmsrrMsK9
4YLiDUivaq8ValbuK/ibFam4VzdGvcNqcSW9aLqLpMh3YCSDKMCFb6r01y6tYsFxkF7mj2gmyh5F
YWMEMpCOfeU783he3wgWGH34cPdcG62NTsDVnoHW6FUOcS0ycbhJqWObBYFvNEhQyjgkNwNeRrp0
nzyBBzvmkwLa2m81wjyf7mpbkawNgmdrD8vJwPq1+z6S9D/ysR0eNxX2DqodqvKJjUMxVTsNTTjW
lt4t82yD9ndJ+j+NoMrBMnvEZNY6EITCPGWtqYN1sUx2f4hWTaZGiLcjbUbXG1Xg3UceUiJRLHCE
SSjUqXfMOn7TdK1YbFeThu1AicOgKYI1l6HPV0RbWOiNhH0GE/5dP0A+QUWahJCdTeGmbzKrZgNZ
ZlVnpmXNHb1xb5gY89ouqfo90PEASTk9S3UK27X7LLbUhkoF7KwAX5hXhZRrp6et7KmwpPL0ArbZ
eicnScLT6isMtrELdIE77zq1CLFKCnXJfI9XHH/XtvxqjNDnvLrUa5+KBNSFds4GLxrH+xIL3gLo
u8hTGB4DF8QSyEQc8c6AvXh3qBlboxcP3JMewKrOVKsNVQEc8e+fcu2zVLl86GIMF4J3j162dTFw
tbJ4hVR6YVc1Ir2Vwomn7hMs3gxautnIysVKOHwKnbNzZnJmbKBzPWp1kxw+IO7FC+Y0wOREzIpF
P3+qAzIIr/hlyLcf+OiPer7gL64qqSjx+5LO3ZvAz+1bKPBRYdgOm+vAVpnkayEq5V64NNbb/2zy
53UWrp4wS9Cpjtw6CCZo1149ql9ZBlQRIUNW2mDIGmyrLfBOsB7Ue8DKLEH4UJoX8tjmlyV1D2ue
ForYHL+6vWc084KfnHnnzVwMm4W+CeK2ldFluGqUbZqRZi3QbT782zeu+4VPNg2kuxuiEcxZL3DW
mRSnfXJEmWP9UUX3ahLvg2c1TCDei1VwIAwOS41YlLUaFY6oObKhfwYBdewm1Pkz+PUgBCLhhNuk
wiFxDI+fVQCbFP2RK9at7pOKGx9pNWICNxUxdNGSPUfoLEVO1exnlFu81b7jzWL1MWHL2vRhW/XV
keljzdnyw8Jj9Y0hvMS52Sqc+4863e/oVTBhqtOEL9FwAgBpCsT3M/OL+vdb0IXCO6J1y8Wk1XKF
ZzTInEHCB0CoYEfPFaE2WjliWRjU34448LWCsYHaFvkJ/WDTAv+9n2hJ11S2lxd7bx50jMvO3FEA
3Pjup3OU6qM32wTZi/LNGbfyzRro8haxmbwxYBlmmCncSBBXn8oSp0WCkH5XP0oW1M44QU+0RkQm
gSSLLGd7jOB5g7um+njFGuUh/2ocXORKd3YWx91czenekrAIaX1nrIvpgPhtGI5WS7SNbgoz+QRi
vde4dEEZyynPSShaOKnSojDrU9xcvA0gRUnlyVpvXCpaqFrh1CtgJqRIFifQrgHElGfkX212yotu
t9HFDoN7mQTzzACFQgVc2cOZcbrpBGUKUUSAXU4kEo6TNrNG5A3FPMG0Yl4VmLcGbek3KQ0J6EWZ
vb/cgGGOnABlm0s1qKmi0D3ODhaMMe07vormJkjYT3luvHoUHobhd17A1VSlohYFSSABo+mVQctL
JuuGTzNYaTT5g0aqrFj2a/GG2yxf0rH//HSq9vx15vH+bv8lsbZYQifOIFQ577GF/wUxhPKTJutp
vP1hpdCVHuYUdeFfUKE+euGtNaQ2OxZMSlJXeZOLF2BalxRInSAZkq760GVGht2719rt5pI6QGzL
rJ4fsFib6mIah2ln2gNhZvALM2uZfU7qusIHM0hwYjt72QpCuGJWYLtsVO+oX7AOtamUZ63Cc/V1
tzVBtFHD+zBm8xOdelct71UxnOoo1db7hrjlsbuH1QYlpcZCV6m0IpanmuHPy3OQ6b9yEVvkd9Cz
iQddR+jijNyIGxoc2cRRrZilj9bSm6iwueexbLwMXSXwCJ+KFsqB0eGxRxGbCft0N9MIYnhLh/UO
VJTd8dGZ5NZUn2hA6gyL1H+LiqzUtrv8dkucn6+jK8gO6f1BtSihZrvtaO1jsXxH464iFrs/nZS/
Y4ksZMRP7WcT4fznTaZs32675xRDC7eWk2lMBm6oOP2JUXUIo6w3UBI19mIMrax8CSlKiMrFt311
dXp3tTxqfbW4tjSZ773APZ0k8qJQBlZu94vie4cqaFC+cm7opWtHk897lN4SXMrUwXAbKD2lQ1oS
WdctDTtuY7D2FyWcvBUy1GTFNz4VZX5vqrsJK8FC20wy7Z93jblcWywX/D62o1LN+gs0kFaZCOMg
twyiyBQxsj1SlQ6PDXcTJDT3CdFSArINkx+sPqIw7jpScS8PV3+4mGfpWJ0pTvBL3HJ+xpuvMpEu
FPFGTSy9MXjLYAaYkOycWXP4a2/RaE2R5oD1vqDqg28JoWgqqZAEs8MLCOs+9ffDq5MfsXKJU1fk
NCl1EPcoTM3DctFYFkt8lEhRLH10H7J4H4i6kxsOtj8vQaOWIvaTIVUeR9LEQQsnZhKgSvSTQZB2
LDdw5Nn4k6wluxoLJ43RUayPhcFuoFUZgRFFO1fDWKr0g2UReiyqkpmIqRnnC4d4DnV5q+ijJ4zd
/teRpDrPcTftDouOr2JkbBQJugHenAXtx4v4H02QXDQ7ZAFYb6Cnaw2aNdOWocoR2iR+4O3xV8pi
+VcWcK4i0ImPc4LWXYdTHG66bPs9qLl+KGPbmUVo9zp36ngLO3gB7PhICXeqBUstnNhi2X8lwx5X
kuTOwjybalP+073RDYMjhER+9LEhjCAuWJi+F5zgJ9eFeNaYqGuFFilIYsDUUUn76MR0bBWtzwtZ
aBDJ9QlXCLOcoH9Hye4Tg8qgvbilwc755NdWHGBDDogkn7Qex78TIpW+DFohdyfIj9EI+bJ9JTB/
pnf4Pw7mIMoIeGX5sIVIYFrjR/PLtu9+BEj9YYypF+gQoq6R4M3z5P3GzE8RWlnLFZyPABY5wFcB
8Pq5Zu9SA/VIR80e8caO0osWh0jXdd9/48MQxW2XeiRv8QymLHJ4N9uui/uHLP/7E//QEwk2eWEF
6a5IW0TPaq62QY6u6EcZUBqSuobng3bMhrdSONNh/t9ueZFn7URGPzAg/zBgmFCn7r1LQhP19nte
P48V73cJhRFq15eWZRTG+5298P+v3kGyYf5WPbaPIYNesvHmABfWEg2YaxEWX10d/UZnBCMrXTrj
ZLmYZ5zcYNwlkjIdkNeVLH8XnTkqipsaNnXqHAcDf92kOWAt6w2sDHHiFqbWzbd4SuBNNueB/AZQ
hPZTOsYBjlybGVa3yTc69fD2P982p8EB4VE7+pZ0BViXO7mLw6cX1y24f6fi0rBY3BOGfZvUG6Zn
7RVeIMRYtSZG9mrGbSf232grDrPwFuxPLdeceSD2mlytAMD06thXHC8eU2lpPaiFKdE3EPQ/O0pv
UDITuI2zBjjF2M2EFTxioWJL15RW1L1RaLNyhGbxeiLTP5be9HXKq65YY7wzJ19FAasUrBu5W8QV
SAaehFphR7mI9ag8Z0PYjYPjtbqsI2LykskvBCFM0pDdQl/oqvyGXhkYip+O+C0FepzhhMnxSslv
2jobc153EIsoHceuHxmwaNrWZruynWs/EVVIUdJkweY75ABxR+xLab7RhIc+e+jZs7M0oIQfOJc6
vBT6/KuxDg6k/2td8lFLg4r8H6ZZrE5uwFRNt2jjxD0FYfPl8E+2lGo2OUNIegAQ623QJTqNH88F
uVRN79HujF/KsIIUxKq8opHwSu5SeHE/Bw/jqTfnHF12GlIxxVwUUZ/Rqi5uXjze8bAkeRXLlCCT
+D2P16Aqd7fTZzhmQyJcl2DiXoZjghWxA2KJj2UoWz5OxoKo8e3jl7OYhoR9wE1aMbv4GhF5I2qG
wWn9dkLGIHwF5cU4p5poVr+e5tEST1FS1z4DjdpedrSdhJTqeeNDhlGQZUXljFMNMOifcDGRC1/o
CrWZimppFlNrhaUIAMRK3ONRFYMhDqos8ooMQBYu9jv4FekXWPFO30R+N+W7troPDfVBBKR/0hq8
9xpuLHpFOn9SJDZf9bpjbYd3z9K8l9ycCpSdB4N7myAj4JImUzC0Rvr9H9ChGU/PK9GtnrlgX5GM
pCdMXqBfBldS4atketyC5tsd9Z41r1tQh/MFLcz3OxJ39wK8X3niU4bLrFeW9l52IThDxRktwh6d
GDcRsQMmn707wpgyb0oEaoWPRy8fIbqJXlI2d1NzhimNeyhmCg+kC5sdaSAwy/2PMIgrMtCrKYZV
2FGi2Mk6y+5T5JDgvQQCJt54eerkwMZh/lvObZ+sZnB0pH0gQs42E25knbbTPbxWHatIV4pwf/5M
+rzj1wa9L7Pw1UDQYqw9ym5YaqUaLwBddGSRYHkUKpf0JPdRto9OJGbtyI6ZGQfHA6knvmlBPmeM
sCLeMI2TgSexVq1IDWbgSJxAQwo3Yd927o+c8SEw3Us18Sz5453ZA9aKzC3dyUIiKdYZSFZTvfFr
OchB63hx/L2I4myM6bMAVxrFKWxKKikQNzj5InehqplSQV1Bh7jvYer/4X3f5nTPYf921Fn2FQmg
okJZ0Ak08CMVp1ZI8b1SDltskGk6hZ3Dy/npNmJp/CdtTiKaKVCON+S1A0t2DPzgaPSwmVOBdIug
AwAOCh+5BQzW1RzPLZf6MpPm+ZEPoFdN3e8KdDANJHcPB9s9SLnePpdUIqaPm2OkxxyAPIDmrNYq
xuBh7Tn+qWnqfRi4cAFC/95xrHcETvofJ/o45yjL3anBO//ucyqT5I7nnsUO2ezztIZPQ15MUGiY
jHXC9q4c2JayZgrZxOPqfIC+u1icSl5KIA5CA+yKT3LwifcUyoKg3kQkxPdpBmCuxxwEWo6tvYUv
CE+7L4qQhgrX9Oen3bRvUazMrREMFD7RJXBvpbI3rvGwa4S3WSGJBGGl23cZfY+j/yc6MZtMUzpw
0Xzpfbywgk915hjULLBRxdcKjM3e1l19AYtfjws9hYhDBZC5J0w0kOpbGqL49mdgIvqqd1YReZij
IzXAbtkS3AH4VgQneo3qwVpK2RhwlZEbsUrPvbtrKzzqR/hoKIk7+vIAhJF/mfhJixMkObZ3kp/n
klGlyO5b4ma7oPtx0eUoU7Pde5jM9TIE76nxhovLKpSmFSE4ROd6bSuXxUTMrHU7bDEPpiRl26O6
9dN6Xm69l29g89k82pCvxpGl2XbS+mgADGy3IaSAaU9XzbNPrY59EBD/ngjBSoq2i9FMogw309lp
xKyHygZ2jJqzIQnyhGZ+fL7TmwH5PKm2FNnXyRfJn2u49US4Y8B+OuUpR5XS2RadbvYHN1uw3znm
a1nSAMc1gZguYMq4mNPgP5cj7ibGzNz9vmd078dyU/Qm0oQYYLlvepZ6Cfp2aaZ6cxcJMOiPS2FJ
f28/dhrl+1pvXKu2GfNY0/DM4l/kJSgAsvEVEmC6e6o/SpCleNWiXkAqA2isxamI3AZ3ycrB6ZlM
BMIahgSOy4GAtMNJGcf/UBqt0P7loUdTUciyvH1ALS277HFdqSsMKOe2S/K/ZfvT4ggM5IywgZ+A
cmOrfVEvFxJjXvFDo/qFMbWsnhYkDIMEe3N5gcQQb/HcJJyk8ZAh+qNusl8xTK73JZ0els612koQ
5Y6T+Hvh59wOyfYn9vgz90qrJN+91Wl9HWGuGC8HKxGJcyLkg+AqwezF96Bs/FRpJeztMaSw/rQO
QrLSIuNDDiQ9KvL/UWnhGx4TH+9CJjUqZtyUdAr34gZPeUilkYmE8/xannBVdh0uFkymrH6GHgjb
oExxBbYawAOtp9idcD+uXIH47sUmWuyQxrly8SAaKPK+ImqShoKC2brIjNDT+sj8cXxOgUuj8Gy9
G5104mUicjMYycUuQHByuj36e7w3mPiUDh/Esd/ylcZHcl/2KqAZK+HgkFEqGpDNsJ+qH1IJ6oXk
8D3UnX21cxioOPWMb4077irtB6+/lRelo1v2QPzTAdrWZCrtIqrj6XTzKBbZZRRiUOF0+LQ3LVQb
9L6YtBgUmyFDQyq8gkW6vCbQ3seoDlQFtYlsbOSnRtGSfi9r1zmYxknYGBk6EYqGDozgGnsOWo3P
qCOMz0Oi+0c0QEFdFBUX6+LEbKmTmOf7tZAVDt4RR04B7NmQSr063OCgY7uZIfNfPEtWSvi1Y6mB
JaFRuH5/WMi6rtjNH14DR9FWnhzTDLE7thB9RZkJZhBVu5S4yHJeb4uFoltKAbeX+nWh8i2aLE1V
PhiWzrK33I/utDcnAd8W8/FRkdZX4CiGquke3rgkLLq9R0f7yINJIW8oB3caaj+/NLNBNx48kIls
MiwHUwZxGQP4W9K0wTSmfKuY9fDSF8VaXJA7Tk1Xwn7Bg6EIw2ebDIBc27ELgUnaCfbGOv+NYx/F
/gqugUMz2uRBiN6V4VA7fJbUSKVG3imlVpMkbREFytNWDDXhUvOrUOjwYO7N8o+qd6rCnP+qH/VW
yEEyCGFQu+5k8Ve3gxY6ndF1VbG3Mqcm9XuOxdYbz6HNRUZrkqWIr0VwzNFcKXneJBNPtaWQULUJ
KESlrHMx2CiY0YG7XQbPmRMLt+dwGSIDbqpkzwb3NjcfC8CL0m5l1+OG6WsK1gjDyLNdL3aN3XXG
V9RWuZlZaZ4cwIZTjmBOYht7rDnyXJ7q/3AzRWy0Bdn7fm0p6QysdELIA0cv2regFilS/E5iiyp8
EWyvm5HuG5borI7aD5fTzHicZM1DDJt3zAa6i3mpyIp+e7LG+xKXD21wyhScE3YIwgMvsJjOTtTp
oEbN/KGsW6KWnve63yeBZPVmI8oxaVFbqClP1EMUVw1aIOXdZG7nnLQLn0uKOE9HEjQqRDrzLXBy
32yt8cjCenalHIuhJ0VNGWI3Wi0yEaDPxGHqlCThUQgWou2qFamq3zEbkxliAC3xpzNVw1EDCbie
bcaHiS0UsosUPrb9GlsYjD8LI7/5B2jrB51tK4I9M6+15yGiyDIBcteIJct3WCHB1YWh5O1mau6Q
PLuOsgp1KhN0VxXep7QFHHgDUA4G+gzq5jziD30V+/PRbhfE11GMNnPeM4tooporFWdXgF0vf/6N
V4qRNvDERJHqKKlFjLNBjohinxcSQroRX1ppkjQyfnqQ1s79LmHRP5U+sy73fRA+PrtMg7rG44oR
6UYn5l2InK1KvW0J2Q+H9moq+pqMmoDkYzzHcM2M3QZrct+zbyBxLnwHWVu4yiqNV6Vm8aXpqqj+
zDo3VGGT8sAuWwzZLK6MpM0a9YR7Gr2JY/XvWCPwkZPejeUahZPwu9acwypElsVfDFMoHN11YyW2
FzKh4ToG4oGI1oGse1jwczuoK3CYzmqLMyXBhRhkkKxz0s1WybUxmI3/2wrXc/0Yl9eHOtaeMadc
YVTyfGd1onuUO1wrurWbD8QLiU5psI2uIkO2NU4jRAg0mDTDhQwrttAood70xfizy2x/ySoAly8A
PaNsRq72OxCHYZia5WwOdp5u6fC0Hlzdgqpq851d+Abr+CU5iRvcz7k/cU7Pd0dvO3PrpJSbyZPC
rCXfClw4YpCNnot/q00uzJyxmdVd7ElI7vf9dNnm1BSWuLGS2kOwAa39EUl6VgS0aY97tQlk+3a7
/fApMSLuBtBHjG6yfvSsc6wZcW27tYGI2eriVpatZrtyVqLoXSOAAJxnsr/hBxmwO6YdnKMOv0w+
3KMeCxjzQeTqt6OE2re3lZSW9xM7GA9wU/wbwVFTmNQNG3Fx7xjqdwU3n0LZXq09O9Ec4uvlJkwQ
yPgV4k3EtE8eKAGsB9Tt20UmCKuEGkKJ0NiHOOPYX+W0E3igvZyQnoRMmmkfX3FMPwMRDfOyj87C
nQYEbWxKSHsLkDCxGPAxKto1SEKJUiDUp+Tzqwv3uNzkNch/r8Va6kBWsze2y7Tbk3owC/1ZdtQk
FXhPqT/6FUwP+Mxztw/ret490U6DzZv4X1aqiDXJU+XG1lfsVHY/PiPCGswmv9UD1rk1fG9MPRep
dN1TfLBF1lHmOv49ge1/cFqBPr7aKq4Z8Aj2FHKDB85QvaE+UkgQoF7PcdOBIf3+uUZEM4lnamp4
Z3gg+9eVPWSfgvHwT2ncadyNXbkh2y5jBFs+amPDHf/vstY3WvKoeJ3ySge2YMPI/HvCI6hFxYMC
cxirdEY2C6IdWQz8zFH6OX56z9/GcaKrE/e7+3hbIrmrmGr+HkHRuYspadMS2cyUp89sbpmojQyg
g1zotimg6j87Pwwt+YG7Y2bTl/6b2CD1gHXVTZLQiXWCvJlDCqFhoS6ClsDcytZm91gqC/dpQNvn
HLLeGA64F2YDRz6ATCAopl8/VKtU5jm3la2QPSjI2B3+dJv9grBzjMUfegqaPTCDFm5Im6hsVl0n
mWVoTLqiigITpaJydhOXrXDCvxlmdqgpzrKbDSlV8kuxTWxz7SursyP014uTwBQqzkL4ZfvFqG6Q
JthXayA0UQFSHi8TQRtqH/NsQw8IeQ7C7y2QDLmr+IhKC5YxeqG2NDqKNwqC17pqaZgcyZ8xsmnn
bMb5t12hqfIr6oh3W8X41qW46yxemOePURN+QBdXCfVk5axCj/YCy+z6E6SjsbyYJMnI0vOBnn90
CJaOjQ1tQi9KaEcNFBAVoJY6js5BBynAqUF4EKDd5c5LvHEhxnS5vtX2fG5XpU9aqfZWiSC6plpn
k7aA+CQoNwQYmfvFmyzRaG9mP+4rDGl9423Pn88J3MDxa61JZ+xbzlJOPpg/wmXuLx7cenBNQGyF
huN7swkK3s11wmkGi1TH/AduhivMreE7FmpxqX1juWg2u4V5Dp+UBljpUQH8qwqM43lIqaDWlnyd
1vPyK+hjVmJAAdOS2bSg8Ni0lg8VrMBc6QhBdgtLsEuZy3vcLjbit1w79ZuOFf+jEH819W/klRlx
XjPlIXbaYsP2X2TwQz+u1vvEkGxKOfCoeFpVsZV3ejDZAxknmSuSW1eV7F1HH6m+1hvWZfFuKyRj
/hGUwppf4Y8v8jnWwDgyYwSIXsxHTQAFv94Sb4AyahHXIM1OX7AS3UbUN1yvT8nHq4OritgFbZyJ
WvQ/JTKDNoiMtuGO4OU2KQDB7TXiQDcNykh7sSc8LY/XzvvU2c9Or+atzeb18JqCEk8EYr6HhbbW
2zNrGMap5zjKM99hUhSUDbVPe5PcUM7IgCz40sDgVOB4ngWqysn4l1LuBLUuwi75K1XC2tgdFwUS
X2EMJbeq9iPhZcqiylISu3bCeFYw2gU8zGq3tQx6W6DWEtNb5RZIdsJ/FmL7o+8w6w1pP7cwHX/u
cABw+wKSWYAGV1jH8I2IAOewaCCcQr5rllpc5Nbq9GuSvyVfk/1dRfwWia9L1rbsHWqi8pJKNmfI
hDnPBZlu8xXSmcX3jmYAyiZR5TEqNAZM7VPRZMOeETwvLGRZ4178zFgHhNII9qjkPPSgkDpnTRBA
r5i345WhWhrk4o0a5dZmeqxQA76rflHM57x35aGhoFjjm/dozVovk9aiyqSZDOb1DcpkrDVRW6Nk
F42jn95AD8iAyPfeavCsVL0fAvdvKtmgl7g/yROfFDUSrvfAFWSFEPxWkRxVofPI3dpWnEZMaZhF
l9ALD8SFcBZHpzEdbdjW85jBNp54Ak2UMmNP49w0zH+qXb+KC2ueYDOTa8ltFknrmCJEWCHysM1v
M6HvfKNOm5SDG8KlBnrqE9uPjcgVTgWF3vURgEJmhsMCgMJ8a7xV3zg/cHct4p3V9bNTKXinefUx
S7aocd3RgYNLxRmYw6U8N8u6GToVVLdQKL633OI/RrgCH1a3ir4GSPQUrRqbq57TQqGfCepi52oL
z5eC6p+Y4o/zVfpq/Byd9ET/oJiEbSsWrnp9Q8lkQY1L1p0eIdBHQsWW+DPJWfzYzILeamFrq3cZ
xXXiAHowtz7d1uMMvmY9wMwrXKwQcoiMU6Iiu6v2MN9uWtL53hSUB/lQcJpzASKuGUfS44lxzuCg
NopIvtQIq/WIPR6MB9QiWZdqjt/IYcxnVVVHffDSOkcpN21ai9l8sCtjEYWZptgBYMnRSQvvcLL4
+Oo9C+OmBH3QU61fivGw9Pza5McK9vRb/cjdJ+8trBuYL+imQr94f4c7QLoTydwGdv6LPYEsRxqQ
hpgUEkunLZF5fnTDHmNaOxnnvBI38f0AZR+cNiAv7V+7whnxOLGtsvqeFa8ACYKNfaSL+HRqdHsM
RAU8iZXpvIYFfc4S9tvDnO3yK4kPTy5EvTel/e9sCAS5GJhltuDixbhK+4+n7CalGBiklbwQ+RKy
e65e/5M5yFSAvxb3/7k7l5YFArYq8yHe0FHzAsxlwhI9PuVMm1IyCk8tdkKYOZBJraGurKoSEXXn
ZXGEyu0DceC3/ffX4VeV+RGJvUc+uf/dwOPp9I0XFAQWenswz5OkzCho4vYOsxsznGGJlFyYn0Jv
c04DbApdT5TWJOMbwlPjs1gFfWCx3ewOd4bl2ZqH8ySt5A4srRBWHFmymZ8PErvSFZj68ISTknyh
eNC8FHiERgx8ZfcJOp0aDT6fFUY/s3EWCYcv6jrBVtkr7++V76C8Tw3Q8vinbACtLQ/Cq46mETQU
+0pGbWNqt2jUaqA4YVFyDq8CqQ9SoYBRlmx9RFPHI/hlHzOm8Nazny3WNr4tpyxNyh3dUQVZWCDT
Jkh9yrfzaSheLxw7GTvtnvNfGywBbE1ya53yRNltmrb/TfLwDAc177CgvqKwH8+Y/1uATtTtrApb
bIyaJmyl+kQXAPwmQ5OTYl5oVNbuCOe9PRQYAAW2HT8aCf9gIdwqEjrLs23Dyz2lGOaCOfaiAuw+
/Hd4UCvikn6ZLWMwke32Sy6kE7D3Jhz27CfxjExHY/Jdm9kXelZTv8yphd/oNfVTkiSIPG6rfFVO
VyopJC8sZf4PJ6hKMyxNOk3j9D2DeSUcShr/M/DLXroDzhiXH7IA9k0HalSxJogVrmTTcqE7FoJI
19CD14pALfkzyOp43d6+uDnNcH7NDBSlQcfmh19Faz6XRvX57RajzM3071OgjS6hicJGtaWmzaV+
mDhvLqkB19SK548XrUeq+hieb4NN8rJXR6tVYSASNES4wZF7GRNObUHRbQn7dfoM6BsyC1woE+F3
1rE5VPtyYkLSNqs4JqxORd37iv8bYh2Z/c1zrkwxrKMleosnAN39o541muZKfdBjxc4sFBJGsI0u
XKQgtyDfTSVnhOKc2b2fnOjJpMSysOHwWjk+aCJbFnnXoEmbpZDRcc2sLrvhW1dGS59Ze+KtYgYJ
QMNrPddWuXQYr1i0pbgRP8BN8bIgNQ0Yylc2ZICFC3u46P+yO8xnSIZHC323vsalNn0dcnAl6bk1
y7HjL0mJB2idE5I+WG2o8ic5KUpLb0T4r31OtP3uxR9qV+bqEz+OFgYAQGYhZgBs5gAM+aKYdOBk
H/GRswRTtaXatFsZcPNDlUIA9HAyUXabDN/Eq6gUSg5NVtzX+1xXke5Qx3nAnVFrzVXoUL+sBpOu
YN1EjP7CkSJUivdN/82KN8qMWNDInW65FLcw718HsJNahyyYC0Ttl/UGFN+T+iujJYRYGG0htR+7
0LFc53jSKgMhxkIbD5ePtnYTt2TA3qHPkPR0/oBZV/Fmrv9ICxZHj/qmSOLwApyBrOEM4f9zOgAq
7sjYulNxZMxYHRDfnCztNOFq/MIskCXbfhOkX6NycygQeuTBX6Iu4V+VO8JOGzQbXQlVCMkOtd7E
UV0dYoeVKVCeMMRQSo0DCGGtgeYO81640n+J49HT9m5oMkmb9u0xTr2xwtrUSGEeau+PSJu8LEnX
AHeuRK7mCr+8qPwmyiflMFfp8aXEcA0dJkSDyozdhX4q924tHtJbYGO2SQ6B7moo4R2/Swi0w7ry
/n73BcHAOJnfyszpyoOo+vMlCrUS1bbMUQwORKGNeTCZErhd7FavsvWKoWexDVs5RcVzkwgFz8jn
TuYMvibrY2ieCiOyioc2ocLJGsqFXHhlYFW0JCtCxluTj6VjVRl/TrQDfwS9iUZmlD9uLSJcN2vY
iIvV+4nM2E9dI2jCywXlSn60L9NTb+6+ZZDYhRl+kil6FZiYqznn0iShQiJ0p/qgJCivRtMZmEpE
1a9AV4kkWTQkIqDtqqtpUeDffV3RO7I2aSCUXy7KEqi0zf/OplNAjlcDRJHPyLUooj2R9w5wt7Ad
o4sLSUDt7KqrgOqZ2s30MtHrDaTY452CxgV3BaWqyfSIIzoWJY9+9PWLA/+mtWMP+PsWGQ42MwHK
t1EPonXxZE8PT2mSqmoSx69xqSGCGfz2eQAl8FmbphHz7bKl9gHm6le9QBL4aC+JzPznW5ey+lDo
0XYN93zyhK6J7O6l8MkzQV15xzbfYqAyYEM4kTeMREGizTJWkDVPeLdhQfkQvxc52ZQB0jib0PZd
xUg98ttkYwVrmj6ogVNH6KyxGU2ACWXh8EgcGaA+OUuVQhUvksJLvuWTL4LSAmr7/fGwiWP+qZWg
4vmnec9aKuwAjq0dVHP5s0SL2gj8RxgSACwi0R/aanX1V8tfc4u8r/sDvD8dEY0jCRxHnYef/0YU
lPuT9+73S6eCwaFJas7Cux5unwKRvDlfPxWb9rqFCIbKi95lvxHDIkLF6VC01XdPSDWWc7qn5ql1
e1QQgR+F60Tuow4k/8yhClF55v75VxOYldbNZHYJUXCr9ve94R0rPc8VGsmykqdVYDkHfft2al+2
8UrsaIkmCJDznx6j7kJxR+r+n4o0HIxeVNJQB3CXZq3vwl6ze7guN3OiDdwiNekizxliKUAipMQw
GzRWW6I54Vxynk8GK6SKcsFCc8BtYhb+7C/0yZUIUN794MvJLTas/H0zMp4H1mKJGJpyQrK/olnB
R6ZN/7JXjAujWAiL3sGedKia65r5fDai7IUAre3JWYaBaqwng5J0cdeUJJL7/6FiEx8la7SdVvXQ
xDEzytGqcvXejpWsJyKjhx+/hc4MY8InwArHoq85shjTbJrQ4tAe5SitAWe5yzCJZ+lFG0MpAyNo
3BQ3lQ7XW76EnZmtpYWAEyzspygWy7Yao+f+U1ybkB97DABIH7oVW5NczWuN+UtNzDOxHJo1hEIV
6h8kJj6u8MmUeUc/svcbhoYnJHcocTCfN0g9ZANDOtoySIrQNi0hjPk5SJnd3KlLQDIcTWNzszTi
qUMn7lHMk/2SYHfR5NPgqlLX70cXREsNStmSlqZpNuN+SB41xOM+XbfsSwY7KCOFxjBe3hiRnYu6
v3kU67kUMf9BjCYeHUfrwcocCunbCbbWy+Wn7fNoolLzViX36klfJGZ9HMP2mS1alDTEq3BPry8q
Q7vNpNpJYSrep7f960Ij4cbOfUJXBjPtOjNIGYuO4V2ZmYQljd2zXIih3GZVw7+XipZfNuaZbx5V
l4uV3cuHyW7OdJ+CXRulN+K2z6OGlreEock4cCBLo98Mk+w3qgytJBHCGvj7+dOxmlgN5W/N92cY
rLEy7ZWtNatXii4nRK+RZMgtUVMmxBH9CIGYrvcV44yyo51dnY9gNgrcoEXQOLb1d9cr7eKia02i
KxYMAKdWGrjFWhJv2o9XV0EMzvhK1wJJlE8TjNODhHQq/JgI8ZmhwJc5ypDQnZqG19GU2O1wihY9
PDzDakqkXqjEqaz9TSSinIkqoqigiROPSR/Pj9OI8FaDrsSwtjPimtGuSgguKEvucCDXwrWYbocX
dmJ5+dFmUN1vRB/qXiANinghxdNwyGyZ9rHtWhgxctCRMObhOEYuYWg45/9W66zW7g3O/C9Ei6Ip
YS5IjpS3kB1erKOjvtLZDvZV2vG6RnUZ5sUUy9RQalzslaWQwMfENJ/KCuWGJ6fJGKT+yx9Gg/gd
M5BUy21nwnArnyhoQkjSN3tuJbcdBM62cAJjASIEJPkCtrsk1WwwSzgkFpcnz1b2h3VB/Wjws++T
Jk83slyBC34b8L4RRJ2tIAHakEMxMI2t0cL2HIVNWXQ2+23mpykZ1IkjXAUJpsnfa4qbiX6FgWaI
SRJoZwnBVas+r2dozXkv2L7pRAvgN/yfg9RxbLVYxHSnuRgjYZrnNu+CjcXx7hDsuBkzdTdTV0Qp
o8frjl0GGkqsH5a8wiZUpgbR72t/wff01ACgeEd6PMwxYPEIzTxklsGNj4qEeY4N3/WgCOskUPDu
nurL4VVyx7jYrUuTp1nosxvGTW8MbhyxzUSzVlbXTGo4Kakm3VcNONxsVWkKU+zaFREHmmHbu4xn
TfWWGyF3dOhJNqO8wLHwr6Ap25vOoMQww7q/zWl8eXWM+z7pm2r5uQjwbPWtQgYV2tNxm01l6aVJ
6bzViK/2c9xR6/Uh9S48oBqHO6rZhqmJQuc2+WyZ5o8Hexwoszps/dQ0/k773n4+NJe2TVH62mVb
G+V0CKYaTFqkIg7E5TtWh/jSRqD2FIUmioxcQkioNWP2+I7HJfuMIErHDieEAo//E8PkkDeiRICh
t6yUC943MvrwRaGGw5rzYdZ4QVA0/QUXpwGXU1wj+hWfONx4QHrAdYMSjSfrAABWY/dLkPFLVa9u
R2ka4NlEe68Yglr+N0FsmiAY0u5yPzaOBHg0qhRja2iE2PctEdneUJyVEpLKYvxOKFlkwbf6A+W3
fKeluuGfQ2/uX+coG5wEaKX7uqRAUMvSDHLiOC2EPIIQl9BR8q8WL6YYUqEGAa8NUDigg31AngCV
NZh5O3T5+tTSgOFJVZ/3tnrYApmawnHuXSiPUIyFaOTWLuzZK3pa31CM5AuYD6eI9siMimZn5PzR
SJ/gmOqG1lE60RWGZpH4ZH1ws6YgcG55yk9LwbdgXFErrixxRDPIJOS91q+hQ3uEN6apqXKdJ5qP
dGgim70agVt+kkVE6RdE8PZ0eKhe3oPJAqN/DiMqnh/opr2wOfHhft51cJn8pBmZbI/rjpzEnhte
e9LVfhIxs5m+6CBjyAKlOnxX43SFrA/eNXh7yJokETWvO1xU26hVfbCWwbor/E764d2avNre8MSd
1G+xN7CeYb+kbN1d6I4Gz2mYRyAIUiFDL5eQ9Uv2D6VHJMGMFAabFF/4mpWvOeZXl6IyxBOD/6D3
EHD3mhfMaor/sL1E+MFxcgjTJz18OYalP9WXhPwX7d+W2ZzQtn1lzRRwYUDbcZ0d42j3sEnws6ri
vpzJ6VuEjGRotl9YvLv/FmEyV5JchBWfvwigpDNb+P4NciwJEtbne7zy+7NDDt6D7RMgBAkZJpoP
mnX2jN8P+9+cYGTbuvwzrp6b1y8RZMMySEHjQjLRheLQjDfeQQ26PKxfnaFiTFp0+fn0lsSsm9Vj
1AmGfrYQRRmCH2C2zjPeSyza6BNYaOPnXYig0XRp8/Da6Pnqamee2dsTlvHPRFvoN4A/Yox3Il9B
LAaUzl2X9SEqV3N9NmG56w/f/lr1TguU5ZFM+f+a4c+h4jWfaeXA/bNPreO/2CfU9iPGmMJGyJv3
TQT64p6wewRKh51K3zk3XOMZkZ3+pRAuMI3PMjHtuy6c4DxqQmn1IhM0O01xikti1GaQHwwj5HwT
Uke5rL81uFoUR45AnBt3iLb7YOADJHYyFIrWjEvSxtcoORYm+86349eRC8eEV30Btg59rIX/nytd
Vb5quUU/F3aEvKWZT1esspkKzwTRixJPYWDU2LSFqhMEwWmexQa+OgHTlBhO0AffztVpaHvYHtAU
GiC7JhucdnlbngufuTM5auG2cNf8J+WlNhr3p/UuFJ+0lWRDRa10gGgLAV1rVkNDq+4V9jJ88erB
KVSNVXmVxumAojuAJ0NLUANZ+FLmaBjfmb59SHYdlDCglxZcUhrnsVs9d4Kp0O2lURZKXfbZu6Z6
oHAWRctYAVcDytVc9xVUT6bsbWKSa9PMSrxFfoiC1xVuqy1PlfGu/MWzW5AGTkIyE7f6IdfhK/0s
YoNPb9X1GNoeVb2CXNbCPBkUYgY7WeF/T/wAczSD+3DSI+bsQONKGRDQMG1fPZycFi9lweKiNov0
zqnmG7fIoL3JeGUFG7KmTkkbvTvZWL/ILb/fOdiI6JJQ/wm4m1Xpi7xbHnSqZZwyIVU01ic85/Vk
uvMNjTTVsho3foLdok+5RmeACjpaVeCbHBEj+lmq2cleinvUa/2OoRrmSEJiClrkfYciXEGwy/et
7po9S62aZy/sX8yO+s5LgEpOhNEuX4K884wIg5Fs9bFUwWEvSo9944l5zD1EscVJoHLbfpJVbtso
jIreclTNKsrjfaVT7xPBWJfGzHMCyCHlmwZDOAjZiyHXk7JhYnpzcFSQfnFWLHrAe+PWkTul6YLE
Qxojm5v9KrI2rgJyp8s5+p85vpXcGBNHp5brKoU2kqdQLA4bUyCxMd7ZNH31DstxvfbzqnBfQkgn
XeaVd3BSu4rUjpBKT6EbwlI+vDDlltCX6AZ2lxQPzQRAzJ0/M/z8lBdt9AQhEk/s9Q9V1Unaw7Ho
RBy+XAhNvNNeXse9tJvq7/xaRjbhCC0TAKc1rnyMj13CUXU/RG5TDbihbp2mxhUQPIAU2phdcM01
JUs6NRAiUs+6P54by5VgssHkNAwhcgArC0MrPSsrEMwckZLxSvbrHKxLuauDugETkrImefuHZEHT
hcq2khznpBIKJXm2+1cihM6UA65VBFVqxuu50EuUXqyzPjsfPKuvJKcg7rqW5iAalQEQG+ms+8Dh
SJyDQkezehQlTpy0p4L2bGOD87JZLP7f3F9lJcHAE78mnuDYSGol2qCV2SeK2Lkx7YxaMow4Phcc
2z33e83jPa/dmS+Wt/qtdKoVbyncesGROiTM3TGA494eOH67JKlyxQ60Ud/2xJB2Fxh+qOVItUUZ
DDlCmsiLqU+A5lMF5/NnGeG75hjws9JpdJ3RwS3m0Q/kLT7xE12CEQoDgw1n1qZM7tkw+LZ8cQqX
GqOdKN7WnNsBtYSLcKkDm0yG/7+zXv9lNoax6koUi63TVdoCHgy2DR/c81NE145yktADVWI2YPcc
raZbMRWz2s8YAmwqG8leHvtcfgBuB2p0aVEl3dizRUsBqdOaiPuYsGKwsHzkKt3aG9vRXvTO971a
1ePaUp1jymGowY7NRmZJD5KlVBTXHQ+2dQSljbnbDn38KfAhVnZXfUUhZRTW9Shg51KnGZRhRwcp
lhdDqinsiP4cBl32xquZq5amV1VVWsbC89Dwj5/FUugQK5pLrCo/kOZ4D/jdAhov3e0SuXxHAGAK
qza4L5pBiToYZCGJ21idvyYO0rsOQomk8NW14Cc3oVh0/EsQdslujC6PE4ao0cHN2A4vJikaWVoY
tBLXD7GW+znu1wUqbTvrOaMOTXZYXK/1lJDz4JAXavd0eX7672e1oRjIHcF1m06XH7TrjEFsIG8D
e7TLYJn2WxsSf1Pne9znT3YvrzluPEiF+rqQL5BaMucmgOZy92ZcPjjpebrhU0I7H44/nez71pCF
RHlm1l0UPyaViofNK/9OEizC2Piukj3i260XcAOr4Bf1qDtqzX2a6ZVu/jXRlr8QoY0PACOBCvXr
jC5UArmyZorJegrhJizR84ktgtAEvBKDiKMjOq+pru9U7mcJpEL4tbFfuajJ5ReiWeVMZG5S0wbt
8fcz02dXgw0hvkKK2xima5Utc1CJvcRR4zjUtJZL7IO131vIJ6CFFtKKmFaFnWo3+3UXHRhkW+zp
Q7XNZyZxNYn2PQzkB4h6Q/phpfeqBEH8znRKlL9LK0BBIuoQ7kBz2Rz+WSMqPaK4WqksNp0gQAfv
cte2M2BfF37hNn21CVyuJe/gpGpxwReeKHq318fexwziwUIVVNgNNciWEIq9cYxlZf2tFGvaiAv2
EkNqc7b5GKcLcEWIvYLFSUAjEI/pJ+zHPG4Jf08MZjFpSvvlAk/uZ0Uyy+JdHKVOQnyPoV8bhVTd
jnuYQDnE5EVAavGiGYyp8ATQfyC3dj6vBrrHiS/VtE58Cfr101Dqt7dQBFT0KWmSpPvYZ3109kE1
KwEHanLJjyeh+YSBZbVql0CDVa/HpnFnJOxcY4+qNF8O1nT0APs0ly4PxkwnGKM0/W6aHGU2bPLZ
+046J/LmDwf4txkWoKVlIlPwtoCZ2QYUthtpJ+CMhrOfJ22wqZKDQ+8qx+VRGVCbQdoiIu9mwT4a
SypvYpOHpaG4yRD1Iq1/CaOI63w2UpXrwZleOJ+ZU3vxB6i4JU8irtHhpRib671aoD8ouhcBAIda
YX3EiXBjOCF+lnObe38MOJk8LuMNokkf2fj6m94OG438+7yM1k+wCKbm+da2aLdD8uqnKleMo1wR
CRzzu6wWh8r1WsHjT8IqyQfFWsNL1LRHTKMuRE3bcbrX3/dJCpDp0gM26UpBCJWI9ZuzaIRI21la
jrYJUnhHXyE5G8LK6Y4g9GUFlbDeoS1hsvFkb22eQFFXJo9Dx3XHoG+5wqBuVmf2FbOxTVwTvQ+d
JUMAst60TTO7sLOX4jti9+aEp+KAug1RD0a9oQKq1rJOQzGfq75lbwp3I/DiFboNTTSf1BmtpSI4
NbwbTUfZDt+Sep54qYjKhZtD9R1G7S4NU3kdRH0nYiZPAV2t2lPhy1yYbPTM47yWSF1xctHY/Byr
L6lTrYPhbXEpV5ue1fkZlVfQrrogLhsOTASL55ldeLxlhwdKREKCFwM4VqH30/tAo7b2vcSDOBDp
hMo0JoPsLLDP8XXhjXZMq0qVpcCY1zHmtZwQbC0IEnAjAmowQbMm+fkeFrS+mX54byeG3nrnC0XO
VuoskEYc/4H4w7U1S/5G3s3GjieHDez31A0fOAerDSpTSZndZdDcPX7Y9a/Txng8+e/CmVCLaa6v
MDmjtgXiuAJa98ATS44Sui+q+86fmhYesidjyMoQnlj0kp2tkMq+M1/2nSKIUv7k5AlBZL1jKBxa
D1CPX+J+ENnjAqSJspzBqjWLh+jAzs2hHm32riwYQO95BEvBF2V5R+BFSeqB9gt/qKA+5kRtJzao
Ksxy3hocEx86nGKR64HdyD9gWTzGQ1D+WsAqhnMJOG6JAx8/yGZbdIdORHBOjc9S83l/iyXUNd7g
If7TIMXSsIeMTZuibwdLl+yfXcyz+Z+g2qgYs/uyxgaQ+azLAKIAPPfnYMw4vmEIv4AZKK+/SfIP
xKvhPReDVRidqesle8DtnhQrFHm2iRKzmgTjdWiJ5GhFVats+IOincP3gdh1MJ12atBirCoqi1PA
55HSDxSpn1+nIYui5xAE0H/yoZGZh3TPslxGv1qGYpVnvWw4NNEV23ga1hbprKbimP7Rq4zt0ONt
2BLTKML3SouPWAgW2bKxIthVZTAq8lWwBNl7NRJH5ess4tiAKSTXL3MmJwz98+VksID+bWXJmfIM
sV23z7KceWGWwEBe2lfrzJUDXTMzaiOiiqBa7BButEV6qbp1G4QVFDGt00IcG7x/o7UPenx/Vwwk
ynS407J+JGVE6TcU/iT94SHr84dW9nTt/l+ohizUzRFuR7B323x5RiaIgMNPXib+alWazo3Zb2Dl
gBD5O5Bteqa6Cgvj9A0UP+PHa1SxDXfX5D03PUeJCWf3jGiQulbkNnjwNSGpcotE4AVtKbO6LN8v
BQRu6l0UZRdLSWMGRJlSaGiSmyCOz43FJcY+asLURaOqe/tbDN6yMD475LDysj2oJRFRv/yzVka/
fJ7qk+ovKeJoNB/l9bxD5JW3qkTYbbGzRWvhmCp0KdmSBfeymDmEqi0Lz1cUCHmTidAjz2Ifh9Fp
vz2IaOTckj7A+98fZJz3HIrpJNIWrcW+VJAoI/yDi8grAX8N2KR/5HDsTzWXZytWyMYuf3g3Zxbk
/YxMXbrGTtI4Btnu4rbPysElXdn/vEu/vxQW+LJpOqMFXNQhkGUH3uQP6jdrWAZCqp4HzBqkCh2a
9wxyp7vB6OF3rnE9NrL/NfKQEq8QxZ+vh9EYlOt6EIJZZnuHqvX3uWgv9a+ZnQquKarjGT4xZGqd
sVqedJX58aqUWToHcGf+wTxWLBzsWqpCh52O2IJ/rgrTVezed3tf1BJXl/bVXxHJE4i75yDBtIiz
0zT5RpMBPxRz+zP7r6zI5w7EB5P4UGguXOI3qfGOeKHDb5GMqoX+iWPemYzDy5gdMP8N8qkryMi8
mloaXGgHKdopdOD4FnDBiRYcnKEYEAMynJlN5oUu7wNkgwZ9I6nF8VWtZMImShQ81+GiwtCo8Slg
Io9sg6v5s66Ebkx7ddvACAR7uVrXDQqht3GaYns8Pwup76e4ftuF3gvbGXX0yXxPYXVheu8ouhzL
2eFTKrU9YVpgk6fclz8JNzwCy550Wmmsx9+QHGJ43ouvazvHl4S9mqf9xciW6Pp8HSqzxXkxD0Eq
6twRFP3EPH5A4ot0KeM+QaFK0m25/ng1zJ5GOr2219tuOy8rCRtMkSBP2rivNMHCaSaebMF9gziG
VwYiT+B0CmSCu6SROQqmaqQcD+tn3WnnGCDEOGvtts8f1LXwj8PV13mJh8wXFl2TStdIXaV5zvMz
3aYeu/sDoM8ooPYmzyqxSA+/9HLbqbNfdck1vxw02JwkPy6/MqF1mdioJnU1FCNUR2dMpuJOzWh+
gZkD9GMLskbfPQNDJu7dZdpKHcKCqEGUZfxQsjum4l1SAz5/a2RMnTXyUtPAocgHb58QE2pLMl+y
b/7JZoA6LgUa5dvhWXJ3Ftke4Sdq644QT1j4a8i8p2SCuCZ3aM5YAojwBC4Fybt7erRJqB72aiNG
HVvgKGnkrg6bh2ZCv560Rf0fzqRdGosrWuDt4/rGe3s+WXuLos6bxmXfHgCV/vR5J/XtOJ7bV41y
zJb2SB0RbBK/QZZGOFKL/xZuI6zcTasRhwjGVifwe6hj13RR3KllbS7PoT0OtUZZJZSHqtz3t2Wh
QUa2VQhJV+YsGK/6dmOEKjUywuWQybn02fVDYqhLwZyjn2IrX8GVncYr0GIiH6yqRtybTu2Zr21U
DmjdYUe43micv58i9i8ZBExWGhxSndRy6luYfj77fZTXvm/pOwqb263HBkWul1GrKtD9goEFeTki
pjRec26/sQmtlCZN/urReGZiTFq6wxy0tJ55JMmM0hZAYi9PeY93Si97fg6eL8xMiyvFU+Z+vXtN
C58PSbRpfcwO4v9PHYS3N2pIK71lfM6ytVejGEHCVe3hbSo1vSZc5bc9BPQrgGtnDHz7DFMKSXMi
wRuDAaG8dR3pRhSeZ9roQ9Yu7qqQPImLjY14DeYFYs9qzNAdDqembH93CH80Aljz/kRzDhfV3pUb
zBpw445tdu9Fn7JML/jpQGzuUObjLrvq9XvvAYAFlzsKwHm5f20wPdUC0t3w/mN2rsIHdYnp517i
nGPlUAHQBvrCzGIuWkkKSRi+jdG1IUDIG0+O3xVO4aJv0DS1S63y3CzUi1/I5I5nUmfj8nGIPuYu
PK6sBFa9GNXvwPycskYzV3YtT+JbAAzFj3lQ0XeM4vIHyEDjkLPHCMW8I80Q60DbPVE2lY7Kpryd
or+8ws4gi3GSgTwUIXSYQhzZyUVM1JO+oU2DGy5q+ztbOR3dRItlGz2a417d36sjuTxL+z7gEdAF
iTlnewo0/bJC7oAeqwRdjbs0Xzkuoep1Bm0bWj+02kAfYZuDEy5gKth4P8+TRIXbrc8VW/CT0NDj
CKilVN9JciJFNbZh7PvjZEKtKdxbibNKdUKWXaLGWz33zqWMdPwWBCKsO5svdJm7S4Tt7Eltm8Q0
eLTyE5S0coSp+B1kKjC1hdKQzGsb3RAsa41nwXFmsUZxuHiSlXaf8CuPzsRZYoGHay/tHy0dZkYc
lbo1HscHgLZLNZoWLyWhh59GZKQhKuyELEuCwyefKdUSxWF8uZHc30B6xZKlL0/5Wmwly7fb6cdF
pVU4tCfS70CWMjVUW77g0YIcFjKtnMmPejEp4UFkdfjPCFpn+Tmtpuew0nXYuTjl8J6Q6NIoim0k
/UE589gbfhOj9eBVL4RbFg3wkZ2cnBUfeepB39bv+EVANUdX8tvPJyzdGA4uC3nMch/ED2Ides6I
c9cP21jEc/zZdxegEZY6nEeuJqnPDOCMh0QuIdTUZZ5Tq4JDWMViRNjnG7W5C1+itpQ9iPmubuIa
nRPwFxbcVzbPXlyQLY4saElRAOb32Nn8Q7CS7f3rgrOuSSj+utLnFK87R45cADv7Hq52yZvv6bO7
mOgp8wbcJ5fAXmKuyKwFZygjtQsKhT58nALA4X+noObAcRnN7ahrcZYtUQt0ndCXhBoKggfqq36b
1YLH1p+XtNUWqNkxngHnlnEhpy4fjaiO7IK03QqUB0jngxrgZ2n9SaiJKyGU3TR0CET7kQtjPx7V
PZGSK2wUNaqF84ngQ2Xf0HjS229HGu7Xu6HDKR24X4kQkWzt+9tcXGGjPtLi11QiEjO8lP8stno+
BvIDjRhEqbfbSJsHA8qjk+0bzV6qpBgvZr3/+u1KUgsa+UL7MHNb86L4IVIrn3TK0VM+XWdtuyNr
R0v/yhccDbonJJS5fqeov0sdXx2iP1c856VpsVTGt1reeNNYpAMXFMbZHgfaawM+wrDMOsm1MnDJ
a8dEUWOrI9DD8nyPl/57TRwqWYg3paTLjDnJU1EuncxVGZouBvlNH2VlfbGN5Yqqu2dweC2yUfKg
A7lMNLEvufXoSHQTTTsuyb+9W2IigkiEsboNF7aPHgha7n4Vk7bw5b1WDZGE1UdMSEx+zdiV3g7L
W9XLMyEYqPHJl4BjlupwTIq4kC7mJHQpMQFBkLkQ9f/pnFEzn4q0q/BbJ9OsGlUZ8EnhV3/T/klX
Usq57+mbr0IhdMSNkfRsr4q8A1Ox345EVS96w3CI/cddJFDVNMhZkk14bd8MGu4e5/unaVu+7LIq
Ih6mcKJq5qolP1llR0aasjkn+g5wJ7PWvo+RgBjDxy/d6tiqUIXiqaQgYQoW3yi8FrW/4MTYCTPI
UbecxiivtfvqwAe+oKyLMj9g7y1EHYHHBBw38WDgoeewjkr8mywp4FLVksIDpWgi8tUtE8X84HTr
/qLMmbdOaleo9XXoghmV7iLq8TG4O7pWDgcllAzRWzd0gpHBTyKLkzgWFRIkp0ry8X4A6eDPHzTY
d3B+vOzeZryTvwu/6EADBWsn6Sd+5BZyV+Sxrh0tQ2FTIUD46Lg/n0Cte5N9ZyIAstVFDIMbHobD
7ulXVDX07D2WsyIwNesRI/C42FPyct1OnUFhRrjubm8l7khTo1sML/mdldEeJEq6rUzd4t0q0O+J
f7gA0ppW5HATOCvLPAFKrAe/lgHOxY7OsnBVT8UppCUQLY9ZWCnNzrTrnj+Xj1td0xsQRv+QvgDd
TzfX9KvV6LWAs7jEqgn94CFYi7veGJDQd61mq6xRPIwXpBiRCP6MJvMIEjlYaTkQIGm4oHpgJpHI
t6+3HytuWTbABWYiYhq9iGWjJt5zwe8DJLtOIoVFQ5nBltP8y/3braYJH+IiLk4KzdqyO4CIUcKQ
Bcjak1fSe7E3COsjrdU+/6MsjG2xDlIx5+FxwcmaisoxX89Ba1Q/27I5n7MP1rb1LAtI/R3s21kO
etV9WMYVx43VdozJVRMVgveOlhv6ntV/KokrJGHewQVjLo8lDLWXliCS0JLw3/hz7VrZVYeYYY02
BzqzR81tptpI62yv1pY5SXJl2hcjAT0vaz/nAXqsEJmOLQC7AGEqUqW5l0PCJAd0twdotrzus3to
ZB0mxCPnzSjLlaaV97+0ZpQ84zS6eG7vhRJoHhxlg3enjKZLGC27abDeKhtbBOrsO5lomUpiW0p8
G5PU+pxl9M1KC603oK6aigLU3hi8MvfLarU1pNmDvJqXZaLzyb+9+vN5wEX8vJBThcEDj1TfWND/
5n7QKf4t89kY5BDHGIvL/TthqcF3A+4VFIyTZ5d6fw1hAPJJaaUmeQjDEJTEql7reDd8lXBn/Th9
ilbwtwCi7ktcjm4yrjwX1NAzNxbbT79O3O3yVD/7UKRgyV/lz/YG5Oj8toQ6AcEqI1FfT4Qz61RS
oOMvD+t71fhwFoSeaB9j5ULKRwA3zleoYgMlAxcEdyvG6f6wrq5iacstSe1uE6WXPPq76ZAOZBdD
BgiVPMwh2bXvseJyj79um8/8ii+wN6tjPqzDBOeZrBWwy9VBGuxFIyjfzIrEZpol3M5GKYgrGJfW
fOcc915O0aZq/t5ut3sXFxZIFVuDiG3B5YN5kPMyfkRJ+9cMwEBMnOJeE3pPsY1e1y5uZcbjKbOT
0Jr3DN/UuH6Wo2rh4raARlwbljmHc740n+52WkSLgOfrxLvhFEYFX4kZ3aOPVx8c5ojjGY6ihE7w
cIHlM4eXVdLccG7mqvwNF4lcSWWC5ppVW2NVThtHRYe3NrLG3M8H5rPrz7gsvE8p1XejOM2I0lkg
4YTPD8y1iPjpH+hC3VtTTCtF0vK0gc/V4MmiRqF04pwPUFCKA1zUQoIGcsZftIy5ZZjyMMNBq+A4
TdRJnOD01HmqKcIZNffSVD8D0jcLWEceWz3b1wbWSB7jwugZ8++6ID/qhO29lDXmiGmTEO3dzkhq
uSjCdrta6e76YfblyKCy2cyB+MzABQIALxdOlr2hsm8mnNNjOy40Ny7L3p1hyXszBs82rZPv4TO3
tuZxzQpi3CuEoPUvtqQi5uOD6nXkZlXafkci5aM4LZU0bqEjFdz+1DjbmIGVmNgkDssKuEmC7T3R
zrxlemO0KtZ7qY/+KWHb9PgMIv+m5xBcm+xZKXnuC6Mk2OZUGvBglflVTVQxyfjsQ6w3rpsiOpEO
t6CU3J5Ms6YDv+/am4+Crnr1i35yg+AnPzLFktpZHd6F4HY1j3MU9oCzuHIOYe5cHf0ZIEUMDCH2
dLCKfpbPzh9jr1MzdPuCUWRob3LwDGBVcVYSIw2kp5etqAcsPP4uFAqPtlaL+Z9ww2+gZo5aKppK
4C4rvnApgjnZfirsCmOqBTrAkL4vssPNgBeLkblh2rAM/lKZ3q9wDKOlMs4hoqWctHYJZSoHfbqf
H1mxkIx0snfl5MK8onyxbt592GP2NRoTxvnC4Go04o9MMtEeNZpLK7H8DAHRboff1/F3vzJGAbYD
F/HuVTC6n1VvLW5Tedg566Q16D56EAIW7alUGvn6OCJhLTHPt8dCoTr5aMiqc73ZsDl9smc7RVRF
byVHFZvRzK2dVy9Q0nDJGULyU6buR+DyW5HerobcSsafpIjM8M6a+St/apfqqJeE1T8I524ClvzG
oQWk4whxCHGLAn2DOUNt1Zer/ffmvcoScU+I96V+DMECGXlouoLdoAJmN2z2shojLK4NJ5OUCcus
h+fFWEDvKeb6xqvf38bjQeuV8u8FwjZyG2860vebY9BpQmSsVI1iczqL9u/bcxqZRgk0qznMg2zV
0P6Lao2E0mvyiVsIuLqKcD46Lh7ll8JkQe3pjKYcLoOBjZhsXtDlKey/Nvw865z/jAOsJVjBXqoq
VoCXtEz4WLdx2sExKQ/b1316/JfVwce0HrIzv4wnzqJuSOM/ywER7F7a5H3gI3r9cOZSCguAUfIz
dqVQcyw0aDFzvv0gG7meH+ey8DRaODMkVtqA8X7GwORrKQO5cNkHImsiM7wKJxEmsGsgfkgsNfSI
DtlVYjDAmD9G2aZIyfkcl+Pzx1qRqNYKkIkCS4gjMacpZhTu/wUT/A2TwEIlYEmvg/H1YmrauhNu
SS7yd+7znGL+tuKE4Gfgc6Zwh7rZJFc+Erys3499BsbVZCd5OuKALvfGbSaIPXWmk7OAPe+XhmSX
glPTlD7CQwqX/h5pdcpHK5Tl9ya3ld2LDht1JW5Zr64XNGcYQzF+o7W5vbPgvK/z4Ts7jc/UWTbU
cfoK0kOIsL/l5bHZoVmfPfE4fziXxVUn5cLeZFhZBzFX2z1qgC/e5dvjeCW+f4fWc4u2xzlilNWw
/oCwB4ah+Z6OIzFz9feE1DJkWNpsVroLBQsh37B9u8uiFyLre7nCwwmQOenJefFqo3q2fHhLEGN6
f5Z37LveFAJajx/uA5wNgpSbAFIuw5QjWaTdYbIpdEGWeyWs4VyC+0Lnmr1xuPgWsiHFqkaSmYaN
NwBM2J6ZJeCrPyeMzOVQ5FKTbxTvnoNcMKIn0pfsPaWzcrpztS5yswYF7GiAtU0ywYvRtJgF/2yp
7o+qMPAOz1Moogx+O2E2aI5wdgPy2DtECUa1jYH4DZUi/J30H+MFVJ+JhRzpc9IkHOYqCy63zrad
b61mMZU7ZNW1058QkC/I3Jfrz1k9PaI42P8W4pNuLuVqH72ztSPrTnZs0roEWn/xQ9OC9IwroXfB
gMHfRVB94deKVc3EnkiMrX+5D5kITchWXLwy1duS59FKXzqwoUq0r10pYafAaOIL9n/3Ff+6l59c
rYlu0YpHKf2MWkBBS2sNjEW83nPCuFVxAeT69wJ6qSr6hxUAa7goFTIgBVN0xA3JeIjwCFG0HmGn
VCZXDCJpjlWWbhRodi1MsrUzUDg2ZTaifG/kLlCq07tNq5PxwhTkV33cotRM+TwYenZ1WohWHLuI
5kvDLHuN/RhwvgDmzUUJApOGFLF7a+hMQN9wH8CTIH8TapSvqJOQlD27Alb6K8JeD/1fc+0h0jKv
HfP7vKDl9NwvPoKsggVLYodg8td4/DdoGf1Hqu+4fleiWU2TrN/B/TYMWPUv0f7EZ8lMMkQHr5e8
Dd0wjnH1thJFUAsqpK1J5iRAOadW1rLPYzJgtfLz0zQojncNRqd3Nm6WbRvTjfQOeCCFgqZpcX6M
uA85aUR/esTloXeJS1RvgRmxi7S77AjzU75eKt+zeiWPGhGzOgRWZJIC+TLUmhl75D0cA40bNDQs
m1oKiUIf0D6XlzdjLjIJlH1HnOFMFvK1/IUxD8zc+FCPSlyTbVkHXEws/6OssdZlwSqswInn5o4z
Wbwj+Y97jsTyI5ZdHaKyiqVLfSDL2QphLSXWvlvhhEpVOuU8BNT8ZqNPbLhVCrrdp4cd7HmbKreG
8Ea4eKlS0B1uMRWtumWiObbMVSewO5rGsNWiGIG1/WE0XxdRHWsKbNa/GU45ORrjj3QX2xYpR4oe
tCBUazsP51CoHVhpfJmpLBwy9zQP8NzuPfSIARzgExIwjfzp6HgUm02Fj+a6bo4/0ERNZKCHadAu
nhQsuTyXp3jxYBfDRtcZSflUHtFEgpGrEIqL5rmyYOvbwwfLs847+p9aR4mwT0k1hljgs0qU5ZXs
gQuwusjBNhguFbKpMD1HjJKlXbBwp2Ty5a+Xvmnosimn/rVhSqmkKPf5ZfNBKaQi4syAdBreJUqE
ph6ierOpCGBbA0RoMaNO16ZlsX1yvNSxderyY6VFoL7S2Dbs9xYRZzfJUozTMS/jBvmopcFdhdoo
eiZGiOuvtjqiw7PkhEae1qpoOEuXB1ipIdR3jrDiiLnkIlnN/kvjZ3RnwQc0W2+WMvrVV24EEp8Y
q6uEHaMNFCZ0u0NjOECvtdRXwyODxVY9Ge43qmazquQDjJstkIDQ1fYmeHW9nCkyNjBS7DH+No8/
fDC6Szl+TvoqAwXwIB2hmZ7XkOjUm4vVCe4YTsuK4KMBz/lqpiALHXd3IF1v4hb0o3sccGjDvShC
jE5L9aJkGo6uLavluP8guZ1Tfv+eYf3fRbTAP95MrhEFc72esT7Q8vHf6nBHNS0MVUJBLiX7J3P4
V9kVUa30XG3nyyP1l6OE9SLmAs1vds4Sie+u1b1dgkvaNSPlvvT923TQm3IiSkFdolv7foDDSN9O
gZrvA7U4N9VjVNRuTO0zuu4A2EOFi1YvkQCqS0wG/bBKSY8PK1z9V7oJluLa7WxKBMuQvRNUryAh
lyGbsZwn4yAM1n8PBHJrPOtK6GmecHOz5aGQga8x3NwsF6rZMnTJxEOdVBSt+XEShgwQLeOacWco
fRxypbaTna+Wh4/Kd8zkHQ0vjnlOde3SojRNU+QySaqMwdnLUpywgZj12sI0XEBfVmIo8za+cjhA
oez167CIUDFe8hPIQ3rbq4wfXEZuiYTjvZi7HChnMoMJb9d7v+gcQSPaffQZU5ifvQb2HXOFUX/D
ZUxjkReTnzM5T25W2pCZrOpLsJb0QXQ4H4zMawO+14GG27/cD3XFV0JmgfzOu6g4neNMRQPmzI3j
Qtv7nVT3sFDVYy/coPZt7+qHdHS0uuKmJpFk0O97J9aNgSJY05qNzNUV1+Kk+4wOd7lvF3xAEKEe
3htzTz2+8Zb7D9ckiE6VaOr6n1o3OOOsmEUWAQLvlhcpqLU+MXhMoRJpCEl7maWrodz0fEE1ce2M
K3IAHAO0A6IH3CzQr/PKNi9SejGrwH/iXUMCUIQL0BcwxSdppq4s3kEBkRYz7i5szmuK0bVFB79p
wGvnNa9omnx95Ct98yggM/sWKx847KOKiekk1KzyYQdHzttI+CtmxqX4mdVCJfot0oyJ+eRIJXkw
KEw3j4R3KPuzBkcS54Zdz3PC50f7JJwCVRD3D2DWrUgswdHfBefKsynlr3XLpRCWS6JcP8HgjFii
9eiNXzAUAII0nh8BCujAXdRwCG1ev4lsh5TA5P5VDK76EUqhsKwKEn8n9Nk4jrjb7uo0UI87F6jq
5by6beveihevoFvcQuIg4Q5v2meaaI3Wb4qFv57nknyx8w6ovqyggsVXAV7dWs5nev76mB4TXA4r
7GxJvLsGStXWyCHPmtvzu2nszP4uBD94jFqAaSrMQalJwhs0o/5OgnbDcZVABjjxRIAuTUhkJ0rl
8R49jWekRKFULbJo339KC63QFOHjGcR+Y+6u2DkhvqTPsO7gSrixzDW5B7ZRAxbp8sYjfVqoptB+
bAJ8fseo1yhRMoeRI02O16U8Wd5s22N/tZ0Nzz9abpFhmsMTPJaUT1IqfFdb3+thTLKI1XJ5yIhX
hbeEsL/0D7ZoA68K9dn6tFbYmasFfXiAsc/eCRy+toKVwgfvIT9bjJtg4lV0T6nBTKbbzp7aOpNV
pHbN/24PpYNrmF6Cd1BJab62J0pA2drYvMog3RkK4wTpl6BhbX0t0KZJWADlNHOtNo2zer2Zt2RH
bVeOYr+QCgORioAi9tBXBN20HbP+jCOsTLENB+gc5ilalKVYGN6/jsVqTQNRrYJp7Tvy9sDiAa4M
7yFk+a58lrQgUky1+ak4xpqgoorC8MJkQiN+5Ev8pRxJ+s2Wx1WRUxCPk9Vzn4dDA9boU1nWdnmJ
kWK+WlSltFs1W/TDbIztHlFlUGGu7LwyXWxW2H0n7fYf8L+kZwDGSuB+GMTc3jF10Eoj54MCfoLp
ZnDIbw43AadFyV/8bfcivLuJGnmPHt78k87uf2M/NHe/vI+LZ1E2H9xxhow8dalZg96NSfNdAIrA
cYxjuDk/tqam7XoJdkoGT7eT9v73QJiTv4GFTtceNKAe2Z25HC7XMMGoYuz0OjQiK1U+VWV21UGa
JbzV4dcsUrn/BDHbRoRj/xA/cCqoRC5RjtBalkCshheGxRvbfEhxZrIiyCRtp0utv51OMs5U/71a
YLcreDotxMRb0Qk/eLsuolf/FRYc6FYcWRAEjN7qDXChdkE+ySvF1ITIbQb7m1+Ob8mZ+WhR2QrQ
JOkdpKJYGYJlLHPzEHdxxYwizAIfrr+ZKht0OVMswWTXbKS9YkBPLsmP5U1uoM6juDNcJ7rBSvtt
HPZNdNrNauL/ME9CAwP6PsbaZriUe7v1FVNx3AwIP3uWIyVO8slOsp6BqHpeivQ84XCEXBIGOfLB
E4kPUewfOC7BcCDR7kQLr4A9K8wgfOKmluUFkVZq7OPOgOYRlXWnjM9qwazIJGMtQZJkc5IErNfH
m2vxernh15BQ4sQgTB6ny0bX+3Q6DcX8+2MmlOWUSbz5BoGXMmDGaN5rKfEhRuo0VG9NYcYSUPsc
/x+kHjLiNMnUymNKA43pS5S7RJfvuhrSb6cGYhn7UGwUOcxHDNY2U2F3FIN1KSFgndPQAlY1Jaix
pIinJZAwjfeU2hml7X47cGLZLHgaJpiQD9nvqBcNX30sGfUeId4KbClvMVviHzC8sHQJykAAIm0f
6J9geFsEW7/Z5dzN7rb5XelLcsfBJYogWaxfuxKXtn/MTrpEQ1oCVJ/UfYHYjDoBd/Fdlc6jKlM9
5Ruy5ra2c7lU8fMLA6irc1j6r1eAM/Wp6dsv2N8f3EfuAfXXZVsqP56VebHAKa9nR+nwMKFKJ2XL
lN9ClsTKTXIL3n7tOuvFTEMNjxtfFJddKNwrWEBDbYi+Lwo5ZhqVTCLdFyRhJL0gWB0q/tgR7FU8
DObWdw6aNAqkseaOn9729Vg3PAvAJ8tfvWXZsFjmOXcEz5l6s2y56yC/CbnAdUroYUXn3M5ZrzwO
3nMZYqNQdhbDmtRE6M/W6ivFYJZNk68A+dV9OP4myq5rkivQzlrKQfTxrHUQw9zJVH/dGmFiWiX/
EXMwp8N1iZQNn7kIpkIFARkL1OP1bmdmv7awVIeSo/C8hJI3Bj7jLUmMPzHSZpfdfNfqJ1w41eSM
FFio8H1Va9ac3hUVAjMcPdph3M2JLz+KXcKKduq0Wrw8YQM7rYAvxmo//LEIE996zR93mJg/0I9E
r68nbsinHap7motuyCNfFxrdycpnL1NutYw1O6n0nyblRE436daorwrpRSnsYHHaE6ae+mRU5zSP
TZYBfZIEoS0RYZG1Djlx+BBKENvhuLBawo4A2lggi8J7xTkSs9hazIIvp0ld/jc8DbT4HtqqBjzz
9hX7hKjSp1VluapElbo9xE6ekQ2ZYdaoHifVwDKloZjcohRygXqdsWnE85WcNq/S8DKbqKuWI9zX
ltI1NpWg+1Joh4x3zYHPXOLjYKQRn3NQQLeDgSNcjiG9awjf3NN8XPrWk/jslptwpkIfUWq0K9/m
n05ySYHOkXRn2Y1SjchFR2ao43pgf56ZL7dc6z0Iwx8joXTKy9BlVwyojLabVnMN56TQPbje15Hq
CUt4WvONELpaLar+c/jxGMwnaS4o//dGILjd2hZ5TNxwUD8kqJQaV1l7N9bKRLR66fDhsC7HyvOm
rcBRluswZ2IUIWpsVWNcsgYSVTw1IE5MRPWPfGCFdx8mvuByRLJD4PG5tQShwnNhC9izGy0+uGi0
ULS5iiY/BRdb/NNby9/XYm9pffNxBJsaAsr5tbJfnRF5bVJFwelVIRr2CeGjATU9/MVlJaNQ+tTm
QRO7fyG/8tbEoY5rbIhfO9OhU+nbMCfjEGfoKqeWVVpm+R/f+UcYGd7G46n9A7GT/I8kfirkH0+Y
xYuXiRdro1oFfAaK9Ez8XE2JbyfgS5RAkvDtqeuRmmprh3rnmvBU0zo8OVCNMySu+J50WAjBNz2E
3e0q9BcNku4HO+TVeeJUkOgqMquMbewDQNikuHCpcBRNwv9uPempi+1On8afAI+nnhHZZiGiMgF/
Q5xEN7ybF8FpoPjiWxYzhz3Ut3JF+03MXbEnoxjERwQu4zIvQW9dcCIy2Xo4KDgOCzgSTcQN+qh2
oIqr/mP58ljfh5dsnn7PLdjSsSOdNy9Kn736ysa2jO5B6/ZmrY0b51VkoTMcQFbVU+0hRIyU+lpt
T01EmXDyhGpKc11qMUntRkrZQCSuyYWhadQ/r+2k4hdrFvMFhGAljHr3FgIib0qLi1oQUJbUtuFs
nghPC0erZwDunc9mq1F8B5mXKKwzvrgPLPtRaAqt4hRGHw1Y4Yiql4Faw7CAFumjimK1JV1097WL
OmexRkrVBa7A8ANHQRN7JKajZngpnOkIeRgSATl2ARP2iCMdy+IpRlxgFXvJThF2Vhfxg8VrAV8U
D7IsW/A7V5Z+c2nF6qWZeIe+TfrfZMjMRJtDGbnM9PwojtMbBh7YX0zC7WYi+i+JTIUppHEKv+QF
iXtsAkDHBl4ANLQSoahjuec6+Sx1Qi5UEOySAAqx8uL86oI4t/uBS+DxJK7UMqMSkg3QpQIxqlHo
Gc2LvF+hHIBI6xLtXJIRuOYFCMIzTtIQ5H4/j3DXTrX+seGWskf3E5NML7117bRfMo1SeWXLblBw
dXvOXkkwOgfsN51cW0gvS0vKwBDNENSc1mnJyDbvZRSUkFzWeqUr3J/V7UCSvtsCdMr3Jmqkcrpj
+kQBs0veGsgRISE4RnSgwojpJMPHUDQMNkQToluonTRp84QwJpkBfxVScjhA8EWVUBcXLGKgorKP
M5lrx63kfF/lMGN/TSHBcpklE2t3P7e+ecpnaa/kxkmD4YthcxomtGbayc9MOHDto8kqczUybr+G
XTfI2tbNrSv+PjoZ7OCOBXgZG3jlFoKGZTSVXdar8Rm7GtUozZ0pq9+/Y0UssYQ8KDrFPrWpZVxZ
jBi31GoxNgESoHy2ETgoC18U3N+fM31F1f/1g4NjBp6JAk9461fbO3Mi4XmEpHwOnR048wGE8Ej5
/u90MzZVNw7n/xhXY3aI7DHQgoaQnBL87LdUtfGxew+zDGU3HQvlx6vWNkllaMyqZ186sm4A/A42
f6AwkTrkfgbYXcvPylfkO+mFy9d8IhTAp7VkOim4tWq4WmrYkYEV89AgPzIdCmrPVfeSkI1HhOxh
ZFqI4gjsH4qBk1ZwWU2U7DvULFgWm94MEUOZMJbujxA4HylmvlXSO13tnaUeH6HhGhiWmqVdbdtv
eQX6Xmcz1BxYrVFGUF6j/KCJs5uYf8OWKzl6Qly/MosVPiIaT7zn/l0kApTNoGlMWqieFBoGOqTg
mXB69m/lzUg/lkJNyie99QUHyKAU4ZTrvcRW3WVM94UlpDBP6S0W3fik43bkEcY0Myt3Rezf+3Xa
qIol84Ee6b9fyo3ghbaAax3nkEhFJ7HrZrMVIdtOvj8YZnwQXVr3R55+p4+sSpkfdN9mhF5f1wkG
oYWMyBv6odCTcYwtFJyp5maGsW2nRFpctZB3RUBJ8EBszJdCIEDJy2B5Jma9tQ5I9dpAY04hhXin
Oq2XAvr+cwWHoKRlHgQg3Q3iTFuXOk7tpQ7zNNd9S3331sKX1W2v4XQLkcnBzBjgBhedTvOobd3x
aeA/FTA+gvXZ0QAlWFO1K733Z5iuFn56Oa+7pAAotktXg026jEkGxnADfI6zhuQufCeV8MQUY6az
Kk+C3foz+6+3miQz/mpklvn3Ap3y3KDX40bGJuGYQ479bRd0rtZf3o+X0Re2mkEflFPEDB52yoYd
iDUTFle+n8SgEQ4226tO9iKPUoiQfsikWEhoKlBGWuVO75F9pgDYOQDakrYWzDEbwHT4TOaoit5r
UU7Lod5gPjQ55npt/Kf6rnvSt+zavpI+oa2Uk3wNlAoEJX/ac4+G0Jfl3LYm0llEga4oB8jgHySd
s7ZdYBsRoixZMRsRKKJ/0kAN4jOPo11d12tmsQv468plN+mVyZ8FOouHZO0C+xkhkYyeGgZB6Gf9
dod3Mf+NSyINd0QN8RZlgZ14a5d01cTNyaS6QD/e7T0xk1d3eWneJsOHFLWqLIibZWDo5RCObstg
DB9uBd9QfLZXvaTlXO4CFSRTxplc5Ke26TBBWN9VdcILKGaKceSpNboDZdV1tInOGM42Squ5UJie
LlE64Kk8lCvAzUvEFFjrwjikqEAQR26UtyIsN7h824QqxbVeUkWhUDeyjqcfNxmoiQcL+ymMqQy7
c7JDKkvdVA/NobCS7Dv9aeHa6XzChuNy3VIIiH76Lb+auPu8jbNrr9Byr/v4KwTDqXMZSLzHg5Mf
bjw73wzb0BwkREN7lI2ykSqYLoc/tXzcOcEqaqHDOIG2EVWVG8G70Nxh1bq56axM/BffBi/Dpm44
zorKhFKguFqEFPtp6+zRvEdZf3UU3E1PtULM+HPOi0p5s8Hg+BL/xm+xTo8JvgtBJkBLtnPwrWqG
8aXIeg40IVhmYU2M8TUpb1fCOqNCEcIh0GVL8mecT/+TQtfR/MUJzgvkXkwHZ0lMi8GrjrbT5uN3
tKoMRku5+xMAiU038D4aVa4rPagCrlj4doLDrdr2CY9BCB4j5ggBRRbzq81VNOXiuqEV75c0MZLb
JxJwLQHvAkUYRWHBiEkclJRKWIIeeNOLw4dB7+9zFUVo6ZM8Oq/RcGf8DED+J8STJnlTIDEuTa+v
NgKPYnNo5pXAEjlHgxrtgNyD3dH4pGabsGAP9Y3IdcoBxY/wwa76zTxtYZSoTJdbQBdVLvrsj6Si
42vtimiWh17QozCmHxSsZoE7nukyIDSqUIu/UkOWm1Xo7Wbk/zC9M/rURvglrdaVVc0zRej8Bqk+
ZvB28/b8LPMI2EitSz6q1jrmyoXrfoxpBdS6qL1sS/ErUYeszpqruB96fuR4oN+DzaZD3vyqbO4e
kYhqUl6bmVAhUy5bbl+adercKSaBQe5vfCWWOA5qEvd2CyqjmsCyGl2JPyZnDOjsHMBOIjbDq//2
pYcqyoBF6JY1C22vgLpmKpRf2/TEUJU3dbSmseWL1BMLlKufrF8CnbyRU8k5zAlxcveF1FLoxGlg
DCXFcqTIGA7vFz3kPzkxei6WFGbmPQuz2PAtV2XWdrYvX6AtaBrLj/dKNQbM9nHQqQ236IchRn6d
a8S4eFQrKiKnkQp0rrTGLeJQWGzs98IGtwzEiE+8uarESuM+yvoEhZApY2fyBuxnlpZ/CADatEXV
vYcHSDPY9o7z75rHOUNnnT5NI3KinXe/WvLN26M5TLEk5WzQHkBc8enMla7323IkE0B7jy8/+NH0
arHFAzdc/e65T4U+eLzsMFXqPRIrl3u6DUkwUlDVeEPVE+nDPgKntJsD7gHstsNHNKCjzxQISoLy
wT5iuhPQotc96hHO5zyGkfYh13pO/aYd5uFXri2TRtNZBc/x/emo5rOoaxeTd8Oms8fQOptbxKOh
gmhZVXuyIO1Ow725epRWhNTsYIrWEGzl2xynAG94T1ygQUyo/ocRHe6U6NxDaBOYhxlQS8FC+Q5T
5ng76/6zoIgPUz50+HCgFBRr4xWS+n5k5/8WRqa6rQzL5V/amEoCV/Dei8rOJsgqMYhTNxFgv26I
v/z7gvHs0G/T2iL2iGXCZc3Z//A23e9JAcSvEK7aw4n36PrYnC+EuyKJDak+5GU5iUO6EH07ExJd
G/g1BjMyd1awH+mmO9I41jI81FdfYxMFqszq8L0kAHSQhL3sn/f/prqIHJm3mOxrSSvAghwadjat
9K7WByHq5IflpLkYl6SmnmKDxb8Dp3Nv4KWL0EKhCFX0NTg3RZgajRus5UCuG7EnHgKZgJUA2hcI
zQWOMcFYlv1GtPz2iOZRvVQzeFz20Vvn/ombjMlAbo58eV6pXHG6uG4nXdIcxnz3yzuEfOZnv98e
Jz66p9OttrcyDYwJL73uJuevVbP9LZtrERVCiIE8aglK1cnh4+/uiateClsRVHwqQP71enPYvCg3
hrQ04AnuzrgWatEB1B5cMRL2mYXWvvAkvaPJUJqxpNWZepYfuFGRLaCj9wZ7azP2R6OC4/6a6OFZ
SkH0o6RvbPTT54zojP48UgHYIaisIFsGxpSyR5WOEsJqzZMMGsEAd4FMuiIU0b81Q4zPUAsYVbHI
MiHAh0JnbpqqbmyoMCNTRIjG2fXqrDIfMo4WLNqVIZZ7eUixW95Bb5DvTvTyOWvJd4Kl2ILWBW+c
SxVFAnsJ8jSb1KX8RoACCxe0M2R8Ucd46trymvODvT7ic/gyE2Okak+dFmSYxtXa/vlTsFgJZa77
oRDH9Ge/Vd5qGueFbb4gYGBJAYRhaYKkZyQZfk+EaTBCSqBRrdkeGoiCgIPFiTiWa7d62W4nmxkS
dPGLbpuycmtRZVeJ2O5MxBE5+xu9Efaz7LsdGekix5Sv2OXDoPjSwDdG5YWp9HiBycaolGQQh++I
IlzuJP0sJq7PSH4zmODQg/BdG12Fyk6/L2NNTRn6aYE3iSwGcWiYZbfLRwchn9cllt/JezUeS/0T
Y6cFZ7ouThLMN64H7Jbf5mHIpdQUoUSRug9hcRpCukHKZXSdpRiciAMu/WtM1MyTlXBKAlXnvpbB
iZFAhNtETlFD2D79Hh6esUoaMhjoEKRSJMJ1TXVSna1sYftyC1e3cqIdKx+xTkuAVvbWcpJbwDrc
x/xMVVXiIVF5+ZRqXRAWZVtNv+Tco44GEI4/B3gbjqwQN4RXb0tO28asDjQcwUAYbwLFqUiDEsoU
PcmM4ByJFNR4xNH/VpmmmqF/vK1L+nE3La1vSATf4H624LEhlxpvbk1lmMKLMcmYEW98EsO4Pfx7
vNN8TEtpSW8IbvRTn3Zu8pY84JXh+zHoKPdXmB/mhh/J0isXQ1qnRiZZgrQUzB1zqG9tLxalDN8o
Ttn6PpVHe/ohA+Q9aqT5QwAuorgblqleoA+a6UM6ZBy4U9Se85NRbttixl9CGHdLI0r0AVhcY/OQ
/735qQsYHoROqy6aOXiCYdatgRj3lcLcKrStEV/vDgvJJ1QtWmznZvp/V+BgbWizka3jrwyl6ATk
+8vLlx0TppWKlpT281QXfaUhD16nf6KMnmgyxZ5OEqPryhgrnYBPj7sFHKz5Kaxe+s08sYSVYwlz
2i6IcblV4IGbM1iqP/lUFn3dKqxYnhT0STem/74TUrHB/7jQg9riLKzc+c9D8zVZElahSSNiOruq
W29ToFLtRvso2B0id1eI4CRhHvFhLHMomOAruYTPL/bR5uQZHQsDXgUw5xJDI4KepU9Vo2fXG2ZB
ezxyK7LkkBX2C55xXzaLysmac0AIxmrdYssjivLbxfu41qQU7vYjc3RnY92hDbznvd1WDDbrIc26
7rkf5IpYYNb6FFdjyDHPAd+0DY/Ne9IuWHpRhbGo3xhWwJ6iw6lwXUkbbU83wlwazroiYaI+w5J4
DjcrG5l1/S83HzOfmGKRgEw1XHQJSrfw144VlHMIgQNfK6PA+2M+0KXRBdt8fJZ5mzHMPyClKrOS
hNeEOvXTXx1q1J3SZSl5tocuFBoK0xbM634R/T7pZC7SqrPTnl4Ne6bZAaVgOvw8mjh1yjqK+XBP
x7nxsdrEufnZUnEMwBAsPpISKrgYS8wvro8w/L30CUwSWF+rWCF4e2TdzTU5Z1nsdlrS2PyzzxXy
V/P6BLB8kBp1LdApZjQjMZCUx6XDesFVg9Qc81ODC1FeUz/kj3TDazAb1M70+qdA7wA1yAsa/qm1
4rY6XS41AGYaOpQahTBT/NS0r1+G1cbZ7dvrKlOxqkYpSSvJfNjc4V+ofuAZB5z3w4hUNs3thlJC
E9gNH6KCV1Na7dxdzihcTk40INr/d0KZW1bIa8vAdGqFW4S5D3h1f1jQRn8YChHJbuWtKWoB/akX
C5lOb1JUKQY5ufLvcTlsIjTcL0Ry+6OgWgk3/Gqi6LsduGhnQAhddQBEcsDP8M+PNH/te8lU/RXJ
Z16y19EtBJEnsylN1iCUKp4uwErgeNebYcKEJus3enLtxeSJox2y7H3m5tyablA3Sx+9k1FCvSrN
iOp7G6vEkqhp0QdM2kP3B9H3UTswZHdcUmaVcB3xDCRPeVatI4rK67QeCw/xbDW0T6QIgGhSSi1E
Bm/thjljxf00dBsyvbOc6YKHGQ6rZiF665bsV7WNcdvG7q4rwge26GFn3Vlmydz/R9Q/G5Lw+6IA
/kFvsp9hzVussYIEbjcpP6+In7+Dv4NteaMfSmsSkuP9wd4xcRRYhquodImO1/ogplxLVZSaUXHH
hkqX5MnRPHXBcwEprZmZFgkB+hJ4wcj9EHudHcF/IQBiQ6FKW3JA1ueeKJOSgEj0EXOc3hHaIMh2
E/praltNcyUH+UKanCHZoTKMM52H3m8NJ12sIW/VOa2H+BOMcHelpf5Crkgqgqmckf1Ko3MALLq1
qPWlYlwpQj775xLe9RaQLEPu8Fi47qoHr/D4eg5lkXbmRUp+d4qNHUTUN9v7mwXqYLqLdDSBbNvD
zZ+uFWGmerb2a3GcBvSB47k5V47ag2aDPip04uOWJEE9hWCUJHF5KxDBPEAgrCcvXQe3SYRrmbVZ
kAN7F9ldjmw6z0MD5WUY4nHkuICCXpQ4ns+iVrhhYIRfovx9UYK8ePg/jsdzkFtBxnQ0jNd9BZ78
XlApDDPlZEg57azItiGjZyG+pCBFS3RUxVWBZg7YauNeNCUK7EeBgZ7CLl3KQxePTVInn47HpI13
EXdLc6uwUh/46DY+pwSKiL8J4lf74mdxRPU341A5WFvaIxF/k9Dn/pwkCWJZbR5SX9wRsoMomJq2
oxUfFNy7XLAdvCNbC5Bo9BT29Dg37TfuLnWwPF4VsgPL3k0zYhXicq268adQfHk3RFEgBi1B2gHL
sRIi9zlatQYVaGoKKZu6W00L/fDCF7MDrzBgChnHAxjUkOgTOyxseIkeh6mXW0dV/b8eZVfEctb8
FanAHEFDImh3vKKi/NfgWKHpdSAEvm/FvLINGu20jHOAY4wtyalKQa7G3NP/qv9egIn9lrSFS/RN
lbwHLoNzd7y1oHf1zklMpl+2ffajUAMkmBaSmKhrK4XqB2MfNOxDnIlaEY+tq2eBLaUwb4RV+XeB
YHk2YG4EYzQqQg5lllfOCpPf0xkbyJYyNDCzL/O9pMyT2wa5HTOa2cXu0wWTDmlJ0Typv7s2dmU3
X5Smcq+hqBeyZMYznkBgDlVTkXqtzXfJ5vkgpBsZcv766nIPvkc32RWRn2YuyBbMcfb6/kPa6p0a
wfveMQbGCnzfRGcJgaqg9cAOOz0lPN6vLSmgD6xaIBDTgQ82fPMLJ2zdzIiG5bcm4YGOx04jtrf3
P1gGwc3qR9tpqUjet3Pa+aljVd398FaVQjtDgTG8YMzL2lCrg6DxVrSFkZKfS4JndHIaVSCZlCZd
R09g72l6P1x7EnuWBEpKqB+Mg4eBen5yGbLClYQRfvjAgedQGUpb/TZ6X3eeXJPgNPYddrPxtVGk
0ayBC014/X2epTkORSyjPiLDpM21MmuHId6ShMA4hQUXp08yBCzuIFOG/bap3ueAaKyhKnlqoqGp
VCJjx9zhp3+P+qo1dz2RARFJmTgYL5qY3maFtXp3GXgtWmXdVJ76nlHzq9ifHAdMISGq7UrsZDTi
/clfxCB0AWZUh050O2bgfx2vCmWRY0rwajnt/BLl2q1ZNXT/UtpZAPdt6jN/KPTvxpz9lokrPrQh
T1lpzzjY+eXucRsRXaNSruyVgFqZdEC48mnykHgdSSjjStujQgMwsH59hlGJaejuzuN3SyxuqDr/
TbnzdaTi47fFdsb0jRVYdFNwl6C9nNISkkjapZsH1rKfy7ESIS8tezy45K8kd2OZwJ8OSgicGxxZ
lkFECkYVBSGsDDtqNYf7vFREggkm5cNPd5ImxEZ9oQ4V4p9/EDGUqWU1MkcMkdEfWa8zSKqdm1dA
KMEfaCJq5PTY1aqhL8458n8ILD3nMR4lm2wbPbEFeBgXO7FUUutn6FT9WsWis3ySJrLPf4zx9Sth
xNXomdU+wlZeQeQ4yb+YfrftCD2QwJBhxk3/OTW6z3CWpYOSbFI6G7WV+qiQvSUg4icmaImq3oYV
EKG504PJ6awvLssf6YmiUknw0g75HItNShSpwqiyLjLVNY2cQBVKAW0YZ9Jm62ASmXAOyczJ1ir4
FondTD2BdDRyXpPGtSH6/3das9E7zyMVlhOkPC2TCCDs2dQ/AWfyCXm8cJMuHXyTcsdhsnXNi1ik
UPrRha+cTq8Qr4fHgagyfMDZmhwQhMRtggiLqCrtuofJgUTB8UiPw0VVRabM3U5r9GcroOYywF82
4Wi4rL6FVBQ+gAaD4o2YQwVjj/tIgFFCC6o5m/fgv74heQfkrCYjnnEU/YDOHArJJ1H7ZWnrzfUg
zW/GAEbTb0ePOsdGDXjpp6Box9l36d5rGsegSBMPSrHyu1I6CnwFZBSEqVaEoRg8Sb0jdNPYeQ8+
rvaLUjm9rkFDH5lKsQ4fAn2jgxRNiMyank4z44d22qU8O158dLFNefIaoEUNpbYLIqPUbWaHI/Vb
9f04gb4zfxNfcruIz0nkCw+JvP9kHxTkmLqP7+G8pPieZJ5CWvlpAvFDn7S1Rf6cX6s7Z1WvOS0d
ARq3jXc7A0jDt1dRQOJf4wKTIZtAP95zS2if94dP8/A8uh31C9p6H60h7FBGJA9H6g3dkDlz+iRz
zCV8uP1tymDSZN/LQYoXtiROca3/CbbNzh4j3TbwooE/QNgWlrhf2xldjcUNLQK53W5tbiPPxClc
3a6fjk7hsbxAD/WQwQ9XUPg9TE+KyQIFWdIkGNYR/UjKbWfK0ISG3d75bhdzBY+6U7tMwSBwIVAv
fKcf5gEP4S0koK9G4JLoLkhfMu+k0GO8MbcspiVfPvP4d3DEJFtclz6OtdRsG8JqfLKB2xN9AFhu
DLJDNEbYVYGB4FdI/LhXZyrKf5zmxzjxn3I2WApZzDu6iHqlBruC0OKDo6MIqO8NC/zbNHC3UuAh
DMrhV2R8N8XGL2aLrQQuBiwLFW6aIm8JyMM0JN08XYkHQDvu6ZAtETr0N8d7dqHiw7QA+bDI7Xz4
BUb4J21SGkJ7qHrLe8qD6bm3oyad/ss+iSA26lN5GBmd0fBISS8KnQrqq486m6fw6yyXWqR3DN1a
nJusobOCrGFnHGpTvTNnwm9HiYC+ib246tHZ2Y7xu7MyYdfTSij3vhvHlWlN3TMD2CU60fbTogca
T3c3Im8bSf9cyxb7kv73tp8uC/A8XvHU+e6OyO3vZQUUWCC26hahtOC4o8bE+hiHiOqiM8hZfIB8
eAEB+XN2JoFIV0KwJHcWt4fbNhKzu6bxELv/8kqdyf6Vgrr7W5U+Ms/UG95efEw+KMcmgjGp+3rM
d/PSZXY3f8l0oUnaKr3cEceMVu5a6yio3RGsFKLJL6inRdqDh6QwOKRLjIypt20l6ljD7Re1t7XA
1YhEwMjTEltzjbLMvP8GzXlBqWE2e4T5NvLWmEhZvmmZ5l+m789yE+wVPQdPkpV+bbW55YbUaNy6
cn4l4RKPZ4St3VEfICmeQ9nNYQSdk9HbmaxvhStBoB5BBeuleH0I+j7m1DTlQ0G8xsJuHqLL8JNN
ahJ8pfZKFznn99M9fMp7x68zgek0jxMdrgZwCBCwClKj7bLszXRBUYf2lXS8AxvPGCiZDqiwOhhm
4CSxzP6VAHxkQXtOnKYErCpasP5w+0igtPpm3luD+tvB3//EXmjEQJ5mtdqLZ6Kvfcytrc+r7vc7
Hm4z6XkHPZo0Psp8d75WPDohaB5pp4CoK8mV8ckAoVijvJTQM76q80tCFtM4uxj65WRSIy4jS+UW
iVQukDfkSIAVDRPVhrQ0W4vNAJi/ihRO6iYcYViKyykJtN+C6fknvHemQkFNmj3rZm0dEQG30joD
fnOs4niNDH9dKnl/g0SI8mr6lAvIdgTtZmKSZKqgQnw2g9RFHJrOZxg+alTzIsQDRZuFlvuH6T/5
AzAdwdG/BXmspz9DvBsS/00odLaRTwagL5DShM2fd2zyGsROuc0y9GzTuLUtsHnsDXdwXxcNpw33
cUY/LpvSke4hG3zQoLAUevVjW5GAu+PvzOPXsL9b8t6cuRFU0sBt3gT2yw1MIeoJ3N7Jc7BfcJ3P
pYgHNpwsIhKLgYpoSeVg+/ahIwEHmqnMYTVdWHpSt6Jbr3IFI7KjhW4/yyn1VWq5LxFG1fOqtDBQ
eQ9pzee50EMJ9E1Y8Wajc5TrZOInttk8yF0rAHPXuTlc7uqESGGELtYnKe5B6kujC8790RSJ3QxD
NH44UrkMxSEVALF8ADez4ynu9hMKAE2gxKn5OWXPC6sDap+Ql7GQnVJhlScbcOfVx/Sm8Z/UB+T6
DM9f4aHaPqLZYK0I+Bah9JxULG4jR+5NKZYL2yv+xhvmtBhCaCn5HDuMIK5R9adFnkxoFAqMzAS5
Y35ys1H2+0W1TosytNcl3b4hhRbkVuMfXSgi1FJtQI9J2wJXjDfFvQUzKpDLt17GOeGUB+e8GXR+
0Bc8KO09R030M9Nh4CSJoTt49ts7ce36oKWvWLyJKbmQBErGhohiobEb7PgmBKmG7HnaELns1M6c
z8CQX8cpgxUDBEZtIQ0kr2tdDmZmd2lQVy6xFdUI5ZivtWnrRqF2IP5BYbpuQeC+rXCSfP9Mg/SF
TJAf0DelOBKx01AHPQgo6wN7hvaCY3RTdsBUTgLuz42xAjbjtnMjV3iBnnUeVh57AjnlqwQz9tU9
2j/bbStCKdnPw9RJBIUIrUGV0bWl7U0DAvO5GI0/wodlBgr35nPThblLQYIVUPsYU+8JuhpZZxai
1ntvPwQTh1FgzRYRL5D29+kfLZCW6SnA0cddTdTm0zP0BbmkXPsgAXvoUvWbO+JB9A+C/y7iK4sm
I+KmD87BXIV/M5pwYQrGt517d2INFoV1rHhWxxCmqpe7EAKsoETG/kNQwMNi1caYTxkHgDl0zVPv
gsGc877yglP77b4k1YtOKzHBaaqQPBKnMoFup9ZHqZZTIhgtXrtw1rbmrujdF6l5j6TRXgkmbSkz
6edDDQIBYfZYKl6MyBctz/vwtwtRzq6i1FHON1YCdy6R3JYiHjuhUclQl4AjwfGDH9k2HdBiwF3+
lQ+ny4E26Hjmt/bRdTQ6iKm2XN5RkN/nY8r6ygcSjQtcVqPUvU2vBnsXoc1dXJpjEFqApAYZlcUw
p117qzWPlgQ8zaq7oS5nkY6Dc/Krky0iGtnxvFLW9qAaW+m3Nb2b/Vowpn4CdBWeOs9pmCVxb07h
wxPi+rATtZSC6UBuyYBD6AZeuUf3++w2uLSD+b5zI7uxcO+fAAYUp2ZRYxo1GsIvOZ1U7//PlhIj
egDXqus7a4hSubjGemluf0CF7Kmc9BT6n2A70UbEn/jpuXsa8v0tkwC06r+LPCM1cFWgdvcWmwxc
kwfn384uDwFKS4hnBVzNy0RAp6s8kqqmSrJlhSOxv1OCoqusvjqiuvpg0KjA1iyAOTg/rSz2MOWO
/Jb60HdveZcYNPkovb+tGTjfqKqW6D8Veaosy+zytmSm90kK0eKjEMXgjVbiNNVBOvBXeNCQL+rx
xHEwYBynhLBe/q0q7ASKz62bw5YaY/peQce96tAOfI94XQfzoGbmXKrEk0c/VXEKTI+dTsDi7FYI
Y+ZwIOfKrEpuoAqfCxqzdYLSQfbzPQyKtannKghatMbhwcG329e3AHhGQDkDxBYq6Rmgp/g1OKC/
vNapDyMvOUCIN/XYzWxN/lQ979thzO3xdPf3n71hjMQQBZ1gEEkbS4/sLPBu7RHXwqgDNtuLjMg0
9RnFGC0Go7phVuP5I/BfZ0cRiJUA2f03rMh6sxBQmyA030GCkIqZAY2VfJNMnaWpWpD0tdOiBBxy
/LP5JKpqe1jYz3CDcqNuls9bHcC/hmBgvL2bPibeFUChLhIJkfo36DtFDsfGqlXOpXqyJglbw9aw
ftKroQnlJwxSl0JArACK8KdEJky+LFiftZd7ZLgymu5gQ/7BEIu8DovKpNFaLyRmkzCBMBeHb5uJ
G+vD9Kd9HYhweQuhPd/TeE1eUCjOsFAfgAuUVNinVLXaf9ac9ZSRM8+MUZWxRMyYHDluX0DxCBKc
A/Nbfg5iRCtFII1ltqpPnXyJOfJKIYP5RmF2n/y6JHdtcyO8qKPMmMr5CqZXEbx9zu1tPeLmCMHr
M5kdbNUuNijXlMz7BtIPFxw+ZZf7LOZ/LIkXNDnPlW4tPeDQbQo2U9t6dU0jpAQiTaiz+6NwN5NI
9883NBLMY4aTL8J1jjKjjPRIab6cV+PGCyU47XqCUAdAbZca8U3DPRTgBn1GkVPW54LwJjY4tf/p
YQ2Hh+oKzs29Hm6IMnpWzwkPY92XxZTbfiovjxyyu3funj3KhwGxIS74NHVa+cOsTQKSadymYuF/
vuX/yjoxpE0Dt1+eSqMEFvOoT9l9SL5/OqK6j/WJpjWDS3T8wm7lpAxWrJa9YKQRq93QbZCFvu2g
hZ+Q3cNrn+q7xMZJlLcpMOK8bfIZwVxoTvi+YOA65XOnnTsOK/iVlXoxUaZvoishIE8q3ouuRpPD
9LxMUKH76cl5YDnTPmAp7wdho5BAOH0X9E2CeDQqsxgqrk56kgcytAgG31BbzJC8ZxI1AoDEFANP
ubLZYcX2qu/dQOxrALxbORjYJoiQTsVCfgKmb2ly7Em742QW1u+EGcNfKA9nFcKzxiMmX1q08Qpp
7/UgcOH1S5j6kXicavkZExvJkOz8oLa9pkyCU7au5EzOgdinzX5XHoDkeyAD9AHRjoo52f6RE9cx
hL4Q2HLqQlX5NAVkTbiLzmhK4FlEk+lrMJkUxz7Phnm/nvpfIZbRyGB4Sq1OA1dV4TO5Dmfchb0O
xAO0QUyjKgsZkFc7HYI9YXbUXRc2R6uUkfp1WTWcaBMJ7AFg9w3es+6Qu0xp8Fq62rpIgbFHNItO
LXkYvSxlBI2bKiKOkd3vNCbhSkimX4Z9ealnEp2O3KNi1+FYOawYVcYh/DG5RV91R/KFa2PdqkO2
c1Ka7OS5r5TVDDKSsimVQUdrzLBRU5H01SeMb9aD3KbyaOtR1JXAPpJV59sAPIY5SUo92R2EnZPX
Zm+iypCu8L61wvSwl8M1yexWiZFcGYpY6rrFc1ecScfnaKq4O6MFEcqKaPl4gVetNtyTgD3Elyxw
9YuBaN44YREudxTRKsnn3mvCUQBjBaVz1V1+hux91MrMgAblmiKmERQ6R/dxXUCyhFfQRpdJq5Pa
akV4lQnnXe04KZdDhLlXY/4osVs6XhCxSk10BzqRyeC4nKKljhSLrs5U0zMT/ak16xOJLjsAx8/r
RiQWYboHrlacn4+s6M/j1Mo4Lf+r4Kjhyy1TZwQaKn+wKZgQ3snse9PXqU1WA5RBwDMyWqsaIKpC
ClsyuJcBOUu/5vUWJsHtIILN6tnN9zYcuBOp7kHEF01ILQ+P69gg3tG/fgQoceXPfSnJV+U6cEll
4yzuVL1EG3/XjUyqqvNvAT+7R0gYYhPq+TLELFSS1WLdkO0Uz57GhnnqfzxSszZ+t8fmCsWC+M1e
rizmbf+5d/L8a6IDyVQt+Onsp7ihcWCYm5Y5cjoOR4X11QOI9MomW3kt4ao8uAeXVBBVfbV2S8Lb
2TSCBdVJRJzZwIugMv/0H8ogt8R7TyAceRG4zSNqMoitF4+QarZT8a7tOFDbSRezKsUJPJWJ9DbZ
cviEVR6M62ARz9JgBZhTvQ43hC1hr9iShcMu2nItQrZWEg+8exwBNA20EBpbhEFcJJgmgqOuqbdu
BV06zruDKHo1glXuogGkZIWTUZT6L3fOpj8egOgpXbW5yi19Z3JrFQvRcRFN0l3GIgNwXR91Gycx
ysVC84ESOnuWBrTPz0Oj3j2ZP06WTWAe7rK/i7wOmotE+1l0ADA/F36eAKr34EUDOXq4LZ5tInBF
8BeyoLeGL4M2aETRUwU1Y8ohhiIX8939iP6aW7u4Qs9rlyUuJO6g8K4CY048SSkhXzOAirpgEBe7
K2vYm+pAZTHbCuFPVi1AelF1XITMJoavmTBhG3DLUEKfVB0iZgCOfVMWkiSU0M/ThZRIynM0JsS2
xf9Bjtvmxg7svckiaYgWoYq3Jj/bDT4jTHve1dy+HQfJ0FFGj7fkAyPWX9gwVgBbjeTo3ILEh0Bj
SYW6JtevEUmdMXZ5cFnYUUzA7oGpGbPCH8OS5CX2E7K9T2SNd72J5gaIWis1tyE3pWzhv447yvWi
FOE/PYbEpENoeBdzLSzdzR+2EB4oO1CXmZF9unsX0Ro6yJo2/qzrWr8J77FRXoklmvBpnoCQwB2f
XfDZSSGq5G5QAh41BPZktG4zFFNkcQhZ7jascmdNo4xvnuZgf30Tuo7Zl4gtykfHVlCJbBmhRBI+
IysdgUv+3hRy0x5myUvssqXPw87cI0WIfizxTS7XoR14Z6nDfNLMypF3FuUw+S31/fGr59fadphF
yIrEZ7VigrwN07XhsHZSU2/xfTK5Rl2N+PwLXgo1EpdI3mONflvvpMxVlyqY00KoUN390wXtSJxF
NXFilzSiJpaSczZTM4muSBuut+ne0CqKbZ3muQqCpl2EjhAnZ0Co9ll8oFQBGaVmCCUlcT6qfZL/
6mf9PeFqAk67tEGo+2PcXoHJ0QKJJYcPhgHW4e7ScCE7sv2iwokLhGvD1UNaGsSy2jKZ7zfQz4rQ
EFtiZiM4chlrD3sofhxG6WVyqbhKYj5xRUzJR8SvCe8LopPZ6hgY1P1+0OH4SVvCQh6j9FPngJW0
gxOliB55jI0nA8ebhvdDRdiSVQUGpHLIVmXcQzmSFSAG0eSIx1EEkAR0ytjQ7hZLIoCDspsVL5Id
tDY4YGP5CyjG2imHBcmZqyGxSmPQC1fExf6/iW6amdWXMAEudAqb43wDHOTcmexw8NBsbyjiA2XH
xRTSwq2ydATlry4+KmFSk644UL6UHd5zPUMnHnGslvx9bYgI6CgyZGa0bLjtfO6XFB1yegwNm1Yx
nMJ/oLe3EEAiVa0y7BEyWgmWnBzIWmmrmXvVS5EBd2q24C6MOO85XsduDEzcE6UgvNfbtqK4FA/Q
KGmJ88mNbk8rKVjKoC8mikbd/qXZbXApiqrpEHJDLqoOPy2wDt060FswA8gG5OfoQQO5fWh8L4qF
pR1tDnStPfa3vVe4b1Rys3uWZz4OYR0utAp9DDbnBvCDLWpAuXq9MszpXskW1mot+ganac6gKZpD
YAyKo+DJD/ufRgFSUG/aTRBzG4q8ucbG4ESvS5L520BhdIDcOHwTLwCMrMlPCapaRvIHnUouIhNN
UkJUXYUujo4AkDwc9+RghYMpo92iqqPolSj0tu7hoa/mi72tY82EY8RhADbQy56SvLngpl2xyLq6
YGCFARLsqyq35BbYzKpxKOCeIfaFtsq8xzgoWeG4Jp/h24bDiynYaObzoFgCuIE+f7L1gqxaQsBU
UWbRARY3xQZIswB2tvf+qExVAQsbNqXNH38EdSIbYPlpc/9kwKAA/A2BnI8TC9aPvm9sjgBkc/2D
hIwPH1biuotq7wwDOtN4wEaT/pPvvFoc8U2FBc+iyqYZkq0eZzS9OcFB94/VUkuHaLoyShQwAoSJ
/qMWijWj4rI11dzC3iIlyS5dclrIu9u1nyqG8eERMATTeIzFXglkZPh31j++qYf4W0eEbE9REezn
3ICmZ+3SHfO9+GX0wHNLmFits/fcCMUa0uUGlAhp9j/wXr8vi+mtdtYE+tGlFgki/42xHE6C9iSz
yMQUSPYY6k2C8EFeZ3aPAqDtidqn1Py8o+udAAvVzWEMLu7NTBgHYmQKZgbA2Sj781yVcrUWUfM5
p+iaT36srpQFPbG3PYv5lukjaGDG9ilS1dTr9IgTQXZwgg+p+Ib8kpcsqJNoIfuFmQEf+yHe+gVG
FZwi7nacj21Z6xZTR5ZBocK9dFWCTV5OjAcFjmiNFvAPIPyybLQeChMAz0/OkvfuexobAeyXQH45
9dJmHyr/ZlflNC5gvhFVRLBjkhTdxbi0Pw6e3neEM5nlyc/v/GUvNwXAQy2taHRB4uLz+o2oj93I
fDRipKqg4V5JqM19Ot2ORHkW8zAfRkwL9asGc+9hnhhdtuD7Uj1h8uKM9Da8BY2NqT3hhQX9bIKj
cnLjn5/9TXXkn0N3f4fPEUQ54gZ4Y6rtQv8z3M0kltbc1KWFruBnsIhy6MZiC6WAvOBvGIH7djl+
l2aGRQG9YnoaXQiJbk+vTRjzCfSZMl+9blfugaecuJ2Qgb7AdpR/CGcKAEi3NXAWoDgd9+Z9QIAX
8umqScKFalfrgOaP1cI85HdCZLoED0wx1vJuaQc6WE0oTyxHot1QwlqlEXWtwCMBBxV767BSArlp
J8bvXokZqQIslh7Td6upUfi53Jcc4WZozhi74Dk8WTCHNUOY65JJPqNQld+KP6EnfYtAQe4iNoCy
Qeo2DQZ4ID5bsGWQ6oI/nRWCGKwYiR+5FwxgtjDJe5G8UXq7ELj5f1wr2dUrZPLvr9VM8EUmSF7k
GrDM94mHmzDn0ojLZYznKToMF0NnSP242xcC7u87r49M/dHRr1bY7TQ0sOulNWbC7Hgtqrx/VVea
1WX3Wp5iAoXA9i8q9y0ZQ9QYlXZAbyKU5WIhZozFkzUDa1+KV4jyQgVc4RZppnHmM0Pe6h6/Vy77
6IUaARXxSBt53iKnG1vgPGQ4tsMOhjGJaknQL3QHfTHuS/jeYf51ka2GIkZENk8tosuRSd2kr/Jj
USR64ofJQI3R027fs7z2a4mInj5n+iFG9JuEi7TEvHXkNUxClPhDn2kcut+W6HCna034DsbJrc7A
Wkzt34m/2ws1J1+gdOzqOjGrc89zqeEO7PL66ITNcmaafJAC3ENsbiuRkil+4qGm31qSUksBFbCf
AGRF1ewjiuGwXv8UXT5jmUZuUj/CR7GclpUOfeWTaf7DopU4156cpJNBhlQ7Hr7NDm8HQqR+KpCU
amKgnmraUCGpsBXbmiD91GEuIXzg+eQZUYpA/DLUommQBYarlhZGr/Eif7poccUiGOv675FekpQW
KKJOkD9zLIoL7O2vxuaJoKOGhwDdYhsFJkiX8oYo1gFBDCDnwxj+A1gdw8M/OJ+oOwdSAg+rpxbu
eon+rSWs98hO66q3zn3rmRxhvYxaBIkUOadqzF9RHrfaKiKCrzYfJ2rv9MDCen3McgOt7Hgojoay
SbwVNyPlJ6ska/IXm/JI7jNUZZkn9gNoaWIOB9tfMrr5ZVhWQoPKYhIGG6+7mmf7/GXjHUmhcOhK
8OqNYY53fl4XUt55G4JJc4uIHDzx4f9elQzkDTvWmRhhhWEZ/4oQe3to7uUACGKIG1wWP3seFGmr
AgK7eCK3wJFcZRk4jko3pfscYVRR6+DScAT7yODUze6klbNyN/umGQmHO/CkSpX5ftgORL+OEUH8
gfVIAB2y6cVzzIodOZRRq9QqvEDVhzk4HhgaXOMoa3T84tAjn07VeENkDjQPYJorBMxEAS2k3G+8
ORukpWuFhhm/Ly39SMQwzTjPB5DUwCzj7jNDCN8dXKApY9TjPYymCwGtOwh7QY/A97Eg5C9lutD3
4SUIk8k8xbAAKJjtpZE0oGl6PLt7vB33pK8N/YN5CEYTskKhXN8fbFWKbQxjhkUNwGIw68t0SiAW
0sEhk+QohSjZi0v3wbfaLcdJqsRNfrqG+DXL1mI3an1ypsNjIsPq/ZNqD5PK8nfAMiBweVNGWCp2
sIuXp/q7pjKczrSk+xDx1sISgU+Jnp77/Lj0Y83DiJ7+7JoBcmTOjZF47ZKkCeVv8IL+T//Rcsap
i+T8OFkwmLSnQ9/QdSco5Y0vw1X1MQHy0Gogxkjy1sCg6q/OKnoLNJzKqNkngr/KnaTjf4xos42V
HYEm/nYy/AYeG5ELKnm2TAt/F0AHuHKE35v/SlaYgH91Fzs3CaXqg5nqQrbFntcrggxiq22qsvjS
mYkglpRcQ+OEUVvAJp74kzKf2Y4KpWgZZkdnjjKBA2tDb9Gbjp1XNQWSPA4FZVk1thHZ1es1BgUU
zGxT3v5rxd9sTCqGjZO30SnhjNoaXvDdWYbR6k6513Q4idWQKMXVVSsZC2R3BXxXxrFDo6AIC4Vb
P2ygYCQDFBDLVa/5mWoxZOHndD5nVfOQsC8184pQav41z4COcXJD9yvTkkHzPNMDsMaKwo7fCoNA
Lf3cMbBCirumI7+8IBOnywSKI/zn9GGAejQ5UmdXc9Mb4UlZjBsm3du3N/iNEXs6U/vLP+mzBd7h
bWtYvuRFJmbPYXjChDhn5jJn/QW9KFUCR+lyu9XKQVQ5zVS6Md/BmepocWIMEEizNu74TfPfzu4Z
WKcDN59MFu81IrSnY1NSpBZPgS9HqLxdrHFsf3axvH1SVvpl1FF/t5q/a9oxjrbeoe4e1gVdBXNz
2A9WY3gcyLYEBPvZexsxqqKJjweaieVWFBZGj34UknVkBKDvjZlfsU4A8oKrpcXUWPOtuK9cmPyt
Y72+EpxyrMZUhQX0fib0TZr289b1rVOagljIwkzdRSYxMBSNAZwaDU0nfxmt9cdOahqbL/+v9NkX
kNlkK0K4YyiD6q/0Zm2gMunTeydPongIEvKi+2OptOu4PbsPBgtm+GNBDSOYY6D2TSca0kNCGTa/
SLJ1hD2iciRYeYqoTOySLaJkvHUzQJvcDi8hLbLc9mc9qUtkrcN5vzdi+BkxgN9KYffy/Un4/x7r
bpKSXT/nLR2Y+kMocRsPuNG1PlgzzO1jQzXkvr1ConGmHxjLqHCCMGCT7S6ZPCNi/ay7DXWcnT3S
3+Otr8x/qFy/9/n9j0FldHEC7VUFWAwczbywqK+1itdleNngMQ3/2FllPmIuDxcEV1/M3Madwj2a
jU3cK6y0QsC1BwP3xgoGwWR8f1BjYIbqUv03uxHNsjnbWRNA8YzaGotyjT0fgxOHduZ80HD1FhcA
rntphq96DVWlTAMxMy3ttCKacG5KuXuYKNdzTJH8JtMI74artPQVhic7rgMMgNCLpPugo9fWKvkO
SgJP36XkWW5BuNE1DR62aS6fnAec8N/OhMz1H1ncqxjyXM0NqRV2FlDp8YwV1C+JRP7UGpC/myu0
zh4VfPnx6q9wPg96etiCclOtY8nTvxR/FGySJr4y+TFzYEfbZa/2fSX3FirVmegyZvcl9WtgjD6U
U7kx6l/zSzfs34NVQB9JcDDQkYPaZTeVW8plsJR+GEgwjx5FMei0VvOQJf3cK2ai9mMuy9Ynnwck
pwjmo9f1QOXIWgWQ1Hve3UD3MYHmTvLXeeDJqCN051RhtTaI7xlDCIgqeblXzUQ4uKe+HQHqEveV
WOnA5yM1pSAYYXES4vCSzfH6F3lEzzPVMRFwgcg1NiAEnYVGUCt3LiUhx4c1z5sA1ZPMq9cZNKqZ
ANcd1JRzJJvTXvAJtEWZ28/quXwWRTidwHmuXknCLzFCuqxICKPdvb+mqXxGX2c4ArsL8skMUBkN
C/TbaHBukvJZ9fTgzBiNruCBjkBtk6/nQdmNmPIMLDzkepujzHCmUZUBuDxWdv/Ws2zQDd+vPMYe
82F61EnSKoFmqGeinbDZ1DgPXnoMZxW7cUjEKsedhognYTBiINZ1MQ8M2yDblrIQ4pafg6ScmmxY
55od6U5PMF7NdUTCwyvpqgozc3kZMuGE7cTbHUaAFeX3Rki9Ef2gOKnBgM+ygz3ZhHxYo8PJ4jqi
8KasKyb5rxXwx0MI3NflkGFuWRYgGdXi/HWbz2BWaovkLDOhG4ApqyYDaYjxabAXVToQEheFHbyR
e1L25WuLK2iaO8q4uGIcjcEBmCnpw+qRo1EXkI4/JagVrz87eIQqNiY1eex2eoiN85g5ww/m9egP
DRwbEBO7+scc0DruVDfh7X26vGc2fGiovGsX09+uuGCitYF6kitxCdNy0bGctOMVRSdA63ofo3X4
uUWyKLiwva5lVux93W0hjFAmcFhUThPVjqY5Xwf4bGiWPyB/5CC9mwwebPY6NkaEbW9JT4XsiPtu
YRqcsqZIK5sl5r4ZqiS044DJNxCIqY9njOp8X7Run0fqX0pipL0SDXaeW3uvTNZH33X/eHDxBkkc
faRnl2Xg7up54kmctlfS3Q2B7lTEYHST2Zo/k97vB6tJJj7MpKDNJVqxJ5b9N8H9uhcC5e3Ln3ZV
xkS6YNlek2jPvaDr0FtdnbpmPrOs+Et33jN6uXbuNXgFyjIydKgAaE4DlIJ2lEtAknaTmIFu+5ma
neRSbj10wR/nwX/hpcFf1KOGeboPxqDejlrU1Upa4JsiM9FgFk8gh9e+e/SV4JHhl/quhVYROffw
QqBBUIBz/alh+eNl3LH6KjZhjHDS1Od2baNshwX5+36MloA54O7uoOHpSjcqRuwExQundNC3d5Ol
KKPZKxvdxOGoVlIeA60dRjwBsYSnNIuqgR0gsgfX+BMGDmWWlBUbwyz0T86HZuIYrwBDBjEStuJE
4I4NneUAvWJ/G8MQWfkfFDBHBKHgFOFNz0FpaArij51xgDdGi9LyfLPXPY/osGoax/IW3MEq1Tr4
J5h6Wga0P+VFXezeQAY+iSHrPqSd9LiHh2VT1p2kPrNata9pMH3g/DsZKZJVMephw28oa+TIFdvA
wpz/llsMNhQgY9y0kBq7Qow4VAQVCHf8jQ/9qzUmQBiqpEhPhk/EvfyIFsuy1KXUk0Zq20Lzjp0f
wwN1PX9/mnVmsKgISm7GimxSxxDQ3c5g5v/BSMna6VfBgI+dPp+e2j1KEptdYz/yfX4Pa1gZNSjq
x6Y472TVynjSXGgbQ+jAR8GIh+KJeY9rARLw0yVpDC6ZFhmJi1iGec7KfKhv7BDwlZVyZE8MlOWm
NMGsMVCGQsb/NHknCwozbQVAnXfm7bSk+KefWeOkhsUsClvilwgxeGJv6HcQpy2MlLypk+fpXzaz
iOcdVnWT6eleFJsveMwsmhjLmgYOTakdF+xleMXpB6lojlOavHIpenp4AqQVU66VxndAlQvWT2bU
uHL7ijn1/8+p2nm6LR0tUWaRyXdrl3ocA04D3AAvaytZSkwVHWfk8AV1UIjGW9QSxvz4lzJrLB5S
xK8CylPPYhSDYPi2BCyzfz/9o9vqhy9FC4qtY3Nv7Hy07wmKN3ZbIyg8RUGUvo/5FnYqqUyWQqAa
PIAY8Uym1m46FQyXeROQYNtbro0ImKOiq8JOpWFp67cvICC5pKRzV5wNXEFi4d/FHFPhIbqt/dQ8
oab45UWajN/5nfsXlG+I8ZK11CU/JRl3MfvhSrrfxMav6L3GuPuGc0bSDxmiaubs/D0JaKiOwQe2
/8P09GKcylxWVHTfZ1bJmQsG9BS624r3TA1DiWVgKJhomoHroyPQ2IjV1kBt1gAXVl72syKaTfaM
e8/uk4Ow3udKozXBhHj664XAsG1DWNBFp8ucc75BU3/2tby3mgUDX0pOTGfzYKFyM5zLXkvyuU92
b5zxaU83K+ZZrtpo4rBEheeI9BpVKIdT1kO3P+gEsFWRNO3Lp9aUIY+L9JF3zWQmoB24Y1a06O9N
zqVBWVKe+fYUhCP32FWvTsaYp4bfLQCAuv/hrPo0lozChBOTRnoW6M0LZMgJ9WNjimkA3sAXWuRR
L0r6wpR1prB9f3qSvUlzJAHNb/4dSvICzLoFcOcg/qdWAFnxhNFyDlSv7G7huVjwFDw4VKsTdlsN
PBh3L8iX7BC6/NXYC0xJFRYBj3WdbG5qRka1Yi8o4L21FFqwNr5CXCeUcpUlxXHC6h+mV3rBNBvF
9TcsKdt3XQY+YjTt4e0rlUKp8EKkrKhS8bf4e+q264P9HLFCstnrK4g3RaxetDW+PNqj2W7Cx4ah
48eVSv5pph0SW+7RjKuEkarY4k95TDudxrykUB+/gB426LF6qJuuwM4o1shlU732ddYEJg0QhIX3
33Z37C81+F1rC8pyCfhUKzQVDEBCo2o3xKP34BU1rRFABmUd9rpM7T3X+lApMePLThEWszupcUvf
euxYVMFhOWjijWnSeE39YrOv1/kJJJ8xn8l2ygKMnTvK3CM+6255NXcO0Yl/xASuA1PZRCQPHwNQ
dPLkx4Z8ryONewkg1cmCma3CsqOLQT5+t22Q6Q0QGH/MJB5VeStOAoyMwUj8ZPP6fed/cNWSNUdA
+9YZU1+H7KOQqrj2q8HV9dCVjGXeHqUHHpa8Tk2JMZIWrZurRGPPd3pj4ln+Dd95q9owmpUxQvo6
NHUvWmZnWB0iohbEBtKpk3yH3I+uGPXVlKjnaezpe616fcTmi9ctY1yXW8FgtxDL8EEzdyaAdB05
AprowTTkcV99htr8QZB8+ggDj2HuMX0Blz1uzX9Bu+ocwOm8e/YPMqEPeoj7ZKS/biMQG/DPPcBo
AgZvzeVPD5esVQYLpC0CrNM4k+E3eNGP1ntnWP5EUDj01cuUdjShjVbIheDSeaFIDcv+4MKcsKYT
deGEyC5nBGYYgbFCzZqk2qJiqvlb0CDdudSy0IEJHNsWbftu5JuzNhkLre6auZZTP3oBVjFY0Ohh
NkptTF5nVMVyCzFSulV4n3sR1MYzxrF6STc7o9n3pvpIL6GwJsYZJhU5khUY/AVflUUwStZpP76c
7wHQb2ZQfxfersT3gYUUIjHvzMY1PMVtPp8BtSyJte9gVwd4MOVGWBjgR5cBYW4e6hdjhaoReYoq
3p+MJsd8Lqqrt42SbawWUoEc6ikHpdHAgSu7/3GLjpsm1VVKpdDHLMHqjpLqJmyTPiscn2Y9c6RU
smO3rXOqflN+Tu1JQZdxmNWBcmmvNlakOMibzA6XFX7KQS5tIF513p7RHSUH+KL5vycHJ/f4oYoh
G7fS/p3h3WIZN1NBf5P6QpNGe/i7ctds36KYUhx6xPgqjdA4E9Njr1C7SIzvboGWuyCfMR/JCcEX
DC48qJ9D2XMbR7TqN3P2G5Rg2+4S/UFYUHN6CDMlESOI0nZU3QtUTClUpWSRj00LKSRKXh5VG8Hc
Rs8wiFQFj82hNm2dPSQ8iw9cG9zyzOGB9X7edUKE+BnsrFbBLVlBf8fmHxwh6bRtrRQRz/IPfVBN
Ocw6AZrLTljwWO/ikXwem7cph5B2rRZhWrRKIzsFhSSFlB4rKYmlHWxy6jOjNSUKQDEgCa/vx5yb
E3c7y7uirs4N1qNE7f0IsewuMrQmyW2HA7pE1a6BBKGJIJBm745qfSGtvRCS75IsIJbLQuCIlhBg
t4p9I7O9Ax9KNXIYxts3arvCCTN1+vLt+INVpiIf6Q4+OWM5M0rNIuYfKZPuahX6vVXu3Q3G265h
VS2IRKYURE0ByBrQj7lEhG9xNBYyrVnPEptAjw2Z1DQihr8k63wP3ojzA+Bbq+z3GW0GoRH4Oca1
wwctGLfb1MbGXqm/aONNZFKdrouLU9z/akDJiqL1N4E5xhuVxfaHREFCLLSaBV5ZFaRJKA/b49Mj
hYDU/UHNkoUXU/28e2vci4sjbRDldy0Y0dud+TdHm46/5VbRDhUTYQVEGMRHq6JyuQzwjQ8auH9H
rramn1RUzNdHfD7TH5eX1YmtYIEG6c8x9r2F5XUW0aHDUFFnhGTWUZG3cczCiEWgV4Gv5Rz0F5Gc
qBE8zARSevXDvbjt56N7FW6jWq0kl8yVqM6oaEoihGbvX0q5uQdBYEIgGu+Dc/tyBg7yiwgrN5wr
g603RIsYnIIF8KU8A1MM9E0DD0+O+qSOX+GaWVJPstMUA7tMSQBjeCZpCCTyC07BvQ80GvpDeRO6
P44b5C2JdewQPleYJqg2beSmWbXAwBGd3Y6SPOqVWuqffzi62NFtQLiKIqzeC1Q3R72tTpRcqx+h
PPp0ak9RTu4J1VDmMrJQPkfNJvSjNhVtAN+PLqvEFk7vyO1hmS/ErOG0tJ5VD2nGiN1et8Q3YUZO
YjY5+Q37oz18habiC4LaULkKSHIYwF+OgmHr8DGx4rYjyG+yBOnx1r/bLWbZPZQU9SnDINYJNEep
9XV6LCawO/P4gkv0irSFlL1/SWBNzgV/u+3FLDX80oJ0xcrOxDNovjL+CtWm+8ecqU5paUfzHG6W
ciQ7K65YalH9/4qZZ6oB+/boGckdiBwFBKSuYt8dwygGa6QKlrNosuC60kyLcGcrHquUJaeTbiHW
bB6I7nzeiSb6eGW/99O91dHh58rTy9ITxr3zfvOknKA8RkomlkbiGUAyuduPa9SmxRQ4pfm6rs9W
2ESAIw77GGLRk/KJncyEIcyZ1q94lcvr0ZGHnJw3FwZ7pXwyS1Y3E/PK9tOhJtECqUVa5wfnDqoJ
+JPqtfPSjTarSF5eOicJU2G6SmzuNqF9vCvLS/29O6sLv2wMuGAnMBSL+IHnbWTWexdBMXZc1NjS
nYctC2GEeQe4w2UST786ZmsFAj6aooXvngJzlt0Ym8xqWnCMBsjrQFt2jcGVoxmnZPs8OZ3GUosI
OY0THBvhA6ginulmH4hYY0xeLkaPwZg4t4wnjMhncOZ60vGBAU09P+cFVoM26uWD16t+wdrrVCkJ
4nEhVXZYmWB476jrQCHGDg9VX85LCPxa1g4yV8tqULlWeDnKnl/Jja7XXQMO1Chz8ulkfGD7LGbU
k8lguhgUK18wWzsH54rg/viDokAJHkyRaqBv13+Gg9TfydOF90DqBQPKxRF/CvrCAcAmvUuvbw8a
yU9NWC8MJgpH3Ba8ium2Zg8bGMPTaRMhwcf5f1UkCSb69f7I/qrOJPX6TbegNEOatREyfiueNa6u
VRDmKzux74Ygj+ni0fAIjuRi0K1TLRVE4iKsNrGBTRG1LbiXQZe2GzsP9HkaOgX/llWQBOcQqOhv
4MT05ZRguUnNcWoU2USOcRSnR+vXFbZ351R/3MhBB2dCr5AevbDDLd0attTtj7oL+XNYIausjZI7
qgNm6k/sjN+NF6a6X4ZqquS1XTa6PjHb8SHb8jhdam1FmJKV978QQ5TCX1+MjNEeGGW40uUswNN6
LfQ6AV1yRCvppYnTRSH5b5ua08bRJ6M2QKCrkX0rhVk8BW597QR5PlIz4Hk2h/YlppjH2MJXmtpY
mffTns2Wi+O355+PD1szc8JijjJC/PlXzXHQ2DoT2I/7nAGfF3Secv2bZorh+nLUbrUiXmP6KvUu
3i1AKspvB1aA7jqWHd8w4cA3dAX7mEalV/FGS2GldF2nOKv8jsLMWb6lLXiDAAu/bobtyaePVIFT
fbxYO8lmR3UBlvmR4XW+tljqUZT29/ludwTQydqQNpsT9ab+Sotw1pE5H5ObfvMJr62rtgnICFY3
VYHI1NrPf3GPOu4J6G/uxC+fK/xNzV7eu4H7A1D3NRtC7W3vxRbdw/tATjZJF4/WLfamkXyFVgSj
tHmvH+le8s4rvLvMZhGnlc9iiw5etdDDTRi8O5VkR4nASLAT8jE5/dzS1U8pb2gBWteIz4rKvy+U
3waRvx2ELrz0/EOOjj2sICDu9h3kyecWE83SYULLvzMR80XvL4w7pnVmtPPbpmByeaJr2axZqkxy
YoZg6wnQ00uURhxyx62Yv1uhZho+keBAaVrgxNLBgZyu3GA+HritdQ3vJirqxvTJU566+xcTJrTZ
F8QAVW0azL/Nh+hAZb6wGOTI04VovNq/MOlDTs4FZgF8CQH9Kcr5ns6cRWBapC8z3wLwS9qNMs2g
0SXZieRyV1CKDayBuLdFBsEFWyZVChyL3L8Vpmn8NO11e8tkfGUIhU6DcLp4bOLEUXzBTUSjdhqx
8lViMd4F6lfPLWB5DrwJNBf9BwOEHt5BLStMVwbliUeMVErBoxhP2wLktO/vRvo2JCwjxFVvQkKN
FhQf+VPlR+F8iXyIvz+Qda4x/lmM1RMs0C1uFz/vr9DCqV70ZubYbUf0N1+MRvJ3+OM9AM724thv
cnBLPrcjaTTTpJQgk7qEY31lJN9Fqtd/AaDziWVVAvyRaFdAQKgHdlODfSmA0+K2ZX4FJS9DxE7Q
Y5H3WN6m4/HWuprfs6km5TmqVwNuQLoYPjEXIodhclw8USwBG7sHZW0Fd2Y7MxtSlI+U/f48QFJj
4jWTzGBOVdjgmXg+1wZxErp+pxnd+WuVDge9v1kfOGBQNQWTxbM4TeFjXcLqSlxP/Fc8qxMZfJiU
YRlPkld+FVhigNucRnAGV5Fj3vSzp9cXpF/ZkuIR93sPf8VEnk4RZIWDpbBsGAldoRbIFSyMOEqy
EemuVCvrGMuqAi51FNVFFtr1zwzmOgL8ba0gPHp+NWOy8G1mFpRQUm0lKZ6EazfsUR4+L5/pVAP6
MIVvCGsBw16pYpVZ9/e12565jmCn9u+utDLvDWstLe8Ido1mzRXQwY7Wdp7H5TslGqwJ71nl44CD
uf6ah7l+zPu/Fl0TStBapELmtcbJyignV2VmvcR1su0/bg2iebCMEkefWDC3utIW25AaSPqYOGel
LCq/XijjVdp8aklSUTNy8LWjeRQNf3nSFSmkqZ4tqmsrtHV6IUtcFOUwPMNEKI+0jprXWwUzlM8d
hbbgdbaXBxTu7jRah04KNTyFZk1/Hd66uL3JLrQyegjCAIkP/FmWH2dgned6tYPXmNIikAPhbUf5
ONO7rrVB4xoc9OKwIZqz32g9cg17Maank8/CUChfc9YB31vSCcTytjYNgo4ah2ZHLE2vADEAwpVs
ssDdJIN9qA6iw9WF84WW9aCWR1pm7sgeM6DsywX/oIySvvRJWoX0K09bD1YHx3T1rimgJXtbo9zR
anBWiaj3FYuvzL/+Vzl32Z/xB75vTLhZBd//AMbyflCADUbbZLVDrLh0R5+IBq3AzGg0wD1h9iXg
rbOpudtMugsc6dn9kWSokk9cxyFpXWuwQ+t+97lXFLoZbtyCUMLLlvgNGQSE+J8H4XoqUhh4NVxi
JN1WkVFR+tdt71F+zAJwx6J01W40dP6oB1ZSiS9ugyMd+aZHEibgmVL4oz9O5uHmKh2ijU8L1WQR
YpXGIllIIrh/bTvRKrFYJmyLHg8T8FRiP24EQWToWUwnTuNRuFqeR315xkDK+MfuxA//fDFd9Jyx
PP61z6/0OmMIyX9SXROMPVBunwWBJq/ybIiigzmK7zvdMhQ1cVb1YinOv3fdgzP7s90wNA/Sifvc
e+oRq37uKZK4otzax4lszugfbDSXYKDyYqkTLwXnCkDCyzIEu1/INmq5uhmD+2S731pwyyQEcTRd
wlMZoLd0jlXeSMjku5+1OJqY/NItBox9wFC5mEaNv3TEchniN1eb5Va8bnEKHTNn//HHJasP6LuM
yucXuISf8EV50anQMhzPXaWF5rUUMOcaCLXTbRINQEqKjRSUzTDPvjU/IAcCDDH9IFUr17ItkUdu
fEY2Poy3fMi02jiSEIy/p7DFTeeLAwoaFrEcLV5qYki865cGdop3Z6DGqSNF+DC1B9kfxGkZIRDp
RG+TOWspjK7hhp62N0+UTLTANvHDm2P27bZOZTFILVvmGhmULbkGVMT7SgABUP0jWmwH1PpqiGXE
+Avs3y/8dM0ikqpXuHvk9lWPuSNAHGqSelyKDPsnGPop7UZ9ROIEsVFOD10tHVdzRBeYR1NRT63Q
8tXp+o3Hf7KMcI8JV7NsiM5JfcwPcYQ1N6Vi4As765SuooiM96h2IGm199orEfSE1d5gzKWeZGpS
ZzveCt6Y60ejjO0zlkBBozfNikpTRMt55JHpq7kGbb04zwRxzxqK9YEw+aKe082n+iqRGA5iTcdd
jFMF4Iue39pZiFXbhECnIIS1YvmDV5R4qlOM0Ep4MweP9YVi2Vl2gG+aHTvLptNUJSWARlo7CH0V
co5ehcIfSqtDCpG+PAmzyP/3kdXPDEjmLA+rs193O4gqf+H3SAs7UnC0HgcI5JLyTOK/6x3SkoRw
GShjOu+8SSHNer0U1V6TnWIJ/E0bR7OmQsHHd+IHw61z4K3yF9cg8fNJr0BebQCB/ZGbJprS3tai
dxZiPf7XI9wc+qtIAFQnUP46gI+hU7YfSrZJsmRnatPtSp/o+xTYuLY/m8l5g5N55HweIsSJSU3P
44jS8NYX1vDwyisojlq3lwIRgSkm+sBsxXrVeMDE2ceLCdSlGVdUrLNodlOr6kN0okUpK7Y2fNWy
IEOt+tOdezkOj2O3Q2XNBpXs/L0tf22ejYMs54rqN2sRBDBYKx0Oie3l7jrzo3i3MPy0Fl62t5c4
p1RgYczK5vB4f3PLrUPzhaSgaR4Dx8Rx1ZH9pffLFfLjsqRQ2hkijFZJbDOJ0/sC6okcl4dA+jt2
h9YbuTmREEc4wTleOygARe5TkRrURV+BWCLrpYS+vE0SDVNeUbFigWSk3aGC9VNm9xQmErG1ttWR
XXQB6KJobL/b3iW9U7Re3RYtBGpqUyotx7xxTjZkUcC9/JRJvS3V5FeOMk+5uYwm/Ltkk4qaclrJ
yrv/VvOIQIrSXnGokGv6cLvmSN07P4s40BLDCRD2sGgzpe0bhEcgNP8Kro/Ahj1AbKKDag5j8wfS
tS3muTYd3en3rFOyGYWHL9mzGuEiPK51T+s4NAxuZpaVj/lCZWcIVQzO1SLN7QMdFEVAnDpxT9E7
nCOfWBtWnyASCf2A61K3WyP7sfYX7DUgQ05nC1+qs7yMaD1VuVLtGztHvogRfJPmksNZ6tlsyFYf
4rTUfwYf+272EFMxUSdt4b6VfMn4PGhZhbTm0cFiF+zKxQXotjRGTu3HlJ9G4Z4SolN9Eqw62xfa
xL8f0pIZmSYkjKaI9c51bV9z0CLs+FF0k7wHtSXvKGuTf8fN5IvmHWqVwd5CerHlppgqGberF5ws
Z/1Iaa9RU/hBpqqdD2DT1PfVowNMMVQ99WZ1gtqVXc6CqdZ6ObfP4WmLK3ORh9rNTySfVGQijAXL
CJcSSYLIUQS15Id4Q4SFv3lbE+mx7F6gwZuxzJfJVvm6dYuqhVBFhMO0KszsjcXTQKaGVyywjjzN
Ie1/lDMXWHsp3xM+3ScMQ+UgpSOwwd6PeIsl2HtKVk8Ch2Z+d2HyUV1cRjbL7gFo8e6/G0HtChGZ
dD6SSYTmcAmN486u1A1u2Khx2x9GMhrs+znfoVPT91wcTI8Z+NH2Og5ch1Ym8Y6ytmOGiAIkl+TL
mP92SnPGERQgIbg2Ji2miavfkgvdjhcKQDqZRL5+GC7z+WBu61jpGWjJkdqTmq805xI1abwa4FjT
Okycs84c7RpwsF5dtSX7AYlPWMZvDK23eQIBDLAvF8QzXlkOkFeH3Aauiwn9crwG9WJRbi1I3H+D
ylVksXb/OyrLk9tVNo/TZgs/oPWbOpBTTMAn2gcNh5htspmibo4vPkyvmOteyxYKi8clbnu+VC5Q
dgrzq9Qkj5DjqWECX67Ur28TNXycz1MXAtX1d62AHkjmYXCX0HflZbIQpXxp/VkONOItEgK9jEMv
n066srq0gquXIpxgrfFdtnxdtF+l7sUeVYoIvUAnNR67vcpco1rjwRnzHXDsgr56EvM4wY0579vB
myaYnL0FcYc1Gj7msRYrASkSqJE6X1bNCa/c+gCOgi+WHVTRukIPnZvNlHiWkKEn3tVKcITEbVfO
SXpY0CeQg8xn3I6Obffand4VLA7Dl25e3OQfhTzOVie4xB/Gd9BCYim+mPYQz8bFkFivE0d4Y+sx
h20EdJ4FuJHEHzq9ZnKi+AqOiCFiT1VaNq64OOPsK2hZuCyJjzAMRlVYQyZmZdWtiGU3/eST090L
OYPYje6NAXO350ea7m0Qg4qQpOxZQwyU1grl5/JRJTdmDc1DTG1Rse1eFjH+Dun2agwR6Wkpk6e1
vD53D3x2ZoWBvwe7940IQac0v6fk+rdpVNac8PbBDGUs6ummvg1WzBcIqwGKRU+ofJWuJXs56//T
j/s1gJYgqCAQgcJMLZMP7wUEhJCJpEzFt2zZN7JvXAqTFcZETtKhMWKwcS1d+yE11BT0KSAnFDdS
KKg+gXZTkjM1ENYQUG1N2+HufW8LleUJ5GiS+kf3A42wYC0VgHSkPd9b0mngnjtGkKuOGnIzj22l
RC8zOwqAmoQ/A3AEb+NjYEIRMnpUv2kAMYSaD9ArmbzkffDYho/XeJbZH2X9Zj3qi1MrJKvLpji5
35tc7A4fngiDNIieQSCFgtv/tTkDgHGig1wSKv6pfZRs3KxqoZinhmN31SCcwMnMgHGPJoAfcz9u
ZtKzKYWzs9xCVtj8p9ja9LxenjrjMME/x1OtVHcfOqFn7BR0Cl6Cw6YRTK3Cjv10s4pk8CndNCsp
k/hAH3yS7kMxCsIcmhO7v6ZDSSjfw7yA/094VXvOQF4M4q0LJnvG9nGxm3yU8cyNNAt7R6hehAzy
gNv9zPlJgqnxbQfMrW6o5htNt+qMUpYDU/LxDzrJGKFyV6rsBDGAEr8AJynb8qxdNbENLunQYThs
P5brP4E+AvsqnsyZtAN9uWZiwj94T8esdIomg8AsAsp1VcQibK2Ok0ukWAZbnuvImgMdcy2F+ajr
TjYqm1mTIttcaNeh34iHcj1UNIYQaHEFcwzHQE9uffxbdVzyTExD9MqOCdjhRJ3ETlSQo5l4DI8z
0I08MaH0YfOJjT6S0lbULRC38OGFGffXMvWloSTp25oULUK6yaxz/wroTW0rFcYeQF95mSY6mOxr
AVopaFzt74WvwcRf4e5DXwWdlEBS54XC2CgCgHbMuPUvN7N/73OD6mID5Tn8BebBGcSqmmCQoDZE
FuKXB+w+oqG3wde+HbtE81CSnGazHsSCOaCwA223fRhMwZs+PbaFN8jAvB1TgpeOpcd4YdhqfKtD
aKRLYbbF1g4SDlH5Qlz/gp7YdNHqyNOSIB0eaJSI0DzX+rY41L8wQQYQ0TQAm+/f0Vfz1ozidnjB
vT5/cTaEnHj9l8BbfOMV7oL6DH9RAJD+VtXiz2PcFq23dldWxnPiXZ/RlSR0TXUFrbo3cogJJIRX
HzZgscwVcuYJgh4oHHzRXgcYpCEVsJGoaU5LyedRm2uvnEYcnnjF+L2vPR5a3oKitvXlWn8Zndyz
EI1vsLbD4DlMCDPKjRP7s5PPsEs+ulfGyF3jSSyOcUyiOUVHqfisOoLFgM8eDmt0+GLHnAVoOvPH
JDjtljn7q120/EjjG5LynaSKOWzahWMjVrr2ChoYXMg30TBGgClgPmM0pq0hoOxCGr83KIoI7vha
ISwQ8BIlevKK6ZzSdsKtMFQ67PP7F8yLfJagupLJCqrp2syWkVNRcpNSc9qNv3zuMFx41eZGynsj
RXRKW5Bd9qjH/nz6MBDk1snKpY1sw0zt9Md/aNqBryYcCtM4pIFPS4HGqnw3/VZ3qAgBXw60CB26
eGKwoP8/p7WNLecAp5BH4wOw14cXNuU8pvhu+Bu0TO5QfL+3VQDOI5OUwteyYVXJQCztICy0nP1s
rlMaD8Eowh4HzA+DXDAZC6T6xTueENbmdifZibWqw7IkotxPSjwRRrU7+qAyBxtiZikDyRebWTXi
BCuvexhoeqKTY2ookJttOWGCIgrsWcqAZ4nQs4S+qoyA5wmN7Hl4Pd3vpB0PosDQk0EMVoB6rXDk
n3y3DDESqmlNsAyT8Kx82voh/acHqc5NlBp10fBi1CU2dQP+MnG0fbkuzsyBu+DjbIs6ROj6Xvk9
4TpxYV21zggQS++MBEzmkF4ap4Bl//7m3VAHyaMxZRInimySi169mvfVwynK+YvYFm9oRh4FhMIG
+G3uTnPlF6j8wCDlHKsNuCbQXZUn8nK3s5gZHhcPRpYqgGLNVVimEb7kPc3Itw+puu3VsuvJ+oy5
u+g7bx5B/P4qQ5n0fFpsbULc0VQlbd0D78VsTVa24/I2yO9UlwawDyqipQ55reXhqAbn7fuFxC6a
ThfL1xpDkABNp0W+z1Su8eWTnSnUEofcaPHZKvOnoavNyAOgpKnG2bfGfmHPCdR2zussQjOAoUyW
gZQkG2feXxouj1Nngv/TSY+zG1hqG+43+dBj9eEUaxNbaLuIeFYYcxboMJan1/0uJvrDBgwmFaXy
OwC/UMY4bAli3K6O/zxHKzqqs0CzRJ1un7mQKeofPirqHFOlnhSU2LtBwHSUYQmBBztW7kq4UyjT
pg7mOZ6XqOfE/rP4L7AfLMsbOU64xChBM48/A39d7A+Q5C9jHyu35S71DS2cvXmFZFAvi/uVxMe0
zpACCM15MBn7FvxaVOh+VbFJzeUwQegN4H/bsGEJRCkkPWeaAt26pDFwOC2osnrTEQXlSCSp3rsW
hPznRTO0CVgk97HZoU62cHjswOegZoVBCnTIZocvhAz5mkbxcQ7ky26dGsQMjBnALfQhQDGVjTEE
fV9uDqfM11jvicyypgEzcRYhTkNfNlNbDD+GePHLG4h8bfu4PYy15KVGhIIjmfNtNmzvglgQw9QI
203fr1etJZhwlaAx2J8/NJMbMVgHn53a/fiu11eosltXOFSlWST8fRBP+fL8htF+DqD3RNd4dmBu
t8EcwtBihV62XJ1W72h+T91HLz0beiOTSYM4YQlzftq/vKwPxUHnoKCsXtK2atZ7GC/pqlnaAyFi
DZxW6C1K6lTZQBgB1f0yletxDU6/h02PpBAuRKqZOmsBoK4xKK3eDnobFLTJDHE8K2oehUZIDM5a
FpHyWcEUJ0gO1Wr9vO/XZFBa5mDGOatkhsLlkuwIEwQ0WgBAUhP42zKLAnRUMiiFLKvI7Heb2dtP
gZ5Ubpf2N6lqy1Vke8UE938Hji4kdWOi+2rEIeHpUEeYK9TDSRhp3vokroJZ8E5mDvlls1/EE51z
LsI2aqv+D5vLH+yOrYf0WocyDLDRig4a6g5aTqKV+T3vfFHoE+c//QkYuLF7Had8GLUB4Xi6kIU+
cR2kT3HGQIGfNg2Ul7NRiXu2ogZWMXR6g11QUUxJHetwV7jeDmxg9Anx6ujJGENZlhgUNallaWgG
JzPwwWW+qQA+ikm9nbPl8Vh9uVHBvFNURfxa/QgPLp2LPOQ4aaLwqzkC4619/OgVsjDMJ/cFAAnP
mZekYCsDppVDL3rcEwpMIDspDu85X+NqHsvFD/mxFqhUl02JwhQhZU6VJZlZOcwckJx2lQeIwLnU
2wqKoYQLLImgB/A6InXARgdesEWRT8pnn6PqlpGJQ6TBip1YyCppW+wf97N5/nmFEf94smb2yH6O
1Jzyio2LczAW8QHC0kz64Vd8tYvAUBbGpqAsk0sBDv7C/XV50dA2p018tleoo6pmKAJxPqxunzRJ
CgwoaqzHA2gfBKkRmWrdvNhmIlpaIFM540dSTvMpzipUWMA88GLd/XM16P8bWb5GbWekFRgKgcBG
WLOFwW3A7VirPzdKPQlOPehmK9oBtR/2v3P9HWlktssmvvUepIvqOT0V46HEOpQWUXD5+IeDO2jw
1gZVkUXk1llmZYwH92PMvfp24lI4cU34/xnkGad558o6oXELh8J6HFf+uPDdF1k5vg4I0kvD4S26
NuRPleYHaoA89dm6K26ovxT2cBFOkTt5VNJ+sr/yEUIAsCIRJb6XzEV+8LJyb4vyrRxcmqjKdhqU
oIdsJ69y4N5UHtrOZ6KqF1gBki5u2c5JARV4fJaH1G9/o+fCrMf015QMiyKO10strI+pbeGg0RXB
SnF3+cjmFbKwHBIh4RO6LNtQJ3il0jR5c0GWq5Pr9bDHOr0KSyo7EVD2F2pkrt3V5Ib0uxtspJV9
MTvL1chcl0sR+uIJh0zjh2yJt4OTpL8C+ewZQuERpqkIJUnw4VCxzneiJs8Asqnl8oBCmr0SLP4s
AVFB6j4prPfOZmzgs3kHvl8yj/dKyM15S4tISdb10KMUAdMEQffskL2HZfJ0CupLuFsCOnRO2moe
/n7R5kV2LQtMhwK7fjdLZOGaFlv7/A9Y/P49spxImYKnD1qExBSM1k2/h507YlgIhnEG19LNv+Y4
Aht1apXqXns/BFyHCR9qAG3ZuvPkUSuOQnjZ+wok8v8/T+fV6cz2OsaY3FXWC6Ce9krKPJmaqE8X
fiCyRh8V05PuOAKe1lhE93jzNNmGFybULdKA6DqzrvQgmuaBbpEFmpG1d2wPgjD5T/mf44//ITeA
gcmgjjXZdpHkjIWPKQn9O6J0pscklBCDbqcQJyWP/xEUqGJIW3Uh39Gms3asZupSfJEw6a/obN/7
8SavHuRuxWN0OC95onInAyt3rCa1k6K3U//kIOAl/GHQLY1rljnhOuszEm6LqtYUqzFVcjrseQ7S
inWrMNPIj2PR0mUOFrXmLYlH+NrPEj2Icd+dhaQMoQGGpltKCL0exgJly+L1pfnhTq2PMoXTLW9z
25zgI4W+Sex9OSnMj5NOtAoFriV1D4VaUXPthLzCnDiVm7AykixLH6ebE+ikUDprvNL9RQn8u4Ih
UyIuUbloSxSVFoR/Q3u/DmmxTAr2yp23gcq2vJRdenlprmce1D5FOwNbrpX3hiT8uAGR4VQO2vKJ
pKgam0vNidptauPS4aeDLWmSWUh5RzdhAUHhI1tinBe38OmKA98rkPL3K/O4SVCna4Vz9t6xzUkv
OEk+EiN1PdmmLqTNsAMQ3p6oC9CpBpUTXO0fK0nLPIma2fBOPJt8DICQ6S5w5A/Sz7unM7MfrO53
zHJGMXlzmC+P82j/Pvc126JB5Oy0B+bvytumvEBIhZ5PniknvioFh+EyJcWTWm1z3ebN0pUc1Haq
UnOv+UvADNmbgDpgRm38DJfEzVYbFWnRH2i66caO+al7HfJXIlHXE8YZn9M/5K54rVFbL80oPHFu
ylGXvvS1/DbI6YVnHVcOGvazHQjeiNmHd3J7hdtzbXI2azghePBfiiEGbmZBR/Z3lisv/DO23XOQ
XQL60LvVWrCi5vBJfhU+j5TV2Pmxzqj5prOe8mA7tB1pEZS0j/2mq/Cdu5GytLdcIVhvhk0v25rn
ainq8HTFs3RvzafDDJ+Av2NpmtZiTdozQqqMAXAWgBMC3Jm1mBGm9LEIJFOibNRHXqmCFP0dmoAE
DJ3cHnCvtcQ0Lsn8x4uDhlu80llizyLMP+eajJ9qG5QvuiwcC4/TusrPRubgnRLl2Ve5wVppEgU2
ZDlqtVoy3xXQe/Y9bNsp5/1TBTpJUyYAld9Q4hxspJi3o110Ut63Q+FF8y1vGujhFoQo9otsLY+l
Z0cTsYHdj4IWaCqFK1Vqnad6/PDjsyfA+JpY+nYmyY4S+8PnHZ0Md8TBfcP3G3MG+iRHRUJvpf8m
AzwlJgdRkLhHkcfZa86OWOQeMjlLXh/qpDQlxSjupladERdLh96IdiO/VfGxF+uW9wyMER93/Lot
NtSm6hgD98uz08IuY+rw2ukdq3Hnvf9LGZk4Q27sExWcu3+WOK9lX2SHVcSmAybf9ye+lBTGHpwN
Rv9VCgyF/vJcsWypBa1fFaeQ7BWn6e96QAcaINWmOSBp6ModnKX4sTdltMeDFrMq3QlxudswAiej
F549QVlsD4mV/0645+NnfH7gHvh9/4FqisIK6uln11pnxybYLmTbg7f1appy2RhBxMv4s05VqQni
Dr5GOwUGJS0HCMqZFRKsqGI6Xu8s++iswWk+Iqy1zD9IqU/6i21KVJlUCozDrZ8Gc/sGG4QoxOcC
uFz4A6XOuCruHrArLzqmhmLmufsPlbd+/zRBgsr4GPoY+VL6MYe30+PT1JEHGItzrky9t5i3YftH
WfYjMD31KDm657GGmRXB/hyYGfiQAQk/+CvCdu1y9u0MvmIlHkbUJDrXZxw0YSlMGfzBwfLe0qvf
cQ6GAocaG7MZZscEt5afwDz65mrGMBXxVPohGdb6hxW8lb8VFVDCRDur+0Hi4QypV2vzDLW5+Eue
EmIHuvAm1U5mSp2yJS0ID3ZdRAozkyZtryOsUcdTq667FUtFYD8/lnT+HxotnXAPlo2Ovt1zE+Jh
YtdeSpXomuhj9XbNQ94dWDlQP8fnzaQPpiw5xa6giMicw4DxQpVSDinjV6oxsZiBVJipiU9ehqLu
ATxzCK2IxYrk8FPVoxxlkPEbLTGw4gVZoYdOmor9Kv23S4xTlAcO318MIQ5E9aeleUbIkLuzH92R
ULa0OgDMkpj2rlCaRLJM+lvwgY8mLN8zcDVyEXXrtZM2HHIab5XPI9aY3/fajJ5lnxcbCY9e+djn
VO4dlxi8elnzyFe8bP9iyx+kUxD0W7DXMPkWeczTha/3FcPlJBr0A+QBUq1ZEk1vqfhttt5T7LnO
zaSRL73qXah6wbpdio8wzQYYU5TMBd64NlfFXw1v3pq9gwdqNv5rZNS3oLLATRz0q6g+ckj+hUKL
uxYCwBVSh2H0MlE/4+5ZuT1CHgIUvDCjRCkaI97ZBFZ3gufMC57tBJONSHBgDUUc3nLewROURpTR
zOvt1lAe0EwCPagsbvqcS+3je3GudMXkKMqwDGfpa5NfvV7kz9rEbErOv5vPZmTykDGHP7hh/ZQA
zVfB1S9Fz/m8kTZ9QKAxol9cOj05WvVOzibWiU127NvqRIUuUFeaBpbr8U82orAidusJZ8hjymtd
/dtYU4SmBZlE78HrAEj55QOYTfKqBPmQ+b3onMqow8Tuighq/RDIIEUl6k7TLt8qGwPRVg0YESk7
5n6LkbOn9+HhXLt8rXKspjUZntzRKvAzfpgWkTwHdk9g4pHJovkjmnT7a4OKDGPDCw8QiGPA87Xh
PTu4B82aEuN5MlQnaYMPaCKEHjFIF6XMPPuUwJuRgKW9w+lteqYTk8AlejA704c7ukAqQP/4gQfo
LvHBHo80eoAnB5/ajJ/+P9h+w4MfcKf1PbF3l4cXuC47Xc4ZMcDaXUDR1KaDGcxeYIS6YqKN9A4Z
2mnV89ZwkybLEqKcTxQ8oAIDW0MIzloI+St7t8lMrerpAomxGw1aO3TZE0oHrQ8IOyRdclEuDC6F
Xb3XNI+ONHPh+bGbJX8VLQ7hZqxf1Yd8pNm1r8pnagIru10QPahKBzsMBy+4CubrKXzfD+tYSB0F
dHL6xQpzusA7jZ3rU36kkPneJpxfewRqET/NEFIxFrlQChabtE36QgabIDhj9ckQ5p5yswuzOCBN
FIHVAW7JVKYSHhmrGnkXhlr8JjgaVpahEtmdnxYyqd90Vxtgw3cwFTJX6M8m73b/uMEQf7cBT12v
b57OKdKMn4Zc5EZ/9OkmALKr+gEtVV+o3MdMSkezFTlHSdNqjjF9i/7gzP2+x8LwGQkjnEq+IU54
/s6Kc/lpcEtm0bhhgmV+kaSjTUVDXxfwR3TxyBJwytd32iB/b1tNxgyjBs3nyz2WuPrvwgheMaob
eQJS8PNAAnDRPpBz3EbthPXv+sXvwfSbzIWfAInHYHjO93eAwRzb//joweLnYWDWAllMJrynVh3n
HmeiDoBETlHglirAM7CYFpjtv2CuIxTo8OjG7p2/OgoZPRQ4zoXZTUoq5hi55FrcFOleu3PK56Uh
8Dvj02pPG5b0G9t9LSgkUIL6aVsHmZNnlzhIbu7TdKY1gc2rqOTIEuw7qpeTCdLAtKTrVk0i0B3E
1QzRUEZ830qASYycp25qZ8IoxVQjYCF3Iy2bd2H3PmkvVMUbraIzth5v27LzDaFbogLYVYD4/ycU
pxA1NSS2OStuTd4clF/HMMpYLRCKu7Uk58fpNQ6Idu5yVbDYlOs1HEc9P2Xakyx7chjm2Nu/0yt4
AaVpkgxKzzgNKkALtDdq5oARdk3a+nOSalsDLDmkzAciLE8BHNKi8BL3MhxsC1azRdAtz2dOz3as
C0JPpFsPKWKSY+iyl6DHheSCB9NJ8oS4wIqdG5tndYqmOYDyX/dOvGyFCPm2Qw5i85Wh8Br9B7va
lCH8o+5wQEJ4GUhdFLmlpxGZCN8dTeNjMRnWscovnLH9ebLKKpbJHw0NNa1jZYfWVMpQBc+6yVV6
N8Ubqi7NHgSJQ5+0xP1EaFjHOFgyAJcJ4ZGH2YxSsbWiMBkeGTqd/74TsZWh8lwscIrmKTraooy1
+vC1lgtXRKnvKJ7GhNYdvH0pdvi6zUp4FKF2ibqvob1I1YLxzw03/mI+137gli70gTJObjd7oRPo
OTjPrvG7rTDh6W1SiqW7fgGowXqchdjAlBi5qKfUURyctAumy3DXXq/siUommLtldBIlpXsteuzl
q8yM+nLTsWkpF5aTh7lVl27nxUbng2/grLKb4cDpxAq3fPlEWmmkhAPbZWXCIcoVuOKZXVTa7ouk
Mi/D1ZlSCPCjvIZwbYj4YnE9RomWg9xhgo7CS7EXG2TDVFf16/Sctho2U05lOWRYM+1l3062BlCt
PnaSNc5+67+Nlvf/mysSNZ2xOyDU5Z4rbgXUsQRCAc00by/83+swXgzXquZe6q4FUmSwzbILyWBp
uL2iTjGe6WH5ricuukQcGPBQJaHQYLdPNRnceGvf5KN0HoSCdRM0MDMRXzxJf9tz/f8+Eo+MPRSI
NjjxkSwGtbx7Jl0fdVZNrG9VOnAN3CjLOBGQPwfqneKU0a+RH+kQmvxDH9rDWErm0AlIXA7I1Nrc
ilgH8F5huSuvaQkW5NS0SntiE05hIXnfOteZ6fRQ6V4wZx+hbnyaaIHISNZcgE7VN51PywTyoXUi
uVcE1JfsExEPwUNuQWdMezgIgQnrinrlTutUW9N5dV5g2xi/oEolmMAk4nAkIxxqo53cM/lj83i0
SoIjYhisTMztOBNXFiVqwLB7B3NOlf5SuTsD+OuFif40kborckQriGTcwQU5T2BDFoD/E50yYDcn
Zq5HtY8ZQsOV0DEk8/VbIEsIjqhoX1RRkF7nH9nrZNgkGkhh8bElmYk/zmNofXcqj6d7z/pim69V
RW/y4eTtOsE9lGWaY+d87VX6Sxuel8zcpWFLHjV1Yobz3pO4uid8Huyz0RDzWqRgIL6+lSLBQ234
HgoU+t6/ejtjJXUOA6v4VtxI8Wcj+trqqHu15rgAXKNvl2915tlehLvB0CbTTMUmU8ln5X3Uts0y
iBku7uvLEqA+g+ied5qmaQ1a1rtb5pjeCs4LI7NR4zHQcdfK7QawEWf8pgreFhbP+QfEOekz2xJX
XXeFl/RswwiUF6IpfKaCG/fruFDiG1VCIsYOFvadIBWWPVZkN1yPi/sz8M47EiIUYe9XBuNi4Jxr
WOkcilMHFwCJnpExVhr+gB2AS6g+MnGsrdvOAnQUho4io2uomIOoi1MMxKBMZaxCQbt/F+oNz7Ua
CjK4j00GWUw2FvSOu/NRwTNOwI/oL5azXYoN15c5VTxnAGWpzbP7hjZVdi76s1asUI95EziJGMfl
qpJbR1r+mcz7lX5fiQuiiOINVpklp7T+3vm6+yLNSaO1k5WOjZcyyn4PDtSRfL4cVcqcJQ4sIlB6
EqQtQ0YdchbY9yQCoPy8zwM9nXD0I+D6pLXgqLbbKdHTqLJJiEWsG2QYkshLfVotJ//QOVP211hv
YL82WS8n11D4jl5VZszxPzRRsFXzHI+IzCzUjYQgpSlS/wYK2DjUS7YuK9aZ4iaxJ63WkgVjRcRv
j1SVBip16z2KO6tGVFR9zr4yVm/9E0zJFaOTSsfb3vaLKWBv3yco3o5B0//ZCPtdvvRNobtFrylu
Gl9R0FGXjKsefcLUnf19lKVXpPWl9dW28UsfYoyLxuP5BpPWiXfAsx8say4lAPyfN8pZhsJNnuoz
Z3Jt0JoMcSK8TQ0ZOYTiI/FYH51XAYoPnDee8izmGqFjJNEuGjLSq7dIy4lV3yKc3HulJC4l5ubp
qgSaCcFz2FNaIZA62GTipVpGsRIRpJxKTq+muirKZAKfG4VIFKvc+l++TjZWtZ9PyFi+PtpYPiYu
PpzTyTWrRn0M6qeCKGiAABTB12Cei3fIXUy9EJ/V0Ay1Bopko1do/oyZg5U4JI7qSai7sgWzsYDx
riG/VGZ/7CJNOvL2oO/hfTWkbV1biGzvNskmkVfN36omw83O3tVaPlvD5TyXpJP5aUvrhzbCUvMU
mJkmMpxM8zKbHXtTvIfkrQ9SogK8+ZgDP2waTDzB4gphFrPivDct1Yi4wDwqv7sWkS+QeM1PJRiM
jfswO70ppZqqCA97hacgPWI3utqEYxsT+DbaCd4tLkeUTjrVxZtOz2g2Qv+YgPzJ3EKwaLD/50Yo
lJnXX+zqgDp0HfWxQEiF7dowTi5eajApG4RtJG4P8HQKZJXzDp+R21b+djD6E968aQMhTZ3hSikE
TShNIunIw4qzR7we88O9o1hcxny4b+eSMS0iBcYZ7EivX6ZTAzXJevqiMF1hcTQ5MvtqXNHaJwaM
Sza1bGoYCZq7UenVYYr5mkbpadZCPED9yajUmjBHgPj/W9NZNBilB0o50PDQ68gkHOvjU7buxtln
WxZLQYQTJOy0KEhb60GsDykYrL3hFvimzknhWzgtDdPdo9R7Ljx13pU6YAzkO2kVliJBa+FLL0dg
cVD/dZddgJ4YDY33xHvB3Iw2bruIid7LlP/GxxiweIdLHXcZ+2TFGnQGvTNb8S/EccMNO7+D0zth
xvFViQgUWbvN6YwxWa5YydRfftngLZg9b1S0vasEz0t9Yk1hJJH7K+Q1CbI8nFbRZkiBZgnGDzV/
kMmKA9aZAVE3iu8zJ9fO7SO+H2ExTvRI8RWtRk9qrJo56nXKQgbEezx5qXnh3PIKAvS3YrgcbR/h
2eeJWT22/yZFx3K72Eh81ESzdSy06qUjFppp93Q3X7j8ErXBwwPo59tXsjXZdqWzoCkCamBbcyz0
JGfOUbN1hPr4+aj6XEX6Q2hFu1GrwsLqLD2vOIVLV0j0YaYtT284mBBNtDCvDSk+KGp41801raSP
uTFS5152Txq9yhXRAziPDbDOsmTndiUnNqVR/5X4BpmwMd2wFVrL+ueJwnfC/6Fs5ND3pwkCwuJ7
eidy3PThnhljxE993uduNOIbkcsPJxbVjMcp7tjhut0PjuFE79TJRAdVebE5o2ycKjZstJVvtxX4
V+CihILfJj5KTkeqacMuK08wrsz/QpcmXjw0Z400SZoAMshbCgmz1XfALh1mad1n+hDF8a8qZUk1
s5NkMlVA7fJmPhwUew0kh4nV7VC2wGF08QEuqP0dBPJPXivi9UkPQ63er5F1tTiYzF7eKaZm9b6K
bi4RcmkYMM25n/kDOSbUDwTc19U=
`pragma protect end_protected


endmodule
