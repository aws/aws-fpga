`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
lcVCgLxPvCiZmApELxUHmOKgmgTW+f/y5aAxdy2VZ3E6BCBh2fiEv95VGXNJZRYjc8qcU2qESHmd
5g2l+ll5wB+W4zguUS1Exw339OQAl4JRx2pPWYEbLDCu6pvIqCqEHTvWsb2uglXQ+sOVfeDOG6Ta
wr0NoQu+kZwIwqRLfIRZCbe6cs4sTn2O9B8xwYAuY3KHTa+SLCzLzy25a0ax3uYDrBYAKMU7vFU2
7CgFaETklfCMc2Iom0yvrdGZ2HZgmIffPLH3wXJ0oGzpXHLcEmcZEVtHIaGN8IZaLrT4CFlrhuqa
1I0Ou02vuWOCvGCvmf9RtPYrA9XEpbEzDvrhYA==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
d86qNH6zuthTZ37fEyg+vQPGq5nmZTUzZi7btKBiZ30p7LxS4kQ5eWi+4SEJpPN5lCEPn3xtPUDp
Rws+vAbWR7geDZhaK1f8Z/7gH3Vk6MYWVmtkTACGG7X27RCiYPK09Onk1fsC4CS33yapwq8yFtPa
Wg5iv3XInC65ti4Qm5g=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
Qv0H3a+/qMbzHXO1s2pPx7A0ByfRYjISt+jTsmq6O91WKxLNnIK5+hDM/PCPbkTe125xuVj2jyUe
+WmdoSf7qBLDFIhquFuZFLx4sXDlh+B7A/LNF2DSCJ6bv+Drpl7kburGvdJQmGUMl4YalLzskiG6
8dQn4LRIK4Y1tVE2Wdw=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 35824)
`pragma protect data_block
qaE0LxXUQSYdG7420ZwfTwEocJPxq5/7Px0dtUCVx+IFRjdSzhB6RpeyMuygullyMyorlsOASCex
i/sY5luzlO6zIjqDmAIeKda9WirXodJzjpfYbBrJGJduq5/yKGb6zAqKlO8c8Pliv9lF4Aq+Qn01
3RZdUEbe+muCGSJ+KAWvMtgPIeyqujsdHgfY2u81XP2urswk3JS15qhHvT6N3A5YqDfBxocPSdbt
F0wrGRPnhwvojlyPAQO+MGW+sKhg5Jpzy7S0sSYSeLIJSvXJIcqvn1BByALY9hieQJZfxf/PAHJm
t76lMe15yIdFRcC66O9RAXlVhjuEtD+K/O3RHRoLYeF3su/FD19e14TFlFzWvlzaZAZTQ+SsOD1k
GgjTbBnBWH3ssGV4iYd5UGJDb0jxHYgZKUpqfkRkbfVpK9OCTlQliaMlDabgxkv8fznVxjOQiTFF
4saTSCHzWKp1O22kSLtFF4FvYivIYYwtCvAWvSoYT2JSXehfmbckMUP3G7MJy2ckUvf2PlDce6F6
aySjlcZ/w7Mkxs8cr2CHAslBqU4iMUUojjEmdpY0FUc17iB3jsRmFl3eK60QdZ4AoKTr0dEKMoSq
+6HZGa7HjzKhXqNhXu5J0SmOIXoZui+Hkl/gHJkZMzwLZddHPg1PDSDLG3qAv7lZ7F5wjEW5UFS5
BcisnWZO+ShvkVdWwnaGxeLD/yn4rOC8t6jMDAKZy6gTaECFEOkOtZSFT6y+10UATUmsURmCm5qA
SotvGBPvH6e3np1qv/ZHWy7VYgIb2txIX/GGXT41Z3vaNqFMQhdtXsdnZWlp47MIChb/mHl3RnF/
xh8WhgUzkjl3NtHAOyoL5ZbB7f2efEUAckGi3ekQtlV7tDcbqP4f+o84RORCqZ7rF/1yP60GtfDC
RrL0vRFOBUfTMAjupUUzLdt34EkIhHkvW6Ng0W2wPZhVayG7LaJJ9CPNWfeqqUTN8znr524J3kHi
EdVSDDV52NdPvnNyYTeMfFBeJECZEnnaHjU251iUyVajx1WP1cjReNhxoI7+iyKWvZKlfk0zkOY0
/RsT/sGYr5i/sNoHrlkMCu2AOZJBG+zlRYe7AzNq/1RfGq5IqiHFdW7kwucOxxQFYT+qyNXBoQoN
7bnoaVYPueOY8l4ZPReqcDT2T7JjMoKyoFYrNaiTayZvKJdHHobKGJFAZ2V6ycX17ywMEaL0czqy
LHMgKeJiRnzRe4pvbeYSwgr4LSgNX3qlC8sSYok78EREKvn29ZqwBd3UCqV7OL5wB2KnWiqt2ET/
Cfn+WLdpYiddI2fFLyemUV/tLp+u0TyNtrhViddpcl635ISwzc8G7LqLv0ArPd+e4PWrbgPyN5QE
S87B6k+ZdlP7yiBE59p2COxhUPiRxD6CrBKma+b53gsDLPwTj4qh+eMt2Y+kAuLjVJwcPzBVubvq
Mq1d7H9wi6bRhjfhjgzTg5DmECWyWJlKxqhM1/OLIbAsPbuUqvgMn/18mTtZyVJcPQ8e/qomQsZy
xzDXCZLm6gZEnrWrPP9qZRpRQ2PXhAdudPBrWDxGv3PIw4YBNW8SPVY+7YEFV2m0Ozh9jqDLxEqB
fyiFyQUCd+BXY16g2FifMCvu7EvrqzoDtT8Q0g1UmtIgT+jD2CrChDLGk9x2V5xkoyNREGmrpod/
8aGx4ZgbAe+7BtJQDflDlGHVawgAs7bhNg6/YP4j4ave8dUJvzXB/o7YWieUWqPd9cQc68/LHp1N
T2r/4ggpcN9IKwJqJubXBexKpIjBeCojoeuODObJjIk/hdXdt6IDLs+GoPcRHhiD21J4m59496w0
YBjBphUv5CETu5wgUwmQYJqjmY6DcMyRxYBFFfgmc8gy2Ivk7UnNglKsgTiGdBS2P95pXzkRklii
HRKRroIu04TBNqkOAznHS5mXZDKmYjSgMPEk0vqdyZM4aWGp4sVYrClcBnYsFkdKmg2SIndpe2iN
goLFZr+3Z3V1wtYpWTTROp0dddWWz/nM5edRvgg9gSFZRhLVijPt3fEMWDDUKefYPv5UR6uena4e
UfNm9NMYsLy7wtZ5M1iZEk/CuyRSoJBEB8luPuFislsPwl1Ohm0OfTw9FKHD7BM3a5BRLpWXk03b
HrxKQIMKXXYZxFIYQ0hd799oCNn2kbv2M94N4kkvo5MrsalM8vTiMn8QxCWfq0gMnKMza3W6GSgw
7jhaNvFAU9lzV5jtJYPiPv9Aq8mrQqOFelrRTdbSeLPKCZzTd+jf93fFAt2DrFTsCJrToggFwkyu
p0+bryqp8TgIl5Mfo0lvmR1iJLKSaF7kZmV4Y7JPw9m94LbS2HyhUe/SVwEe1eS9IaPJcdRU9Bc6
HXtcc9Tw6XQkCOzINLeUUuh4jNx7DRtRgC9JHv3hc2ztgxel8Lhh1SfJ0/vA+KVD9gmE2nFwdZuV
AEFW+SfygLxhWUD5MqAweSmZSBm8ka1BUobbiSkoE98znOfbE2cX396eYvCwfMCdTKAChh4K+YN6
lz9hXEzcWoA3yPLAPw7TleeJN/ZYYu/hoEFI9el2oXb7r0nRIzhxvtQw/xfo+U93j5Djvb4bdzBK
uuW6bDcl4o1fzCrK5wPAsLy+RPlv/dvvPu4ACsMZ/LCzMmyCb6d98VusmB9ogJnKI4O/yDMRGNLV
KZxnxoLftEChyKacAi3sUzFZL8RU+h9rsN3VBze93LbJNTkzLkaE/psuQ9U0PQ3FmQxhoKQCa8wO
ocTHPGfEX7dvCeSs9mpWHJNQAUw3bqBN3u1a7fz3SW0aq8frbsY0RqEmdyMQUU0177V6c8jMCYdZ
i0jZXKXxhhrNB957b0vcku4iVjWw8PtsWH8piFEfH+lyoExjA8BEu0F44BdUgSHxAsK5IC6eMIbA
QgOID09NYMlNbKF843fw91NAIdhfDE0qgGg2TyRv7PyUG/Z8wm3FTH8cAij6HG7FBPb03hLNT0r7
N+tXSHRFwaOtHtKjVNG5ER1jChsq1Bj0+Shqkkyxu95hpzWh9ORzB5IO7wzcCb6NjsLdBtVQ7XEQ
rQeDIL1QtCPLi4Rzg2MLeUw9emvuJtOJxDxgmLrDxpZlCxUbldQt0TwsY4kUx9bSAcxwRCmdTzVo
gedVNV2VOBz8ijWrdDIQes1d2i647Zu7ouZJdUMRuqg64KXxbb41BVSe9WAgRaVQziBiWr7LH1ZZ
rcPZXY11qBBwXN75V9njUe7lap9FDtm4jzFtwEi9LL4b1zTpKTkJf+u08ezeuvdsG/MBJAlO3x0C
/3hvkGSQUSFAezOGlT4maY2xRBLM8wSdL6XWKmw/Plr+GT2T2NGgZFJyvwhagsHtKXWp9edKimok
66zN22RcK3uoze9nDEWKfI87QsiRvHHrSPWI0TYqoQKQPWgXOSCD7wNOIp5JegJxyjGkgCrD3R6h
7qMqvGfRNnfYOWR3EPB3x0JvU60mcP0QcmYcO/iEJLeKf41PWTVYmzx2rT+CiihSiEvJq2dqFLeR
eEm8a6+R/R7C8Eaj2VcL8p9tMtxeCogdvZVv+f8E5zZhj5SR1EiAgv7GEBOifmEx/G8eKgx7vQpE
pHbhOH2ztXqhgjgBsdSdkFTG9sRIka1RGzNDfklnaY/jRPJhxlqkcs7uFFMF3CDNtMwMze/64knm
ErZ8xVEJ2s9mFeEwHIH2gTLeUACOI4bEuwgPkL7WD6sEIXqGOm0odLrFi2bSX/QuIB47QTTYVsU/
ADcVonLyp6NBea10EO/6aMv7DWiUnyHX1s3z4LU33xQpyPyGJrI2BpkSxp77NDCz1290fAteYkgA
0O7eIRkyJ58aUOdN2R1ENxhKuwwW0rmafYevaV8eotL3WEiLpcRXC/FvHX4/zYefxHx5hfHcMdC+
nJ2DnVeXCLDTYx20WsT2P/L5x0ismKN4vI7jDhn9fU+qpG6VQq+kZ7npsh1l2U6nYtiqbdurrCbF
c/wCCbjqSSUkcb5Ky6vw34Ce1cwzft7TI+PszPG2FfhgwQhN6S683rBv5HB36Ufd0zAkp8NP2di3
B4WUIT4ZSCgGGkvbNvaB3+m5V03DEiXAluxY5RwQy5kWUUApmvHdZKLUa94c0XGswn2OE4pqSMmX
SFB+Ai3VYSOdoBlklybiDKApOOUUFfGLHsFr4oEDj4Pre65T6rCYeMx1ShxNOw1MCplqd9LWNyev
pI0+UiyRFt6f/vAUlhqDK/GoxDXR3UmQd3RjQMZEI5hbEzoFuCQmxWKLxKj/bO/bJvfZVGBfQcVt
tgKfTz5rd6qb9P6F/Mh3doCsOy4rtnPLNLGqv0w8lpJrgSJQQ6JXcJ9pKGyX2uAAHtGatLzDhI0o
Pd3NLBM/i5OyoNvwHhtUQq5QBkd8T/KWEp0v2Wl4zfefbeDtkwRDkismdiKF5daXt0S2w86qhpx/
PeTDgz2dUQUU/nl+oQqI5OZq+s0a8asWD7lTrajQq3/fzoVC9csykEDWZiAB8RvKLK/yRAEJgJc5
jrhmGubUwMLafMi6+RdYQaWFCeqIL5SwFDaXrH//Qw/dSYStRvGOzsh5kX9ZOVaxp52eNAs0b6cQ
e3k2KkJ0Zt0wDsHwq62R+at6IPoDdgMuwIWeYG3MVdOsRFfk72XwkWl6shXoqYHJNa2AOibbSrGQ
lle0CAEgHE+nJCPLYxmvRTjWhjICO2wUlbWecpAmHyeA8WYkl9fOCUx0YlcCqgdgUGhvHRvsDCIT
uJYWX695stiTXFpSQ+WW1CgHDK/97MvKqvDXoDSZWwSlsh6gl3onmEwpklEXYDUtxJwBhQOqzF9C
+wu+ay63e9FD+1UkmBXUbB8NzInVMSDWwm211MbApVZA4s/1HGNwvXKYJA8QMpKNcZwxAGumVpFe
OWyWjM+pvi/M5RaEWaqZUiNrVfFCE7jNgWACe9G4R6sbXqCJj2DTROFo4ZXlu2EMr8/jPiC4Y44N
2iBBTA8EiTX/DC/ZP5tDB90FrfN8szLLptwQWLDNARwmyZr0S5+jwUBGkIZTLuNXsAJh/QuBtVCj
sAZdyqTh63t2VPLtSK+e5wI4U60s7dUc/lW9HCMaMRyDxRJ2jduTUpnWA5xtFKGKK+2XfVx0ZkDJ
aojA8kLTfqEs7xdpbarUHl5E0ueeEaSUHXEyh5PsrzLflKeVtcTiuuCH5OVBCRWE1e4rCSme3VNv
Taq+Y0+wbMEhu3B0F0ukELxjROrZmr9rXe/xaEBa4BNEDSjnh11vKOz+vt79lcB1bJkSHWwk3azv
lsZ6IfGVPj//RgSNHqzpzeHzufA1v6eQ+3dstt/NtbfwKcUupdrvDnrq3Z3QXELBMo/u3Oe38L4m
RyZ7mDe2z5+C+xlSZpnwehngkT2MfHsNDOTj2s6/WyKyBacmYoNs+n0Gtlvf0qhCRwsWY6F8FeAu
a17NsL3nFUA3Pei0QDQQKT2HQENRZMCEcpcgOmMopxwVqrUSacIhJPBl5gN3DQ9szM8Qh6a7uPEV
bX/cXheREuSaeq9AOYrVkusK88X+ta6dpjmOBzQXiDdrglO85Gcb9opLkBEib3BbDMgSyqCkfGI6
vfkoc3zxDJeg6qitZmbGG3z0j4v13mLtAdSnME/SXTP1+X8cneXjEq1Yqn9b3qjMSEyyq55bc9KM
XZ/+grbCEAoB5EK43uyb6S4CcojC9Bvmb6Brg7xWqaiPFdNzr2MqsB4s/jii+FiT24RZPI7iTChg
QKrmtgP7pjla5lONPCDv7iOmyChmPl0ZYbUXmaS1XGkpgti4E/18lRWpvn2fdsb5d5+1cXLTwxD7
bX/7ayRZVgH/gH6gII+B+LI25Dpx9rvya3akBqt2kQ/cnSGzHt2iZjQP7wEBiKIyo1q1rHs3e5HL
u4uOEHc+d8Sbhl8lxK3DU3J3VhaE//T40bmzNF2ZQ3Qu7/jDmw4hSQ6Pzr2maCrXp1ljHzVrliNE
8lgdMP3yAV2QVPLreKStjJlNsMDvHQ0Nn3RFOyu1AxB50cW8iSHZBz3C5h+tjZ1ciN/h449Ne4JA
BM9UOli5vHGF8Y3E5XGi3Qv8LI0CYbLYLaeV7rueBhELz+SamJ935mx6aR5ZBVmlkXx0xTuxtLF/
RoIDwdJTCQKGARaFRNDYQ+meR1GaE4fI4CoCQIqSiLmrSFCB+wfLbaxYO9HT27uR5erWHMg+GI89
VVuS84YIQPr4ocEXtOIZDfZaPbNFAXQ/aVc47GYbMqE7mnhTiWSGlyeT6PoVrTbKpIfyj4KhRnUN
fSoDNw+n7m8vWl3dYGY23r8q0l7y3jPy561mLsXCfcG7sJymBFnAUtEQ3Ky1LwXI/gtD7Ljvi9du
yrOhXJrAjgp39hHPVZ8XmULjbikCDW3aTVcx7QdIzn1b+oxdChlX3V6/Tpq8e6wYgHfGTBj08Hvq
SSHE3yKnkOwbEUtRP49bDt26tuYBqmfqrZFaDFVfbxuQH/6RRcgZIJgPn/l7lqHEOcDUQJxcvvsS
ghMS/OykkFiE7PJsNTO30ua4+NrmhaXYjgnHfmNXpjf0NIZkTnA/wRQgsGCvmM7q7RXXXmao2s6C
5tMIY3HGia6glE3i806QYz8KNQnRJiY7xe5+qDPArMmpYsLIRot0+EbTT6r2zh+0ync86pDnnUQf
6QHoDIosvvTCvR/RSKnsWDhlyC6h1d9O/yBHvGfGUOP80ZJtxG66v6oDqDh+oM7P9qWUZqxICpfr
MySz4rLtZ6+FoHNbs5HY/9x2oyjuaiCAF/J/u5+iYWs4ObeQCQ9UU1az3fNsQDRgYfOZk/s3D5o+
pZXd4NynpoQLb4vk2W1I4HDYulNwdcdLHV4sNDcKhBCSaaUUzFiDqi1fnYU8X/3ISQpGGbpfqrz0
3tWf6CPmupaMw1Go7656RPYHy+GZ4+rfdaIZhGNx8UZjjKnvvO49/AU0IHB5vL1yUQgRmeFgOhhu
d+qOHtKkwDhclUMPc0ArCD4FgnRl27JBM3U7T5DAeh1V5auzEqepbme0+XSgi3A5X9wrSBp0zMQM
N4Yb1kRBFlR+3z201Cn5/Xx0ZqKyeWG7rfzaBjZofrkLywxHnC4+8ASKve6tVegyb81MI+jiUbxS
lE1XE0vkpv9P4z9CZ0BYWBW+w4rax530+r2dnQam3MRK3xj5EI1/rXEj92j5JQskWtp/nL7Hk7nm
CYw+Rp8yFNFFc0m9gedqxpcHtXgJUdCX9dhCglFqjEb45a99L0gLDlvHNMtZlX+NL9UU6y4nTQDl
w6LwXUVgv1DCkvIWU8fU9jmF5gcF8XH8+UklRaMJFSlqhhQf2hgk7mymQ9JXvhNDnsb1iovCIWeE
Lab662v/jLr9nYfwnVyKsaLExg9rp01q8qffUlonNzdOHKN1Tzx+suEFubVARZ8IFfHtk7H1Ou0C
73pm97Q61JkrXDcDUvOr/V2+job+WDsuX4r8jWFzn3cLh5DjNjD8zqXh1Fh2SBvgW+Mispgat+L/
txeSk9YIDgR/2jKh1Lg0YaqOaiOQXs38nGe8BrdHtlQjem4s4Efwvo1imJy3fm7IzNczQuOPnwUN
pCVWmkgunBpKcLjb3Kw5dzyfACp3LS/UJ6/71d8rbi7aReb5R88Tu+6sS73yYpKsOSlE6x4qkmaP
/PaZi8lpHB9rug+pjstxn5oVOIp/+aBK/fe5NNW+n9Obd8W0cA5WMAPBNfPJUf76ERgqbZmnQSDq
Bs2CzLC5lK3pWL6rRjQp1EKh79Vfvsi434LQ5LzrEAPtru1mVZB6Nwe/LWCt9q2jRypAooFvTOSZ
KKl9hKFXOnaix0Rv0GlI5FtFbrm8i6jgtqruVa0/oGy93amBsX4TfirfKQU8cG6yuDUWxUegete2
KIeZHTPsKa7zBe3eTeEVcI3PXWPFIWfyDWvpniQXYKRawZ7rqjnUYXljPr7VGPBSpY0Apxme+cRw
ADqYiFNzGYqHcrwidIxX/rMzqNrrCgqozjuvaK1kPQvasHQusqYSVlfa4R9iDHV4E4CLve4C9x0p
c/elEd3g7a65k3ZhnAEP2ryu62osK8wTFeR4ZhZbnWrPwBI1xhJOUSbmzDNsB8Cm29TDJHmplNef
d7s4333AlkKhib/OS/AXlsrztw8ka1w4xRyVCt+oE2/WjN1nJoEdF8tqQhayM2mjPVMAl89ymWJX
gS6JGoY1VGcRNwq8XIee6/rT7UdRaA6dQr1YXG9FcnhqkeFb6764r09ZNJnbHioKjEx51p9rWUht
QuUgF3uyDBR8xv+t9Ext9FJnUa2tPcpVIdnv+dpZdBQZ2k521Zjl0WHeQ+/B3B7+9qF9NeDG9tp9
ZPcNg0x6SIAzwjOHGnwaqd4tbihEiLgm/qUwK54xSHexWK3/BmQqhmh02yO6JWn02SbrM72FAhcg
M869SG4hooGkT91oGwMFYPpQPqecyBBCCaWWwUHiMG45WU8NjuuvVaDI+kdCLKETmm9sT7z+8e4x
EDACv8cKix/FR6YkC9Hg/LX4Cs2B/7H3sCZvgfZ9gaQWts91YpEIcBWkcoJ1Q93pDo7bzXiJulYf
ivoG2R4zrQ2uj5ajJ5LgH7ZTZyXESLGfkhk5PV0qrO+BIp1/FVZEcaTDySs/NBWlOEtW5hklKrmN
h4FIo5ciDTRb9YfyW2FUWIc25Cd/G2HNLLK0xBelKL2h4DnFnfoXybcHtdbMdTtEt3Vu3AHM365i
MVCgQbl+XAJt3FsLtvInRIwQ6yU/adHSQ8E0dkMwWn8llHqqUqBBH/pY5796GbhIKrgp94o6q7Ak
zuZiXYPsy41dc2EMosxYeNJOVgp79SMjPhhSpzYszIN5awSzdD3fOlcTNtk/oBbqz466lG5i/1Q0
FCAGVdscatAXxBUGgvbieW95Yzi3x4t2yklGMOBsa4nGb+337JdRP575jjJ0ddRA1UQEVJNwyCQQ
eOSHvlJdN2Pkow++fT3SXVkBFYNKONNIJJ8cLXVlVvVzoqX+pJlFigsrl0MmEqz8SCNlyiR+RhcH
35H/3YpGlEMVeedO/CcYo8EUBDFdLt90QSfu8Uqo7uO73dv++W+16hJ2wFviz0Q8FHEvWWmnvbeb
+MfALudvVuu7EFjgs+LntOOxgSb1X1BGN0Z4MX/A+fDa2olV4sv/FG/2rFN+3Okm1OauDXwsVxhi
NFS7SnYhfB+Djmj2OiVK+RAe5dmsqhu7KOJyRsicpBCDIZ5ymYcWLPnLn2qge/bj1OZwzyjNYUQ7
DC43ef+ilmppIrE1a8K+ouZnv5+g6E1UkEe8/NPkidb4z3JwHFaYVkWjWNaZ3zSlKHkZnEWHRaz6
wP1Glu1gz2GSA+W90rgh58Cnb/zxQqWVMAYO4X2NKoOJOk/mIyKUHLJQe6XoQQZceNfeHPbF0Sa+
hwvJg4estSzVAmL6f2bI1pM/4e9QbSFrpI8r0eYO1w9CNC0DgTGG/FNBxLyP3EX0kreionNiFcdc
Ag/F7krd3p+DGmKo1wdJxHTAlZeFL+G1BwPT6E9ygH9Q+SGXpyS4JJtlFgf8xCJJ3ZljjsbBEtPs
0R75cnj3Q7n5+if2DUcdogSnTyT2+Wb2rZ3PFWAcQ6KIg31EmwLCFA8hs+a0Lj1B+D2Zyc+iQ7RU
ia7Cxb14k+Rx1KNfDcV8wg/m7+ZyzF+qQCxBrpa+ESADhF/z8j6zIW1EleJB+G9WiqGC5uaIDpM3
01GWw5vqbHX5/PbRCLDfajh44AJzb+Z3y1X1OHNccfacngyDIL3pvWmA6hJ0OsJE5OR/8FWmg9cC
QJZkS+j8AYGKs+p9ci73KxYwcsrHrHxQZxLm92Jx2KdOBb1OWabNuIXvEI88nXE9r5VYpGRD8Yzc
1VCiV6dLqXVqdrl9C3FmXVo0/7Sf7jPYO4udVQ3BcvNaQkyMHdfFlme3L95qWjsEiOMZPBIs5v0G
ho4jlqgl0L0FKRVTdgk3yPWqkgiKEmgE1XWderLlxCb5+2QpskgpZkjAjF1aQayHNELb7WteG996
1AU2vSVvoPIttLiDloaEbEurmNpIF0kbI0+mJ02cOcdFEkhUW6WQxOR7vEYX+gVWuX4TArjbF0m1
Ap935KJ/jLottbdonJGPymE46FQTCkRSyOSCeQJaCOT5YieM4RWQyzqbabXS23gBS7dVLIiQ9NcW
dmpH/j5ZJo6bny+qn+lBiKWERb9xrnGKm2ul5l4tdVu9DTklerLWEx6WujCyS1TJkluWZ5s2kK55
IBFHI6IyrQ77AQ9MHguAc0o59KqjRXH2kU4Uz9NnY55jB7LxYs1JWA0pZkPVa/gcjjnrrFJkywAq
89GS4bbd8pFMC65abA/BC53sieStVGV7dNgSNa3FGxtfnIqe4smjxY2MURVloxYZjEQiKblmt8Q+
0CepDPPSEJWx/7coEU+AsmyaIGWtp744YFpwoHYXVzd1KuXR+bFRe0E240Id1ezx97EhlzSzfLIE
8ue46d1zf4Qa2+oHEpUgtAF2Fle5RnkrZTseBFy2gHduU03Va1lCkRePrPMG31fTyS65Y6N2gaXN
iJtYs55bfS5iI5K4BHOK3OImUws9KPwcrdOTmsI9LaEuQNVqoKmT32qUYKBncamx/xs1ACAjjdwe
tfXkTNav6C0k9jkcf4b0VhdzL2Ci8Pf4di88TQjxM8YP63qPtTGay/rwzRE450EKb7dYeUJGQy5V
i5zyoV4bVlhJ3QW4UErnFEegkDAJZNs6nIwJQNYCju/nZbWnPy1/liWl/ARczHqMKBgcQK8+vAla
4FcwJW/3gClSlhT1jwrdXWUhJFX+77j30R3eh9hFjkClvvNWB7+5+G9/11cf7GCh3WeVTGX2nqfr
XRntzA6SrxS0Qsu+0E3nPkHLUITbw1CnmbRxto+48dwPCRzJ51Yz8q9Jc8MYkVsbpOySr8/RqQqq
H0P3qLOiGVCGRqOwNy2JOyH6OXwvCfaz0DG/fS6eWoy6i75x/8dGe9FbJEktKf0hm4PbjgC94R9V
eDqy4MGT6QTYpB2xkkyL8FfFL7aVOvmbVD4GOqKG0iRx2meolveNNEldwhs5I+3m09FDW186HdKT
rFPU0ggevU7F6o++ulZW2p8nrLdyIQyby8blJ+1uvn2wvlzB+xs+L6CuzywkKGBIB5SNbeeopjoj
vwmijPu4rUNgr0ZppMoJX2UZWVBoQhBbV+zBUqPxMhK2CnLdzuq1C/kR/tk8ENQuSo5CcV3w5KmK
62QrKzX/X9j4YgfTqua3FQJ2uIvoMIbddvPDzbiS4j8ndLBmWw7GXv/ERvBA8L2DTGZcqibheIGt
rJFqt2zlWVDeDR/Qf+MHcljVu3MKBMGjBNNszGSjGqyW9KnKaD9oU54BQxvf+kE/Uc4VLIbspUVH
URzX1vo7okVmQXImXRadJiFniTiQWJfdYqnUM+pyklB3qdTQHj39Wp3WAOr2SLAMrV7Rm6QLuwvq
plizxg6Nf+UJbKbRAZpU3dTBS8Caf2Vi3bqfPgMLbIaKCSkbCKRUd61yEZQNKNgy98eu9+s0CDTc
d3Jf1OYMQAHRyiWRZIP89gecHDgLzSpqiY3x+dPY0dRzH6mTocn2VeHIy/njqwNvSeIYOMaiqNPy
+pDuVtiBF4rkOGtShQL/EWioDNLO90LXXirlKIo9aPE2TMIOsfyDhIrIQiBLDkgrw1BWhytli8ZO
9pLmm2BngUqNI2jVjT66kfVJAmnkzRdKQqp5A+fdRY/X1WiHPrnzC9MVnO67411mcaCCPKZYffCu
W0BKwEe55YMMHnN0+HTZzkD4zP+g+N33k6toW+PoUz03MO0GkWLvUefAy00+q2PfbOiD+bhho0Nm
TZ5eSQVxHaSwRQILsmwgx5KPTUehWR3BhvC13p8GlY07ZWqK3IM1UVQ8B01gV8TZVL7bovKAN6LA
Phi1iHTIeljNYFyBAasygMkLc2u03VsM7daAQquXJGiV9WwxkBjxh5ziQf8ojMY/F74WoET9c17c
lMDKq0WZzUw23UjaMGCivcszEKQg7mGyEJLJRv256X6f+JWSIsm04fcvM4YM6i5JdNuurpTs6zMg
HNwYbSetQzp3nxpNKWihklwfgziYSO44sVvyYAJWqo6aL0QzMr9mUQlyj01EljMDZXnSMcot5Oxw
v1DwZoUmNkYULqOGFYGDKm5d+XoXGejP8gqPWURB6AVuxWt9lPG8as8B3PWmy7iJdgQvYz5h+DVv
VeptuYB4p18REBW8CV92k/5lXsg4qNaUwt2TRtqQz1gNT6Vu7YiB/B7dBlczRvUuRmsg3m37i6zI
GdtrrRQXm+RzBga/09M/M1hy9qgM9lyzSJ3wJkimRRn5t7jdVSaLdAOIJk1IMkg738LPRi6Yd92j
fVXDc+FoBNnKphbwA7PQf7tx9sTznQ47R9dmpueLiN+86C5Tg4/bXqw5LGo/DUAKwEFvTqXvjWEA
CTRORLnYVdqbhVD6o8Y8hIFH0GCrhHjYGrE1SLINB2ALLVds9jgE9+ze3+LqEPj6TXziGqxK6WRg
7cEpCEtkuFV5wqsQ8KgfzHWLRr8BYISCle/2HdwgBP4hkkM/l4X6Dt+Ts4qWyTNg9dgmv5ve3W0o
E5LXJYiNCNyCRGtF4Uu8a5IuxgA57iEuj6hkfOq/bIFIQXBIvjZxVcvGsWmGroyZh9zcPRtqFGsl
hoPmFl4MjJ8xohUNL1GXbFoc+vt5cwt8RqtsmzO2Nbdrx+PjHVqAxc8oo/7AcPYXhZGD18rQW9e+
Dd7Wv9VfmCk3HVCo1lm5Xw3OgjXQqzsjJ5vCzp5hbYUNvu4ZdIcOr8CYvGCFG+pcMRZdXafpO74c
Ucyi4nAsEOoxPaPWOCoZpE4zewQVWWZambma5OacRQVktCleGR97uGKef6LCnPsRAd4jsE7tJg/0
3iBF1MjdT1cAFO0se0HB2AL9ZFeyVgNg08WWkTmTjMx8LAl5ydb2n0zXaQ6NQrIFBfEqyh0HeOqt
5lq23SkQZHz9sLnfrDfSBI4DV/Y3cDJq0p2jyDq5xL9n+Pl2hAIbKEWQfNqQ/O2wHtfD8o1bcV/q
tZfgXzNTiaDUvMNoQhfuGghFMObcnz4a2jaAFLY+hCFNKO7GEMrs6hqjPwWokfDa0wfIzyMzM5IR
D9V3RSSrMPxe747U8DT7y5DbR4pFRTj7z+phlO5dPd04bplxAp/Lz5+huWhq2iQ70Fa8QTdKkGjR
mTj701NC1x2sWju9O25hN8RYJtvTsuCI53tBefmeL5FHs6WJbADn+1KNXxi0gk9xzigd+OhaqQJB
aEQmQQQKS7b0dJjlUOUmBowpWLx0PbqlagBq3FpxPNR6VkEO4c4PiSFFxGnsN6X75krviV8RBZJj
qzln1XWtJUqBvnhQXppz2aBOi4Y9NKJSz+yx0zpmvoiDwByJH0eTgYc9HrcT6rdQy4SZ7tQUwPku
pVS4fTUEL/eBe4nfQnfRTY7oVYl6lZkSCQqzIoD9rovqSHd4KeNsod+2s2x282CXOarxAaPDyERF
aBusLz8et0Vhkb51Co0YVJavbWYlPN78Y3AsNhPI1p/QuFLdUaKTcQHuyrlu3IOi1UmkBtBY3FKs
OD4N6JoNfUpv4n7KLzxwo21YWR5bbiECpoW6cT+pAyUmqAkr0GWgPyUwT/+0BwMfhLYAenMA5GNX
FsbDWv21IZRetci8Il3sNGzjGPsq1to7deDWCN2U3refr4aL69tEj15pTivaBl/SOUMRvU3W7TF1
shtB/f11VB/Aqnc7J3E2RbRFcqyzzQg4bvReuZswKA5SrgD78XMyvgYzFlIrWf5Tq8S6M9rodFVr
ojrZ41/8a292vmQ737GhbShYDZkQmm4DHworLccjrB22JRdAx++/kYTnVZiB1LLWVQM3aP8EZLFR
d82HZzZg1oaeDi57RrFQoVpoUTkVHYjc/FqfEb1LGbLsn0/y5X0GFtrufpz9oxLV63ihaOa5IWq3
XT0zta5Z3dxA5uvTJLw7w9wtwMLgPEhEg8fRhy5hOAmK121X6v9+Lb47inNJ68Cb1+/F0r2LICv2
a2qxWKO9pJ0pN+mIrRzbTFjCq22DdS0ohbQWlMdpOScydXbCaK+4av4tshotKWaIiAxrn02//se7
r1bumycFx6omjJPl9PQn59TyRGiIIRVGIHyZihcnanXL/tUad2bce8I2VSY4olDYmY0eNzXsq5S9
HFwnEJ0CsblOSrQsKiXr96RIAta5Mle3kLB/j6Gms4MCDFLc/z+XO3CwAzhp/92+8CCjPCyzOHPC
zxAJCPgQ57Lq0eTBG+78pddhIz/BKfO10TtvRYTncvfhETEgbi6qxQ3PZ4BAMp6gDUuuMUcHdwzD
95DC/B0gJ2WatSROtmY8yQcccu3ORrHrQdwnr9D7lPzBfITaDP8pU4batJBDq7b1HNVbhh38bGtV
1jboVtxXB2WkLsUL6GfKAnBd71zFOk4ghFnilifksEyXSLjuP0SGZ7GDa4tFA+MME90TIZtwIuhf
gCceZobiIrcDet2OYYiBXdtHnjHUOWjaEJUjJG8M4PG4633so/6H/iQ3JY0HTEOdzq4jupReqKin
yaBQmivtoTWJrG8vkqa9mbnodFSkdG0CNIUNPOaqx6BhSmm50omVCTxnXQAf79zcflkTsZElpZIp
npVj4R2M1FV77Lt/X85CWvh3dEBvEbktoC8vQI7BQZycJZPpI3Qte7MVG8eYkLBG6ESjnR3in63n
MCz5BSQR3OA5WnDxw7xrAZI/z6JYJCaTOotYcUPBClad2Soqa75J0EzpYaJqSrvzBpUg+qyu5Ns+
Wq8/uuol+3GgayOnHxfhYJPQYRlStUfTvbjfHGJG/T2XpJPz22fm1+RCRCRTueUX20L394nCPVT/
ge3H2nuMwmleRefjQG0pOW7Di+296nkpB8VNo44ztPj+NTUgZdTyuTmShe0H6qQ6edgJRJYsQkLZ
KIyspkwwqQxLQEeE49ddvnVcz2qkoNi9lTUjiEEXrk7A9v9iHj8ql//gjRyK2epxfBcMgoRYZADu
UwG9iJuXHiLq5Lu++QmZMQRD39ggt1Ep0LYfRbsGPize0M5kS3TckxD1mdt6tJNbeWaCeVbdb2ah
gFg/Kw2EJHCzpdhOk0K8FfOeo0JPsZfQrPmk2APF+eIe14oF4P3o4XIw5C9JUZY3n1YnAAyGVN1E
8gJUjIP0KZPYmIUhRtNF8EymmUvKJj42VxKIi2M+JhEdAimdmTNKWERUGGAdaWn+oV1P2XyKeJ9/
zvSbkGK3iEQEO7mo/4uvkzHBehmh8krl07znt9ITAT9K071W/xpMFrDQBRHnlG9KPL7i2WSE32Wo
DIiiwkXzclc6opcCjWgnDQRxQcd4dqamYlr9UpINudf2+XJWsIL/QkArnOdJvMzkF2viYHBsLc1+
BQTlAuw7kpdYDUMiCM6k72v3BUHLP5i50x6ZOt4xr/1Nhz6Nsv8tmlLXu7dSepXe6wd3GRJCg+M1
pvXcYFA4oHHM6XZErRYa3s/grdedkG142N+H8k8mXgL8YZqpGgBUPPcu9hhGLJA5fhceaQi9JegL
As9LzjBq088NH6EeSm/sRhBuSEm/ns2USKNBS4LFF0EPFs9XOmR/q7wnHiDRYD6/MLE334aKTDtO
zMslT8EyNHBiPt61z0EYmiOGt4DYTCNsiPoNpeDJFPI6K9fS0y+sIETh2yfeq424f+coMtuWYTUb
i3tgaO7xNr1Wws9nDqU094et3dxo9ZBN4zRkkpkFIDWNfXyly/5RprG2qAiYZTnKf6M3Wh5M9ud+
JKmJdLpg0eQcFP4eX43z5dgvFn4xVSqN05ZgY7Ohp+ZWYyzu0JOmlh+s/zHc+GH3Knohd5x0TLff
yS0h5gMYkBBMLhwjgyvF2MbHBP7m7Dgl/mHc33SmSF2RAsdTeJ3I4v0+ebk3EBL/jKsvYJcaoteE
bZzkSwOWECdzfMaQBbMRKRgG+hSNdIrx9cg9F5SbEfiq/IWJRuaOd2sKNBIgFFes25NXAnb9QOHH
GbJmq4qhrMQ4jHLteH+1SPHiHHmdQcPbQLDguLTKlYMPc8TLtNlYCS6A/QJGjXyw4r6HBTfrqce6
BwFJDltBwaqyIWfbOr5dtXTMPXCIPEUwK4AkqPn94RAz1T0AphnvMYhC+CVijjpkiIUKRybnV3JG
6F9Hung/u3+/OI42ScIBxqE1RZMR/MKHCY8R+YnvCBP40fAZ3UdFQYtOUWD897LHf4IdIi8nsEI9
hhzm8egoahxdgeK0xQzzr7HDb0uxskYcgKz8xoxeiqlr6LBUarID31UsWWx1k/mkC0PQg/8Y/bAe
eSeiN28pdGh4tGJPmGSl/P4xmyfKg6o9TmCkNEhnVBRW59yq2chg6ys2Ag3xK+/0cCA7omn49riC
90GMDT/B7eH157sXbrQd5SBvwW4oxtKEbhlo0U0RopQtsJX5cNpe9/7483ajYmCv/DOqysULY5ki
ZSFjyOhm065qKcwwtc4MicsEaM8mbl5UxLK8gVX/pbO60FvwfPBIGDprMCXDQUUeLtgfFh8DTNU8
8Oy+sJWBHy7NtN0+wIIl1wmaR9Xp23mV165cqjnFTMZjzTMguBvjVVLIC43qCL7IH19SLBzCV8zd
9nuLBwFOS9eiN65RGYNe777w1AHy3XN0LI9ZQgMYGr5PPWloTDH0IFG4vKcL+0n06cj2ETWEWhhR
Af05GyXf2V0tjvZLJzlwriP6zAEuBIJA335ripYFMSX6jLG+A2S44TqkrfpXpcDBx1RydLC7LzML
qPyHcxW3xBb0KTtGDaEJUV+FHsntJe+otwa8I4QDOPxTEC8hZhesFVgjWIEDt08dUreXRqfEllE6
XI3A7Pk4L9bjJiRJtxremsK6vQA7+Fvb3LrYrLxSdKxSI2Z05ygg9ju4mkC8QzLWxS/kvVpSrTdF
FodxkbZpE+SbML6zkMiJ1TJ3OXhw/oejMcB75KQSEUA2EIIEsVbnbUJwqU9Iao+AjFZ52Iw+c/k0
QPVVtS8jj2lVS/+49qEPB4/CV5Qx1rsH9DycahpvpzDw9/3ylO63lNKkXmcP7s4OyEjZU/6NiNy2
wVb0QKbklejTzxPp/wzCimp9RG4/84PU95qsLVNQgOO14lnqLkvzjn8NqiGWNpE9wDhBnF6Pdv7p
YY2EC1p57gVmMjPxdjNi1jYKLJVsVGLFDO48n/pAeGSuNAhP0GyziNn00jLvRh4youuXQk/nAYvN
4spF+K+tJULmp/ANEiSJZ3CMeJeu415yIVopJac2fXkccUl70HnnWCw4tmc6qPO6jzFeLGZaYzHR
N0+q0cU/K5gbffua0aWg/fuklyu5KWTj30zUzsjJ0aKnAn9o1c1QOD+wbn/M2Iv4/OCfdwRbcd4C
M9/zoKnVGlNTKW0PepeRg3SWoZv7cHG+NjER9zidzNumDBk7yKwwPoLIw2ebaIIExUcXRBwEdjyZ
S7ClS7xYsZczqjrDj+VuY1x8Phn9UoQyi6fTXGIxLd0LPJLSZuJL0Xl+bsiq1H9aurCLKwxFfR6K
DXu0RBxBail6HpG48KRRnr+IxR0/9B5bFgx22WixcA4U7/IstXykd+re79SIFF0vp5O85KGa3yMv
P2JrhNseOlqehPDeMExAzgE+eh+fbDR4tDH4FBJ+w3PkXvCql1sqIO84yIk1OEAdofy5mKKv0grM
QDx5VdzhIJOfCNg73vSDhHBrn7NMbUvEakTKTBvhg65xyCrdpUfaZN9lnAwgGZc4F5yqXkHaMrIi
IHieN7Qqm9QBPyh24aqDYb8VB1vaZNyVryPzmjhIfycsweYnsYQh26UeC2AoBqgTC/fxIuRsXZbl
RG7jTxglwQjEQTFCaOhKz/eL/oah9JIgqZFehW4BDg4DihepSO0mS6rA3SJ4sLN2l8h+MaCFqiNv
ie/lq/rVMSjyvrE0ncAbXuDf6YhzEGHvPd5zOxZjk08iXRbZ65yLNxZaFqy/xXeTnlxs9KckGX1M
vizBlq1K9SAhLZIoDX+9UpSG80X33PMbIKGGCn5Nml4HufAglD42um0gSdlVEGxwlUYH94nOxzcf
FQRtzxlzrVT59EtKY3hNV8/byrBYv3RpWw82qMqb28abd7qONEdwtcCem62Td7o6vSajIstR463w
R18/9k1h8b/puKgaUmVcEJgSyiR+OP8xnugKQfKvWeLwHxsRUwqntNYV9SXLXXsUOvc95Fe2EaCU
c3SBTSl9OILABAGPk4l1nyGLgliptG2gvUwNRvNUz6uqtGKdQ7KH8skLjmsm26CdahKKR00m33A/
Rq9uBbwRjTrB3aolGrnSMtE2AVukxN2FUbL6tXpIPsTFdO2J6fXN8eyrRATVYdTvltHKJqzniAMN
Q3bQXejkmukoz42OZFQFvLnX1r/dglCxKtzux9hHHcKYAsPD/m4oji8d/2f0TI2fM+P1DfuhTcsE
vUBJ6pKnxh/UmUu/WRPk+hnY9FpWgEQAsHFI1Wqx0Fy+GZR6m2I5rDaLdBy9w9Q1ByTp4GBlMV+X
6zd30VBlNWjvyyG3ny0BBN8ET84H1xh80PWVtZtRpRiBuV8dUy8GU7PXiZIpI/WnndYvCrbvavGy
Xc66FzLUzLGV8Tg6epITiL5+4GzTtSPdMCCf4WOBMuFgywXqt7WB0L/vJngmi9qbbv6RqeYoe/4M
Fx64ig834kq+ej/FdpjQ6k3F1g4lNCRw+upAAdmzKRTtbXEilQJPpjXksr7O589kCEAYe5XkvG++
hYRPqFHdO33Gg8XfnAc+TVDZVJYxFC7zcoV6P4sgvlR25zZQxpaZbC3SIV0TlHopBrF+ktBScrBq
W3c0jYY6UPF6R63Tu/qsRkoKYKyc1/zs8HDfwxxnuEPD0D3szlTnkZuckNVZkYroZKAbfLaIxi8a
RjmGP1EJKX2GI/LEXI2GZhoaGbou7Q8oCwnPqZJNDocZeZWkHdLiASswg3vvQYKk2c6FsaFrOORy
xaatsSdculz7j1XkS39LkBKKJstmZ/3o/c8D8iiz4+ShCPViB94CpuFPeVtD3MfgfoR5YKZvH+Z9
YTWUyz23WDr8MQVZoc0OSRUwUn9bgUH4xiIBZGZqdJJOMmhZVj33v9L8F+Ue6r7g3N68pQKF+n5Z
dIz04Ae9pGw1vUAg4htRr29qO8iiZHRYtP02x1A+4njWSbkL8+WC1mhVlk5d08GnWecb9Vhv7jUH
wEP4JJDRVpO3D1+SlYRGht3OcUmCqSvoyHakspwKbNLx/mYZXC+rZw7QTSp/yGvGQ08eHgyGvWUN
Uvqnc7lTCDHbmneG1CIz2eycQdu0rV7hkUcaSrhxbSQrrCVNwWtA7uqF/YHUINv6QY+4f+elYynS
2XQNKcmU4qLRfQSaNUN7+q8SRYxEzyE2zPTErc90KWHe0O9PuGB0G7vDnzEDUUENKvRArHHDNE26
cve8XAy+tON2+VV0ieGwqup+G0qp6iCIuqEmBEGlsUbjyM2shrYaN9XD4jSFg8Ktc58G61qJtSPe
3quXhl1qfA58NYac9O2wqIa7H6lCb2DjOWjk48TWefRCkgtcialUh9RJLPIV4ptEn7APt5DxCK4u
rExY6khymafnNqgVvccuPun+ijY9U9Md2vEpMVdc25rj2uz3Ts/W6GDnv4va4HJemL62Hfkq51dD
NfgmpfbwawFKeZ0NsieVWQlsRxWQ73WW7nWK40RSSFvW9pLWgWYejOcm9CRqjexcnNyDFIs/SnMe
GjKwfMlVECVLq7bTg8MhJ12sUrhEOzDuvqCGRymSW4K632yA0D6BVex4cWZEexHs3yAwRRr79Aru
74dEnymvpSYiE4qnZbmN4zA14Z+TXlRTfwnganoxQgLbpyDrRUVqUulF+DflqR7q0t2CbsaBYFxo
ffBSYpHBVIKtpUQRyUzsY7HLQt8vv1fwCnO5477IBfFyWP+vfAZan9lyfZyp6FXQUPZr9rjHczv4
stxKeMyycanuHeud3LwhZqyHup1dh/+tEg28CviC2gIzZUSSarlh/GHR7pzXXh9vo5b8ntRYpoE5
7SnFbgZt/SzkK3rlfGvPq9EaMIaQloYH5bScE2Ed8EeJcuaBR0tDzM6IF/keF0Z3Snho5M4jvag0
YkAjb5H0GHZcK4XAqg9xguvX6TsadM8L9Tjd0xBb6FazPy8xxMr4IifBQ3iYd41PjXckEXB77/fk
t8QJLWR6G6ip7Npg8z7ARzdvLw0m5q42MgngpH1iGp6K6Gu8jekU40Gc9P7BkNyRWK7+/uAA16M+
4rP9nakR5PLJsBiGmeU5rGvGACDd8EEodEMGAt6w1dWAdphKh1FrHYi8hlWoQHg91CBLcXMvMZ8o
ZEAJnckGAvg0WoikPVhO4UzqzdYJlIQYAaIF2Sx3dPxrXvFBX1ta4ZzU2R2G3iE1nKBqWCuLKcCv
s3b1KJzOvPy4VinEY6FGL8TnAOXkK3muIu988A9xDLe72oQzn9vIc5vqtGiPfl6Kb/wuytZRzJvF
vF96GdpiqP8LWnwNIYmKltcQuidB7QVawAnZNqN25U7oLv2vWKJAnFV9KlG6GOQ+FjNic7QIB90O
gSXAMQSvypIC0PFoqM4nimDWR0wJxfTY/eP/Wr6ZLhPh2xNISKPpr7JP9OtSyhIWRzp6CQSS3hjX
/5iadGxdAjDMMul9I1/EHaCxkMKBg7pgKpgfSC8XG1v6nrUw2PlN/5FB/jh3pfqewcBZiBI1Q8Of
gFIybzVuDoFGCEnYOa3gqwpjdCIokrOcIvXfSrzn1wWFlg94IssmGoKbHQD5B5SHcqZO3Kgejehb
ExeQVdpSm9kzjUysKs36CS1N+ZaB1unWqW3I2j16e1/c4uY4YxfBfSqOKYRw+1+IrBQxTlfhke06
KnPWJfjU38N0CuVTSRO2JZ/eTql9fxkNrdIUl1wYFOottYgditj/oOf0pI8+JvIRftWPKpxSEXQe
IofgAvo1VskjRPD60iCejM8tHaUQbq79xyYjVB0pECSSE/Gg5g2rv7F3DMGqqNiw4OsPaR/vtvEV
SZ6+ygUr4+i8n2tPn9Tid1/eon7fRD77XDN3Kjm2tomFKYzjGIHMvJEdi9yojNhBBuZ+3ZAklMKQ
5YAnnrrvVz1iL6EwQszdWHG7+76+SPUzgGIy13U66vgmZourbanjlaRA+w1H1MfpgdiX0yAB3445
qAW/aXl7CyDaL+bNQ9VkHDaGoTMNFa+uBWScqwV2lP5Cl/g5291zLApbzeGdLwSsqxholTdXjeXr
/pBJxCRDDiSmPqRHU7jRgU3Ypdr7PgHy+bQoJrLuMP/Gnc9TGATy4iiDiHiNW4UMiJMT3q93m9B+
CeVbbQvS9qaEU0LZTaJOX7AsgagT8FO+GIFff6IflSJE5lTsBT5jkYUEqFLOQrSBdZMznXCTL7xu
Wisl1tt288u9t/fkuUhiNz0Xdh0KnpKPmqkjqKAVZnydv2lxuWOEhKxfHRJNKcMuANrDD5s+KEAd
jz7A0HVjjsc0cgbp4XQuRfuA7zULq9b1a/yxQU078z5vHQLKOYpjsjO9x9Rl8Ih4A4hRqw1FUp4t
llRRYuDIAR8c3A1HxMdI0qZdpa9OhER4bllVWqazqPv3h55HwwUbtBOrfFIl5isf9C05RFMyBBxK
3YX5icUrM0r92RQf+V9ZB9zNrEhyhuyfZ9TM5r3SMNGhClE2urhswfZTy7cTtPtrDGnWuPw4+fb/
K5hho0DECUZQZeVBtS5nq5CQhKQ+0IV4/YYF1on2g3NIOK2UVrXY85WFlChZEDSA2vW3Z0M3vw8C
gldM0lUj2Jf8Q9hUJxASJ/cZv7DVVTwedlD0q+hLEH/twEHI3JEvg3pwMy0LLPrnHRL5x/lnsMwL
eHPD2ZyO5wKBCUP8kixkfGcS01soGHhJNwxaAixjSgCY7j/l/Fu/gb6814YPUdMKTStFQIJVJwE5
cpVbZSeAy5fNAs9rZGYkAvQ/pExqD7fCg0iy2BpZgAlq3pybLBTKUjnJmKdwPTW0c+iOWCmjsJmE
c6rTyUZguaD7/lMpDB38vqxfZ8covqeLhUQ/vecFGLjbKQQWXGMTJM13sqxSAtn2oIlBK5zqg8E7
TuU6smPUXlJ4TORfm8GWvWRey/M72IkykRrGdDzv/0IjUc7YbIozhxfVGfZ/19KBBZ2/kSSj9U5A
DBvCzVza+6/evUphJCJ72Sy1TMX37lXugovPnNMR1O5s1u+896JwkyPV92cQdHLDUwdOFOEKpqkn
HePYp2cc7WH4JMQzMvEtbbujSsNjaSplElkU6+ta7l6nx4OAxBH+q8S2qlEaGign4j6nIEL/1iap
h40RqvPDiKrHiisr+k4IqUPRi8SRmDpluRynSHBjBi58N4X03dBjpi5bKAvf8jGnuG8WhRNdS6bx
UMy9RqcQLPwFdn/5/iuS5ODjmzN80l2Js9PH2z2q9ey6gOnvIXBllHYCfV8newyIM95/jHOcbaUE
1gPZrYR16z52eLqkPitFsWcOjQsh8lvQ+nNbSmoji7g4xqTVDafuZz9MUQxD/Sz/sKZVQ5zxWeJP
56ps5reN9QpfikVuP4a7UKp585dYf4xqiJnIKUzIldlpFwFFxFAIFy9V6k2vzbEMimNmB8oAT3wK
27+1UigTxS54lYiqOcvyiKcDZVbTkhXkcn+uAPIST/APSJyiHKfjc/jr+lwGEpQY4SvmZCv4Kmw1
Ll18Z4x0dCJM2LrKNsixGW3mG7Kn9c7Efmr8oTooCduGrGHTYmmiNrDExQHS/RCsFaKtWGjE/PaQ
4Z0/G4n5AAA2jguv2sKdphC0xmGlnJPN2FXfxMsj/jQ2QYznvhs38/XVe43NDkgSI9i20jMuXEqO
zrdZx/xcGdncz2WatzC52psAOp92UVR/Jlfv3UqlOTKq9Fj8TSBOXX1Tk8w/HC9pOJj3gdt/1XmY
3AOfyKCMdvtDrVExSrmvwqn5VUDMdopEtvpRr9rbcyJ27g3yyvo13PFoZcHdivDiztNYTHE/CJt8
UBAXFSejVabAzZnHTCOmNwczsYi9M+uBI+0cmg3CWGf31SHeQIkL7cglfunRAAoEB3wJNHvV2Dzu
kO+OJuK5hxRNUSmtidKMrJtEC1YNE8cFPFICbOMm4jszcXnOB7hgSVe4ilUGhm4eHh/2AaadSMTk
9jC/WEkuELs5Dr9nNyekfZdr7Gl6hDoo3ELWsIzjfdk6xE31SXlf8Nu3J14AuHoB72qCjPMvECIY
98jR4GP9vAqN70jq/zjHAY+pPdziCHzUrJjHgc0Xow9DghPIqKJ6OdkKM3KRuxnreDJR9qnj+qC6
Vc4EgnATUz+E8YdrZuCX/mTYMC07aXY81eo87Xf9NdcVSoktnRwoqzM3+BNJ05Lx/LbmvEN7pxpc
PAVJUQzsYg6k4lerLxm2Iotk/yQD84f1h+6RT7OJJEpjXA4qQ2tSpc2i4gACKJNFCSY8N/Y3EyjF
1sjoV2uZ5gi3nYqGRLdpPt3/lvSWTDnvNpyGBndcmAbX15UBM6IgBRv1EQJBsuU3doxV45u8VLMY
7hGyp3gJ6drHuAXT80L4PrpSzXhqb+qYfcyL9AoGT03R+vo1YuIF9mJq9kPJF3/7CNIbI7ePLr+l
VQYTrXxU1ux33+bln9MNcfeOxVpF0lE52geTxlkgiqn+v/hoivEKvqAtFFg2X4PcsU0yvCWkEDdN
UKXnM8tO9Bm6ieYNyjoWp5fIYllH9+QZUI0QOo7wmhpQY22prwYLeUh6uDSZ06s/NqwG05iwO12z
LEMNhHQ5hUJ8m6OORXozaEz1VsPMbfBhqfblXFeOsKcbqA77qa3QwIfFP/XEF2ljkHTyZrsA8sJA
DbFZVWpCmAvp3xvzI8OjG4ZxjFVND7dfHj7m2m9QvEPplfEyXu0cuTIw26B8SGDmnS9f02xZuKwZ
/xRnmTkn/8hRck6V0Gau04GeW6JEJk2Jdu5WZ0bhrtQMsb8eV0Fk1uUD+YBbBsSLJupjsPfY0LPf
BKHHeCAZ9hSbdBd0DynHOBEWprcnGlxEKYx0Rpjkf0CtrtJOZZX/ZvnBwDaEGpZm6At4/bG1DKu2
a0yxx+quVoOSGmsmz5B8yhxypd2I2xl0+ii7ryTsprkOuexUExPl55SWe7CMD5+MrIBd7n1zru0J
kPnpX0/u/mFvRsvFvPlcvwopNBlkU5cbXRf6YmIoLtJNuygRDoN4Xl82Ghbvyr0nhC8ikuXIiEkf
Syn20uC+t/s8icfcIX9niH11m/kLpKbmxZqP0vg+GmXcefnGcNQ1XvTtWkbDBvQ9Lozk2C2io72m
sm5a1rRln2IyfMtnbGhYb2s9S8AshF8V1m1hunldH1Zjx+gmuvcXAazMF4BtCYUFAftcOd6Jjs/x
dl+rS2jf8TYhITuPk0L7bE7784BFY70VvyVK/FIRWDKe0S73ZNX1afMGzEK0exOIQg7ePc9FBtLT
Vde0QHA14CGVIs96hdIKO2pjQGoHwgflq9rAm7hmi/AQel2bF8nEFnGyjVrcblttdfBg1Ws17Xhh
5xpIA6IbC8et6A4TLzC6f+8/MmbUn9isLm+tPa2vxpbACTAHykkQlaLQY6wQoA7x+hehWDoxcZIa
ercJPVlANlUmKi4gbtc1ZImK3BSKE8afh+DD1sM9TYfQmmBcSmu1qlUODfK03TUKCnkstQCEXbqg
QlRBGppBos9TOML03Ea0PXny1QDkhDQ91C3mtBvev3DIKWmnG1eMX338pyqBNq6XVMCRfrWbz5cG
idhL7W1JBtnX23fH2UrDVU73ElD37MorM4D3Se+shfGKHZYZNLGkrhxClGU8NsuFN3mxbtUBG7/B
3hohlMSMFXOgj25BYl+dODQNoaCAwjWYekpSM+9eYB0Npxsa+XAZR4zsPptDCg5aQ6GLaScLQSmS
mdK9Dw6pHqwxJt5S4FjOB+GAUDVR1WJaU+9IciAsPCQfHc2Aagjj136jmq3uOsQqWN/fXtvyj9My
7uHe2cAn9xzRYeKcJhcP1pDpygGRzXNP41+uSKe5267g0dVouoW626FSENYuf11aHGHGBVSCL9BN
OBwoQkE8ugFQN+bd2BTnMnDeukjAQcbTAya3ezp8CZCb/xH7JLlJIPYIo7Ri/t7PXTae+7mn8c1N
0a36iWfJhE/SVU+yvkR/9SnnpbR0UA/sL3k9d7yCgHbb263DVtU9kXt8CQxjeOudsmLl5HR/RVak
MIUl/nehime13NKzvn9Dae7Ma9Y5rJgpIRzI7lZxfKMDUDq90kp29oEVG92huCCQo7Z5ddLxEI+M
Gg6rynbbmmDp+OklaaHFiMzWjiyxPv6OLithbp93KlWdCqWaFDno4cx3Reqfx9Uwn0XJzuydFid/
b+acXPfdNQhm5RHNkceonqE2lslgCH46n8ppTCjnK3s2xrZAGaSmVYTdcPczf7JperifkjbXvoEf
3KrhQeekphnHa5wwXyxpevaTViDqD/MbvBQ9M2t218HRwzCZbEWac5J3jtSQ+ggP6HhK0b+nRSk0
WPBz9vEY9HhiNpD2RIH9M+peWcZeR4HPfl0qIfH4Z54gxCapHLPNrJVgofrVMly/uWYe3saFPjDm
XAqVJB1cEEJ0Grq6sL3TEI1e/hp/mZcrj8tYthDEA3QYH2FgqvInzJvrAjltUgebxmr9QSMpNOou
7Ypeq2BcXmYaGlIED9zf5h7WwWHe8VtxYwspVxjHNo9FP7COa2690JDXUftip9mYBobtbuW4ldhu
314yBIVuI4ryqIaWaYVJ9nbQ4dYUYuZ9pTCLmiI/9eK4/qU946priKUbigpayF4Opk/cbximJNN4
bKpQTvLDT7mev28jLciU3Z2R/VRwwDSznNEEgtYMFVHCeS9aTloSj/NSqIXvrW9N19bbG0vOR2Df
kZyxJnZHTZZxGcaixrDgRwsYkYAPxTkJyPm0Yd2gN8iwF1vmyVZGfU/O8Poas1fhaUezoV5PZJEw
Pe7V17QhZYJVureUsbZWxPI6/YD9AEQcoabcycmAAWTOdwQzlzAMGJtUJXS197tt9D4JuhyAPQmJ
KAW42acLWJDbVWd6j0GkdG4eZu6eWLrEi90pt7V6SUZSlp6f8pv7yCHTMsUvS30bNnKOvHbvf7mJ
sU74cRUBUssiwY3bOi2bFS+zKttRZSFT9hQm9oJ74mPkMmbbQxfR9FY0aUwTA5LUK2lDDZpd7gwD
/rCgzQiXjdicAAVcs2tFu0TEt4MuaL8CTJNZyktnRoXWJnL94TI7KtmNYgXvPMOmmpWjWl4XwvNy
6jbrH0YR+ti7aiCuNbQFth4vBdq1GHCB0Zjug9+mOKUnh+NKVzQmyG8F6excGVYpwIigI0CqsKkb
2bWHiqYo+Jz1YaCQVbMUcXPdIDkWIM5rS/4NLELyb8unGkRxG85/va5Cr1BEn03uEIHokomEaUH+
+8Wbarce0vgNXnXTTfQOHn940h7HGKauH4HOdqUjk0Gmn4BkpY2UxlhpHZZNyuSvO3MHEMC9yLTA
VCMx9Hx50lqKNLcHb8AXqWCTtGqdiym36LFbDhqidsZybNCxN5d94e7bLenI6B6+Aigs/5Kxa3aw
XXT0wCI8CJIXrt85pdZb/1H+SQSp2lgRvxQ8Og3o+R3rAj6qcr9+ApDYdD+Y/CqZM61m5PVuZNVb
UZ3YMGsG2T1DOUItHGKrJe8pV1kI/bxa7pRqDIzqvCZl9penwY9IShUfZLXSthESu5ux00Mkxz+d
JeHi/7TaTbsSZmaSyv4Exy9zRr2n+CmdQsByhnUluwlM9VFE8MNKZxSLxFidyaugUNgormCMw/0q
z7t3v1yCHUvjaT5biB3zM4fOEBc+Kr7NKtjXq92UwI5fRWkS7Ig3MBwz73pBXy4WaONjvUxUTCxe
O5ceoRQ+QjiaEeE9l/fkrWOnKm4ph58zLkuoA4GiY25nldSunuE57SdEvjAVPqYAa2C1SzJcJC3K
uFOTKaXcp7pJ8iBf5qllbc3ZDg0OYuNUuoZYOJZ5hChOmEWLqfpNULMkVQNl49xGAl1ou9iTbLkW
qHiWmhmYQ7Gs0Ytq2/CLLTRev3dHZNmSbly5RsNINI3jEd1DuSZEiH9w7887UC3wyPHU2kRNWqRk
TJYuNuYIgkzgCp5VAhgMvgg3Knmjc8rohiHTipKjqgQj8mmeJSlnjBBZSCOuikVwqsICDsCQXrT8
DuN6EbKXpSc5c1uJWKpCAwqw7sKBrzZZXXdE2HZyo7hfo0vcp8jPTR+z+V8hi6rD1v0rw1VYiWFQ
Eh2K3E53h7IbY+vAD7oKi1AObtMqYKqeppO3RGyPx7jAPw2KBziFdDoFx3/dE5pOuuS51Hwdc9rc
Nl/5MuSV07rV0x86JW+d/0W8xPUYq3KJU1K65kjDcPWFWBNQ3VZOcW8zFId/CKdBXa8XiuE+yzu+
mLlRw1BKEh9nMXkrMu3P5iiQKn0m+t6jQF9mp5+tpYAbBFPo6JAbZ09EJ+I0gT/oj9cJIcimjNzJ
TmJlfs6G7ff2CgozR59cGTj2leGzOsUM316tyr3wYZKpniaHczCAdt1QCkQU/IsMoFHY5F/PdpQH
tjL1Jpc1o4EJPjS+OiY8SYcNAkv8WHPh0gG7TTCWxJgjYFBWSVrtaXOtgZmK+YBEqzWYE6kMx9vs
1V1uqW+M0NtK3jdNWhQaqW30xQUh93b9e3BAnML45+cBYBmXnUHk1PuTcgu232tpUeQSv+6cBQuK
UT9QH8FFNxAGmpbV32A/P3+mGcw1xAlQB9KuQ1UKnlZZLePm0l8K5D+kRM7Xf3AdGjG7u9ZkC4T3
tu+avvhjnkfiDEBtm+EKEI1otv0XsdH5YcNls5pEfo1eGp6zBqwInwxcMgpUdRU4ZVLVCvBzEsqX
UQRsl78s9HvQql9bMV+D4kO2FLVCADPsoyx+Duf9JAw4Wmj3nNew+GDQyxeG7Bzxgv7z8VzGAFrv
iYWktLkEmx8C3co3O3Zqe+Jl0XVrS0uGmvLOgDwe8N8hwP/6acXAOY3y2sCg/zSeifYAU8olAdzu
GsPxH3mSiQ9r5x8gT8xink0BwxptszeIkyqeQlur4+kqluwMDVFpJzERSozMxzuBTNwx+3eL/IMW
2/SydhP6svfLhvBeXlH9gjholH0Wu6kF55N/YEBMam9unW7zBKUNdB5tFWc8DFpaqYAmGHqv1148
iTx0pkmjNkJ2Ifk1BwPravU7zt6sgcLT7Ri13wPS2jZ0V+1CtrZKh3x9/NsukFWF+YaFhmpvQ+Na
yaJiGoOIt2CDNskmLYdSWu9RzB7MIrbM3X8oCJ+sQLNE3Dc2NbTTfbUCiyAv7AJd91WBoToqyuOV
DEJu4Ubr6nP606o7JIb/Vezb4S+eMUrDDfBi7EeDsUUafkBdSiU5Zb9Can1Jr/lJqec3i4DxLCsI
IJVPYkHai//NgBBmfln9ueClMleVzkiIZ0u6zyReK9916DRQxxqR2o1gFaCQMvfhEmLQvt9/A9oL
xvpfSb/eeEr9z2WXcz5yOPfSGL2ckHs7NuQxmifXKIO1+zAiEZ/K5d9UQxI8tM+//wCdhCh4Jugi
cnHFtJxGUmex7TqkIrAgbgKShD/kl6EgTgm9HNz0jWHB0cuNDTEYDheh1ZH4MjAOLbPnCfqFi9Wj
UKdY4r4CxJMR0oFG8u4QT2BiRorJglHGPyE+nln5KDbiPiiD0tkZWr7SP4Xri7onsbiFkntpYoGP
9Rsl2NE7t5852pgGEmMYd8N3KtTcBqB8B6CEWANIB0XZl7pkFAh0A5av12e57msTIpSuX8lpWvI8
q8Rnfa6xVMSz4UAN+SwFLn5FUq52HK667RlSwaUbAGtwnCRvwZMOO2ue+KjjtczxsT+RN9Rrptqh
UgKpJV3nzV3USZdYNXbWNxJlvD76fTUwud+Ley0PXXkqdIIlW9IWOrI3aZ172Y2d5F6PWzRssBv5
VwjCvYUp1ar3Nkb8893Z+6fSkj7++jLIFAjkhNVUSkNUdTFynoSPY7/MRBkwFeH2q4qznGKDKzCL
tbMO3WhOovDDPeOP8pIi/0j46QxQfCvT+t3B73hLe9Ys+bvIEAXNtbbQ4ctZIwCGlrjh86bNqXFt
dkeiY4D9psbQANH041/tolN0wTZBe2U/QXJrUJBFXGI2/BtLPTkega3B6iiBxcKOZM4E03N0SnpS
7cCt3kk6ucU6NoTf/wT50uWDNXibKKRc10ms0nz7NiYsEZtJs5b9/gWw5cwR28ML72dQOEO5PsA2
ifKelveC9ezFaaE0dJCERld9lNb6SL8ASsus7yvjEFH+Wbj3IH8BjA6boKbZ1kjgReI3mec0wQKw
/azjrDi/i05KsO8ASHRANa6sEWxQl75TJdgSZU8TgPPROYG9c73OsdhATXzG9jutvp62TLAwCqmQ
ktX59Qw5LsNtsaLNlhlnxxtuT8crAOrKFVrYQINoER08aVQnnh8gDFHsUJE3E12kjtVlfZkkBY+G
QVo6LSJ7C3zpoazz+dZC4U1eO0AGO78NZM/s1CmnPFeU1VJGNyZ/dkFVjMkiebkKiLIaI4MLQY4f
59UGtAoHn7+GOveA1Rit2DsyixUgLuNR0MIHdPyfwPRbRCKOyKWXX13G8QlqgDGzRx+DJOdSGZb6
EOc4M1LkO8nlh4jaqt14ar5sY90y02ZHeWs0XgCc1Xz8J9yrPkJq1XQLDXgt8UyM3Wnp/ScCExBs
pyBS1Knb6WJtYAidL3Ww3P96HJIROAeMyGgJL6fSioR/r4e8s9x/51tUAbbYClaJKqpBaY6ASBoZ
ghzj8hhHCja4kySVkhQIdz7CoOXFuxDQK8o3K5n5NdmTFpDeZxzyH/iuwLXczGl+PYVTLS2s7sc2
jXLXSgZ6KqChm8hXNHGiwBHjCtQFucX5hY/Ya2zfWCbeHY7ka3qu3Na2StkxvSVLd77Xavdl+sKc
GO1dkwwICqLs6U/rqE1KhActBrPAZQpmUK2txzE/iNw4pUNGZrSyRrIGLQurIAXw/8j4+W7NbWva
QZHIBPYWkL8pwPO6nZ/tdeeW/o6J3IzZ1sfKVEQLIr37scxGIE8Rwx18n3LCweA2mQY8nUg1vJ6D
HzIr2EJhwHJ/vf9rle2FTV5oKnDjeiGx4iEThLVhSPcfDWVJy+xNx9Payl2dbxJP2AbbPhrniIUm
TrA429P/T0hCSAWersVyKh60mDHspTH3TIp5nUDVtzi/9GHl1a6xOnBWLRI1AEC2hgH70ukyUty4
NLDNRkyCHeuBxgfx8+ExaAFvYb9kt4w21UehtVU+EGw7+w7GPNXerOVSx2ucd3RKlxEX/SxJMI1S
w9Iz/Wa8cKQxJchFgNRSouWZL8KzYxfuC/fRM3w6WNBLg9Y8czMgMOY0Tu6SQXbxrQ1FcgNG6p45
oUT31lIr6Ao3Fybyz0MJr2oFkd9hf4GaXejY51743jq0GS7RJSHvfRKeEceJLC3O1xCUHd0GsHdN
Pd1ljEWDXGCG4BK81pwM51KlN6w4Vx2IDw2rtn6L8znZBTk7Nx0R52Lgo1KY77Ift0DjarIR2KDE
SRvp5H0qBscLRpayNC9YDqzTLR/5PGPuhMGhlVgQzhRTjrKI8pA20ftpTVpzEqfKpqjmSMIUoRVm
Edbm5VF2X8M0hxKjoFPHhQ9akfkeap3cmB7bCX1Qyc5TRLYm6FcIwlcGIjuKieOsB2vVFIOEirki
bGd6MKqKd25gRb5YY+ioLDEWrwsqqlsdK5x21RcHk/55baLIDg8jptrURlLnEbV4lziyheoLPenH
zEM8wrViDxFGzG2XdKqbeQ/ZDRjbb6yOeNPgxBKz52lZEj66bnkOO6uilLwDXUYgtun6pm/rP6Sf
EOwNfeG/Dn8cKNdPwcNDWsJgq3xbqa/aNXIVgxe6JIr2RyfVEvmIZ+82w7LwBGgm7GMlPuHU4bE+
QSyES1cdwPiwzWeN/E8BFaMIWIJbR0IDGoYcr7mfQyfR+OC82BrzBgiEv/AYr8pvpnb/wV0ZSW1E
g9KUSA7PhiHt5Lj07CYNrsM9lkQbbFkPVIXOfuLdxwmUAFsqEv8ywu4nQpvXFQJ0XYqfLCBMBySP
ztCC7jM1K0O+TEEvufqSdZWUeIvLMdzoE33/E/JSJBJH4+qafN0Ts8h45b6dFKpGI1u3nOPYP3ir
plfYYqxu1cjKrnq3xAPLnxL+fkdQ4ar8XdOsDNmWDe6DpcOTw4Gi+K1QjLdyutHCGl+HGPNaTwrb
NvlTRz1eqDo5PwjwB/UpoiWWsrkvteg4XuK1IYgN/p9chb5tyfYYST34Im8mEY/uAJvDndPr3JRJ
ERfeIp+QRtY2a48tLA7a46+toozAbuN9a3/ygoZmHde1uCPLHkASTzfMoq1xMyq3Z6BJBmLoMfNQ
OVFzfzsc6OtymaCkz+i2SY77ujivK+8qYHHwORTvAfK84svWD+6JmYT0K/mGlN3TIPyDCzbb1UdT
fxfM+iVR+JOdt7I9vgwVG4pTytrwCukg1K6GAHzEIS7sW/81wtl0p/nTvLjSIUtMN3OpZk5xoffa
NSbFeR8f6E4nC6qbYggnmQ7igohV7w45Dg1YwJGfgzP4w/VgOUdUwq8yLgVStNE3t7SvCT54u391
59tujlqKJKczwW4z233Pe3HciiS/SlLnnyjIWOcOCyXB8pyCXgttgvFstkcm2lhdnPHI2enuDF0B
5FFJ2L6QM3210zFJFoKWwo86GkE8TOxbYD4AiRhucA1MNbtQZkUBYZCvZ5DFt+lxULqLwfjr/nEc
YqsszLkcgBdYd99D6hLH4UEpAFa7shrCpbeEXmRwGF5KithIZLJgAXBjaUhvDJMIK90NML47UgeT
IBJj9hLVPkIl/dwe+C5lOPmIXjVamMiNsGkh8w1gH6g1FWEcV6HdZUDSb6ATNli5o0qYRTz5akbV
+YAfK1MPg/4fmlY8za9udq3q1sYlrLXeoO+DD1v1NbiTkA4CuHHWGIxxTMr2rM0E+Kai0vYxQxu8
B0mwlKkBfWb9M1CK2G2FjChaJ5cSmwqpKYYvf1ttA/f2mYl0kzR86okkxswYTE+GquvUuUp1GI1D
m7Ws+s6FByH+F9la0toj+ETgDTjjo/iNU0UnPUbeZr8A+6J+1wQ0pIHiSqQX7TOwcUROpqdiiHlS
NsOt4ORkCrcfpz8iXmMUupeu3yONhtGuXQahXu5iq7cHTs9M9mNn6qKQyx613X0WEj/xQXxcLz4J
5nf5J0suVNYEWq5jELuKjdcYQZwM4/6y6HF00G0AoZni9wUAbZVXx1UetNKGhI0emMuZgtCCbjDF
X31eGXOpuWKlYPgg40VcvI3pRhn6SwaDHLy/rWUouVOK/oDwcXg3ppIR65yWydAfIUFS//V5cKLv
wxyW1ipUTuO5yyj+g3//kFYgw+UWG65j/nplDEsUJZtYYhy+9X55dquOGhpXB2bKNuDicTGNOYA1
Qne+4RTMXIcpIKcKXpjr/Aqj7AzryW/dWR/SdwqnmpQ+qsjNxFlZydUitNfG/aydAGbeSFgPtQVZ
7EFbt6XZX1xDw9gNeWGQ7HbMhkb25heaGPob0yT0yUvmE8kDPF2KB/Rm1kpKSu2pNcQItkNBblCb
a9ixwEXiUe91kJP0LMPELo1IIPt2BMLzgXpW1qCCJXHeU//i3vldF1r/gOtLfQexBx81wBd22Uev
qtkjFJXaIG86hHfjOc65LLBddffaBfkusB4uEnZPujrU111Ua7+B0ajWbMu/lQMFFj389sJn3hB2
H5iB5bGZEAnUl99IVdwY2KBg2xrKPwJQUlbXy0xyS6igoicJLbOnQEX7D/leQlAhSNcg4GCoamlo
6vrc+iU7HxHju1/b9tPZJYAbWLeKTZu6kxiJOXXctEAdA4UcE16TfKgp4pAvmQZxDpR3kaQbVO3j
1H8vhKRwi7dCiXAFen2obRT7RNafcEv6uk3iaTVSJI6E3iOaBGV6smdM8rvxi+ejjvWSXqHej4m/
+qoD2jdJ+QRGY2CMt01QsDiKa9M0te1h+7NyH/TwzabL5589j0+TmfxCkejcyOcEwCWKxibViRZ4
CBPPdN1cxj1WxZSlhsyNb3Uo98+Il3gX7+Xe5cjNjjWK4TzGa2v/DYX7+H8F/B/S1EWEaj6AVf/4
pzFVZO+UlIwMbUjTuOlaIDI4+FFJbM0CHN/KKNiFTYHBEtcHB2UH364LT54V7Caosl8uH4oOjwIZ
dDFE1Jg02lRbNahAON96z3D2tzFTcqtbvv1n7cTy4mGtoZWD7bpK0/43GbJT1+88LBFOY1OPkmL5
R4XbnQ7A8W0N4reeS5EzfR6M2rrIFnwmjEh+aGChGiqNwBVgvyz4uUzxpXtZYpkIIWM2FzFrkkOH
KDOsC+GLxoXn8CRYSf+zTHAdq6Z8qPnKja88EAIN8P9YIW9BUGw0VFngTK6PvTGwEMUSQUscIP3+
EGNTkJwDRXoykTVY8akNhUYdS8m3N4fgsXuBzBaKePym/Ab/7Ho+bz5W36Gk3BkjePT3AF3/4QQh
g0qAa9TJjCfoex8KxXSxJnwn7D8yE/tAObeXVrjl21qjmNdovnDJj2fbssyAanBtsPOnydfUlW8q
AppOQ6PUb43ZoUFZLc3Cec9TP8H5KRmgbHPzN+31kELkZ+yiS5IlmEHNSXS4lqW5Rln9+FRCzYgl
2Idu0A5V859ybKVB7wl6QK5pAUcS0mRHKlC+yCAyN8UFpuufq5BZPGhkxCduoMTBbhhT2qTiCdbq
zrfpGHJvYi1ki9VdZykxWCpZHOZZkCQ8bVfS+dhKfsJ48w7MNyEi88Q0fIzhmrGtaCqJWTR+4zZV
wTwdOtE553mwA2yC3tkCCoeaa6y2rdqG+sYgFB04CNzrktgnh2A2TdYbMhEw4qmS8HlteqAMDb7a
3dbn/flN/CGaNnTpXC2D8ETmsB5zESNFqH+Z8Uca8NMQHpdjg+b/S8gnpgAPNMGjpY+aS2tAuhPj
8EPipq9WjfaEKau8hrkfhp9WSU3eanNxMa5XSq5q569xRmgBhPZBxWtDd0N/SUIbFz0df8jPFyl6
5UsxOK20qW58uU8RfJoy6ht9z+6Dw6FmxG8L0Q5VFs7geRjONlieWl8HnRTaZQFWEu9HuT9pRdoO
CY8Fy2iRdx/7hH/SRWfXLMsoN1rfsz0pIlrNKxyy7pDxNpD3sg4LhBLT5ML5pAq59myFaYO0cOGN
40uD2kGjmz9V2Gt5IRinInlhjJrIgOr0xisjZ+nLgpcT3ePzf0ICPYBFHNbnZHpFqrKaxoiDC2B9
SMpEalvC3hkum29t0YDVQf67w/QO2l98LxVtiDvdvV9vunzNofrsrkbyfEsP5jyw4AD9oEJABBBZ
h7iEQHW9FYHb9fU3D6RHPWFhOH09JdImtaIoL0BK/0INlD6fie94WiM4sidD7ZpTsia2h7drdl/B
ZENyU8z0biRbSEgS+y5P7J4FIfy5FqdDuKU9f7IBmc7i9rzW7sr/MAMRVctUd34fEQkB+f3K+aBo
Ump2h39nomcZAMs17j+woUqxQqkkoiLs2WEM6R1UJZRmOyfar+Rd1MqopqpztMYdQ26W9DsBnkLd
J590j+8XigW9Zc6ek1gC8PfEXzxNGCDVZbDEajk7lLVICeB4U6dCFZnXoTEpZ2WOysHq9CiveIy/
AZL31d6mTl9BpDhijgdN5rYBNvv34fYq6Hw4anGdwkpnvcFJPPY1/YRoUhXI28W16m9vb6llaWzR
UzzI92dEPCiIsy0L3lIpQjDLROqJ148DFCMnylMWmiw+kOtj5N/bj9ARmxSOY3pD1LHQDNPYfoFa
ClgAmDkugBIbxU3CzNvr7AivUeX+XC9fSTlfmaRJEUNHCsv1pyTe2uoeTmH7FIX2H6hAtG5/yfWR
/hnL75uuccjePn5Nva6R8PQMwgSE+KHcjEM5d0CKlsa+VOSCmPSML16oinTmuF1PXV1vCv6pn3ht
bYQxciy9g4FFr8O4dR3kQT6617A0v+sXC0Ghg1UgPR2jALeRppMTsrRHght4BJoUh8zyxUoeczMr
Nc16twzWLV8CleXORpawoYgPCGmFEjEhERFbpu13XRp4mgjjP8CaaAjMtrX+Ynf5wxGOJDcmx5gX
/e79bQ+f0Uh2WxQ08cBphd2iW5F6Cc3kCIJdfnu/covAlSnRlOs3I5XwYKx97nq+k52u+9AgrqXX
jZPpWyZxh7GZW4dYw22ZgOUFc9ybt8Nhb4W6CWlwa2OHS6X5yZfrkHOzkoh7UKVdlwH504bvaH4K
9xvZf51bN5yvy9Fz1LAFRlWLupSFcvh7P/rUJfzA65cHtEMAhmFbMGCl0+O1RzEHmUuk64+nbX5Q
Faz9y/0lOTd9UdcXkbynUqo057CzltVQCjiw6S3N+w1GF13ZDz3oAwfjbeL5RIIHg57JaEQIb9e0
6wO/jO4uwFZ2robs5BlWlOwpUpYYC16kH83drqFuEKKbJKbNIVBIJMzW6qy9oUFagFKXlEgpKmNL
KxGLR9bTVtl0sYfYnV+b0lRVN/Q48uzkKoCPcr8sf1Re6eU+nhNsAc4gkDS97xUR90Mp4tHOEQ93
Ymj0VRDUUGZNlFO3CGAsDSmzAbZcaNc99TTlMmbTSdFMlFKHD6uo2Az14eBIcv7YnBO5qZu1HZCR
uSjb6oDFluTx3JalJ+qDvoIA43uctW3FteeREB4atZqGVizzl5InDLImB0Hu+TUtaykeXFrFft4t
s0tTN0/29ADThlm8+FBgbLF9ZHT+1NC7LGDS/Ao/4mJevALwSlnZcHtivzgRIHP3V7DRkWaO31hR
3RmTDkpr2zYeTuRoMmQifzFLTW/BycxJx7Ccm+O9WdHGt7/LjkVamjjBg8xuo6QxTTrqVUd1q5VB
8gU1RnVq6/PhaZPIBQm10GE2BUUWEpCUk/dIfDAJv4JikAPzGEIYmBYRzs9dUs8C7U35nm2ZVsdq
sDjWXBH93NCve13OhdG2UDOWGWSfiskl0kY+hksQqbeemNLfo8BB8GXKs7ea59bZv4WGpVx+/+pQ
NmWjyF7ovPg1RA/pEc7b0Fd7Bci0JrQJj1R8KvpizPaQqV7HBstsXPH2mfKSJNr38CjURGIO/hnf
M12/np0Ijg78b1J3W95Pu2UXt5Uh+9HHZ43wv7ga+rCoRjg2OYU1TGqBRrUZr0y1wd2Ajw5lEYJt
H8GRQRxUqhOzx+ut8oNS34ft1pR7OAbQkuzEJp6rY5PUiNHHhAPwCWQFuDf6py5q2g1mZGYxMH0y
Es1asp0lg40ry9vcLB5frmt/T3bWXDt1b+jW7RAkPSdc0ccLO6rK0qHPuUIyrnKvO0zxQJ5OOrDe
M7YB48L7mxcTQWzNS/NMnN5ZIf8pnnNKl9+ywA287CaKZ7j/qoaNiz1HPxhyDVsy06tUNM5JHyEm
XAgaq9YWY/fC3EjtNLl/Hdmj2HWTJVG6XyyX24Uf7wmC+9p7S3qqfhpujN82eI6JGFSfVIr2d9Nz
paCbH45NAhVZwEX8BBie0g/BJSwLaAbrHtt+VSxVjm+H43MvjDUXAZ9W8/07JVMEoUFf3tw4W9ud
IgXua0+KfcckEKDUOdLa6drWqphILAmkqkboeGLvpJD2WYgfTAJQhtIgYa24qOnDtuH1PLyAS/Wj
484F3ya/9gbm+xJC4xqxrQ12vIJaNZNcIuiTLaPT/pYZamMu2Lal6cgYCXP/RgLtwUvJModq4Kna
kWZADsb/lHT7+RM52v9xIFuZoftOJe3UykYZlZzD3XynZQC3VA5suibjpidRC8kv8So3CrS88/D/
yCzirdNR1L6XUA8Roja6b7EwTxxaBTIBZKxCY4A1vfqiApEMUKXOGnvQrqkkx+5+bEdOWrj7cVY6
FqilrupSkgNnZY9zYR526I9uiAhnE/0xObaZX24wRCjMM89+A862OIoFZhsYGPd/Hltz9PvQ4AgX
wJQMfRRQBOIDSTIWlYm4wfyvsJkMIgLXqcDZwKz7qsmtYWWeAVhOYccZ3uAbc/YzKLf13eFFU5sy
GcTAlUt8IP5xMYJ6v2cDFR2+bVjRZJvAFePi68kTomRGcs4jT3IwjFf6Jo9ne0UK5XX5aFcjHvdN
c2q+ccP4R/x4xSfk+46Cnu9KxKpOOIxFug9n0v0u3yrAoCyALl52x5qGbSphMQuCR9tOvf8cJSxp
yR4woa2sOkym+H1PvjpRLil2L25ZOg8Ryt6iSx7HuJsgceXD+zJzqK2io+eU5CdnmRl9KAGQIXEI
rQAR3gSgPammOEgwpfVRe0F9KKpJIWWJa/k1LtqJUAYj+p0NjOqydri2SGueHqw7QDUj6zQnxGu8
8Dh9Ph3ydOcEjujPtbnjsOqQNOxBRzxO70XAnBHMOXm90XBD+rTVbL7+LsuBSK0RzwOhQLj0EinW
mA2DmiP05neJKFlpoNphzKsuWQv0MibnZarwWS6DZcSia1NJc6NkLykL6hSG+BiEeAMqEWwf+lG0
75ttdWlZ5WQNS0Ko5twLbb1ldRtiaBo6NwVYK6r2lOsADdLxoVYdyasMBNa4Ynh4jaZdLnC/xFFa
nqist0kYavlhGOrcN2tPqvNsj1NKto6qbaH+iq5gcz7mXpuXJMsH6ma6uEKuK2JI2Y0kNss8T0LK
YLvK4sAa9ojLof0D2zyOrRivIdHFSaCz0zxn1v3So4hgGwAP21k+wWChbEq0Zjqrx3uP/tshdV+9
omlVRcqNSpmT3bhWyXR5FvyfJzZjsuR2hHBJip5s9UONBRlZWXQ2A4h91IwjlR+wQM8CjxBeEsxU
MuvUbHfwq6uIndpvZzMM88Sq9yl274xSDA4crCKRpCVUAW7wMpNIl4QcvlPICJ/otiAr21rv13+7
TI+OMMGGAs35RYWsKmuylsAroCaTDGaJu8F8bSmXFktp1c52pKusJe3O0sC/rnUG4WrPE98EDGFd
PXWHqcoJtQk/QT+izIBXbyHO2metVMP137/4J86sZZhG+w3q0oI/th31Si481gbzqi3g1QXVfkH7
Os8hQkr8lZ78Ddui2rPxjHM+SUHEL/AikmygCML4W+dGBHfUE5+DAeus5e2I/MzLNBSRG4JTUsgE
xvBoC8OakrRjXZwl/2opP42Tg3ItqF6nZEcB9DyvbXTU/7yhcBkG+5VtCEhu6W5an+UxPkln4ypv
Cx+WCsv4XqEU/7rxkWN3IhecgodsypRK6o0mMc/HHzarwTclMqf4acztHMWEakda+tK/FrkE0gpn
tOFpqFzsl83xUve12n9y+p0NQReZ09zORhgzp1VF5J0xj1XeLmsc9msKmyfY4454q1DqS1kmS79I
KUE6dDZX4aeNAEdYpo+rMNanVS44IAV7aex0v6OIKR2GbKUTxcGJft+4NUJcalXeSaO8Spd7SK0K
vviEaRhWo9ybK6a5neGpUVNA9FMNDRZd8ormClRo4b7kGSGxNCmxB6zCuMMvyxkCnjp/5JqoD2t1
LY7P7NjL7gk7weanGC4kr32mTp6veImMVPJ7cNjs4il0A9C4ivt0dBoKqr78aENkLujn9cyfDQnn
e93WK5WFKpY8T8wStr1CeFtixpeu3hG/xm5m8ceE4nWkTGzHBrWCGugH26wQXILom8UygHHTbfd1
BYoEpRdOmrqNSsWflHOXMxFVGu5AkMk/WpVaEflHzs8eYasu5CJfGXNyI7p9Qt/AbMXHbfIEGiUB
p/5J1s3HVtEVhJW52Tpjz81NQVVReC5VvY7VZCtCaCDD/pasokCwJo5fFxjq/seomTvuRBrMzzeR
zcCRPIQdKIsYfs/LBcwHudkfHy+L4HWVzICLQPJLZlL5SHYTxTrDdVlZw/+4eQ8YNba6LB+LXvS2
XHrrghGP81+rkQi4ZFgAe4cO7Dj1u9IWJ9vPwCVswJqu7cXCxeTqP/nWzTt2+CF+3+txGQ1q+or7
ERX2qo+tw21o9/alfjRPRkxBOeQ0kIifsmkgVVuVlUPINJ5JGNEriVnbpkKOhSR80wjrNGJahAT+
y9VbrLxCNVi29dde6pbomPjvhFZ99QwCEpKa9D5rmh800Sq2VC575+vRfbQNUA24VVdJ7XKZsjA1
rbk+MBEWdvTF9M3KHZD/24ogMcFok+MV0fKSdW6C/Cr8uORZlT8ZMdhu30mI7iQs1bwE1wbf9cuB
V0yvtdKuJwQQOJmUKld9L4WfFZZo3z4rz6TmQN4RlpnWw2seddiuClII2GydxkXFvMZxk+DW4kus
qvx0Q6RSfo9gwtLaD34KCnBqGV8MAIuyLBZaQIsLMLCUeQY4e/FC9MtTvrPReaLfzZsYPZS8v/lI
1/zMOnyHEGLWgsMdOSrnxTMod551bSVJbbhhjInx3KZ7AhwDWbrN+7awmDMGiKr+gLoDnkHvIlxa
V4Bn7KtEj/T8e65zIaHDbkPk4d19JF6VjqYzsxxycq89E/FzlfcAEHBQ3vl5naWtYOtkx4wSWkdY
+v7a3Y+lGKksoMucU1F7zJpPDtaS1xwMOOEcuKTfu5GdjZ8wHQRHfRwcs7TIWIocdx4P143OTvMf
W1oady6oNi4AEdxZkxF/EVuu7mFMO4HFYxvx0OejRjKTO0+uY6WyO2FZi7AM1xrndjvorhqlq3oc
OzfvE3Yw2NAOB2j0TXnMvA/FHaSmZiat4zIvf+/Nt0RqerLLfEZDhJ8H9y4QmMqXFsPAKRPO+oyv
z0i1ynKsXeppq1KfnN0iSIfMGbE/9IzXvHoqy356wlrvfEXC+lOANVY62NHDeyhbBVt4JxPK88YW
ZcnQEQ8kEX5OXkDYEp40LF+2ccFUk3yM89OQUmS7oeoD+ibmMzpegoyi1In3wSVhgp/USbgXObtC
rdmY4muVMqIufQUmUlsrUZ4zpEyfm0pTdm3VQkIPSZtjDxXO+e0jcfSHaaPkwpFCF1M/gzcgUWdY
Mp5VGJHKehSCRp90BZzQRmUq0FyckN/W0JTh9KrjOUIr1hnTR8wh+CjQ7tXLsUZMDkPCrNaGLv/w
Kc9IGwiy7DkV/IvC3sQVbn8c76rNtGZ7T5dmdy58xZSgR6dfPZN9l+cSM7VaSIXkbF2M/p6vEClc
/XtapJKo/LjA2msJU2cslQxnp81y3T/hhVPMtLtSQUNK/zUOODiE09BMdWUKCYQ7LInhnGLmOMiE
GHWc9CaCe9bhP/PvmLsoejKw1SAw0sSOxV/4GHE+Rxzv10WPyhp8DB1Q4GS+fFoaUPoE6m/W2bRi
UR3aWT20FsjLVxWwGbe74VMJJy1+NQJ3ijr6MHOTR4QYYhf1+z9oozXP85b2GmR5kao54bDyArCk
cyGGxmyJnMW9WdY0qS8IAbW4sRDaJfnEq+1Fv16fNd36nuqPJUNd6w06N7qHnq/H1ydy6EKUOHdA
FmYUvurEX3sjdScZYPRjdsPu5oTWWAYGWCs6pKuD6PNKAqAdRsGdap5bd7b7C/T+aZCkzAGnj5u9
+A+5ZPmJEs8cyIzJjRhC4b0v9+IpMvB7kPTDZR+ktXDTs19sDf6Pe7kndw1bfUyW+A3JJNPW/9FD
bUPW+ol+TCf8Rhqzr5POQN6+My+/UC5pnNLc+dQGeFmjEQdgC64dQVklHEksH8Uz7N13z0/b/Gyb
5XSt8z/2IQv3Neu6sUuDkrpWghpRjIMoBld6ysilkezTATop545VNZL1N1NxjZgMgYiQtoiTxytX
JWcD6HKMNCtewthqWkXsZZr+ef/TtpJMCkAWoZg46kMelfTUmIAsLasJxckfGQmQ6wBkX5VcTpCo
xUyoWOPs9+a/266hcotzVUzU+yIhoZF2kvnAwz0kicxSb7Z9yomhZcC7JpgafETUGNbgtaJ0NUA/
94tJg2oNQgHJF0Hx0o6blFx+AK9VhIyMPiWUysRc+F1SXY9PC7l88rQ0oUeefbiFCQCWVuELBuga
WkzP2LClpT8qqtT8PCNrXXgctYguS8Wf6EfyvMMpA1yiC8cWoi6+Q2rqJm2STdgyzFemO96vflhl
OJgT8K+6iKCQ1Wqez8LaUvnC57lFRNQF22OEvCXHNxl133pX7XslbFUrgOFE2hcnIgWBnwud/bcH
tHvOqo/ZtnppuB2yTIaKGieQY6PeQFFtrXPw1hPcw6YHIbiQNgneOCYVioVOvBi12dJl005xOvJQ
sb1bRC3pHdpQ8Tyy9xBWSCJUbaJt4VcsgET1SelhlQpCLzB0DFoFIeS85d5KoQm0I+NX/3poSYUX
X0BJBELcOTTBUrc5RuyqCXA3Xfes3rngUYmmi0VZbZoETV5XqnEhClXEuV/4O0a7Qi4XpJaKNgKI
YKezaFIFkpUJqH3/TfMt0qe5eeFhmNtDhuL09sjF1iF0AYJ8BHU0B96X9QjgKdPpQyvqBvibGEi9
hiFiWdO09UA9ZeUAgDz3M+k4KQun1jUbrlKcS6CL8L6ji1J5KnOfrrzoc2HbmoSNW6PIvXhIQu1/
5eKLrgDOLZa73j0+79Ex/LRK4AtyUlJ4N8P4UWkV/QXiqZpAnH+XvPWeYk9ESrvO3Fp6ECkXpdV9
QOFdmFSEiZ/1AKi9OPQgl0cL8J8c2YTMitVpu0j3fEU2ARDhEDsmA9nFnX5gzU0P5H8y7FVg0Htf
abdJHp6m6n74lOMxmxQDDjXu2GtKFRzaaaY5M2ovKdTMH5jF6seWoqfy7fLleyWGSBaoFyUNGBmo
ZKUdfy+muI9n6RnRSDQytPeYsXpNulQFe6aTjao3RI7pUJ/+VVTn4dr9QuVBVWvdtQ0Gll5mIdKg
1y5pgbY1v6THPO5CvkXbyAYHgRAcVmpIC9s94TKve7wtdAQSAfcjPR2NA1UTfz5Pzl2Y2Ts/xYB4
q0eLDX4ZjJVWQ/HZTp0T+fBpOd7kZc8XDrD2Vazdm0pDV2tfTegcLeIZuofVCBB5MEB+i94Uq/RL
qV/t+eYC0LFZ855eA+TIs7eQHeJqAZ6zFtHwSUkUVuoZEQecKnL6hD9TT+kI2cU9vbi9l4GGA7py
kg/QWwT1ysnknkwsgwpLMQlwWAv7WGRuTj5gE+bM/GpbRQQOcyCwD9CBERQ4ycDI+o5whHJc9T4L
ifn8tKcLIYS7Pw2UNrMVQ8E8yVh2oRb7ntxgWGVoKIChsv0texh4SEvxvRVuzBK38UwesNMMjEsK
BisXEhXNE4OR61rUg5u1HBshtQkGbKUEHxcYHo8pkh+keD3fuBAS74zZORvOFCUWwd0vgvSX+Zw8
q5M7jnWhnQOySP5Zr4vi3u5bq+BdrhbN1er4AdiCee95jtwVcn5IENFg/rXYmEbQg1Qr4WQDBhmB
W+YIKPxzKxReslcxUYqdvc6Lu5gxAzTqmNM1H/j5uWS2wQJOlLnh0lgxPQaI4/OF53SE6BnRjMUN
IXCqBlmaaw2Z3hdcL/jGyUCPa4plVPdcV48pp7bZ2dDzJoiLcIKtMCqAJ/JHDJo+K8Ckr6ui1oKN
9ik1bXyFHD829UwyWusAsajxnLH2CWbRI3r6PbP4JEcNXIk563JL2jxa7cgNGmvyAhLYenLq9eiz
GuXYRjMJrQKcTQWr3ZdoT9E0mBZlEHKEhJ+T3dBdBtmM4oAKyYbrvbxOdFHZvJFGFgiYfPPb88YK
uW9Vbb2aUuiXAgnR7Dl1nlrqp+QYeJ/CHs/kloYClngL2Oa1TR0uonki9wK/vLvCOYvU2RfSFsx5
0GdWF/mc0p4eDJ+acMVk+iSsqM8cHeQu65EQPPQBs8YEJgmHIeisbX9FTuNAgGTi60cjFElXnW+3
0n1WDQGe7PlhaE+5BTEFxlFOSGfvPNkFcun54tJoJl539hSZs/Yh8/gPtbmRy3oQMr3yD3e55nSp
6+l9BOxD6g/Jr0/iFup8x8PzDx3axwJYqaU71ZPbjXRqqkHSCVSVN4fVNUyTSm2o2bUdKfnSeV9W
PExyShws13NYFb6vYaEQFw13G9x4WfouzXfulq4h7Pn7B/kmvdeD97nmrhaLyTokldWnCmyuNJ04
8CficiW/46Zc1jQ9K9msg0hLyxOFrhRR6Ni76lBOZ/2AUlscog9C91rP66fLPzlm1tMFy4K5tlLJ
w3GbqOUzW2qLybVkoxE8Gv3In4O/4Mqk9LnwMfJkjwo6HHk716gdPMWQd7ohgx1TGpIW3a4Keqfr
1wNab/p7LLqD8SdGYf+J7eD6xayRGMVnTNvqoC7O08ve0ulMajE//PJLs3tbZNS/raVuWaEN67E0
cWYbi7Is/O7V4Nr4hvwCsOmJANUl5pDlMKAoiVJVUis4hKZ15B0SZXhK4dTJfcLZM5mLJXjBdeOi
J6D1jGUC7r0qgfOv2vnZUfT+KC+Bi3irZfMX7ryPbbMWuiYj6cREov+ktlr8pgOGh9K9uK/KLbYr
Ysgsxctr6KkawaplCl5rsqznW5OOuI7QkIyXMmzaMuB6G+AqUniw+jHoHx+7hCAI2wQ3Gy31o6yX
BvjPuZhfmo0yTNyZQEyZfAg8GCy738uU4piXwvXT1C4fU72g7t57hc0jCiCgzZMzlHFbvtR8Y18P
P42wuem7Fjm24giyQP45MBSQI0k/L+ucgaehmQ0byT65AbWcg3eNDeO+FQM5jFMnmI6Q6F1dVj9i
FaiVnV8iHsGMtySvf6kTGGlMvfwwMFunLk68nz33JvwCz3cwj95KOPgRwPhI5u9LRBEfZUbT79XN
+iQedqM6SDxKV6yHs7aGz3PbYQ5YZncSAm/ljtHu5FrYkwGn8BTurzHOIuOTPnllmNHOLVxuIQdU
OGxmLpEKdKkU/kawwhn+sr/VyqY3U2HeJLYA4pcdXm2cR9TvFQTXLaDGIBgnE8WNPW75Zf5177Jm
e9ecUWTtGvcA/bLSpPFuGqplaLQT2syv37/qV8Bopzg3VqIJ7+NwjJFZWBzgph9JLZdhqJFQQCvE
a6IbvvEB3Ov5WTDzoYAdEk51l1htBZEDdpBO4aoEflu3T70vp8IZKGxvXSlWMURsJV97eLFdwa1G
eg60wekDqED0HxwKiJJPxr8ScK/P+VeGm/vvuJwl3jxwXpu5lpa8Dn3l7B5Q8TAD/SNOuK947+WO
NNkWNXsI3qJ11zyraVNugv94+Nq+yIP38RJaoz9VVLtUSWXFJlP9P/gsKUb0y25rOwpwob3ti5NJ
8sRCr6tpUn0LpQjsSi0anSbaUSa4qqkXbgEQl1kKQNGPWqTTmPIpyR20k/zUOMa6ZWZw8GNdctrg
AyeAmIIN5HZML3+XlP4IuM9sN3bN5y1Y8znmJ0C7UQxv5E2r6Il6i7g+Om4tCLFou/Lclq/mwFOz
l4oDgeT0DrrLfBBTPEfvWFiOnNNEVeFuxOlFRx6KU/SsATY8zx45O5mr19hnsrM0nOV76HAiYEnE
Pl8rzkxNQrpx224PI9qnDEHG+YjYH3LvRdqHIR1RW8dtgJhB5DNZSulcw53WCtJC91GIRKmrKaTM
qgsem5SLaUNfJiWLT/aT4K1/7JLsSChnBwI8aRTP6H1RhapqyGhdKJIM6ZleJsd8+kivtRmMDgBX
j1XBFNnRkeo1DxB9s8AkHna2zTNe30Y5aPBi/Nzq7ewkxbk6sMDwT73Gs2dRiLuiJlSxb84Re+gS
Qk0GKkisvE+KATUjIMX3qejiBwBj8e2/HtBXvx/k2z3bixxr2MumKvZUFn6wf50kXpbmZMDp8yMr
kL4S0L4ABAAX03pSPhBYFrFnVP9u1wB9z+rHK4xOrpsykjCvS1UxbiaZZQ9UOAm9qxpZuFcHkI+Y
i4XKTr1ytm7wI6vRC2T0bPCdek6vt+6Ps3N21+56rLZ2cZ+JcR+pZxe+ycY7CzUziQq4RpJ/oaet
kLLbnPGFJ0o/d47Fv3iRs05F/xmIddOesHPuN9k56XxK76md/X2fMkkrdotpaRHuM9QadQmBHiuK
nGpk306P5loNR4XI2v7HksYVrv2HdcWPlSoKNivZG6spPPJ7dsv70S0tkKGwNn3QyO+KygJxrqw/
iF3qJnkb36yE6HlQI/fdOe5+hEBFQnSsdZCHPL9clCTDgU9Xw50F9+YYw+A50JSmK6ocJqeD0pFx
mDfUct0TzwIZzwpjqkSc60uRJkS14+7edDdWWmaYTJz2HoGfK7xt5zUpy/mtgcErMj5xD8uG37XX
AS7pEX3xOl+X0k2TplWoJnQbNxFn10PrbNV1HRjJxTVoIWmxX4qKmqHUTHonYY3JFRaBjfUFUyz6
EL+dUP0N5S5H0zJTWw3EKr9Gjn1uP6j+vUrsHCjDBbvhUX20WJPLFPD3lKWTMHAbM+TysQdiHOsU
vbW/0i9leb+zqs2Q2YffvUtyuZz5sIhPf1pR+hQ9ep4RDgUniedzgMk9z+XPSCqHpUxKcZ+o0U9y
JeXcXQOry8IWtn1NESwyePR01BLAaXkkagyoMRwAvwAqyEDvCKgMnn1p2GaxkLa04AWmo3DOzibu
pRQbFx8Jx0B3qQh7+hjZIMPiMN8XUVFUGLRdLYy2en7OKmwEqeZQE3FyA+6r93RAk/nGJPbZXggw
GdHJLCbfqAoka/MVEO7Q4VsMgbMgKlQkiuEJBZqtP815EqwPMgATct71QvXGS1MQ0H4sgRFrympE
u74dJsw4kNkTdcGTBF6zSUrgijAHHngZ1/jJ4LjUeU2B4B6/Q8eNn6FNSJk/9MB8oktOSpYVAUO3
dfhuP+zD1oXoTtRS4JyllVh7fDh7uoobhxRaEiy/F0ywttSMLwTxYHueEBbja+JPy+0JP7M3XDRc
VplcdY/IexYajQ0B+veacN8hdg8krhYmgntcxmJzN1p3PLwN+5QQ1drDkw7z7h8it0/7RnZaUixt
jwtUNuqHB5PgbS3O9btkQA4iA3rC1h0TLDrXcmced4YezZ9eDNz/gj3qZieIuszh0i+CS1A7u7vz
jrFtoEErXnK/KThVNtOyDmJ3JHBt6PzWuW8WU3QjlCkpLJnC4JXJ1HLI0U0VrTm0slHGPl7MFG7Z
ktVhe5I853jGtRjcZQyS/4xLE8iyx6PMVc+2VFyk6GPTRyMvL1dsC1zKLu8QtTHga5TR8k+6C2R3
4yrVoYGGycWB9VUoRHxUexZyKJo4AKq74I15EqHnDkSH+tgc/8COS6FkIjHF4g2zgeLbwUU/SrHq
OSx5enou0kCSeUusSQFxvvxc0xEtLOQiO94XnpWcutcd++HmJWo112AFgz3lCdqTYRZ47Y0MERvY
HHrmNejyLwGF+FCwFLb4ek/e2TiWSfv8hJ/J+UIL549nN5SrNEUHsn/lqxOz3hkYZ8iF2ZVhG6Hu
GAx94RhRCZLOhRDaiYhSyyin4BULxB07OilQYy3Jv0dV/nnSRCFKlI1Q13vrdTbcgIbx/Shz+EY+
OksTa319dMnum5z9pTg/f9V4KVQ7oGDkoDPUL8Q6YN9u+hDAtyQWg13ytdBjAmbyl6vVVYEDp4Rm
uswOylELOuvLeor+gqfxFww2rDZ4iIsqzH6JPO0/5T02F1BuEauyI4/KBatNeMAP4Lhr9HNsYHm/
Qz+dSzidTC2WGwTygD0suBjjBc/9hrYdI1dvPE5G4ks0ccASvMTE31XxFqxRvDlEEBYwBMyAEmiu
3xkP6PYYWfFcjDXsrHYwuyX5Exh81EwRhG1QyYwcybV0znrTWt29M7nE2nW+jzPRSGX6HX90qI+0
Fn0BchuGs0MrZQcQ++T7btOT8zt88iWFGh72Cw8CEdEwqW4n1TrvSmIPDEv8fok3SVg4+UnTPczZ
vXqd5+8DtZr0XEIGHa9/fGRs9YA+47hFA29r/XrZgXyqTfo16XtSAXqGGnDG+idXh5ve/UX3vVq0
8DwOXOe6wdUGWE/njJYobjWqEK5j/EgLfr/n/WZT+qJfgIJ7SwNmWYcjrQffiXEow47UmtIHunzd
29fyHxkfrB0HMde2CvRW47Ruq1noTkW/rMFifp2Q6Pis9lOHA+xysA/I46EmeoSHwgS3XJk188KD
o1yPwkACc9OND4k7A8GBKVocxtcKW7YQZF/2QM+12gq8K1hS/pCUF65XV5xE7uLLVUFipDAoSudj
nUuAe+ufbwvR1Ov53fC5Zp/mLiOemjjLEpke6aBVigoVQAqfsIBxM/RULFKjKRxDipWN1qpSpQK5
wC+h3J+VQEOnVi9pI2+jzutCL2Nv3SQatNhU+edm8b3PQk337fPfjjYVyvvY7RbIkI8kHrVdmovK
GsmXGx7TuX/2rW7cYJrVQ52jhcq5Ln2EHuUKyALTlTXHmAibVTHMsziT3CYQruY+kyPJa1SGMCtN
r6/99G0MyotYiAIKyDozciQTQCQhcqyrkUb0LJ72NsoowGZjV1CvKaxOavk/3qkDL6xWpM7hQuin
l9iQw4JVOT2AqfHEeIHgjZK8vJE3r0FleLpORyqg62bWfgoCTncfeYt81bLTJt68dS8i5VB4pqEb
RvvtRF2zzAtHfTrF05TPO4f56M138QwuG6Kb9hx3+qiQOw5GQBBKsG83541M2Cb52MGYrD0qBqd6
8pZfs3udlRx/kFpznjHMXjsOo8gTrL16189+kT56eQjwuIeBrKCoGsKxw4/GwSpQ8KOSBt2xAl6w
5SvKdihV9JVw5MwMtz6qL5nWfNpU8HxSow5s2ifpp7ZS3NSlpvblEjl7S0BeKUNiSAhO/EfVOSUB
rQGewoGA7kCkZ5qD3h0/BaxnEU6DbLApFycT3DyZsBlfz4lZ+pnW7DC+LhiaU8y6XYemtU676EOi
HrY4PriI1wjKRWyRctMJdBg0mmSrOh3rrIpt7RUkGJVGepyIxgi5dA0PG127sqDhjsXBLRs79lSO
xcbKeNdUdIjBHcUeyYrnyCpYMoHarXTpT6w9h4sgErk1yYIdtRFqh4KLTYyjOKvkef/ahTqe+IjK
UhwcQWx+qZ0sGu6OFj0RzClITPAaSoII4bhjzA==
`pragma protect end_protected
