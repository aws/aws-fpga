`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
neUIhZqZp+LplbPVVCNO72IPwEJjtV3I9aRgqKJNrANLD4arTN0ixDQdP/y9N8lqJ9vhPep+jTUJ
M7UsyDqbZxo8J1IRSIhFppEq6ThM+8szI79ZLj8xg/4tTuYoBnPQfW2yg6XMMECoDQYvAgBDYamT
baMIIq8TIeCow7F3nKdxm95vlWfidnGwpc1V75BoeES5s/zp3/CHiIyGY856dHq6gzVNGUzVhlY9
NGMMsY6M89ko6dmv8rpYb8qYU0D1ZqgDijhGZjsjg92iqcTwR6rvfBO4WpbRQtme+iK5Ks0PzRQC
XhIEAit21Ordh+O9QCKxxlPR7oJ2A4pZQ5dzUg==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
DJXKCL5wZhdj5E5WknL3LpdU9sk2QG9PAOdCsihOwWEahMzZSsxDL7BN/USz3jqJipZxLatJnLJD
7ksMgrMp1S6gopRPxm9UTcZR0omv0hcX/G80cnhOss/bR+dAJTMM0DxnJC7TU9dtDffMm4BbLQnb
Cqy2ZeX7mCC+b8U5fTk=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
hoW0x4nv5zPyv6I80P1ONoMjBsCBdQvJ4X68ovBAYK56BC3ZriQOsrBbi2dFP3T6NJfics+gkkD2
yiMA0wBydA8cYNL2K5lxFWHhJ4mK2k8QZ2EYcRKpzL3pgX9dWmiyHe3pQu4f3Zrf7rjgOWKJalyJ
S9W+UMu0SwBALB/XwjY=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 17568)
`pragma protect data_block
bj+prNInKSUYsz1WB2pq592dNw+5+uiJCYazjLPjcP4SOrDW9MciDkTQ0vogWXUoqj9E/maEDWh+
lvVpoSw+tN1tGBT3eJzFdVRWw1ZdjL25Y6kRembEZkdkZjaWMw9aQo4AkZPaORmgSaaLpfNf6ezR
SmxFPylEW3I6cZLBBz/fh6mUBxHbXi0zgi2HC8Ra0UfTBw9BaBThDIYle+daogjle9HosgMk6fSQ
yBsj5XO40ozBOMrOB8Mu4KmzsxT6R4O6re40NMmtAAphGtzA9TqCqMJHhvIHmLC5b4iCCu7KSWso
KTJ/v8E0/Y2kIkncRthdQY6kUN0kJ3gjn2LVJYGt7ec9a8NiQQh4Xttuf9JrpW2ExyvT+v++ziBA
KIcuS7XUMDnIvItK4Zq1sz3EiN9T0T0MNPlb2SMNOqHdDwlUBRK4rovJZKXh2jou5gh6Zi8a7iZQ
0zS9nhDKEf7+d6Os/nGx6jFvG0Ijk2Pe/WDmNAboYEuqn+lMSsDkUcQDFPhdtCefX0h2IEbfYrGx
vuKQpfWd6zIQZKiI+tDL0VpXUzdDIw8Siqihb3eQyXPJaXfEiYJ1amT6Dcp0TWVGCXZCrhW9KY1T
+19lnsVA9Dr87I7+TH9IobrjDpSh/f11m6CWTM3b7WB/8sq0v7Euft9JmHSQ/a/Jc444EknlxmbM
6G5tbEb6myGvaYnzoLFns59DoDCIXVYyeeJr9VoGcmBcwXQ+F6GgImaG1UTILCna+aKEJoDWPTvl
SfBdoXQ0PqBOfhZDoGg4rrTWEsJWJZhcmTFz/yUpTho+l+HA8If610oSr8U7LDPlxQcKuloaM49D
EbA4+xSGn3MXEAF/xdN4lAJihNwlPoYxm0PNi/7UcZvE96zGQ+eLHzC6RLtb43xVgkClYJcQJEJa
btN7GL40ZrSA0Zlgtmoky+OchHT2UDR9n0vjGOsJmf1sgCN5ldIOkssNldAzfE+OFVoWaF6LcdXg
jqINbOgYXjC/BBD4/YjMlv3ix4m1Ea0p+csSd4VkmCEmU3UEyS7r2USdk+6vGbxPFwx35fwM/sH8
uxF3wsrIIQn5gCDqXALhLHq4vjk/CmT0o2hNyGGwjYLs2bsIrdRz6cvfA2EKq2vSuzUWCI0p9CV1
0oPH1Qcv6OG6ZMzHkBk0l+7J1DpVFdhfwc3jYc1xMyCOx3aTD3X1U/3Iqkulsmjmy63HgF7x0PZ/
ldcH/+uEEa4uronmkisLgWvW8MHc7nflPmb7ehO0mm5P9MElZrTQuFEmljkBaczzGQnTtMUCh2nI
9N8pBIsdW5B817nP/2G2MXdPm/Ln5S0oEF0+/TkN+uPkBrxJxvwOLBdjm47ldCq5xwsjaC7v+2lO
Z+74O2T3lEryb/2GQ0hjH8KQOQVZB8c255eFKqSui4Bwto0Jp+Ck6Gym5cpso1Ew4nBLuJiBYEo0
1VQevJ8HcJaQthHNx5vV60NWCw2+oFWEH0HTuZu+SStsaxCXJykDnWWXV8GhM83DEf/edvCAAynN
kPcryVnDYnJCzZOyomgEx6vU0vzlFEu6nvZ7k61gcAN55Z9Sdd7TkRJqzfOds8iH4nK3IIpzNP1r
yYHfME1+sfl62oLAYx4EovJSMRD8maT9Bc4XPQTNiW46I+Ae8vNQ2KKhoKI3RZyPUS3S3VC+7gPY
eRQNoVpfCxF+5xhYTAZFKeXvt7LqMl/lesTNaS1Tj08sHt5yhawC1FwsJ+T8+6NrPeOpysN6ZwXe
z3Lip59lNRKpf+ip0sX9rgMVCvRU+r68Y85459ukV7zG3ZrIDrbC7pIp8ofW9LJDHTxJyZ8S6ACG
3dpr+ICIcagYDJkp/jDnF0m23VkIex9xylRLvfj2Z68Bq7IH4o/LZtfGPZT4zYzTlxwc5lfhwIfl
t9ZsR/5Mn6tsiDepOAGNRbK3XPhlQTEsYZKi6T3zZ11Ugk5uQ1TiH/e7J6PEA5iVaMqKCLvrSeSJ
vEIl1rzVWqAr2RqAFqIFIejhNcI8yPeQLq1VjCdkkJHhlReTWsT2oiTpkp1UXlEEA9Gn1pSLTWcj
2qiGORc4oWNPcJCtRG83eoAFL7qr+PW9QZgnvgcexkVCjCLmO9AVa8s3rMUSp+JpsGeZAdCkhiwa
IPwL2cJfWgrAx8oUaZXYCRHHBKPyEhrtVMFjg4jQ5qBgo97gFL9rMTdqlGXWB/bPuiy/5q1lEc/t
lkw3xG66RsQZpdKZfowVRPIJdCNpRtp5UNPkQLAsR2wn66FOKR0b3AwCbegeIj0EqWA39XFihIWi
o+ezJn4qtrtUQ3ebdEA3GRrQQ17qbs8fqidz5vczBlVskyC0TJAIM5LGU8VmBYkeXi3JVW3MpdlB
v4zg2WqGoREefsrWs6f2f8l1ppXuor0+q6Fb0RqSkjDHehjKfpafl8EdrnrAYleZt7He7TeaOnFp
624v/lkwTfYlmY5mos3Y9VSOBTZb5pVD1/T8FfA7mPWJGBDGoKBuu1zJFxrRLMGP/9Fw2gWUA3kw
MZ06LKOJSTErIBPyhXQ/D3DBStffL4QmlX2q48vZa+GCEv7DbRjpmarMX+jQG/Fs8/fG88LCGfHe
wP4rl5GL92nnMINZeRGuCk88j62VEz4hia6GyEe/OdUqiBNPWveGYZIgl8YRA1X3zF/10xGghkkr
5Z812dBZ2wwUm2ERCx65HfQ/F7wTrKP2QMSjXAEzSYPgo8hBL50OofkdJiQeZ1meaFvKxhQqobCJ
9YrJVb02/RiEny9Dz0ZNWUG2EzwXPTUOGPpCWcHRRDMXJ9uJ2stPTN61LsDcox/WjvVetI81PL8k
vHIOyeKFozyY50/1YLER9I8yzzTyRyAZYGDwyMsTEjnmzWMnTEsXi/eiKwguEya5coAPuOz3ggpY
pWZjiTFZzxOuuUAhiMyFdPMlJXXos7/YEgsDbgber6SNBQkUtsjf9RnqlRZhgruyu1RzkwWCwKmu
WOPlagDww6P5JqTsnpMn5bqNv5GqRRw/5j5kBJJgaAbESlPGcEyjTFryhaMDdtFfWAmeCRuBDpE/
bGDpzXAweyIihBy+mERXAMOPwOj4EBDrm3+Tw+ki43x2ca/IQTMwu9JIutY70z5pmIMGtevjFtAK
tSDUGEy+ETwfiq4VB2jCRErc8echpj5xP8f7nn9zTuWi+EDLLN7OWLs2P3fJCQh8P3RYPHxgO90B
v+cwu3OaGINvtqFhx/b7ttkXQ0FufLK4jgVF1e/K4Db0/sdYm8+h6RRfl5MASArpFB++OVzThIbr
i146L6X+9rDAsc4bW/pj13AegUmb96vvzzscfCRPqPyAsWL9XHHB5JQFtMIXrk3JYKUpEjtmzzp1
VqeKgrA8M3QDOiIAoZYplxp5OhfAzOUHCnoF7ZxEi8gQAczyHyYxfdho68p4Aetji3v1iQS2Mgad
0Jc2xbNi4MYujb4KZXmMcBPwQNO26JrUlIj5/VYOm/KulM4IprTYDnzTrirmzMERMnJhcuBaj+hD
6lXPKvbZYHhy6hZh839psWFscVTcvKO2apoOGWsCJDLdxG+FH0PrAGyZO1frLvtUdsrmdvwEDfLg
k3DgFr7kdk6ilOv6qvqjYQTTwOrcY4MkLuaoevbA04Wo9rs08GhHOJGvjiBQA0TnCvMwzTasqr0U
GNDjKHdYzH+zTdfLKF/x9kFfKaIvJ4+UmVXjPOLPkEg0Di2vezLJ8MA9QwCzt4PxU6I5MgHas/xb
s+qcKtANaCcy+xI/I6qoAvhWY2Ci+icF/L+4U0wK91i8mCBYjT5XCqZNftXPai5luUuzlLzWTNaA
FPciqm6gZqEEacw0/Xh0NDoIX8xw8GQ/AnaWjL6FbMrOexbzhYypZ4qR9GrnLNo/wMQYNg7wTU7g
IE/iB5JxS9luia0a5y3bI7boUxn7XC7Uhl45WBdZeeiCdK2YvQkYJ6t/STRYNmt8u822OhqQnjfn
+jSkVENX9Bi+uBA7cjBovqXa/PTBHntvUoN2N+WTehsCJ08ztv28gQKZdK6fRI2IhCqj9JEbOPjk
2cul8iEtQ5WMWWuvYhBeuJ6o3kIpm7aId42bA3Q2zC5M4nvD7VfBnCShW6R8xVaBXjElcruuuBsY
mLPMa4rTIMPsIcBoxHQUrYUzOau4UaImd91SyyobtVDMUBDGFT+zyrVs7koieU4XQVdVQJ6SPJeU
H4tc/8z0mW1/1NAfme0OF9mCHxX+lF/RmccDuEHVAycOoZeojSYwbF9RkJoYINNituFFTiHpMtop
4eBVM4VNf7KBkkIz6gPkxATsHsHSw3nxP5qxPFh8hydD5dxvUD9i00dLoWCkC5q/USUZZaS74W2W
JEdU8tDwwbMgTvWXfvvAat/cuNcwiimXtRXeIFFXnoCJT0Ru3EBs+vgsx9H/KRSOQW/R9QFnFd14
ZFA1DoiGlSy2RwEEvrySJ1k4N0AA75qPBnT4V/fhegxXfv+UZtbqvIY0xfDA/0DC20b4bdSUUiSS
n80Qnls30R5icnlJBaNwTPZ9tGPyXsfWyuILigWsylDd7kzPNTyUt+9ggbg59AfBQEvSt7S6HQc4
LwViQFn23C6SCFf0LbAD7TXh+xlrPr7vnebkgciQ4mQOfv8HnNr2tfe8DjdeSLmglFoRaMRNEAtl
a3CDkaIeZHxGM7DQvWQzZkN7S5aYrGyHQ+2RIHIeFrmrtP+izhITamA5AEMmK0kv66z6Mw0LbrEP
R2VhvPMCPPgBiwyyZUL54rKqu4+zZkLud4BnwsbpELDaDcBzLnAn2+7Zm0in/S9Qpwgis+IK3A7N
6Vjv8AWwhPy7OFlNHdPvcT2M3TBGKzcG/8Rax8SshSi4MqATA0l5/oFggtqcl65crqoN0Obn9IPh
uz+13TIa8U6y58gNN9q+ZWv7UQ75jY9F0PPJC5VVlaLnr9t0MgzsA3VgIdVGFUKrS8TjXuF/VnFE
2qziwwjraqVgkX418dzXKMJknPPx9sXkPFeQMxkQP0+wIqBwZomSGSh9PcbGgHSn/mdUji6gvURa
ly5P0wcmg6u7yRQ2V9JEItArQ2SyXLjSTxEul5WVGo1QbCzdaf6e8ZmyFLaLNkBe4yFBd2bzVMv2
D+etOMspdEwCsdmwpK+uU1o7Ns0dRwSp84OgHB7WQpk29EHaJLpBVJ7jwN10UsVj5MpsqH+mlYel
MJ40Qss2tGJTTlwnheewlhzpHSzhdTMicy8DECkvWgCxvRzLnsBAx2k3wgpbdfuiVw6hQhaFArHE
Pq694d2W4mPtu7GrLCL1ISrMK1neNwJYxCc+9XtCHJ+07q6PqMj8LX7W+20fyhL4tqgPzDHUp4Vl
i27nBS/WH3QlzV1MuUSHCF85trbHKa8yMNBWOHlKyibwTgH7uDEdUxSDetq+4v7o+8vpob+QcKgr
/0m0VjyutxJ1jT0yiNZQ3QufhjCXvXWExZbOGzIwtDzNFPmpziaqjZ44GLzAKqo4PwbYMzkDAwJ7
qZMnQWVRvPo5H5T/CA24d9JDc1lyaGOxvzRpo6JEKyQ5SoU2OzgoQEWIYjz8r9IHPZWFzed4g6+s
q5QIBlBWJAuyBFajOtnST6rIMVZ4a3ph93vlaq2kJI+QvA040tSByYXIQwOeuKj/HKS42CPu+P/1
ts74Ehqt3Smvte9vXi1EpXGY0PDR7AIaOjDolhSNnm/+bE3QnC6iVDmHzPFxts0rsrmI98R6HHAs
+cbVUOa03GBKMkBVVxj7rP5RlddamEKTZMSD1VEHNbvgny3QKvcoS0geaU+x5IFeyZXWVQfQriut
+j6U46Fo+KzCrgWcTM+f4jPjEOKL79xKU8aA1xyVszz6pXNW/fbWH/8oyUKAPvQKEuLS1KYxb8Is
giWwiapJaivrGpR9awps+uvNovnyy9EV1bv/73A69XaQGAe1k6UdWJ2viaRWY6YQzLavPCqDGwwq
VvrkAnsiZW+hQC0IhLigweDrSN5jixTtTgGzAcC0cSmv0N+MNJpjVhTgbWVKvd2ky+STpr2/1RPU
O/88whj6HmheHy//XgScRLG1wrhveIDTwYcJN46Pu7KhSKqu5aLTHn18Js/+L0qo1WnMXp0FYJdb
g8fcOsV1N63/uJdwwrMb7QxNQcUC7GQnKCW9684B4R7mpq2AqkTyfVuS3368Lj3DUGcks+ICz/+3
FSppLhq2fpu3iRzbJ8svEmozL1apbigNXJ77yFaWUcJGD4EyqPjhZw7fsOnKYSaKtK3GJppKj/y+
hlEjjD2SCqf89Ysu5SCkleHPATu+C6DrL2fQUUeWa8pLxMTlRSKJo0vKgbBgqIogpplEGa0b830C
1EbMMoTSMt6vtviw/wsh+exf+xjcknFbLxIBWdgwpBaD4wLNODOabEisVAxnzmkfdLKgQ6I0mBpC
cvBVfnmcMgiiYiFrAvEa2qSq9bdLSMdVV2VqOtTuGzYq8ljvSYV94tdMjgL/l4M5O9cIvzv74YrK
07QFWq+/flGyzWWL7pd6a3/ax/ZdiN1Bfo20Hpdvo7dcy7gNvQ6JdthuxBV9VbM27q3RYvwCrlU9
OYrGeAS+W2qyliSiFWvApin6/nhlqXNojKfGpcGO7MYxgmExiJZ8j45r243FPE+7ZMrfoW1il2wY
K6ZSSn/dHOw3zqt/XBitl1puIPvhPggFcQNjhSFC97maGG3kmrg/dfLl+f4mKD9+OxQceJjQ7mfb
TtLnsd9sMcPn8+kG66pncjRHKHU5KYH7dxzIIiG8QQ3QOoaHe+tUZrarynvGJJQzK88EtdcGCBsO
14beIISeQQ4lpgkklZbn8hw/aKWrG9rZiW+MKypjGNtiLIRs1WfVVQ+zLz3hGAIRBJ0uKCyD0mC8
o4z+I7k8NpLB0nE7aEF/2EOCpxnmkvGZpkCKKbcBHH/9t9YjbZYjHc03bCtmEndFKUbYrdePdj5y
Re4LbeSDq6m6LjQtFtLPml8ZSskaLsWcyHCi0DlTjgXVPJ15k8czn/aCAZBFoDtp90lReowMNgCk
XaSLaosDoJ/9jcV1qiwfuEDzTO6EVKCDvOqouFUox9IhTBp5auYCEOHJUh7ELSrnsqdUruAOz4Bn
DvmOTt2Bhi9G28iOPEzDULxCrpg+iU5v1402CoqwNNjrT0Zy/3bf1fQtDeZ0Tbf4ieprNFN+wb0L
rxNGYLX4ac1wM6dtKoRLcBRgZP8aUHTPvJCPHYO1JdHKz/pKRY5GFsDEpTVhL4afcSf7P11uyRVk
2z3AcJ47TA21lh8IdPOTOUhED4Ks0z38D4IkaPVucJAZ7LEU6OgsC6KYQlsp5bX1u2L5ZfRWkVAb
HNZ60cwAbXvNleM2kSoRmgadHLn4CHooXYPWyFnHXvRxO5fDYvlEssq0mLvE+Y6wvnp4mvU3GTfH
yHFaA8Y5D8EBywi+yi/3X5Unmxe9OxYH1fvoEHn0U8lOwboBBNetbOXmSqxW/+RqKPpjgUK/3BjH
cFZOD3EdW0NXXtVUJlUdqfkOvYf0pPL1cmRTuzc3KJpyKqbhsHxpw9nXafofbbKod8prnwsrirwz
o6Uw0f1r2HykmxgC0y4FbSCtJHC1zMHv08G9L+FWgmgRfI5npfmOIg04uYSNf40geU04/2WWxV1H
+pZbtDEC3VnJJcgRIGyQvMVQWgEDGKoNfNB/Bc9sTKP8PGiDZwZzgkbbkKwfK93olFH1cVMruTt5
mCEAt3aq0AvcwwRFCTD5w4ZTdy5w2gBM/fvV4/GrqxBpOFQxzll/n4dPeTGVsdQG4n9NjO8t76K6
7MlQDsbK5rmmoRyP2ksaWKiDrfSJFcbtF3MG2hXc6MXAs8WSXAWtoYa3hVc17SnYMtlaQMMhs/g1
vBIIp3wyTAEuvZs5twOahc8iq/v8zulLqK8aHEx6ofd5BTLmr7v4JGZU9cMXdlCyxVaAB1quvHmT
2jspvtui0MQYpS0mtXGX4EuVwuuZZcRPkqyhm+r9VhCa6J7av03OAd6GymvZEWr04I/CrdYAi53Q
IYYVJ69OT9qlr/sDRohh8faMAHdeGYBgZWFRld5ojF4mdGHLunjXtYmaiFowftvUFt1dQ7ovNMMJ
mo1giUdbWe2fBwDGk42um3gIIQHC0K/l0LlVxXHHATFydC6KiFAGoujsE+ffBAPvT2P9zLIM59xo
yRk1pNlbORWnTf6Jv9ZhIUlUE0pkvR5nJFyF/JfrWsdcFFDBf6YF1Qp2gWCe9ccCfm4+asiXSDHp
oqQiGijBLO/cLUMHgtRX2YZu2fsWMXuQ3U6e5w274ukkmicUsGH1ZDbB8Qy5Bg1V1g82s1jNa/sz
+YIB5L428R0LcvC0mJjybThB00euLURLwLfiDMHG28csLOcdcuvNeOuTKFrg6fmCRqkTR6fgoupS
konqlLWG5yduHWF5NIvPr4UuNdBtRlWME2bL2jEr8FCtp7o3wdvvawkzoMOqqO8BbbNzhSfa0w48
Rj+U7i/ZxA1Mq+W2VKzCzBEbq3Uwf0J1xBEEZ9F+0+ei9nxsrLUNOd+otaDdVZ4k4OMwctNdtTlZ
H5lbfmlb7Da9Crq0ZTd3w5BOfkXs7I305QGlbUp8iS1eL7/mgNGoohDUa9wQTtbyF1SHLfgTEUG/
f+Grs1+eVoSqnv4DBlqqnnYK1qIMaS/tGg0/0ld6xfqlxhi97otKL5+OxIxIZFkATSEDrsuK6CW2
E7o/YbeBMYyROzMKeS5nZGfQi3t3Qd1wItyV9UTp6niLh6EANZ/bjOiYhRH8h1WBYTN1Q5p3qAuf
LImR7Un7zH+XhfgbxFeYmkCq5rx/ubNwspghwnhCWfjPp2LyjeHYG7WOct7UPu5YRw4S/v8husHJ
NffRGnpj8Un+5h1r/RwV25JUEyk3JdqJMO9VKQi9eYW29Rj6JCSKwUsE7gr8FNJQCE1v+6ocTeEH
6blT4S8Q8kFb77JD93VLOze8ZLEBIprs8lZk3I/9HoQgJpE3vNEyz9E7DU2ynPb8hGD/g4hi2iTs
v3Ns/oq+lS/nrRPDn8OMHzInTsSww2IUhNoY3wUwGWp1a2tvHEY8n+kssaqJNwr17JkxFiz82qee
IvgOQ1oU+4DbzuvZZZNML/++qVEfYLBkYedOzIklbsSTRpi0xjVA22FjzOdC05vTrtlpX7pdAZCk
kuG8HfApojRQ/E4QCLYmfEMUmREcn75ZnLVrTpLuBQGwNweSLpMhJlWAdmOTBY3W7ENf2ppZAJRm
mZSbv1eCUsV6YniJ6xPD6wuMxkPwTDgGU9riQ9gzLxSoRsgL3kFaI+nf5synzhlQYu9hWr8F5Wwq
y+5PWX9rcnI/OcW6ZmlXcv9Hn0O4uB3OKwATptduPDav4KfaIfLAUH4ZpqEGdPkYTciZW+V5qgW+
ECZOWesQiQ61nojULP4aNBxDJ9f/+XISI+PVTcNeWlz1HAECeYJAVljquNJLXsZZovmRIbkvplw+
UX1vXTXGXPGGVBL7qtvg4pJX9gmIvePtFGixn2ok97XyM6MelO2bm+a9BFS8abadV5GkNrKbpDw5
yL2WkGRpQ45xdD4J4XIwOETUQgq1oKmUxpxYQOB3fomBMj1C9TGwilGOoNdh/ZLFJxAiq14P234X
Pino5fwDeU61cuaktfsqpiRlSi5MVGSb7IsBTVgU5/PIS6NK8sTeK4SyhNlYk4smkXdn19TVoW9a
JWQv+f3FhEKTOcSdEBnjvnETX9qPCS7+VyUBROeDa53hc7HnkecvElzYfuKWyWJZxSj+FAupAeWu
rYJPYFA2uTPqDApeQoNFUIQtZpPNqzbNoC5cS5AnsOa5TBczisDkhzQBFge5grlZuKLdq4wkl7da
XxOssUXAbznuPEF4kKXtd4YK/oyeq42ioU8pZ0/B8g52CPMWBUk29xOgUeLTKuFIULGALroSIPXR
4vAq1gfMM1HJn8vElW9YNxQMY8tOFmWPoB4XNKW52sOLlP4czpZBFfP/9FpbFCY7vYFEGNysHE+V
DBKb2bpSIU1uD+vOlPDYj0V3ESB9gf6h2A6r4CiuHB5ZtJBcGTlg+Kv/gHNQaCsQkbvLXymMpH+4
W2izmSkahrhbmGZqIzspE+pR2GVIwxhliORL0sKrm71OGXCTPlTI0YZcPRbkmvfbekhQ5v1J8HVu
6Yju2W8fvWniTH1+L6cgLKD/W17fVb6XZRIH4nWOi+b7MPA777qL71jdbJ6Qljzfc7VatJhxwVBe
EkGP21gm57qLvL0+4NAxvCcbCqDDIR1B7d1kARzL1fcw/WMgvw4N17CriCsZCUU2gLyn0O4t4Aor
pF3osqdd+Y0W/0li+BBWiPvjWmC1WvrgFHPsbDo5sYQ32vZv90omh0Awl3XIcnvl6NcFP4qgFPSI
3Ts0w70mC/LDFtxerBg8sw52nzpLhGxPemqk/PsfTmdHd21MRpmXZdQbgNdu7c6KjEIDbH7fFJnp
XoJGBxQjkCJ1+BnOyaErYP2sEcENdSKdXVRhWJj0o1YXwiCZteRvWMAoLq9bIbuxTnS44yzf/n44
qTeZDV9ueh3QCZfmiWPB8rFbhF7ZNfotvMkts9JJVuVBzriRsWicgZXCPGu9RuKmcc9Wj41UYgdj
EtZzYvSmRAIPumN8DuVAajtLgYUuNF+Vh4DyIojKE/wUHNRFnOl7FC+jq29y7/1DA66mEHxVbWQC
GbJh9MXI62MT2Exw9IqMbtoIaV30d6DDa83w1UVsBvY9nSm6vCLvmAeyMr3DJbi0zax2gIgcquCK
FIFT7jZixGB6r6KLTOngTb2O8xeoGq+DFHndrA7hqVVlSEv7IcoQQRj/SDu92CZYxcZhlUTLDeLQ
suGMORrIN2n1ViAvJbPq1bqYTnCPVgvVhCwPXE57CHF7g7REv1ceSyYckzZ1kX1DiFchvyfMprEq
i80dJTRZ/t9aV/GSmALhSkX6HsLMRzaMKvMykLRCzcZnjSV6a4skMQphHeS+fSbT+8OfB8iIO85f
r7auF2B2ug236je7+MLzurDT50jOmJPqqz7vNqoKdDt+o+0m92SQ/WsNtmgHRaA4ONcWPi6FtfOy
VmEMwgdPQoEwDYbEXrKx/ttgCbiqyVay7FhX5vOxEl5UDehdaYQMy9cfERMq32sRDJIYg0c4WtzS
1hsCIvdWIIPpIQYSwIiheIIFbf9yuubA0y/zGOFUk6ZPB9TifaUlWRDUfa77GkksT1uavyuTAjjl
wNllOcCt+7ZYl8BoPymo6orhesZmA65DlDcJE7Wpjz4AU4uRuaGdd1xyiZdntlHzVk3Pdaa4xEOS
qZiHTSuoGf0ifD3cU8+10sOcI4ej/EHfLGgyXUnZEXGbQ6xu+ej06l4VjgM5jEvVzXyAsaQHEHmi
Cerd3TJX/X5IQvMa6tdx14m8guLPkJ1GQrm9Y0WshkQxPhGRRF5MTYMF438uxgAgGpioyY38+BBC
U100yIsV6+92zTLW92WEi4nrAWrMUPboqfDqgoi1MOUtxIy2ia6yCR9gjFw9XUsQ3lUiPcQC7/TN
n5oopfhBVvoNGKZmgOKc191ZhgvsxWY3ViYhegK2UV+TCx3dattsyQ5+xDyMte3Ah01sHD6QDMAf
mG3LxbyH4AdMvOWGyOVc+DbZkRWG3qwyNlJCicFUU5K/oHMQC++lztt3BoLu+adgp9fCcLJvqlP1
yJUlcSYunf5aIl4i5XN6Ty1n8kg3bKRiNBtNKDDmIzHc/x7A905YgUAZL5tVfWyhO1oxFhZPuWec
G9pFBVJ+XpDNzUkxxuCthTfBb43s5nPdaSg/RMyTO1utM+FGt81dJOvDeXa+ov/VONzgqsgr/LZr
gNgzBB4Omm6tuQf+MJq0hK+v3QZsx6JRJOOdl9M8bToAUcDbVTm8u1Yuf0hgtpT7G1DyqRFH8qR7
c1HEqUURt0h2fCfwVIU8x/V3S9xBufbjk9zi2fs9Zj+nX5NPu/5PdpfGDFA99RfyYPgekBJ3MNEK
GspfkCcLV+Xy4zE93LPwdarm4bSIPIR1SqJl05ZrEXtmeo/fdxm9wKhyi1LgZPR382b6EBBYb2zI
8lnHRzpqnvAOCyCUBZ68xk/wNXzxjnHC15iNZubgsq+kAA3OMIwqjKvYdTuJcrV8i6AAk0rAz00I
aX3JLD1AnVs2Gn3LiU2P8bbhexRSYc8/1uhPUpBR1IYDwsuaFde8tKuAVZMcRPtPkqZTny+Hy9jD
qUcPxmOWCQGXJwPll5SnccRJddA9lP6ePA+Ax8m/37CXAmMROkwEPoOX0bmDBl25DmrXmAL9gXTL
kxZe6cMByC7YS8eWC2F+3nVYN6x3DGCviLFOHOeFF9DtNkc8g1qra2n6iM3QgchGvnMnePTDW2xC
49S8gaPbs9VqIvypyN/tz3t/ArlQDhynRyvqsnrMS8rZNiZCNLjlzIW50zT3U7eDMLWqKCQ9Tghp
Y+HPJSR2Wy0hcTlhOaCfIaEhSk9278SWXu8HWlsOykn8MIgs2vF4cQ2Q4vwabTveWihjkVEEcFeI
hQNQGximhlVcMXRU+zUcXxsaP6SX1uLg/jA2RkATKJSBLuJLKbMPLeTD6JbtU5MG5DHeRNANAsok
al8+BJfK/5jPn0UWisSCuoqd31k+t6WznqDPsPxkf8ricgcZyjQFg29u0LnduUZN37TTGaO9PF7c
8yTXV0ZY/Bb6f37XpWlO4BhxeFFj6DK4WSUw6PJeh2cRKHoRXE9x1DmyCudPxR8zbaOc0Pbd+VAq
4rCOQKyo8thlJk8RatLpqN95tQPjT5OSwmbaTXbW0ZIvyMYPx7JezbYFSzPY48VLbWVM1J9qtMl4
nimi0Y4X+//1WfViyWfMiAP58GZDDcZmM6KDOxbc1ysaPMct6HZ5wKJfHXs2Hc1AWYPivgB7zmVu
J1gfdjuFWkJDxyT/lpU/BRko8I6dFcdBpxaOcEfq+s7/lZP6jMtksNI/+gLra+JI1dP13hWo/x54
692/cbRejw3/rTSLeAMdtlDXsOjqmHmiNrgXyw9q7P7+XGfDryz244CjrIFWZnbWk0lIgKvpeoU2
sTE76Z+9QOecmBjepHOewQWgX5KiVBwJLN9uK0/lBCjy8c0wMcMmIC3vMYp9vrQtky1vpBihL7jS
AoIG9XbSUdt5UEoUdwFK23oWZQQs4zw4GVcEnk5KGP3nGdmrfrewxfTxoJmSuGNHGi1vj7NiGE7d
LDFU3yRdb9fPzmpAzDyl12xlu8UfgDWP+0sn1qFarFkfMUPWsHMRkZ3Nk+OFpmt37oEuvj/H3sel
SPnexlps0PjRm4aGApWM1cpqgkIn+s7BerLYyqsbA9jkpce5fngwQcwi/3C+MVEBfvfsu4Cbw+g5
auUbfXUhNiHjND3XIK1iAajVPhjwExfP81gnMb8a6c0QMngi5zvWfFrYsNsa4aRpxRhqCQc/gNv2
g7UgJ7YcoWsTwRmqe7gd/rJ+2gp76ov1N8CU8XR39fgf6taMUFaZA2PSLY5jRv2sXwaGM7dS1aoZ
6SqolIBfOnsHW2I3U6PvBkvoSIJ9mGqCF+KB7N+abeOnimNHzj969HRHR4AdvOG/iS6VzIr+EknQ
Le3JOxm0u5cpgcBckBfUVjoGgjNMIqSuXJu6uy1RRNpiIo7V+h3ygzWTNzAS0YP7KkIJLc1LXOSq
jgUFkJWK/z5/H184Yy3m4o2TQmxLg7X9nztl6823dvtuhy8b5TQbrnzw4mm2aYFMX0K7hCtvSojz
Aj0+SB9YjmtcGOGsqTU7GdNS6wU7n8FavcrzieOI+i6QUyTDi9Zq2Rf4XGKBg+6R9HVaFuUq6gTC
J8o4Kr3RrEGY5am0c2A5jcSELrocqTI0JUzasndi7mGLymp70IstF8W0vDd1Ln8rf6o8eHHShC/N
nmCsKTtgwZV9cXJBu7R5rWzCgWGMkhJIK571kRZ/qFZLj+x3ZSnzu6iC4wcH77XY+E0GuHpAHY/q
RWn+SHS1a8NVhnGA50hB6/2ABU9YSvtFT9UShc1qSmVwoZQP8kvmOV7GejtOikiPg8q6r7Xu8ZVb
MYKXAF+8BbeglTdXjp6gTT0AXvqL4/W51DHAeh5X/mXRicXbNQ9PraCNr2qr+4PKpg/D2nb1ul7c
6PsUytg6Y+IvyVLb1qLvf76f5vVTMiNSOrrO8V3SDoUr5CjzVT2GCLZleKUYd/WT223y0k0ajWxJ
4cRXXxEaCw/TTiDCmNgRYShTHAhn/24DMYthzLm+BfWGjahrYPUxL+ev02KgUmhBWus99NOnIP9C
+jDa0VrpMVyaZxCGgjcjATMbro+GxL1wSSOIodb1Cue3MYxEXOR7WGWxcVGbomRHwcOd0vQb0pUx
Q+I4jGPM8YP/2+ewRXmE38SRE2N+jUksTUUiND7/Xkf6tfVE5apOJh58+X8ChE9ZZ/ZiuyZlMEbh
T0mSvUTuMf0MpfkwCciqlmvsNXM58yUAnsURAQC+pkhzGOiJrqvq2e51dNDzSCwHaaxVBGIWaNwO
AEAtUobpQrUmEsYVwDg0vQyIad5SoVLp+LPZ/YuzKvns/4rKQC2FKWmHUf1QClR1dQUOquA8GVj5
nQ96rVLOf3+E4BqDAqMaM8ciBkKJKq1F6pWnbtzQe8j44M3FTMDjKlJzLZmCK0CwKYqyh8P/135l
hxvEBh00WPjEV5X/7bp4kGo6UP5i6mGCFLF2CIwz82mKnPkIUz77FU7VzMslsdanVNcNpQicxHA6
OblD8h7+HjrZ8v4J3O602AuLDILyeIps84vwIeWSvv68VhOzfQIt+FClmGSH1hdblTWb1l+z4ttg
upzBmpal3AI0dlDe7CSHs6IVgXUu2qzbych+9Tw1lKWh8SHpHZeCAYbKAiySXYTSVuT92yPVgnbH
Ubmq3bjHj3k7OnbWp+tSqujN6xeC/8C0Lk9EgS3ounH1m5kp9qlK5tqvqq+6M+UQoF3ylbwvPIMn
H1crjQ42ALpgIhfjlZ3N5jkvWNShrzUEjUuJ6vittqXCxFf7OUzVFHR1pOpztnoFB3QoEegB3XM7
XLPWlQ5OW39IY0Uj425ZYAXHmnlqwTV7ihmpBGE6UYZDKdQYp22g7a9b3gew+bFnFsWTLJqc87fb
uUL460F8N2WQuIEp9chVS1orSvmjOsXttSDtPGICrJqXBNTxz43URT5qD4safBEdC7xzf5Tp1tD6
gIjjgPocEo/0OExjzA+eChJGiyn4dy6sIlfH1ve1dWPV2+NO9/SCc+K1CNGOVV4fWD3uLvMQtAS4
iwwUjOKujCKh7+Z2w2PgzFCA5cKN+3M8v+CxYDaA2oWNbyBZVvyg1NvkcMle88Gtfid4wFCSUrUF
oF6QGVBmKNkwLjNNdelMFU0ZU91uPlCpJGiDCU51aRZsAfbjMBQgAfSN2A7CcV0xzEMgc39MwZsD
EvEyN/zQpuL8IRcVNgVArkUu5vM2eIAWg1/GOoNA2f2Q2E2QacoShNE97vdykYsdvpFJDEhNtStN
+h351qVTYSL4eHpTBonaas+mdLS+tKy5ADCJRyvnjIB7BoXSRyMmhC02psX50VuWj0raQCN7whrw
KvYelU37aW4coIZfF9bj3m9TMYTk/eIPh10bVnqzqEDoLhU9hFjH6/390Yy4JoJ6WZLwlZfifdC3
EsbmWt/Eoczdl7RgSxqsZIfNFzKEkUixws2dpt7yjGBmxn9AyZXZmBqwia+n9qd3uBZ/pw30MTMZ
/v+8dUhemqfjXir41tRdEb5igzKShnvehdNeoMRkm1NQ6PplJJCSdeHP93vbY+OMQOnnSc9IWwJ/
12OGApXfch9/o/RcZ71uXyPJFsGygxeLiBIE1gPLueAXQGWrCYiTriHgpGV50zhe9y4PL0v+70Iv
cj9DjyfPbYIxg/B45g2mE8tb6Sz+8J1F2TriHOY9HhY+sqAOj1MynYf85Yg445vHcZ+No0FBwVb8
YrpFSnoXly9+etdpmt22IsoDf8p7SrAx6es364OjaoodpMT1qfsFuDosXQPLeBnirKhoi26vx3Nh
kZ5EWoYvHWJKwNkQxXdT9jeHDjpAIuPw3+uApOqNehUoCmgNQH4gBRZBujf99Nba//7rvNtSBpdN
HR+UeSufSb9bDvLxqMjFSk6i7Kwi8CYufnSsXrNdSRgE4QQKm5yDRxkqiWItjNoYEBxoqzwxJj1z
5bklbjl0z9+dbojN+tFBBF/FtTdgMK2TaRs2kSakG7M+cUFGtCKpaP979fxPYNEPwMTBYIPvUTcz
gTuLCnmGBX4GDvzkJMV5CrU7mEYfVA956ahn9rhBEI11wAOyHjmpW89qcKnl+M6SVVtPnB3o2Mab
of4gv4V8H5Bht9ZwzoHXKG2YInzo2mcTtUyILNelkeEuEGlhNaNYcq2sPtRAUcF/0kN3N3MvtXr+
R2l/T3mMxwguQVj9S/EiP09H8w9ldJ/zjZ2fhctFdaVko0FDBZA33Zq1/uLTLoxWYWhkzanNAl6+
laxGP46/WFwD03Kpxt7sq1u8ma8MB7srE/yjmPBgDy5Ha9NTbXoOddp9bNWJadBKkT1B82JgaLVC
WoFvUCtNAVN3RLJ3zvgV4Vg0fEdJ7T7ezubbfLDt0Y93wTin/rd0u2nNqAYXVvhZypL9UZ0BpuhW
8MSu+FdZDAzan+u+rEncu24ypAtsXW6nui1fceyRmCJbN1OKQpQE/KI0RqweQ7rVj/ivDP8jt+Xd
Op3zPzXh9VrvgQmHET/YH0GKOuy0SunswB/tTBsA6AYKHvi3B5ABx3MWnoXnE06VEAXl+ehT84M3
AnQiII6p8BVgmUwTM5vZEWGhkXO6dzRpPa6h+GcX6YVgkwozKtx/Wd5X/Dl0Ndo532Zk1BwQPd5S
0i4PNxDIG5QZx9qApqZx7nlKgROQ5AeUMRBJMN42qcl3sWbjF9yOk3pTEbe+2QhBH4v3pKyMMci+
ESHv+HCtipztWfhaXawn18q8+mFSoWnO/qaGjlZb9Y+YteUnUbVrSvBruao5cNSylyqH2CwWr0t3
Wc5aJz44x7riBL/WCCSf6XRXcGBmvOfBtkkW/rA/pCxwPwm8WeMcwoTmAZAdvE/hBMZbRDRDqnHy
iJxEH3uae+Z37CFJ31yZoyXtF253ywK9Fl+UCNMzrYqvVoY5X+KxHLFa26bSe81X1DxOxwH1V7fo
Wnn1oOOBR/Vcu4Y2mqwauzQi3FsP41nXdxr6GSLAreXO2JUWSjw7/3fL7+7XiWB21f3Tw3dxiQL6
xUk3aC15xHFtGQmHM5yIfeIc2+XxDGUCjfJvhXkvHliKNgtR6HvN75sARqscCjz9VSWauBu77TX6
GohGQZOJLDjbjA7rmhzin9fbXVutSbxFgQZeSE+WYY1U3/vTJvvEZuEAQNNhrGF52Nxt8Uw+x6R0
rlrZjqWdIqhPDXXbeFvbYL1x9JqJp3IGZlTSvJPzyuQ6e4GHZsQ0FuuCilEsJiGia1CVcENs8TKF
ruNhZDJonJ//I1B5ijLYyga1+WGVAJ8e+EsFxgXSLzM0+v7VTZEnz6xT3SQHWyVfmSxeBrRMSsww
mGMK5eJLNd36lQiwHAco3Xg0hEfZpHalX3VyKc/+5925cPUlQqJdccY6M1/A4wl5oud7E1bi0Qmo
XeZAuW8OrFu/rMLCNVx5Y0Qr6vWmWFWCMuEBLAXoLyI+HaEZhz4/f/3LfjDtkOUPE/3+ZQ315s/P
89s/wJVnN6ErmDmlQ5cvw+eCoFg1gckGvPDVSVJ+b6B1Vb+hk0z0Eg6w6lQF/yj6Y5PMQcS+VjLh
YE8NTkCntLa1PTOryT0K8mXIx13EICO2Ib8j70buM6cV0PxoSf4NE6m96lNHA70oJvoR0YzObqrA
nbVOwb4Mry5wpphzohuGQInH94BypQRjW44rUVFq4jW9DMI5e0GTA0C1rvPoAlci9Ut0YuQ28FcF
JjRvZWLsFQn1IOQGe9Vu3EiX805IwbfTIxw+x/vd1F6x5OJ87xGLYI+G9hRVVw5bgAz56UpB3oNd
onMcD4SSs/iDxROhDC9Dw5lvK/FLn47jEjTlLLg8UqJasnA/twv5I8C2SV5MT3y3ZR9/eUEla95U
WPOMyDn1pSs/svyxKkjIkeGWQiuJPBpW5qNzxwsQ4vsCi+7EdFa6RyzFfQxfFG7pN6I1oXgis8gv
mSgBOsp6JoT/QRH0LmAew93amd+C10tqMThoV/G8dCB905I8lL6tZKyfukQy5mm5niACpMPOgL7h
oWabHq0Ut28ubugviHUFvl/P8ulqIhiFFrHKss+p7HT9/X4AIEUHwQGKHzaHF7cWxtHjPO7lpHlw
6WMJbnrljS3xwQNZCkpvdpCGHdjwEJoqZ8jr2p9dC6coTetajJ2kWkyPjW9ncF781XYVgFx0A16k
pHpHpYaN9tZ6/SLIAi+Fz5pnXMf22pCHy/akKkGl0LRrdxJYgwfsgZz3WU/1Wss334K+LwlUxVxl
6s1oUiRWLba1VbdG5foU33W4pva/nHa3Gwf8SnllNXL6fXFzyReEMbvm2JNgCv6nCwLhGS4qqmHh
fT3R4w9MkaZhk9AGPB5VtQfI7YEOCLtgxSwuxdnMlVjcExXdu+Tx6M1OWBlwdwLBCnQsVf8Fybvx
dCCjicxXcevRdauEptdL/dS8pDR4YLmsk5jfDLqr/C5XvRL78aZ+2eTxA3pN5LydRFueYBktSBO+
8Ij3DwW1eJw1FsPJDOsPj+L0UVfz0b4rgTMmVTxLZl7PcCjHqjT9Ta2x9W7Ev9odyw/OJ/nRqniw
NVYZKtzzhdqlROMvL7BpoOq0xD++tmKMNAkyU0MDCDyTt7ZCEmXUKX0k8RF1Dt/1vb1UUP5bKI7k
wT5QVn2B1X64oNYobTlTjErb/FOuddEaafyQpp6gTPIx6/VC+BpTgywX+VfyvBoTdC5b0VPMAlji
virRTWYfYYN8ZSgOzofPB7Q6BHayVD6FDwUNaOYvJMYaxfdV7kkhct/zPyA8IgFlux4BvkQku874
YLDbznZD6dlyj9NGKJ4UKKitATxVggNjzzJ8y5SMettFnusjO5dTYz2AgiyaPK9/mYBP7+KYxLEd
/qL12ceG6lhUuYh5CqTlFYI+JJPMb+iijvA1MDx4zHzVc4S7mfMaTizvfGjkZT4hratghzxfAPaX
rEWfD4dOzY99Xa26JCl1ebo3MgnoIDBJwwOtbq9pKavzW2L2GESwbVo3DDxQxBXp20DN2ZROHeAB
LZhK4YK2k3Q+wdLrNshwUhXdTtiRn0vywvAMIWV6kIQjPnhqoY41+a2LnfO4GXmSlqVwP2gs2+zh
rp0TMuyxONn9KOPxS80eF3z2rEzNY9I4yvMVuZyPRhx17xOD6Fi1DmQtxr7iJBPh3J3dtV2NlRgT
25o6wdkOkrG79cK4SnuMIp6QlrJhdZNFTg5LkWJLyz2bycLtzh0a6P9PA6yPKvO28E5fSrlGV+Et
6JDeQrY8fqSfAm1fLIgug8INmEoAL66Q1h2WLDaS3wKNjW2Yab03gJSmS1OTM9XQUEUXNzpLdMjw
iFN4oYnUYn5TotivLutBOTfIuCVohKJmG3mnOANpKiZupB1W7SCn2S0+A2T/L6/jt8+hzsuhUnYi
sgsfdWuQJ7qWQqqIGQgqxX3Q+RD2wKEYf5iFGDY2JyQNM7fORMowSFqm8WMWSryDLa/aZloUa8GX
YvKy44M4hD6xIky0ma9ERP6XHYyndf6ozmcQ5mPvaYUlg0uxVnOm3Qg2IBati4iH/XbQvaAN9alt
zmNgmU/rbWdOinHnMnPGwYMELJkAGhhCEMIFelB73FO1tTL/5Gy9yqrxGZKDbs5ZgFz95WkQ95w1
vY2LOmbbiplaAsjBYpQ4DnxEKml01eJ8FGn8++4xdDU23aWU/UxP/QcTWRy4xPPYVONeg3Y5CVOD
0/3tf8k8gfiC69jgP4VxcuiJ/UhsVN0oKVwWEJ82f3QcH8i2zsq/eq1XXoG9Ig6CjL/w1rmv/YCl
fbGC4AjCuoSMgmVoeiDEGb6NnwFQFj4YDpIDJyF6yjOZo33wIPV005/vwm9KWkhFxDUVeat19Bcq
IIYW1B/qWCQj6nnQGRCHI8cwwcuY+4v+PYDogw0bZma9kbf4gexdzA4mJ1oezH7PCHwsSE96u2IC
7VOf8afU/IQ9xa+0aNUZ6Bd7H7WWkVJuJpcPCMenIeged8Yl6Pdv6Kh9efzVOB05NOmyc9WK67QZ
TyNTJ/vQFpTW9Y/DUxIZvIBcITMlq+icLqmrZdi44ItUufrJR9DDD2snTEcBTld26WuYk3ss0w6d
aGLxW9kUI6SXxpyYFkB6ZCTmthNi0f10whLv37wVeUHBWObvM17fnGAvRq4lLaT+UdTKz4DUHbSw
5Mi8SEkps0tkVlES/IbAivf1D83hGrQtItdhI8CBPIYX0/iv/LPArcEqpBeSCAvYmmOLAnvNvA9k
O8I/sCvwQn+xnzovqgo5QyGpmxVN6pOclNusET51VjdjTZIlAj3fD7ankZdWIR079Jlfj7Gna3ng
ciken3XaEXqmqVZLwsnbQ8pXuQUwD49uIKA8O6vLTl25YAlRMiLR+x9LS2Mege8nL3/J9LydeT7G
pxPu7Fls31+3MVj4/DeWPTzypkMKyjsjUvV8SJXWn/USwBHV67nmjVKEVjwU1fXgeBDqAotqQaFt
JpQL449CTn61C2tW1uXWDTfU2DrmakIFlaQ5grgzdLMCveT9zxTKjsEeMvzCAffeZB6593D9/fp9
4zdJVOlwMUDSTAGZruM7UVMC7iEkmwX//BosmpjxoorL95sa3vMGlZTQl6Wxaj7r6fWChPIbu+xd
EIFuOSS0WZDqi7Oi2/9Bnh/HbHjz0wTpsdRO+6X2kuiF3jbTLzwMCAeQGHtuQckSZe354GgUKz2v
khFJnvEjw53INgisrAvo3h9MELyYEj0MwaarKVXNEQJ2aQl6KTvYGPqDIVOmevWBJ46Eo5xy8xAf
Dw/8cnTXQct4KSrO3EXCzZncAaGxSO+UjuXA9H498Cvss+m2w4o8Dz22DlLAQ22A+BQlivcKeM0H
t97OIzIxpxZEw/0NRJ7TKyk+ZkpSERT9+lbGLGLJYeRVwbNNBNsU1POmQAR6oRtMHxVx1Y0+B84N
6Co03Y0SChjpxqcr10rJRJNYugOR5Y624a087wnsYmoC+jiHYvi+O0/4iSiGGWBGuUhIZVai/Bct
wlIXIB6b1AQA9kjzTZSp3SUj1NxcCuq53EBZ3SNqJJRLSSL5eJjd72pYEoCPZprHBZWB3ee5G6Ze
rziyWtpHAK5iDGgI/4Qyt6CCawE+gnnWdZg/NgcTOSC8OdsvQHOkfgZs9JCt7nwxRjXBQbTru1aR
KKhW5pNzG2wLIT6IW6Kl13tSQw2s8v9Vnt782rOuIAulnpnmhPZObhxNmpGrVyIoLopZgodbmrZV
rCydQ+VMuqRWli4n5yVpwZ64+lQa/XOMJUTEZcJOaWRRg2KdKmOgOdB8JqXHB0y1t1Wl+sve1aQN
vkZkfIo7K/19anxT6yi1LhwtJiay6lt8doKzhLQK4sh1opfry6U197rJ1ZjS2Dl0lR9s7mlcwPZB
lBOxSVv+Uwu+fSrrMy+LgL1+ze/icn3muyOc2xZRKljTNLqRtZKd8Tvs7aRZuf8QI8shOhp0/yaO
BcjnJJULhMIq7Udi/wy2F1fhXyRqWuVKqC61cGk8lLUXN2T6FHA5x0kgHS+KpNYVTRrf9oXxhH2j
j8zf50yQZKL4kMIJmy53DOLZn+BTiI1Xtjj/TYtJJn6YpQynLvwG0qyVwTvKgFt0Rqh3Ae7c8H4v
LKP/Sos8ds1ndDfivl7PxQ6NYSMjQjPc7MoPPwAHn1x6pN+3178VhAH2llTcguGpmQrDTxNp2yPU
AQUFrv2OIIRuahYAoZHvBrVIaI2X5VfZFFTu5mdS8K7kg7CUGwgtGCFOdHLvMqMUttEPWXqHlKDJ
prTS5Tv1aOpvMy+BSJ/XuZYfnmTuTkDeGdnP37Gllc0UI4MuXAmK4ZbWcxkAZV4h1HjRyMTKABQF
ifyoP86YS6jqlU+JUZAcTje+FvlKC1/RdmhExpCNZ5DpoVq6tJxxYTQK7oV6hJRwXhZZQeSYMtf+
2Kh6+xQwL8OH6bTHgfTfWDghWpYEU08OquZn8RzH8ZDay1srXxGZgLTJl7nLoWRoA4Fymg4CFYd3
Pfaf//m20yhX9Y3sMks9JohyxLS10PYJ4+loM9eTCoGgkGsczYHS/P9RN255D/Hv4men0J1aCTYX
h1xnXptWNGmqf1DBBDvPuXUoZ4hvK7/8aO/grRN5cjch47GjPGdpsjvKfSJk18z7dDn4Lg9V3QpL
P9qN4OeXbWZfmgdMw4gMsaiiIVXmlYY23G+OmzPp23fBDHOiBHE3uxHg3GRh+tudsN7oyl9oPpES
kVsc07I3G3oEWEaZx+pENxkiBfci9vS6PKTC6aA5QqBo1mm6b48koKRYHS+BoiGrMTfyRCALEvTB
Bq29EikRRhkXp3dq6drsKXs6wWmvQrOcOvgno4uqQ55ulQiPoVgs9ZTeYlzP+DK5EiFHSRpIUXSh
3Ut72Q9GZR/vAfo2JgjTk5miKPPnhMFqP6UKYjTaq4VDdTnLYm6sidP18utKVBi9fK3Q412ozCRj
D2D1FgI6yNFt6OVNdY9kR8hQYQq9Mo89qd2Y+eXUbsH+s+UOFgR7gOi4OIezapAIFYzPFbS10keR
b0mHKLemNOMxgtlaUJHc/WDVdyYYMghXtlftMOoAJfWgAxIcp984CXwANJAXVa/My7/bSlbZGsTC
9N5nJgHsX+pvoZapDbzEa9+cJTAmgmfl0RyJeF2cjBkDmnxk7+eV+YmdKpxnYQdMFtQFMSxjoQjY
H1D8GE9p9wgt5nnfh5AQg/ClwqjHLGglLRCdeiizWKUKRdALW4ljYupL3nahJzuqkjqYUZNlBs5g
EgOio8Ja8rMTFXtKURnjsGQueOf8A2S+MbannXLcZxQbwOQcqijnhWoki0wttqbR536BaFK1uLo4
hZXj5lqbHsxWudOriAjwp1unjcQFkzFsGQVbdsp7ZhelEXpqCfJ+83Smi2o/FFQOkMTjNgxkAyjV
Gu5wrsp8AfPR7NF1QngbWlQzN3V86Njc1GjE4Icz4+4vS7krZZbwaCJZ24KUKIFJvnvlPBSg7a3B
LHqEgz2VC0xdHwfUIdmqVIocXYTYbSBwp/HQkDGPJ5k0RSsg5AN30+7EedjZgzQb7PIGu3S/ywrc
x+89TPolLDR/R0+35BTBwCkd5q1XWMLXACL//gKUwYvCwJcDBDeaJMA9pH4CuMhI2trohB990cEd
gR398mc2t0qngPobQe/LwknaS3axNOa+GV3xBw+CX7nks2dlm/QUuoPmZ0VuKCgfL0qfcvq4ke0L
QiF2Zc9J0GwyE0e7dkniMyO9X2IwItyL9cmhWbSMaxQ103EzeKIOtAaR++411FuNWwhoMrU9AKlG
Q/gpNGT6kTf7bBqr
`pragma protect end_protected
