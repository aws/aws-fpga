`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2016_05", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
b6/iPm/PagUA1S2gcC/eMz+hfa3UjJ6vkYH0IMCBmSMVhTfSztfyG/07hW5Ml2QckTFWlGcI/9lT
e9/vrO9azXoKJUkzn73rBX/Gxtkey7kdujuvsIBwmoJQHKzi9UauwpacJgTp/8N1qXBBkm8yvJ0D
UQckfPGUBPiddTUYZvJM3HgMPjLbFoVcMBGBFn3GXRKV/PaIDynD3PEqC2sN+LpjNeJ6BV3Fchx9
w+++dPRXTrqGBi8tkEbKSXualQKH4uaw7QDqAODexH+EPQ/N+LMDP5CKD2MPUGwfsGpJ9kH8A70D
Ez9CCa0YXj2VoanpvGNUiG41OErUODZ+PWWWHw==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
25ZUOAXa+uPlTFgvJA51/iLSfG5qjbB1Qd12/0j7T6ApdQq60EtsVvONTBQ2vpbpCMEbtq5wQzT6
hfugWH0KT7pmKUKR8xw5rWJq6T4/9dTwqssP0f268iwTLvpybQdQM4oyO4rEXiIaGL41E+fvTzQd
iyzCe9BPG95+FKQ4tmw=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
pZbfPK638zf3+Jv0LCF9IXEH5TL7FMv1+TmPmSwa5dBDk51A7alF1NhjrBlGe5FpnqTSMPzrXeFm
O5XNj/IFH/CFU7uApGU2q94hbSz9vVBePD28ZRCUYjLDopPupyX3UpdYW8akCjVrFGaOGwjqNtzb
F3+oTz7fb2dGtdfTW34=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3056)
`pragma protect data_block
Xc7qgPxhHmoRmZVCek0U7skjsGLiGk+BWBGEBOOZC1ukfCPNKz70MnHMwCIYNjA/XlV05fN6O2fj
TQMA2hqssysBDOGN5lfosKU05Ze52l+nXMoNPMddebaeDRFrTSp1LNZkhUsEtdApfR5BOnoJFO9a
DQBZTcxzvcZbu5KSWz0nVvOfOXn7moMISF90E8QsmGt9Sq6y4MgqjcNVboLb8lcTC1aU1jEGRBhb
GwV5+crw0GEATK2h1apyvHc4/bS46F6RRzNdC1Vmsca8FnzWj8rdbFzvcFp/TPe+u7eIFl2oDwcK
pV3M2oM3Ja3qnyZw8F2cRCuXAE1oduTMYG0bMvXpOC3Ef/Tv9r+EiIoNqZWXnqP+qtbe4qiqJzAX
VR1MRCQfVjtVqRNDuy0ShXCD2DR/y2DtoERk9SioVzdNNq01Ni1kvTlJln4c3Lc8z38d5PdSK7l0
mG7+ursd4riSnO2rXbAzckVsK+6XcWoR4PWcNN14SZuHJHUzVGfq0Q1d8irZAVEWahIbCvtkqNc6
EWG/FIg0yeYqnuMDtntec29abkPSmtTyI6ebtKoHXuIggdMn8sJk/dwFlwovM8FOgRh+0FKl0saZ
8HSnpK0YeNzO3C1iR54J95ins1Fb7oWMakBk6VCIrkvFZS14x4W2p6TqHni6rtL8k66fKG6JgzDo
gGMWQ3y3xgEBej6q8Ad9rNwivxgwCWCYslIouo99bsr/Qcrux0qBZLBqxXMrlYq4GRshE3BhJEgT
iG1yk6Bf5IJeoATHiL+Gs+yMFQYBvqWugIPcaCWH5bUgB7n8ULCElVqNtveb8lop+XyaZ7Ity3LP
P4oXOhsWNPaNPrEvB4bgVeBmTiCjtDon6gYrm7uLy4BvG5QDxyD26c2oUcQM3YubjfwM3BspXrbn
Fl5Dyo/JJ2kiiPIamzKbTFlV6zFXzTEatacW07WF/vzMOYGtl5crKkcSRmUJRb8snCV58USxe+a0
v2OCh4QysLxKcT0PuJSM93i8JImgtJkexSDe0aibHGYy8+hH76Vrl5gP5BUi+5aiJRP/XzR5RXcn
XZGweY2yrgwxRvky6J5g4Xv9TrAwimP+cYUj635GlIEGIPTEzJ83I0inEVOupwspQMnftXdrV1t4
1r5PUXsx2DQCKRdT4eaABqqFeH01WM+htMWnXqYIDSqFp685Kb3ohX9lrNfOuWNeGVvTDrU6HKMB
lmWFg3iJv0c9ACW2sMrvs6wyysSrlL/+C+h8gymqZY6zRNHLrPAIWzT0obINqjEnivyYNEFzJ8Mb
8/QUhptdnthF88v0SrAAa5ggru/ZUXRjqbe/QuPo3oP7viyz79ojtrdjR7m6oMuNmG/ajLz7u5oh
EGlU/eQr5KAKrlkF5cXTHCdeB6H+r1fw1IFMJWLBDL9yzARhWKxN0oWwmeBvlFAHJQWba9EqIGR5
PX9cbBnxOInGZI64S8GXwY6dExkUHiWcYc9LBVvBZjMBxhHL9cBrWdJqclFrcBVt8ovpcM6KkqhQ
TwsBV+qEb2/aFR/TjNqmNnlPxtoU0b8lBljyraLnj98QhvKRTZckNfqvT5K9DiAhvejE/c4H4wZU
7OjqrUROg1hu6BZn8HB9Db+Yn8q7zJLn1zWkPWOT48bUDVbBk7vP8zabcleFgAaLZtp6kExhp6Uk
aIGzy144VSMzbnlZNeVmzBOx1PS4syAEKOhQLkELyAiiQd2qN7XWuQbf7WEztZW5VZxJdoxKhsUe
nDbNgomglDVFvF33JkPAxZelRitdBG6LD+xUR6l+gLZlbF5cAx85S30cEaOlglRMqROjTw9Bh/k1
nkim2Emfo9X7btpm5RElDoOsKp9jFMUr7+2rH97gZLzzk8/9vygWpXdiAC5CerIQQL87cHwJjub3
C5y6GDLVtgW2dErNjpx8hvnw4SmjdStToPRzD9rZvdJOKRPgnYIkForas1YakiX/cYSbi23tSm9J
yjrE5rq8v4JjNjI5jfJk3cfy4Cl+/RQriqzsye1K64R9uXuj38JUVbRVEZelfUaggbYncwFCgf4h
ocCqC1Qbhyit8WL0gnPBIVThNn/vsQ1WTo1vico4RO4lBeH+uurGj+wXevWlNeq/DgC9INvEtisp
QbWfn8HejRJCnDdhUIOUkzZMoyo6ZfA8sjWwd69torLnnuFKB/zbrJlMEy2D0Bwz5p+eBpcF7rnl
1WEVn/JJ7C8FbCR71va/5yoP+Zijpumkg3ZiStd0Pp8n7vexbHeqp1hil3iTDMCxV84U6rVQrjVV
nuc7ZSRM8XYHnRFEiYT2kfLftOEUu3PIp/igcHr1OaU5jstqGXgprPp1c35g95+bXUrR8ZTO7d2D
kW0Ak7mxIozmiWrXQN+2/EaJL1NL5sG0MN6ulbTqStK8IZhzKIRxW9HKAeLS5TyfD1d0AMdwtsu7
Q3bzSob6mBCYX7jHS221LkQ2vhmNbtZVycSU92VVdi7oy4JNIQo71UZPf+DkgwIlp0tldQeTfDb7
vLus7xxfHR0m61IW8sCt6n2Z6VXDvUxbdBMEcR7zZq3EjOdKyUnghxV9H8ZKJnC/VuluH97aEoQL
04cY51tnKxPnPvL+Z69ggnuNpJ5Xq0BW3zgzQaS8WX3Fi3OQYoSpLhIhlepSDPTAS4ZQD/zNRpvx
mMvN+4JTtoaOhBxAl4T1RCFyRYE1KXttJg/eCQmnbIQrP6sQYJ9X+MW1IYbNrhvweLl800jwwY9H
mdz841/pgpEstz9cCQSAARnWzOjX8cgWwPRMj3xCXLB5AMnpxyTc2geGJCw+gJdBLN4SLb8mUJMe
P2Fr2Gbs2l2yi5PLH0tC79D0sD40azWZ68IyR29xNFTlYTZK6rUOmUwdW7PAmwCWbk9H44vA9XrL
5f2G2T8f3lumuTHO83QU/NzzoHi6+wS/KRxcvdXmz6KhE3AswfbssjtFAWcsUE6BJlEa2p86Jqsq
5/uTyKFKYSe8LZs1UrDVmGtpwDgk2SEI+L1vJT4mYlFheTFEbEXTvn30fd1igUS/jzzeNSqhIGOB
e9qT7yyUT1HeTORwJPFWSWRxfvQrHsH8UPDWkpvR3xN2eE4JAYi20PxJUBqzvATX57ovJ8CJ1qvs
1GtWDpGSqSL1GJrGB5+s3K2x8kci+2tWkhVvP9PV65PkDHJWb5p42XDxnldCouv/apqrYVf+yuvn
tJ2EBcWtSG2tCYZVxYUnwqJhbSbRe9Ou4HN+OXA10kJqFZtllZbKvgoPHYWbUJxXg3Vw9TzO/1En
t3tZ7JH60OahQCePOrAkQfHHfPil9GoQkSUTFP+ZE6qj36r6axE0nqw9N8v28t3i75qYQeLzhq6/
hhtIzkBv5omCLE9d81SMr6Aub3K+bXn3uD66dZPVkFKUxWcCnugOQKn6fgVD+8MIsdGFbSRfZ7VO
8nNO00Eol5HH8EHh4vGkmU8K66sUwUTSPGXwfwriOu2fHDEcHz8gSyNPeQJi6hHPR+dJ12sV19y/
gYeG8vr1JFp6FyvF65gOGe3zaeJm3bHL78Z6SL1fAZjHcOqdc0L+xkCWluvpofUjFuIq3UsKTj98
4yYHiIT4/HXWKQOGH0pMCguayoK7HnstTDiifnkVB16lpOhVK24zzjTJFYaPwb1r3L4GMZeCPs2h
64pq18obuwketMzEnqV/1ggHwUxlg1suBD9ieAhLSdXseXfE9t6R7PXy5YDT+IzslONCG9uU9T2r
3+20sMFB37ZbAqGjBfj7pOkJQ4SRcxEqgZHppeLakJONODK1tycFHK8udqIifWoyJWdeUUDPMRK4
2sYscYOAupJmnhw8IScaYD8Z3+RiGv/Dncjq1Uzq2jDEk8zFZiQvrD2hF+CchNFb9J2VONrA7Zea
cw2CISWrzgT5EYPaNRr37ziorEO8sT6LbJMcAQSeEHa4j86MZerDFIkC2/yqCFvAReqCTw/K7Khx
c1Je1G2gBPKWtq0omqG0+JOMqWMsV3M/RuNeJ8hFnaCSoGn93g+mZM6CC+Qtm7tCruq3mbHnnq59
59d/ccSSRXBRdjrz1V5/TZBb5kJkrekqUwry3o5QmVwNX1E=
`pragma protect end_protected
