// Amazon FPGA Hardware Development Kit
//
// Copyright 2016 Amazon.com, Inc. or its affiliates. All Rights Reserved.
//
// Licensed under the Amazon Software License (the "License"). You may not use
// this file except in compliance with the License. A copy of the License is
// located at
//
//    http://aws.amazon.com/asl/
//
// or in the "license" file accompanying this file. This file is distributed on
// an "AS IS" BASIS, WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, express or
// implied. See the License for the specific language governing permissions and
// limitations under the License.

// SHA: bddf8457046b3a64e63d28d7e334020b6f1d09ee
// =============================================================================
// Restricted NDA Material
// =============================================================================

module sh_ddr #( parameter DDR_A_PRESENT = 1,
                 parameter DDR_B_PRESENT = 1,
                 parameter DDR_D_PRESENT = 1,

                 //NOTE TO CL DEVELOPERS: 
                 // The below two parameters should not be changed.
                 // Changing these parameters will cause place errors for DDR_A and DDR_D pins.
                 // When set to 1, they will ensure that DDR_A/D IO buffers are correctly instanced
                 parameter DDR_A_IO = 1, 
                 parameter DDR_D_IO = 1

)
   (

   //---------------------------
   // Main clock/reset
   //---------------------------
   input clk,
   input rst_n,

   input stat_clk,                           //Stats interface clock
   input stat_rst_n,

   //--------------------------
   // DDR Physical Interface
   //--------------------------

// ------------------- DDR4 x72 RDIMM 2100 Interface A ----------------------------------
    input                CLK_300M_DIMM0_DP,
    input                CLK_300M_DIMM0_DN,
    output logic         M_A_ACT_N,
    output logic[16:0]   M_A_MA,
    output logic[1:0]    M_A_BA,
    output logic[1:0]    M_A_BG,
    output logic[0:0]    M_A_CKE,
    output logic[0:0]    M_A_ODT,
    output logic[0:0]    M_A_CS_N,
    output logic[0:0]    M_A_CLK_DN,
    output logic[0:0]    M_A_CLK_DP,
    output logic         M_A_PAR,
    inout  [63:0]        M_A_DQ,
    inout  [7:0]         M_A_ECC,
    inout  [17:0]        M_A_DQS_DP,
    inout  [17:0]        M_A_DQS_DN,
    output logic cl_RST_DIMM_A_N,

// ------------------- DDR4 x72 RDIMM 2100 Interface B ----------------------------------
    input                CLK_300M_DIMM1_DP,
    input                CLK_300M_DIMM1_DN,
    output logic         M_B_ACT_N,
    output logic[16:0]   M_B_MA,
    output logic[1:0]    M_B_BA,
    output logic[1:0]    M_B_BG,
    output logic[0:0]    M_B_CKE,
    output logic[0:0]    M_B_ODT,
    output logic[0:0]    M_B_CS_N,
    output logic[0:0]    M_B_CLK_DN,
    output logic[0:0]    M_B_CLK_DP,
    output logic         M_B_PAR,
    inout  [63:0]        M_B_DQ,
    inout  [7:0]         M_B_ECC,
    inout  [17:0]        M_B_DQS_DP,
    inout  [17:0]        M_B_DQS_DN,
    output logic cl_RST_DIMM_B_N,

// ------------------- DDR4 x72 RDIMM 2100 Interface D ----------------------------------
    input                CLK_300M_DIMM3_DP,
    input                CLK_300M_DIMM3_DN,
    output logic         M_D_ACT_N,
    output logic[16:0]   M_D_MA,
    output logic[1:0]    M_D_BA,
    output logic[1:0]    M_D_BG,
    output logic[0:0]    M_D_CKE,
    output logic[0:0]    M_D_ODT,
    output logic[0:0]    M_D_CS_N,
    output logic[0:0]    M_D_CLK_DN,
    output logic[0:0]    M_D_CLK_DP,
    output logic         M_D_PAR,
    inout  [63:0]        M_D_DQ,
    inout  [7:0]         M_D_ECC,
    inout  [17:0]        M_D_DQS_DP,
    inout  [17:0]        M_D_DQS_DN,
    output logic cl_RST_DIMM_D_N,


   //------------------------------------------------------
   // DDR-4 Interface from CL (AXI-4)
   //------------------------------------------------------
   input[15:0] cl_sh_ddr_awid[2:0],
   input[63:0] cl_sh_ddr_awaddr[2:0],
   input[7:0] cl_sh_ddr_awlen[2:0],
   input[2:0] cl_sh_ddr_awsize[2:0],
   input[1:0] cl_sh_ddr_awburst[2:0],        //Note only INCR/WRAP supported.  If un-supported mode on this signal, will default to INCR
   //input[10:0] cl_sh_ddr_awuser[2:0],
   input cl_sh_ddr_awvalid[2:0],
   output logic[2:0] sh_cl_ddr_awready,

   input[15:0] cl_sh_ddr_wid[2:0],
   input[511:0] cl_sh_ddr_wdata[2:0],
   input[63:0] cl_sh_ddr_wstrb[2:0],
   input[2:0] cl_sh_ddr_wlast,
   input[2:0] cl_sh_ddr_wvalid,
   output logic[2:0] sh_cl_ddr_wready,

   output logic[15:0] sh_cl_ddr_bid[2:0],
   output logic[1:0] sh_cl_ddr_bresp[2:0],
   output logic[2:0] sh_cl_ddr_bvalid,
   input[2:0] cl_sh_ddr_bready,

   input[15:0] cl_sh_ddr_arid[2:0],
   input[63:0] cl_sh_ddr_araddr[2:0],
   input[7:0] cl_sh_ddr_arlen[2:0],
   input[2:0] cl_sh_ddr_arsize[2:0],
   //input[10:0] cl_sh_ddr_aruser[2:0],
   input[1:0] cl_sh_ddr_arburst[2:0],     //Note only INCR/WRAP supported.  If un-supported mode on this signal, will default to INCR
   input[2:0] cl_sh_ddr_arvalid,
   output logic[2:0] sh_cl_ddr_arready,

   output logic[15:0] sh_cl_ddr_rid[2:0],
   output logic[511:0] sh_cl_ddr_rdata[2:0],
   output logic[1:0] sh_cl_ddr_rresp[2:0],
   output logic[2:0] sh_cl_ddr_rlast,
   output logic[2:0] sh_cl_ddr_rvalid,
   input[2:0] cl_sh_ddr_rready,

   output logic[2:0] sh_cl_ddr_is_ready,

   input[7:0] sh_ddr_stat_addr0,
   input sh_ddr_stat_wr0,
   input sh_ddr_stat_rd0,
   input[31:0] sh_ddr_stat_wdata0,

   output logic ddr_sh_stat_ack0,
   output logic[31:0] ddr_sh_stat_rdata0,
   output logic[7:0] ddr_sh_stat_int0,

   input[7:0] sh_ddr_stat_addr1,
   input sh_ddr_stat_wr1,
   input sh_ddr_stat_rd1,
   input[31:0] sh_ddr_stat_wdata1,

   output logic ddr_sh_stat_ack1,
   output logic[31:0] ddr_sh_stat_rdata1,
   output logic[7:0] ddr_sh_stat_int1,

   input[7:0] sh_ddr_stat_addr2,
   input sh_ddr_stat_wr2,
   input sh_ddr_stat_rd2,
   input[31:0] sh_ddr_stat_wdata2,

   output logic ddr_sh_stat_ack2,
   output logic[31:0] ddr_sh_stat_rdata2,
   output logic[7:0] ddr_sh_stat_int2



   );

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
k3CtFsv52ABnOwZWNULUFvc5cJ1cECbxHWQHOSGT0XG3S68i1O2GF7DV+yMBf2SVFSrqg4HmMHCQ
jfdfbje073XEtCppB7i/sec3CWfrfRZalkbRwbPj4MQtDJ4m7AcBWqtY+eDE833b/vdZi5ht17np
QNqaSIYCyMjoUMXuzYShAt/EbIi4pHOiWgCU1UKgP/+XnFnzqgZnKMgEZPEwpCN5f12eYlchSnr1
VRK7pIVe3beSF/pINTDNo1gd2yS8u9sWJAwIkTD7hefGW/7Cz6Ct6gNHztU1kYzW+aSBQF8N0mw+
GKFL5GpNj5yAIVk5TscqNo6bJGh4vunBrVfZWA==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
KIetJ9KEOHucJU8T0PCD1jv8Idyt0JXtK3hdCZJ266nBpquheVvRu4IHzqqwUfHbWZOxQ4B9R53v
uIN7sjnk2Tj48hy1VpOWC8Z9jUy/W6Ehthcf/fQBh29OgCkeXVUuxO7xXlAFRRZ0uB0xW8eAR9ci
k6n7bqNU53/CsMDuBng=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
UvXkCu/3ZNbQxp2u2yO/2n+h5iPF0laeBP/3sK4l5Jjf7XcFTY6A3RuI37f+m3k3FWJRq2RQ6Ugm
3uZtGOLn68rnUQ2GSvjSu1txUWJLE9O3/XlB7zUxw976NNkha2yNMBoFh6OdkUDb3u22MIb9dFU0
xP1Bstz2DzKNdtaSxqk=

`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
YVyFZ8tAKPNd3r4BjZ8w16+ZZ4yYTbdHXUkKbtss5xb0Sd0a9MJipUobgvWhvYG5BtSVDfeOf8QT
pj5mtf4ngA==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 72800)
`pragma protect data_block
y0b1nRf/WJxBxtuO56oD/KaLCFKnYe8z2rsxphoJv9HHXoQbfii3G7vp0lBAqz2VUChLJLCMVGMa
lYZ/Psoy1irpDgT1yP+72AwYswrndMSkdsXzvB6sXTqp38UCf+yr9Nr8LvDcNK0GqetEw9f7Ca+J
Ou4S3kAnXhaI142n49mcGTDQWRKgyLLKZqOscUUoTmvzQDR3nbiePT1kCY/Fycqsx0csM1Jx2nL7
FGmFoNqMSqOrStWEpwII3YrqIL6LC3ZL8d9+ZEAc5+bBmihzcXLIbRUKM9zMqvbEO9RnbZwOxWuT
6i6QVTmbNbEeROEQOuDgrZFWFYNjOmxriaCrG5j+8lNFq7n7eRFI2Oa+U1zSuVPdAiwpHfj6s45v
2TtyTf2GahlMzt6M4vhe/lmOHbpqH9Iqm6TbOvpLOOCR6N7KOiwEfWNqUQWUq3yHfYcg16LDJ8/0
09+xWl2KDMPwO1Deyv1+MgBeDK6Qy8G4UjFZuTeOsGVy9YXj1RfakOI9e++IHHq56kQuzWTShzMn
vTjt5WJGZAY2zSpMgW6eWtybWID+F4qilFDWorqjJIfLkGRQDVzIovv2VR++Rcu0bNeSwKZjC4XI
AW/9kUURBIqzXOTqEkaurRfvoQ+yT5dwAHxC0DW9c59rKxHrktfKAdk4ATUNekQWgMaoo9Ho0Go8
oq/3aVFyASSJ02s74Lv8uBjYmIRstn0Rp03uE6vf932rh4MjvRmbrN/uI51K0/4FlCEnwYB8aBUj
i1whcfFF9bjJgimmeTRfrHKKTpnlydJZOyRw5wJCkPBwQ7yG85HIqTPKoeQQXLMgLXpgQgvBbkvg
skMF4oeZQmROvvyWnxiCH2Cwii6+lLJGLzcE9cjsljCsKzT2HDKpIPtyXo8BW1QdENAAiIzX03Nq
VGJmmKcWc1vO3FEIBFJjt6Dr1ZvmXw5MOIDWPyvh0SI76u5wYe5Q8Vgok02noBADMTHuC4tm1yIb
46DpKRQpZQt/HMePNlU00fSiH/b/YBW5VwrFoLb9N5Q2ZpfiAwvd3Yw5VD+6ZkVgW9FBUWuUwjVD
Yctirstdw+QgFSzA1x+LrSKUVNBDU2nN4A0zi+C3qklt+axX/aNrXAZmlLMP/zUE22S7kOKp5vFp
1jLsm+BK0u2YKUIcIyY06aVNa/rjXSgwZpegSXo5uvTEpK7XdglaIYHWnO0bc/vCyiI46xoaZCMs
LF4DMN+a4aRSiQ9ibSUroxZLkHE5CdXMyaBxOEDgf3gEwU2/Xe+yyvc8oi3YqJ7bRsfJKmIkFhHZ
p/LTxErkPAc0dE3zTDnPY5B2hJQu7Nzoxzlq5QyGJOebFd8fzLAuiIMrAa0O8lrDIE9ZANhRlpwM
ZXFDvn1orhgiapre6MY79aC+8K5OIctw6H3PJIQDHQLLyeY1GC1fqcPukvJ9YQXc72l+RqE4/wiH
2YzMGEPVrGIi317ncx+iHcxPHLs8cLIQli60pgXBaIQBj5mD8iyEgO73/vC7s6u/bPABOaSk0OTA
3b30BWJACq1qXkiwM2kC3RXHe9xuZqIby7Mrg2gpFUwgIoho1S/Vrfi7nnEACkzInZmKqVG8koNC
pnn2/ErfyIS/ku6Jq7takEHHyybRZAy3nvDVxUQG/UiJsyLNsCWKd3AGpjyDkBsPqktJU+O6Kr33
x94OrBulTHdt/jPYzFtdatCTB4qiGvpbLqiV2NoUtGmI4uFBvzPSwRHZiuONoe3pGJUkszSCD2Ob
n+y+wCsoyGqrE7VxPXng0ejHGMepFEkiTcMpcoajkfI3iUorjKyH72MLYfuQ/Zer1CWuLLJr6lmH
FdAPuvqqGOY2daz3nKxkWW9fYdmTzMU6uP2FVilbtLf/eICLvzCSmGc+EJUrABnIwEeh0qHb6cTf
Int6xfmlNDq6xqidZ9KOf7zBnTVtb3aVshl63LNaBA+qfktCJ6F4G/OXhT9DlkdKuQ1Tt/zGCW83
St8z+U26hd9LozUMBiNWMtlemNSMBqHxw4fY66MoZ0rjpbAIYkPrfepIOrtX/u7b6Yl0EgrblkPx
rSqEm8Z/lsdc+e5oHTXPGyNtOo+L+BElqkx7GEhmx/x8OMGwFe5G+Hg4WmZYYeuU9rkZ56aCD66G
Z6pnGafSW0kN25cAkur/D0vdjdtGTUxEjwf6Cq5nyjtozby2osz5BKr9kAhBexq7I5ZOdwiG1Bwi
vBmZTDig4BuNWQz3CB1xSnodFPiyiZbBAfBdnZJhlJeJEpEWf/qvZlG7W3sTlqXyjwq5s8AUCA0V
BhJaTPAXv3zXOX+jk4d2dav12tyz1N6kOd55lnGApSCYVfBnImHGEkgtpJzJ5XpTsvAA5NMkYK6t
Xr84eKOlIacdKz7xAns8J0fAMHR7h/oddeKHu3mn36hQ4yPJhrvtb0BcjUcG5UscxQ8j3UYUScQr
Uf+reUeEgRbymka7DpV/cClWIC381eAYTncyvYKLO/7LaESlZAWjiTxRN+OXt8ri+hBQ0Ezx2boZ
beoSBTvwiD10AAThnMeUN7wHUXLXvHe4jGrn+jMrYyGMGoH8sOTpnenRqenSIuErTNCZMnhhPM/L
rzYVpjKqm16GYX5vMd3btUhyFXPPdWJGTtx4dTlEybuJe9qlGvZgCAuXQkecJ9vKY6Li8T9fdRW6
dOiJaq0FJzbSzBOkjcZG60fM8mrRFjDNp2laqQCiSs3BnH5JMZd/ce8bowS9lpoxc+slrWaq+IVr
QGZbvQx2kycnt7i+QFxIn9mZ6kAItc6vYOsFSzzh1sFsWIpwUHoUNrSOz2IzMoZt67lG4R7d7I9D
AxuClBt/R/YfDVfHxrVfNIN1SUlMTgdY9mQtagfVbOLEDUw8afWySazr8n/gwMQNX95bTKGvvdCW
tYUy6FBLxNcH7BoW3KyI+ae0FzXpDZbuhpby1wM8TG3YyuCUgWctpp+XX7Ym4vy4RKe2w2rm54Qw
tPLOOQQn4kmzQJ9yxmtHcNOrWClIFUbmHTrLODrY1dCST8YtbLxR6tkMMckUGLhQYjKedmyRXdxZ
UsNHzIIaoNlQW4WX/u+A8dSJhHMn2dI7LK+rAnUxiDrBjYem2sa3waRHfSvErzPvHBWewGu0z1EB
B3rnJTrNdI7KzGWadZgFqp6Akx+8k/XV/Nap+syoWn92IMlpBsH4c8kYYk2KIfRxET29Y0mm3vc7
WS2pojTvqPaj7FuCcRW/VYvC2f7p0rrfSpkT3KDRUXv2ZIP3IufSLxHrxBHu3mhW6tJZ2hvbdpTX
jG9EK1PzfWNxvaqwLJ4TqcuajLT0qWu3vVS9Onay2nzM+SejmTUn4L2O4fHMJsytoQpBwULJl7rE
WAdf3OI0ZjpXZEpCDt6OeqGlVJdCWBfRXqm8x5IYDjAQNBGEQCo7Edigkow/jTe9bMnVpqe5P/CS
2IfeC4C445pfQtte7nt4L6YYa37/cVl350FLCZhdeC3ERzW1emY5dlXGAwjLrwEgkP0ms8TS1plb
d7Ia9rIcgyioi4WpoPVJclk4+ddd1z/m/3PYIEt6qpM4Jmwc5/rhydAe1qEzbPArHSYt2UVjVI4O
I1Ny+OGC3amSj/zYIBka9rlj9glpOv/EUHg5jiDjJ6++Z6kSfoulKKqM6M4XufpnqHnAEaf++O2s
Op3B2Svmi5hLxStdLnIJj4RMcNOsPdbkajsuLarltC/zlA5fiHYqkfa/Y0+NYUAigWmKgrpH2R0T
eNx/z16LpdCbXUJIDEQLMU166eI6ZDYOpQIvbQQBDUAlIqPNiHXjNQ2rKnzGXYrdmrmxhnrub2BK
G+qoswJtSfBorDbFV7RuilRwd2FNy9OAo9FQMqaaM4Sd9xETNEWWFueKMgyb3KdCXZ/Op+5FbZms
c6fZCAAMaaTsceDC0h/PuC3AXBuw2GgA8SbBI0b0oqXWnOQDeTSjXqPWwEmEoxhfj2StDvIG743E
fBIlmUKwmBijJb7T8JXqHkZkWAvCmoF+ezvKv7c/NznQdNwmoEhy8Z6npXVtM5DSM9bq1NdFxYTZ
Chc3EyfUYrQJ03b9bRjhBXrKOxG52oVYwE16vexI1chgnbaFaedFNW9b+2cSZvM6DwHCSDkwryuf
AySQbfGEAfsQGA9NCSLp061upxbuEUQn5FxlY6hFyI+gMSbkrzmUej/gCA/zB3cGEDve4LB3pWIx
qFTsjBzq2fhiTfPLN3mzYtMXDZH2fwTbngXjXi1VzlGCwe8n4FK76/Znw5LwwxQuUYzZlCpWW6lD
C3WOdEiAlj+nC24tfQerdt1VRIBX48dR6l8JDAACts3h7y44liEVbPTep8W+XSL86uGLluLxMA0T
/nJRKvd59mLpt/idq0vNlgxaaFyfS6gz1fYBXSqkyX4pMe1sR1OIRG+FB1FELjkr9KTG3puPuyHP
Bl7+1um5wjZr0B3Reimkc14To9HLtDuR+K7GsxIPUtftmuZd2HTdXAcX4CCIS9bOouJmRrLjeFNx
iut5EZLnyHXeU1J9tGyPqpaNIROO8R3afbY0rTBCPImghMsUht7AcuYGg+Na+TvuM+pJowPYKlac
5bMecCPxwO1HL8juebgmDHV8nTYA3IACQpIuMDl8lEFYBBu1EHCM/o26Bst+0feg86QTeLcze39R
wPNYnPi+xb2KwoyTDpcL8afpSnIq8x4SOUDtcLwCaUH5Kl+vOSOTzGEJI+8jOATor8ZKl3CW61EM
7Rdw0nwc+cqNQGa6iBKzWqsoFcNusF/bo77dR/b/+bs/CH2maAWDQSg9hadfFBE5Zhm2pHAyNpOP
Y5q1hA+y4h31HuaUdmNDJKQIGIoUCY2CV6C7LDokpqFkea5UGm7CY2VHJibFgKXrn3OIwSuulqil
efXLQi+xAHZY1siLZXDU0zXw9s68FdaVWn/H3RXioDoPxKN3pisINKhX+hXz66RoN0YzlW1ZkFoO
3px8w77WTry7l49qmYgfV55G8vXsZUDMENKAXxB1RN8G1hJKNfldmpCLe+8ebh083njdAD1yNHed
o+I+aSg9Ct0syyjWMTfmY+a3it+yv+bJEgO5yZA56GCPASqc2zDkOlmXTqp5kZo8jwHTIl2Eg3is
+BIwoTtrKmF9/cEWh4sK9VWI5vDKLgceMXFykYlO5a+vUfZtinH8czDkyZQcQV9QLdghO+N0HZzY
44DT/Urh2FH9HmLTs5qpgZ5Qv7ei/ubbAtdPQJS9HLoqPUMWs3CQP+3GTXHVXG7F6nHzgYj34RMo
FiM7RaIqzd9sW3LiM63Lc4LvNozydk8AbyA4hMKb6pr14FQ2BiUxDkKTEigc3FTMQ/1K4MZMAV0A
3kjiqK4B0MOjDdTMSHEnX/2+RzgyIMnthC8Yd2iZyxqUIhkT42nTbT+VFIGU4s+/55iI1glhyRW6
M33RxjCgMJ+oqSiL+hNcVAQe7OU72YDBDX4HWpJsYMZQqxdBypb7iUIkgxb81V96FgvsC45EfiEA
S282pYdCUkLPlRmaIoiv3SIaaq+xSeZjBnvLcT96hffjZPBmiUWIqsNyylBZbN0rw5Q4QuWg2kdi
WJuWGrWGl+6+ilVOSMLsSYtFtxmQlpaG3S95YBlBvpbdev+Ek5dPhYQ9bRmylIsOpARtQkN2lvoy
IPYmuS8kKPWLYRbEnQRxZH5LEo2z5E5Qc6EGQv4ewQNwhE7SNQXc8MBSxftIoDdEPaF19/nK+qiG
BYxDCotCVa7FbMutvVNPBpRomY7k4Tg6H5vW9KrNrpoX7hkEmCxMwAdZd+bWEdmiWKUfdkKuwzAk
TYvWSKkaMBxgiUeRTv/hffQPz093TnXXAC8tf0/KjVT2/NsvEN/+7w+aoDb60WG1dPm+U6ozj99p
bdCKRalCIbVz/6DAv2i3AO3/AWI6cJq0+lzsZtKK4i0xEGay7YzWp+zRVJAUuYw2KBZUez/lSX6W
dUpo6hMQAArps8sQdqbM0nAxuMd1EY7EPGbuiBHFuLP5ejzvCQKV7DvA+yggqIPo7V4I0DzB0jYV
7aCOZ3eFIDT1+UqD4uBRk6gJ1A0kMSv1RnvBDcsJkl4rD0+tVXkXGY5cfXgQZ1hT4DQywzbaE2nU
xw/GGCqps4o7m8FWWIREZmRYDKdL5cU1g4Uj5/Pok125xf9Q9XHKeQJzDephGLsFL39Q224TLQrL
B7/FX7/ukpI2HSHnWt9q7S7Ckk0pPm0ijtOFLy2BC5AVmzU2ETAfGPISp8TwudAAufCqtFKeS3my
gDi7V+IUcP/im0BMRUbmrTjAtZT40py8sMgmJU0ncEB0gvwsolkE91u2vpk4G9I4k89bf+SwpnXN
r3hRdWo22KcB+mLHMKcJApeAkkwbKHKhs8KGmf84vg9Yx564ZvBv82erfRufvk5SuKe8qruGHZuj
RPJA7y9NPF+yppRnuixtezSa00L/Li6rjNRli3Qi7gNSYSO5MCnwoaYDL1WVE6gdlpOjxEq+gkyb
EWp+yHmXD2I1Y9Rci1sLPedfnafm9o5KIPl6jCqUqGCvSqJqgchLdKYh3v/TkClJkRGSmL3zGex3
nJoBOkQhzjlGXR9NSF/Y8Km08h/9ijf+C2dSHeo4kMGi99wTDpzx7e/1slBls9b9ODMIc/JWh4b2
AqwSULleWLOedC4HFRa/GdEGWxrXGzc7LgCYe8l/v9Eh6Qin5pp8pKPxXEkb6FwZ19Ay8dGCKghj
idUbpA15VhwXECh9iwO6xy8ZKKq8jeTQq6i+yQxIvcA0rY66fMtzJMxK3nBmQvI0ik5nyRsx39xN
keRzxCsQY1uv7GY1Q1P4DqLk/MWcdUkdR9HakYDumq5J+BIpSJqJPnj8aJ6t2C2M6If8Pw9m/WSW
QJ259tnb4d1X5VXQX+8A9kxtdo4XP8wGZ9YiI/9Z3dUwOwVuPnJH3LfuezIAjFwVLzDG+oP88eCl
zXOhGUFTUfiWao4hXK9eEk4uBwcYFH6CPrm0/mrVxAwhATfjHfSYbrpa0ayUYl+rYCX9D1amy7bq
0d/ePBvyKB90WM95KdIZPu2AH1brH0bcpwrbAXUMgTC669ZxI/hR8EWn4jeySeE7SiylZZie2Q48
Zgxw4f7OJkcKJxTRjIJBL9XH597xrykA3pErzA7irQj37Ak4sXRQ+vwj2vtwI8YwoR99UquPwLb3
GiX9z4DS++pFNetZScibpiTuIDTvqkbIQ9/D+6E/9Jt4rEmLmmJYKNzboFuG4xmu0ooOXDB7S23z
SengUfoKO/ncVOPAvu/Ab+QCyFj3oGQelof2+cjL57IfosZFvqSlUaNMfvRoXsUgb+CZ166hlQkp
pb4TJxT4nmNNgPVWm4WqT1ryVkMvUXHUOVH2pkGnYu3nMzYMCveMFs2ABGJ0QoQFitvV5D2QTEB+
iJyRkXtCguu4U+QHjKzPwe5DDp8J1uCuusEqand141VUtOiXcRiKwmVuOzDY+V6tEBegGO+m4nfn
Xsj67RRP8Q1I9pXVUlesP9okB/ebS77E4dCWdRo5BEhJzuZUSt7WPn/vMeeLApm9iJif1naPWMF5
qzYvl2mae+b8PHvKRsW0qYc5nwYl0ZFpCaoV2bUM/RDepfMVCy7X9eVEdvrAxW3WXkNla7P/atzI
Od6iG5ZI+/6nUMmpi8bWtDRQsEFKmnGgfqnN12MxBgBh8KuPlWmGSeFxNubVSP+7jKNo4CyQqKyY
knZ+lY5rHtjwWgeosO7EPZqfVAVETUodFY/ZV1CfaNRb2Nn4FzDvKCnc7y/DxYwTiy7MAIjgdg5N
9wfv1b+Gd3NPkvDS2iB2Odd4C7MfZGweUn8rwlpYw+KvMdb9eNAkEaN3IRujYLhnAC8UTRAjWoIF
MZt/x3CHGklOqQNNFGmpWCn3kS3z56SmWxFzXWTy8yPOCYekRMP7HYt3JO0qvcR406kUlauoKFwG
TU8BHmXl7xAHX7ZlaGyYjU6sPaHNvpkH/E9vxt2Ef0kvk72L5oc31MgaUtvQfhBGKL4Omq9nPh+Y
jFfG4qFUoZRb5CZwqqEQRJOlQizoEvCDFBrq/amkgiax2fSPtpuSl6vcvODvWnZyxYUTNAqr2irR
kV/rWR66NYEKk3ZOHYWxfsBxULJxeeLaZlCf1rhznAyKdx9JC5HR47HqoKQ8ODs0zhJD8i0GKjXe
mSBKDvM5jokmOX6dhRpEO38gb4BnDLyj8aKeAxxzKsNlm563+YjB59fk8RXnfJ13tufiua8L1/zY
xH7lFshaa+6pajubiLmFwQpf16WDSSREYcmw5k8IxbYlTGmK14yBGwzVCTBewcq+/dInjpSNBUlI
Inklg1THlxiTJRQUWyDdzpTUAIzydJrr60rvMFkd2XS0JN7kT0OwqAmC6xvviiF5nTswQxtqleDu
i1NtNnBlOuKOqvvIkZ+IyidIr5hio6Gdy4iZF3opO+cdzfldp5pZ/2XeBzXp8zq5mwXxslUau3uH
zRFkypx5tXmd41CdbKr0rMj95jvrXRDygoysbkleCCx/QNrQrvvIDKsONpmYXilp34uE3Rrw2lrX
2Xqv37NzQouiEO4ZiTlsRXdwhYJXxDAgTSdO6rPuFIvVT5r0gav5gpNViuzaRF9wkwjaWdjK82YH
MSZlbasQlQhkuQT9BkB04LfyvYtUIU994ENNPTVgBrNAi+JleIQA6yOKKc/yt8By/5LF0lHbbuix
P8v4Wc+NCnVBW+DwvR5dtcRPmLkaNfSVgcd+a4ZLgQKfRZIMFN361B5AgOAcRqNVvzIQfG0a9EmN
ZS047XN+hOVEg48GMtN28Nr7uLwsR+d5zBF+qOcxp9wzBee9h8SRNy3ZWUooYbFRYfvydS38x9c/
RHz4yrSsc7a6L6o9ONO83juch5OyrTKbbfaxHqH1RrvWTtlTCfQuT/Bgkpz1QY/0deEQnD3AUjje
xSK5MacDxwA3yPDzl3KcHo6sBQfRCLGBtFf722uaaoRENMSCayp8KzHOA8r96Chqaj8hl3yNR8nL
7j+lHyG1B1B4hLBiu7LHlGdW+Wx8viQCv+GscXLPt4zHOTFKPBrmnWPaix0P0LVg8AvbpaCfA4Pf
uPtvmjsTco4Lng10pSEZekTWnW9QbhWNVAcVzT708UyFnrtq2Hy//9ApMUciR0w8o1twDfnAj6iz
ET8/sqCI2Rht9ZySoYp2b6mJFJYpjn42rLDJ3JBDMt6wBZYDV7p9RnXP6/B8F38iUDvk7DPZTmJu
sJ2qV6nMBO7ODLxU0x5XQXnFsbD0iNsOU41kqPKn5VAQndiECi6qqRSeWJBrSsku5aUUuFHXSJyR
F2n2WaagSDMmsyypRP20wOHYZEnyZ30fltty1FIGMgkl1i5kgoEk0eMj9ZFViXHFbSD0ZFPp7pVz
A/A3cRGBT0F8f7My7kX1T+9tCFgFd4zYu2+cLHNa5VOy06sjxQiWXEsFLIJlANjnjk47TMLA+TV3
XNV+9AZZpD+fRsQgQLdhvMTvL5SaUBdLRFJlG3sJWMze9aRLvuCRhSNZud2WcBVN/kttI+kbPPpa
mswUsiV6ZcQyPrOJMwT4l1AI6Qu5pPSkqB/JiTLMnHA83C0wYVm3a7LbR06wLTw2o8QU0dBT1v/7
LfCDTNu8HlVq67oFd9ww7fXbamKalXDTe4Koo0tZuTz7x1ajitn1UkTLqvONAsfhohCCApeC0wPl
MbQRQ7RgJLp8gwAXw9j9vxyXXVMiqxo2afHe/c8jYmnN9l0ErdFxYbsBA9A6vWgzDysNmshoCZGe
qSZMK8QWwWeeku7Wy83DEmLYm/rGcR5KnqR2QN7GPFCid9874PR7s/NMNiZ+H/DdLyg4FCfW0vFC
v9FoGxOOGXVkLyX67M79yigdfRQWJ7ABLHS6LqoxdumwHHjfeiOFNoqJTjRkPTWj6BylxIxmU73r
k33yXJATHVmfSPcKKLPJzb3fdMR9h3uYJDuI8PX2lu4f2WHiJInfczkgFt4jOcTKBJ7gpuf6HUNO
a6NZInVZNpLXpzwlSXNS+gn/W+nHy6VYdtVmpVd/VV4e2sJuy0e8GUiaT6cbhJBxNwUNPDFg4rOF
+gaBpj5BL6Gu8G+Jq/X7Q1h4cQ9AZLwLTsKrzcMk31pQdd9eTR8V0QqpN8PtTPPmo1eehRWGe3Z2
CLFkoF2YjCldtj0HGvl2agAX9A2cK70xJziL9NZwXl1vu/2Jr9FsZEsnJGnmgryGMPHjQEQiX8YB
McFap6f8jPKf1k3uupkuqTeBdTwHbBMtGxqJS3hSQGOoxEMiqpP5TvFWNORU7dxZFAaS5QlaI0hI
cDq3dc0nB5Fr5S37CqbgsOGx9gnH7fpQaWaCVPQfBU99HFx2wdvi1durK5oSOQcQtNKdWLSzujr3
6XqhecSph1GYkzh2aIw51lHK9oGMqMPNLFaz4ghHWd9P5NVTY2Gw8GC39LEG/OXA82Ub4Ts0XZ33
fJdaCh6FvkLuL/dIArU3jDnzzOzVxXF/fJ530kOVAOcptAnyeQClyH/ZxjaiVQ8+y+od+U+e+Uil
VHmN2fgXtA4gal3PquW6LCrEP/wnyBFJn6P5SRLAVlsHR8IA+p+6Hpp9o8lKN35mzS+ftUL/fpE2
Pb9F0qeVcauTCEANKbRnih2F+Sx21URlwdi0o0wi+gKPL/6UmAirFziZm21uXmT+2auYjo9oyCjL
AubnQ3uyJmS9WQeHWIdLsjW++HjyESu7gUctmAj44E+wtiq98nr67ZnmsPkUog9rfMUOPjET23Sp
DYbUi0h2Gh0DJOyfDnw3SWrrNI7UhdQ8OjBK+KD4r8ph+zu/Zom7bD08Mv1bKQ8Uj5a0b14Xd8PF
1v+lp5nWX/HRg//hI5t7hMGJPU+COe8GtxUE+AVVEzgGz/O/0xn7PJPESZHG2EbobZIYFc5Ce0ZT
joqXHN5Lu3/V0ywFAIoLStyH0ieC0R3AMdvHqO90H3mlSB0Q73sPYOZbt9eNpSG7lvxstZ3Aio8b
ctQXPFoOiiRCkMYGfagUMYoPvYyiW23d8kOc3PJQICpmN5oxczz402e6NFvTyoI8gdOs+oI7a+nS
AGjbLIIVCBM0i5YCTGhJDDA0eBSbfgKhjhveIKc2UwerfQbPomTz5rcQcv72zn3sLO1S3uQQ7+Zh
p4CZojypFXH3f0Y7OlTHGKMiKzfcQcQDx2K0dWYWUNIIrU/7nxunM2QFiZUvA91HmY0aBOLUqPNh
ODTk9PhHfneoDX9rgYSz03/3Zp4Dof5PM+a0G9grgvhTOoG5oXXM7pfiUBcsshYRo8h1jiuneWrc
mI/1+ALvtesUhG+dXEgtPX/qaaQVyEkDLztML4N/RhkG28WQxDLIBxq4kkZJ2vMC586zqtA0sPKV
Mc7MgH68czrjnlYo8Z3MZn2811jUBjsmnsw6YUKgkpXD6FdCHi1N1ddCzLAgUn14Xc1tka2zlntZ
T040gHYFlbv/zoHcSk8m/az1M6RkntlMNv/d3czJjUY07WlAwtJLlQPx9l+rnsz9bd1KwBUorwmu
hiRw8k9iwQuL6Tp4qTSLQk/ohROyBs5Gc98onQmeV/HhuiYnKCVxQUATVAdTM7yPyT6bziuDEyCd
1Vhhgi29rj/+UHNN/8kxvMuzgpeWJNmKLYrlOIVDYefrshD2viBSIshEw6Chx7+3rkxnMK0r2F9n
kkfUNe3KfAB3ACJLTDEJv9tPV7KYmI7POYC3wuw1wKx1Ik+k19xb6cFAlumaLqa6RCX4IHApt8DB
E0Lf2Yc3xaL8jBdVnjH4ipPDZwDec4DsYH1GXiJHOHGI5lzwyHs7NsJazhUq98HJ/421+Qze6qA1
RzlpGxAIRaEZdQqikRTTDGNwWP28+nTneR2545qNEcbg6OTVKZR6qK2r/A27qBxTsdpJpzV84CdK
np5woNjwutgBJ/otT4D/qwQXAq3kQQw3gT9SGBMdPC+fIa/ZYeVyMMBFJxL1cW/0frr8LJYA5V1y
rPMkqGFahCAQfL/io1H4sN9oygGoJFZU+PLI+syrM8ed31lZI9LRyGJ+6DAvPp2sVdA4f2P6oQfN
sTx1CD+bldwW4LhVNaFv2RaNWtX2iU9uSPBw3xZdsxsnExdbK/mOBN2fXBnKUNgWSzY/ib/58tsU
6eFUsAYkGhUQEfltxzMJ2mlPHiwP2zZP0rf1lTkgxhFHoK2mDcwInyJGbyPXEz5NZoJt34/a0DTj
sag9VrFJ/qp6sUFMtDl3jFnb6gzNGbBFul7wgcaWxsEnOxA1mMThZQjIAZAS1A62LOafVzzul8KD
H2GSQ0tqYycrVAlOBdeLRsz4Vtrj378N5htHiKFgHhgUrPTy4XjkBknUiCYoNr5GzTMkbdGRuOyf
FzYSUk+76UlPyupYPwETe4R/aElnslGwolOmQhGu6GtWkbXXI0/JZ9LPzSQAN8SDY1qpKYDOk0e5
mbeJ7BFyq+UsSRempv02gRNJZFcBOvb8L98zpS/SdPNEN0venQVlbMAHj15obLof6JKgcCUKmc5k
F0ASyP8cfnxZpn+4rHtVgHxSXd9Y9mOPNC3agpyAAycTEArAit7x0A2Y0fnUVAo+GhOA5YO3tcqT
xAfknu3M8j4bi7bpNrkuVJPHmM8wJVry/2LCl6QTkZIJxvps7bZcTLTGeuoR071jkWo1VYS829sl
4yVOFRUSDeJ8MrKx/AdEpJLdsBaT0IpZegMG31MQKiRAVhl2qSxMl+vWIi3DB34y5pWVtuSvPyHf
AwFMB6jK0FdeSncKZy1mdNxly0fDxmrCytdESkmy4QblphFCYINHLEW7MKque41Z4ATsQRnFRIWv
chFC58gA6xITTjDjiEQVKsGyQWBOQHzZa86o9/dpp9lgV2fjgnBIfYa+vCMnPa2ZWII4YQhewJFL
Pl9ylPdrf8THqlJwzOeeGXl+yxhLL4ZlbB0vuoZqzvvLceXQGC8vskkHSd6zZPEr/60Wdx1QtjxQ
hv+cvv/a5trXLRlzlWNkNzmhcb054bc7ZUMNSpZeNIw2dhdrIJJpudp2edWH3SXU8SgYiTF3LS94
nRlUqdBzaCxuKFOU1UzW+NC8cJ7faBL8nX+5CZn7FKOnBsecmXMsaO7flMgSCj2qfFUOt6nkjy7v
nwJ7/WcpaLphLpIpRA0MWYUfY9xy5Mwf2Q27fuBjH/Wtx30EMTYN5/vRfgpiQWo/l531Wq0aV//a
XOeJTlM0m5UCg/L0m0cPsj91wI/qIZx9F52lhdRH8Qt2pLzy7Dcqo3gusR0ylbi7nwEbYm9OsnNG
b2SEDkICHoUV3H8bb4G84K4o9eIre0RvQ4vsy3/q4/Fxzs9/FGE/ms55+jHuZYucPNk+YkXOxgaE
w0r5g/TGYc9mWlXwYcylAdi65K9QCNrq8d1vOVdjlNXbmoW7kTJW+CoBu1GNdRy2CqurZGf6XdAS
xBvTB8UQIzresXqNs1E1mK3gBgpC15F7hCthdp+EOte1ab/2PiyBPfvSv+8SFfTu0R5NyCXq3sDu
pYLlRQcFJKAlR5CA2FbyzNYq+kVivvXHv2OSPo/XTjBhhQqzH4/N4S4uF2aDXQ8qYWauiS7uilJ9
k0OogOijADe21RcFEl3qPITDKZ7v9DXPYiO1lHEMtBDQBUFqUj2+a89ZAcXIuWS0hkKcgakUFQsz
5tLai96dShbN0ETTT6SmT2IeseskDX1NO0IDyZ/FeA66nYau14vz695V14oGRzUzb04S0upR2j8r
+bGseUlYSFcKyqxgEsxHeBrWQwbr6IRZwVrJJPHgJP/XbUW+CK07C5TNHiXWTpcD9kt3Sh+Nrrtl
1fA1XGhQ+ApJwPL8y7lKjhBn2z2nP5xH60bC4CL1jZEqewHixvMxHEzxtOY1mkQkVvXI1+vYoWsp
KJVFtnQeczQOkN62j73IeOsfk/dV+smyFl+ojFnbTheEO+FmRkPSx3ZfN68DZr/A965RObPAJAll
wsbUcM48dk3HbHLldohi31Cgnkj6uogVs9PMWxY1C4VKgtzg3fyHcW5NZ4IQl133qD9+a3BvOL1i
9+zWb8mS8bms6+ovWLr9M8RUrBfs6f+wjTzp/DUcfM48rPNfEhA+0z5phCrDWO3IBBPgmNXF4fNl
hkobDXo1C8NyjKGSq3oNdKlb7vshjAf8+USEqtiSE4ZeAIOBgIAtJB3uLBmLSRSR/NklR7gYv22X
/Z57Wih6xz2UnpXifRfTbNIoeN0IqjELC/aymUc1W8Cc1DwAeUvffJJ4gCNBaGWYv2SP/q0QMV66
gXlhKMsW3KmtxJC7vwb7uPfXcsUNBpZlghVLL+lLuIdDabrzqP4dAEWrsvvISm/2hS54d1j3WCN+
iAqC+DgMX5XsnJ93YDnH4d+jV9LzxZhMOMLdUIhW8WTyOIJcLUCX4RtB3JZY7hrHGL2BHhg9s8KF
cPQ+ynD6mLpF6yQIlGz3JLJ2z0NGU6hN8f5ywfxcNhlrEyrUgmTOWWlQsvWhBcwXSBseR7dHSCJx
zbgDqRU0uouqQCrvuqnUmuLI6oWlhOA2YgV4wl1dGBd5rlXCfMBWenlYKYRLn0kckpHAXizUS0f9
WxtyLQW83h599k/hgsAnRDAMnAXNgzanMcZYToxJB/Ws6PGJp908+Vz1au7yQiun6rbVjJARAWJh
Ps9sC0iSwYcKkMJEXB7neTFBmqN0lbhOV0Y/LR4amd24XgGRNDYpj1KxdOk7JOu7Al+xgLEYqci1
Ia9jDjMpaUMHlfqhXSzM/Ra+yZZYCx8OdCJk8/a4xatfApQNtPBBWKkrnfsSBl3xILPZh6V/dYML
4dSKD+Kn959kpoYZ5KbKniZdzAI95hjyuejlECy9tCrthP6AzjvmWjL+zgNER+8+i3Agrifd1KDl
cCO3QjMhuF/1mN4Y6t+U/ToyEwO4Vg9NTWcaFE42QihHudqAMW1ehbiIyzKX0JkwB7aULHhYMBBn
LMBbvhVMc71VzSZoQBual9ildGD1zfXEgViNcpGfOyorsykgUPtRGnrH3hKW6Iv+gqw40Q1YsQNZ
zzdBwUbuLm+aQbQG/+4+Yi5X07XD3y6Mivl6RevoP8bM1LSV3bM2zPREwXqput1FWZwJ45MwykOo
X195/ilIKk7ScDTJAADkJGCH1B8sbM/J8z7Zw3ebBbiXmnDsRzict1z04UPpdrWegPEhKAA2SNyv
nnA/XWVMJDtxmBwfR21WXXH11QEjPzx5AqUbP77zZSMPIscip4M4aU2/jq8RJyEGhAyWegla3rwK
MjhsRhQ72gQQ9nFJSb3yViJy/F8bOibslV+6hWpu4C2mX5wwHUg9tOe14XRDXtNIV8nkTEi+0J+d
8hCYCBmk9+yhhFKfGpHinONOsFM7F81gWtX3XvLBSTbAz1hzCTKvlNghLCjCofaLNLYuVhlLN1Pz
foIQ+hRtkBUG26OmUG4hDWUKoFPcxuy9PK7ZJ8mlNxo1CeUWz9vKDA9IHMXLLp6TKNt+CvF3bBCV
fAV388dlNg0VB5meMH+zrzKxKmKBqqIl/q27Xcos/xaxiW3UIWjdWLOG45G9mYPsCjOzoVwTXAH0
G0vkFl1+ax1qJagabcqCZg/sVQQOvgaueea0n0QPrwSmg1JqYoxrKynnCui4vSoGOOcD0quaBXBh
9aD+grVSW5OedcO3VrfbkwWIr6DvCDgoSoK8YJKdBsNGIZMn+sAeJh7w+mWPaSvxGXExSZADIR3W
kUzP1Q0xvQT2dAtrqm5Z47GN2enXDjA/Br/NnNUwLN/3mbYQ3hzTUhDgkiTso7E+X5+PlrliV64h
dg479VaHxwi8iRddIyKPlRmjuG14Qw04JOZPrTKBP87Z83METExtek83BpgFnwk1XIjLnJspvlML
+DlXq6BKaYNDZhhLmlMcd+vnIxRPvEzVibfSvvaDoG/kzfkUZ8AnYWyz7PsxYQt0TOiia0HwUsLd
V54MmpcVRVsJV89JWFbK7wqAsbu6HFUFZFh9NFguoUMoCb7ZOAfc/H4Y6vddqK/c7yTj9IvWmXEL
8l/PiDoRxbAkIrIr15zMLghaLDEDT1jlcPTSIeZjddekpM+EYtSyRzs7Zdw8QFq+kEWehAvVv1sr
Lq7ABoGVs8vZBVHX4CSc0T2hjiilog6uqhEmXF6abho3Ogh9K8JHMLBU1wY8M99W8SpGzQ0njr/Q
8z+5TeJWzvU5Mo2l6ytF7T8ESqB0712FsB4BquLzRnZ8blDBHuQxVBuLLK8Qrpzs+/JyaZM5/r95
c85Rk67RaI/FfMNzVM+8LrwAhhKqDF60zLmblLXJ0AfykGbabElbpFDIcJpIbRT6QoLfahgWW/9n
V7BiO07+ucJ0SamRFNRQh6mcSM83sqf/ZYCdFdd5CsmTsVfT20UtO2mqGYkGvKi0Gb50gGtyUWIh
hbvHBWq+/86Me2WucRobOwE4W9pxFFhJUwYWUPYS+dtJO0chYinzv/TDM7m92+PkxHGBQxy+URuY
60JOlLFHfRnyu+wUnMt/2xi500wcmR4uui6T0qKrNCLZRZQaCz+lK7crwIcAOMXC9muvMRcyyuM2
h+rHeOipEo7oLAuDoZoiJqOju7LEGmiCtBhRW8EQ7Hvfm4cqIFvPMf9ZSMtSNmJHmg7C67pnKUEZ
Lr75/nCcAYPczbf73jZYrSuRjtHGlusQCcjOMkHsKpoQ/Ejzvpf6IVFtf4QDtZ/Ot4g1dNSO+F3r
PYgX5o7/ICkG15FQECKGEHGziYU3Isqaig0gBDWbvJakZbmpChFvmdcC7lw2HxaXA5+Fyz2BDK/L
+A6iyO46+4Ncicgd/jSg9QJUrgP+bsDx6Scwxe2qXw7BSRwtTdAusslkWv4+Jg7AjTWKkim0K6Nt
A5TaJrFFWHtkcobwEPQ1wG5sycvw0JYWL1Qd6nRcs6YLHFEErviD+iV+RfzWdduIt4ERhiY/LZ2A
o3FmkdoVgneOwz0TIqO75oYCyu1YkSZkKdnMbIxJPG2YGdGo8JySRkbgxZ9oHD1Clkg18f8ABrEq
l15ZZfCfjd2JW1WJWaYtgpDJTve/TGduDgPWPVCBp6iPiCCPa1eS/Wy5W7LVXROERQhjGlw8rEC+
Q5hJNWlE0/o2s3Sr2+QDG+6nY5stAt/HzvAsLY83PObVmGT6og+gxxQqoSTbcJgJRT3lhUgc7pkV
Kdp5xCFJWEmWgM6pj4TeuOfq1NW9l3zPhIrO12PWtxcNuCPoMM4/JGQObG4NY/0W2KYjb9Sy2Tz0
m/yofPHd92TjnNpWeiS9WLn0PTIfT2x6/jAUOpp4HPxKodaCPzHrg58/51/kHzUPX7QeVD8Pfax1
Ar7vcimiCErGPJ8CXB0ugB5A8brs0iohsqxQiDCTKXZUgp+Eo/oZ2RpEiDCsUw6ls0qUwc5uFSMW
+Y9bL/j+DApQdiBtGHMx9BfsfXrQW/W9mQbjBfwsZC4mpT1JU8DyH6MMY7XA2nEbus35qleFm1Mw
0xPJeMIGjUc+17ONRnSpoFKiwpGaxCD3za2K6QFqaQv/+4oC/pDlk0HOsbncSZOMcusDuxZ3sJc8
szcdI6fUJfZOiq3FGDphiAhtYxEUHiQ4kp/fo1jOKz/PIro7iifF+HmJvn7XvD1++RW691GElYiW
jhYRFTt7LaCKK+Vz+C4azDi/wK1OMYpN/1C1xqZDfyGXWW3bwnKMF+lvAyN9/cXDyK7iLIHU3XaY
6J/fTlLbiHKaf0mBbF1/SoUMbZFVLiL7eAylscpejPd95XCmA78LguopHlKdeLTXNOhPdN4zsnOJ
x1L6+Oc4JPwFntajgMpGg0044nKp5Vdzha83ZjZ1YkN4jiuvy9RFWlL2r9rffLiDoEZhyTZunntW
iqJWXYmpdVQ0KzFrdDWr3r3/ZYocFHZ7XW+nveRs7AB4/3CPEgjbL9HAGnsTNCoy1wkAu3r4dwLw
hpuV8vTdop2kemX4ezqLMHkP2X/SMhPiCBQ+dftl3akR7Fq1xxCX5eP3Am8+z0MCY1Vs0PfGw4q5
ZwQW3VNbboe12SlT++InDeFaAlt8rm6EOU7coDPLMfnJg4KRXYj0mF6n4i7+nPspmXh9+kiTiWuK
lLWymMxUrnuUmauKH/5Av0sc/bp935KJ3tdvYbzUx5WNv2FS5dOXf0Sc8C0lPXeMfw/5OxVrOLrx
P0LQUt5DmmLc9wdnaJxVa23SoVPWbW7QpdoNl8nucne90tmLAgqwDMo29WQ25XdJeJKWsdfbOTDt
C43c66fXomuuj8bT64s0xwi02cRX/ddxJ8a6jyzj9Qej6JtKWr11ml37kCUMGItCxmkdOun8div9
vhIszPX0hoL3+dC6SXmwfjoLPGa0ZIYorplIhL06/CYzjaR4JiQuCYMk1+HDfSMxrPUSCstqVg9W
cmOIjuuh6Qoiq+jSOzYpFEo0YVLzMtrgYe3w49OD9wyzulkygBImTawgNqNsj7O4Fn5qkldjxCP3
APh6zBJs+0HtDkTAXIAjAGDP5FuiqaifImfI09ccT0QnIpVhA0hjTFaNfJ0a6QYq9GokxsKTxNE/
TPtuFlaxcRE2tg6VhC0B8R2FKzxTXXb8zJZxi/gNplqCUMEUPnonMWaxaJ4AyP+4Y9/PObrucO0Y
73jVTbXo6MaRTfiHb+IlYMvP0s8hbhPGVY4rWc3b2vAf4vBBI+mqM3TAVpfUZjOGouI1J6z9AWGk
xs3rM9VVIlXEo4SwThntY/DTG3xbyKY6uuJnksF4SSd2OSjMZSxKyZq5WdCP7RbqCoCQs8cLWAYa
Kyj1u/Ql85nOKTUXF4tKMBLdy48wBWcBbKgeY2dx0pliIe9rYHfzlHLPUFqYuR+CgX+YhLirw1Y+
MBH+R91pfQyqsRacj/+9y2G/eGPSSSxFRap1W8DhQeFrwy+8eP1jSANvWrl3z3Cj1iR4yVHRTGcx
3Qvz4hv4SrETC78fw27XZqeZpSDli9FaU3yDoZjsr8ogSDeuzJuc1/2zIsXbEJm+awe9N9HGVi1Q
sLY9wFgn/BhtXrPZp9AQazLC+N/wMLQ4fck1HZ8blJhZPRSh7dTA5/FzxvnWpKS7EjAyN9W+TA68
vDtm4jJtM9qFY3/s6dWlygqdAAG/WBA55sxWLI/WIJYmfh3t9EYbKXd7aLOiKmyTCvG0GTWaXmSM
nLenqewAz+k928Ey/NfOvqW6Yvdt5nGFU1lJDBdqLoK/96TFJ9KbTMOD2lHI77RzZmJ9RzOImIAj
czch29TOM+xXrePdC+xZEpYMFr4oRy4zxx8R88mVXMzJ2IvjmBAKulgcX2hnXZFGpmU+jCz1BCrp
Jwc35jKQ1BoKXaJz2yTINeVPVQVH5cg8jiuqj9ejGWM1EqA6XlUYW4D5SPoNIokQUsqHnRKbYDCp
VEcMqZ4s+x0ncX5CsH937MjX2wCtjXAhwZhe9qIqp1QoqBVtQR2VXicpC0LlyHayE+GZ/GxfzYfG
hp0CNHj0IfPYT5UsJ7Xn/1pQZQ7116Vj1jyBVMCr3b8sHS+NpFE3v+Ebp93bMF5oiRc0nhyYk9Oi
ZDkUjnZBmSApn8JtiHr5ZxtX+A/jKtbfYfU08JP6g9rRCbMQ4Hpds4hhK/qtrkoAhzVpArINtwDT
7slxsxw6QQ94XZV9z4N4PqsfMZ3gla7mooLkGL4MkI17KmUDQcUlPIdzGiNcDdYP2n25WVGHlfy3
flSgR2Q7NgBJQXuOcTSpwzAHbzQ35ASuf990IW1QFCQ8nMdt/X7rmhrOrDAzqPsFyPiWwJItQcn8
cFhA+RqLHwRFB2EJDXtv24SGMG6mB53SvmNEOcEJoP6NbSHIO/t1urXvgsPztcXMcPAqJ8PX7FP1
gOHVDKU2QgGQHNPRhNvFfYawVaYDCTcD4SPP8LOdTTPlb9JxhcU16oBdTow3wd+ptcwVFDjNo5Bx
Gi7oIwdfY4VdOwvUknvk+VmIhcYihAytyCTulEm+u+um1qeMbUXtpkb9dDgsRBf1ZNis1boT9J1w
wQt1EpKF7iAjBSZgF3csZyaq3MGSM0oueonCJRc+Yo36mXMsK9wy1FayPUNHtplwP8Uohd0KTnUf
T+Nm8BAaX6EFnY9DDkSA7ytxr2j/IZTiQgz2mEZwsXwfLlxTkM66lKWWTNcwvaZFH9rEbenszkT7
RfEeNy1h3mweQudyMnUND/505XyV3eYBnrsfI2e1Rc07hwdIYdnLhD6sjawZAxIARrW8HWYVJwfV
ZY70IVAgo4v1VKkWhHx5FBPuMEryKFpJCkOD4JJ4GgVEtukijrejU3lhu//6iO1mS0327oeAlwdy
Fq0hJifLGoQFftsFx5PzIWhSrKg7MXZTdSAOEh5d3VistGJdGsrdP504K8PWM1wBahUGwb1CUDgd
wmMSlUskHMpEW9RDIRfZlr4dMWQOD5gpp7dqQqGk/UjC2PycisaHWUfU3MEdDVstVDL+4KHB9axI
CQwcFEmyvkOcnI0GPLsu52H+2sKON9LaXfZSMkQFiLH2Ix1cFzuV4aN+AuXY6wMBQ6dnFIICD/CR
1EfD+e+9dIELH4QKLST3TkVNkTuk9pX5m0g6S5NmFhqAjpEpHi3dKSVSb+gfIPhyheS3OWt2YH/W
/iExCSQFRjRR/TGxJgQtYbAjvfJRhHZBqU9l5gVXzF/7vt2FvpqJqtzqAaat5S40E8YfgTTZtG/z
8YqCSW9DPnVf/VrjVHnZ3tgI/8WV136QwHdn8GyWU2/4eOPZCo+rMDAcYeLKdRDkv3C2YkzwsCfU
JFCBimA6Oq3+8lr7cWV8qgQndPaptWVCXDwKs6Bl2rcuFJNmda+chxTZ21xKQM1oLKPdJXOJE9OM
BSLMbh4zBo0hwyPVxR1UE3ivWsDgXTUToKR5ZvBOEZDRFiK5GVKidZfovXe1WtbYFYUpAK1CYk56
vs+FfT0UVMYQQNrz0bOg8nwwbCQThkHRuqHFLbs1vR7vAJiMDLvz0F29baMt8RgK0Ug4sXxCHEOV
oRGmplS8vNUUur44krFJlO1es0uGhYt23/yxCcCzg7E8M2uzJuQ3qM9I42F6G8pDI+VXa+XWaYE+
cEL0GhO0JM1jJSOMiVp39K6Y1asa15KvmY5PUedpuwVd4i9uI2DqKkZZzq8p80RVhABUdv7ld32z
CD2pg/hN6DLX8XjctZHPXTQJBOaj+TmXIBqZX403SwbyfK1uRxyWKlIZ7a8Cz/E6EUyZu35BwAqC
2J/bppc/QbIGR1vNjKUkLZ1paIAWEfiJdUIjTEPwTrvRa0KKZBP2GpzxOjEH4+R4oLXe2vQPyp4b
bYMMfmuqMPzwZ5TM4MmBxpUuMNzcF6htHyAEuHVZmhntQ88/Ml5fgq5EKl9ZcC4Xa5jpfDLT0HJM
54YWqdSGMZKl218pb9e5h7vzUMMC4d8397zpnNUBdN2Vl6nkBacRvZ+6aGzVQE4ZwAuOZOZ8/x/a
L3Ivm38bHLqFUM/ZW58pJlLplQB7rX5O2EUBojO202u7J054dDpBu1bNV2XNtUuoyYJmYQtaPwlN
Y02p4eyOWw++gMpnIQpOvSmbcLawmmXwKqPzbZDU/rTb9DiRVtQQbMj1EBebo/30/gvnSAb0G7WE
6VprY13o2Cz7jH2BBKjwBl9aeHHIg/RItvaE6dIkqfSM9cqdfwCuO2/TqKJGeGxznfn+b0jYk4Hr
LpdK8jeYVLsMOSm5YVyo5OPX5ULcR+4+wDzRnFDTfx2z+kM3yLR+mSWNdrKxfzQBrn8Fmt6F6c3J
Vt1lccGT/TewO0FB2Mrqdw6nVexctiTfDcc28FAcIQ/Eo+9nRnrjJYrI0/UjDVxi2Fj6Gx5O2FKw
JKo8FJ6XfIuIBp/WcALFOHvOpPV+zeNA1EEMJvmt8n50qOJKusGOe3jAzmtkLVbl1lzddb3xbtjt
HswQTUPUAPWB4kbRVlxOX8i7YvUYKa/eDjyFZtTijHpxEYyPc1Sx8c1Getgw4tn/olXiQPKrpkt4
4r92boVU0uD4qWzzkIzaQEEi4fSu8Oa/pb+yCoztG1KoTyZa/wSuyOEW7hgyjEJWI4dWsUWCSEti
g9fdbsLrW3T5YfdK15z3BWbOFRdNIvUPVB43McNerl7QY78FpQUns5qcV8O/IVteHtLOzZZV0RQn
9W9mdsftqpQvwI+nbbqSMEb1qvTTqGuwcthdYvGj7JyRo6sj3PfZ6lPYr/fSPZ30BIqlfD5/BV4I
wDx51rP3mkHKuEGlCSa9krMJDCxN92BT8kgtr/zXuDHpycfusYqDH0Uh6FWAmX8Ib0u7efqLahm+
3CLiFEAAD0UYCjeqKOSJqRRqrzKIR2wP4l2dyiQCmvJ/kZa8le+eWXlweofRG2Xv7R7W3u3AxiQF
UPVd65ise+d6fhEbI339Sd7gESSnjOtlzjiL2oNaPlJdFxQHwcorpGukop0XfNF4ILitcgPYzf6E
C0tSFkDDEatvolyc/BXLyznZAs458TliZmqDtgept95SeEX18wZPISxADqbKV3SQmKk1frN25AzE
iSPb2e6foQJ34mEDex00XO+Mt78vLrr7M8M+ToZTGvzuC1U1mZrJ/kewuNKWRwdW+/VPmBPlW7un
aiPevbCrVvgMafPmd1t+ad/6E/lb7kAb+528O6YQL6zWGE8QhH7k/YsoPOEi9D4qNWZSSWv1qDVj
eaOeHhvj5C1VmUinQ+D0idwqj0NnqsT2KEvpefrVqjVucuPHfBn7q6+iL50wJmeoDM+Dcp7N3hbB
kUY3Wz5eOoD7rxDcc02PQXTVGHHHEFWG/kxEmWlnJrkyRF1nLhGs5QfV8+M9W+X/psBT+Gw+G+S8
S1vod2qJlSdcjsxFjIkk90di5KUs2aVoLZJOJZG5zn1gt98d0Cnima5SrQoiMVvMFJIE6l/6ywif
5yhTXdM9kBymmSvt38H6uKNMIyDp3DKYFeVzgIjQaZHZQnv/pBmHj+/YLlJIEX/GLLmvA4BE7aO9
PDH+GH3r0XrdVSmQvlKf+sAtrOcXDIqnqy/OSfMkIFKJwQNS3F88wrHjn3t3+93q3hmQH8pkxCBM
RgcEVbYDEhWnoAnaMf/NTKNMNUqS/7P8Ftmhg+tcr2LQ8A2agIkla6zzfm0CZE7Wyj6WKpX07OTw
VcpB9kexOTBK195KfH8+2Ecm9l0Kg/TimU8/Ft6DZxlCliRBRz+Gu0aZ5xw2Ud1WDZIQguUtM2wE
eSnpRKuer4cGHzhG/Gi2NIBurVIiUR5/BNEjnRCu3kuDJoTE8fDzwxXz5TEJtQDUSkL/+ssf2+92
EO/u6RuxsXuWOJN20RIs6bWaZxngOEOLiTvAOYYzZzkHMPXnRTqFe9ddrERVUVrvr8GuGg3ypAJB
7lKcXA5SmLSzR4EozUYkft7N+i6dSI8EbJf1VLTU1QlnrDXK43PDtxtCYYBrRCjWSI044c9ooV7l
MbCHeGqVqCZ/fpP2zHIwH3YX5+Tf0L4NdT4H++jG/oDBchG+wsjNuY9QJCP6AM7fr8yhkqV6mKdL
rSdHyoUQjx6tAQ+XYhAYErcaRV8fbXo5lyjLOXOnwm1QIFWv7RPRoYZQG8BcBIyuKODvq+iygTaB
AENMkRjR5DbjaGZHs9nvj8FChVx3lBUo84C0CBB13Rl/EfMnaNUWprL4DHh1adw8v4z/6MlRfS07
MmrR6LSIHsuXNv8s/hznwoKUMMia0rnrVMUK6tzQ3smekBAR3o/5G8a+WhthojEFrdtEFR0ZLZ5A
89rbiPIaUqedYAtQEo4Wnkc6plTYxL07qioxDbfw4IQ5wUTnP6llphXDjS6oMlCVvIl8/McBsKJl
q7pQBzMuH1giJxlAjmz8Gb8thKS3K87Jkm8iwit/unJHQar3JqhcxgxK3jCh6HE03nxruIosfgIq
mNf6X5yZXlo6u4x6HcBc8VTi5LXUS9NlKZBjQ/cMCyTUT2JGQ/AfpyKgJQmQxfiD7MFJK0bZtVXF
puj/qz5Th5plRY5Hp1SvxcpMObIHu7NUOfxmyUhpVdaQCSwqiGk+WbqZb6PLaFGm+60triyUSyLX
5ZnUs/cUS9Q94ZtIwFBulwvOQqtkXqEPKEWdWErPuEWyNFHIGMYg7grW8kYvqY8RhkMjLJ2gyfid
v7y1jm0n1OjXgNEyUgo1InuWe+oDsa6vzxo7IsZsYpCFsGwRZfUH767BBRhanWkbInC6UYgX4Wq0
3Hrc3AZSckofs1cemGYd7lsn3BXJB0/Speopnv3sbJg4z8TAtAjwy1ieS6Id6vFosbbcQ0lHX/ro
LQkGbnNtjYLb8dGtNkHOKfgXFtah7aodtuPgcIv2fNGlZfiB41ZmHw2ZYkdcW3ZzIJ8k8BckSMXD
prcj3qqk6Azl2KVETMF5M5qGtVYClEIQSWwUdUADpT2xIqUif07NZRLOg/VvYPgzrrI3iX6Kb+Gj
ZHZFTnQzmHNmJcNk5KPTp6hqWhScIY/wcF/MnrBT9gZCl2XGX7TZcDeBaCp40fgREY1v76dvrlIV
i4fH0SfZg/IUCTONmOsmGcnBsPXRJfFXTkfgi7FImIgjm054K+oYjI7WtILRscF/X9UxUgXRrqNa
WEF/TIX3T2iEu2p/rrW5oMYgPNfXOpWnDOi5yWJ2FTo+IOQ89c4TUxdVsMDvwJi+DOzPTbGU3QWz
+uE2mGkGCJNcizjArGVC6QO7r4NlgHiTkS7arGzWePdi3IAwg/vUZkB4jUJv/29GJTP/8BXsN9q1
WlsPe/jhZhHq/bLn2LAnMExKvZIFVa2Olo15ztMgVy9eH8iZieycA3xFQAW+5qubbi83KNA7OByY
wZnHIYeOrE0uV/FDXFBuwjJV7ISjfQzmVNStmyuzB3HQMSttl7k/rFwSSedkJIiOqpAzove0Yy/j
NP1GRwlu9UJ+3tD1Dp0XOsUdEt5GU7HNBvhpJm+a0BGyJTOoVFzplVfBRJDZ4kl68QZV3nZ1nZuA
mD7/dEOpsf42+7WSbugk/bNYODyXf2OF+zcg2upesteafxRbMbkHpUE/klC/2MSasvVlIwHgVpvQ
FlpPvCwvA56sWkt0rxCNfxp9ud9cspz7kfaaiUSVWYzEsjmBzzAVBM1Ztn4ElKzoWT+mDOBGlbzX
jb0nNanlcXvr2FdqEdnAq8y0euD7alhrFJp4tSw6h8zB5NVe0fR/PFe6j0XI3TgtXDW2yMYBU4AB
UnkgiEO/1xFQsfL4WlTDoTgFlaqYQ9bJctFFcC30L8NuB2gP121RoPCGtv24oDOIm67uQ92OIqLG
DdPUiyRxMcyMlG2FhWQe/MEUWj6YJXvNkmsKZMvlNaedc9DkXB4BdO97I0yGMKB+MdK1ID4Mi+GW
yhw/j+Nk5qx0oijEr/LkDnIBfGADn5BvpwsGUr+ImkFJhUBXS4+To7NIyT8zRf+VGc3rwdokk3V6
Y15UhRZbZvW851yNGhO7Tbg/AFQfRT6WU7H6uTcxuAOSBfx4I/XuD2C0oJ/jlDsXKWysgkQwPO4C
uc3QfJsSHIH48duGlorPhuf/dI+MRPZynfeXn0D+8dcyMRwybAwmnpsE9riSjqR+5bWLr1FYxIQe
dYX08LUOt+m8Jy7VX+vT+TovzNO+ZKlwPOrQ0VwfJESYfi2P+do7cpp+/LFdFc9uO0gYsieLPZMy
IQ5T/J8n/7ovn4Bap+GkdLWW3640b7eMEgZB7tIYUmjI4u3E9nqnKHVf4u3zvZdYND2ow4O6R6qf
6CiP+tAzdF9g7M4O9fNFXTOsOQoXY9pR7HqvremiT+zoRDyG4z0OTTRVDki6CCTs/eVbqnJ9aT92
XmrRf5yL/Z/NawslO0qw/VIfTNCQ91HNHIp2l4tGSB7tag3kWF2fOAkNkSCPw0ywzUEA4SBloVgc
I+Wx7odidU/YmWmDC+qgGnIxkd0/gdjv0ATQqqneDaTCV27tpwiEuN+yrxMw9AoOXympQ4AWtXJi
6vuUZHDNqbU+e7xj3YMTzVHpLa/qzN27ZvNjOYGYTLfksNwQJXz+PF86SWqu39ZpVfcGe/UTXrg9
+2RxeK1aK3esLa+DwhEb1b0+MsFMRh6caRmcogpUTC26f0G1H9d4PzQrpMGU/nuX8hD1UyaHbWxe
XN2Rr5N/7lhnxNfOEwN2jGJBUguUd/6fBwggw2RG78qq7OxPJ5cGWEaxX/YVnyN8IbSSdPeQUxjv
d4GwveZDm8b+tW0KGYpgM01i4WOS0MszFlCoFnHiuvVNufEvx140KH3u8Llo5Ka6Zj/9LxApylXJ
+ozWiEc1Kj/DOzq23bbCVNm80X4yeJ+Vfi3LBDn7CHxOKoAz/QVHvCdEtopBDwyBTGVOnrMKYafc
g9Dp6WzGzXg+vi0o0FlsMarMM6Gs9745uTz1mg9D2FHh6dvrl7sPXkYBZtOnCA6RInk8lmgnJYSx
nHexFzS/EuRtLFkku08+aYLG5tuWEkAw4al2/9E4p0C0MI6wXSTBPTnAIMKFAQp3GyrvMeBHhWVS
GyLj4SpOHK6tzFr5uzQd9myjvDpTCJd15Fh8t/KJ/UadTM4IXhtZBQt5Q29j8UeX3jO1vkxjIWx4
g5WEulLMb4gxOt1TQX9wpptIqGtYpf9bx3bByhnLqEcJ7bcq1nMKlwan9lxQJ5aiCix5bn0Yij2y
42GYnK1qI+tcm8gsTFdMNdFsyV4DDbr1ywdKh5GM9VKbFsTF0pUZ8YFjTCma4bge20dwmlMoxZK9
DtB855rQJqLy8aGaXgTrC8A9q2NyFr4TGAcjS4wdxbg4o8G06K4oN/JwIqgTovxCVr44FfypeiMB
FAUYwg+bSaBAD0XAcjI4QlreqmNYxT3uM7JYvwb82gI/etoseUoPQPSbOkrg7p7/8HHAEanz9qE8
Dt3KjBeqp1NcYuswdl4X/rL3jU0bT/Jeunq41nB0Hz+ADUEJgFud9VE1mnUs2XBB/KzyWA0el56X
nEWzIFVChrGilMXOkVcXjDcjURotAh8GYL79gvAU9/LKScqoUwt8TuoN2+98cqrOcXsSFE0J19aC
w6FEA4lNELWW254SOkY1yry7AD4iKOxtYXTYDRtvXaLey0975qbrIkejrm9QA/MPd8q5Fk9NRYRO
IPAKMZEAP7USi8kFCKcdZXwU5lIEnziEXIO2ystk9LhNLxJMcds0lfhiBAB31j/8OQQIRUdHQ7pF
qtSXea7nogSHyQaYKpnZOXwFhfZ/c66+07eobkazmt5xuwMe99Sl2URfzKyJKQ4WVc3VCBSgwSti
lIh9CcoAZDx7KP5aCFOKsCTj8S6q3+vGSd8v4yu/qcGMfb0F3kq2AUN6s1pK0T7W3yQH2Z5xXCHq
thHHljNhhKYh5EbKYBGa4gSmObrZCpTVpZ3QLMFWSfkmlwHpD6M84lroKjU97mtEmtqQm4uCDdQo
jaP1BZge3bqDVZkiEdcfUYz72tJ3ETuz6xIJT0/1SExjQ6o5jDWqkxHOVGSgLWVGg+t4LFOvrY1u
XyNBZU1NO9VOQhD9aBMk0VkdZubB4sljvwyUfb9w945DrfZViAvMuXzasf7RzEO+BcBsuDu7QkBk
mvvhwm79R41lDk1nU5y7oZT7Zyd+6TlhJrZLgajpiHkO7tzrdzkGYbTUM9slb2V7Z1Wg9zcNc9KW
YPs4FgjsfJFImP7+I/MYVzKrJ50Moy2ACUW17m51LKngZa2Wbp8d7K/dVguYT6c2Y1EIdRX/dYD2
RPQF2VV+Th5Y3lWOA7mErsS/Dbo5mD9OBOl2ygpfbItwGoPmRonKHm3atPd7w+D7YMnCmrxJPefF
9lbBjn5xRAMatjnlAtcHIvMycVRm0aMYVDNUiyySrDaccmdqyrDIYYpSUOttz+wxpbGWZ7ctc7OR
UUjIzn39KeE/JOBEztvBTZstVMBvEVijp8GGwdfGPQCyj660lITpEy0tuv7nGIZfjNYUH1qttbXv
KuMyS02cKVSX/+f3GXNbq8C9kmQV7+CV2bc+2pFJuxcInwU9CGtD9+hRyvp79T2pjSnSF1R0cOTq
MDwl1Gk1YUUvyilK5UsvJtADJByH37+vOPbtgkckxs0/u0M4eIJB/KSv0OZICVZCF7Pj/TOcjNE6
v+nf69IZaBcqqWa/pzEFCb1Wgc6V20X4HV/8SZXYQ2mdSReAOCpUaRouEQraYkyWUGhiR9kH/KoT
Ghj1cXgwtvWhZ9p31nDQQpMi2GwWWAnfJqdmeFNW8EzLsfw35oYIObKYn3j7R6mxHoQ/mYkWieD9
7BZ2o376G6mZ0+ts4iwc+36etiOHXDkGD9Y1qbzHwYtQkk99QFUHNTPGngO9v7LXkomPMdTn7OMk
QaCD38EnlX82uuqOBtKbFiPpm+Mu+zXtIPUaPZ8YSrGVsgpjfxaBMm89pLikdzNqIj9u3rzIfofY
uGBC33RzrD6mRRRXhj+AWBITFJNUVNWXBC+3zDIG8ZLlVhYZhk6JQoKfaMaiZJTRxwgEzkErL3D3
CDbCrJ6M/qNBgBtWMMqPtFLBpmSOsmEQQLoVeBbhIJ8+Yj+Rs3U4erUn7ItNUKndXe2YBT8mNmsM
1TIrMKEOCUkbw81jlPiovEUTfqcoijumQdl3hjTrEyjSxUGQa3FfvKgl1DwIdvsJTmQlrG06zhtr
nOP2ZNjtDsIE/KtZngT7ugZW5N3s7FSoJPjMWYVbbMtvXIZeN8+59bypcaJyJ2G8dRrmz+npzwnP
jK8gdp+/pf68sh9e1chGxjGgA9ty9xb2Elk30DniaTq+WWABm9BFZWAY2AuzMMyLzRogIKpgG3ki
RjrBaIg3enT8UD+4tGh/lKhYfeQfP1xDQgYyOBgzlxUjQCJPi493lApveSoFQK4pobtuQl/c2Np9
ZdEteaZkREoGVzRlInCxAfBon9pRW9n4E8SMLeBGpGhXmX0p/oGcscelsMLoEJQaY94DPxh1kb/M
GFKjt8zvRRmX1VPfd6nJpH3wsT8fZwdEnG1pdBkyd1tKRhM64APZ71cVbn+/Wnf2mAppTXVxPNDG
wJ8nXdBsRIdqu8/Uer4ry6Te3r8jj9nByCeiKwGhsNpjMMOp15QF+wnslkdWJ7mPbDcPwzBLDW5b
IySI58xn/2Iw4r6fWXl6YYwfklWdQwuOanM2WF0mSLJyEOzuIxuR+20XHslhBfbJHr4yjbZrxr1B
gwziEcJXRtOPJkWtQkxxTvHpQIZNMye+7jqfx4dGFChKVBQI00ECh+F3CD+WRn5sQBb+SgJd+CeU
wdqd7YL6Xgi1+zrZCT29fqBUqoFSxf9iAoZ0a1JdZbbq1R34Y57u1dvMp0JMUVhwJD+udFynLChC
qewVDoacUMbWWXN8fKM+AfDUcguhbGGN1ZXT0CszrOhHGprxwO+5vCQ6w8NiuKV6GbS7Nir2HkMF
QoXB+RN6yFc5Ws0vKGa4ggUSMZuPSFUVzoR0vqXfTjEBN+3SlWeVJJ5xoDRzk6WFleeFLMp+vcum
NKfwPCrA6etn/qcfQMUs9MAg08GigJjwIq+Up5jGXzr34yTrEOlB6O2ZU/Y4ela3C94yarhWudsK
JoWcsA6eu+/B21bJhQweWqIZMFPH5yzg0UMtlOyK/B3PQ02th5zz2V/gdC83I8XH6dd2V4e2HIpe
0VtNjvrI7RtCRFAM+1vu8A26MBfONQaSA+qepsgtWdc6wCuapwpMBaRlxmp4AZCPqneKN36Y6G71
eB6gbFT0Is6j/l5OJ2MUfoy/zCXCpwgzKm7GiUrRstSSHBH7vpX6eX/HX15srUiAbU7OTwDdcw3W
VwO73/S1kj6G4I9E8JQGjbA970EHgxudfCyaXCpxjGzI88C7AKUwqZsyAXRsFrxGC8nq5M06lzmS
fWjgUGEknHDbCZig1AHRHti8p455hWi+eN/+iMhfe2XQsTwhQt0yZd5lrqkZVLaNB2hMGDxVhvED
QSVPf0lnUtDGTYYcxSqIYJ9WBmGGfKZnAxctSvWcXXExmxqVsMXrFdbMN2OPnWcANQN7ik81P4It
fPxW5bjRAalZMe5OHE/vQRGYr7cPuI8H8cpYSRksh5kVuHx/YLRxFji6QYoFXjKCFmvjAylp9gXc
KAdqCegp63RY0C4mim4jmiYONJUiRWOetP55EMmvHQklpvlColWcEGN4JaM1w/h1qIcgNmwC/Aa0
WqzjQ96eo4Coq9CGuJScFjvBWEoGH2EvCtGsyE1EmjhNqEz8hE4pJgtxA9rFVabNpkaadjXWXHEV
7jYAXWuiNhiLDmxBqnvTdjEOn/qJJQsD5V/Wn1hhZTeZdLbLgwTWxV6jUSuYp4NlrMHqc7PBGSof
voUv/38+IvMISiBr4BIG20W+BGlM6wFb475RBPlfTIyFGzFJHu9oE0ovKcSPzG44ldVP8JtkVxbw
vvwhyHET/+wVLD4cYWpVGKCeDtaRqSowT2YLz6vSft8UHkwl+7XqrJxTbV+Wp5lJca6u7OaHibD4
qe7DCZcjCdCTEzyo7BYyis3pknvSI+8frpwsVy9nGn7JzWqYVhz+Rcv3EhE2bfgS44q1tjYtKqeU
NXzqTQlvT1JuT6CvCirIOD36x9BdNk/2dGn9sJQpooS3vWpOMNxlDDZdjhofa/L3YfUdJC63bchM
iRtc8d02yZuWXm7SO+ejON5gSkQeIB71ALO46qYktKuYUjEc6A3lQF2C0fK1ycMDeKEQCIB1uVey
YrYYkZ1Ub56Sx4TU85Is3g3SZmHW8AaxmR7AScp9w6fXSOOQLGCID1x5FptAq9H4lznSrb0i2cz/
tVFUQ/DY6z7iq+umY+3q3xZyOxTLL8Z0QhnoLFuDgt6axy9NKdPA+v+Hs/Q2rySVWT18shmZCohx
7GkOJoVbg6pWoMJNqQbOc4h1BljsSdDHlE2XLfWenZk7pLR/jdF3Za5lX5qGWZvIp9pziYW/K6H5
1sfuOmQanV8pF57qKkHNOlX64KRyVXisbEmXX4nKoZljQjMsnrw8ZEPuSnJ0HG8cdwmNoSCQOPU1
+s5OQoNWEFgSm4A3WugsNp2ur4CXS4wkqQank3OYb7zulJnTRUfm1mMia9yrWk6frMk7Y1EWB2k9
3DOg2aabXw2L8leGyD8mf+Q0Ta/1Ug8vVp7wDLdUS553s0zTBOqpMcSwulPCYlbpQhzgxYuyrlRV
2wN2VRcj0oDhmQuxpyq1B7T7S0ueGZohdsmVa9T6ggceC6Y9gnzsuMkJvspmie0qYcxtgi/ab7+d
SfGcImk8npQu1EvjuimzQUDmNN04Mvb6YqMaoxffzaM0AdyWKehJ8ST/viZdxyKXL6ctLDXYY0mZ
jOdGsW0FKhPt7booFOc6HAI2JezyJebvNU/+wvAo8tJny0yMQjUqAykSLbvFPO/rG2WXF3LatFp3
6yTwXoU69rDfGhABe/4kUvTqd2SuoxwWVMeMQhrVkxNvVdMgq3ifj+6zj1lonYQE8z6ORGV9xCz9
cPFk2U4sgdmkyVHYVFqXOhmIam6GvaNCwVIg/b6k1sZbP6ixzT8cOa4BlNLLy3E2mmbHzmBV9wJN
K9bo4iDXU4XV/nhMpU4IVyJ4N8H44Glq8ADVkZ3g02dFprrciyVsGTB6YWnfjim77zbDmAFNg3dE
k/SCX8CjYiGct3eQZwbo5yGKQw9Bhp6C4/OD671MfpZhb7nwqENyq63RnhuFWjmpsOn8uwIDIzH9
a5teHzh/YgzJEs/j/c8Qk9pAvnHhW0cuI7RO9RoERlAqd/KyTR0h6Xbj0+kedkybqqbwIxpW/VMS
qiyAwOAOp4OdbqJvRWEuZNxIbmckwpSmyHd8WtXDa+SzW5KCSIwFEZqNY1tEEVmV3yf+0CsTsjQ0
qwcFRvdI4CEe1ez0pZ9yUF7unEAM97x8sRtrIJ/DSm6ueKssoE/skGS2r2gbocerig/zUlV7QIEi
XG1mrvTpf9rF66StBSNQzbTt8UQW+bnwoJSMThnAtyAHybWSVBe7zMhWC3kO2/8rtMRo+Dh8vtr7
L6RfW3SJ3hJtnp36TY/p0Bcfs/COxCu1k9yImJtdPinweD0UaAqonNqTmVf4AcElzAyoB5btLnVK
b7fEA09jw5HEhsOD8ApH4BRBHjKWnsrvt2mb7V43kSXiBmtf8VxC6jEqyAWyNulbU168gOubOQ8B
jqz4CfIrf5BoboGoeOcQOf2Q+WZYVVy888PAYFkQ/LXBKcaxhOZrE7l0Ir7omsXsfmfdft2eqv2F
Yp44qcLz5YKAVTCeUOW7wpehv1vNBJ3f8qMnsnmw25NXQ/Pqt3/BBspcUITbMT3m7r9pJHsevgrA
/nhAXWHQXnHLKWOkgCVlLnsv9mnzeRvfDLir6ew/XPEN51VHtYp9I43Z4VpwiRoyH3M51280X6zm
MCpkGmBnKyXGpriGDEhv9cj4fVt+0Y3flJwPEKiM/+sN1HTLf/HZZrrRUDZ3gTzc2I+3ujwckaYQ
a4W+C1JxBC9HYRJBX0+m9ozClOAsf/2A5Ef9hSSL4Hhp9gIihdLO1Pdp/Oqyxeq2zfrUmT5l0Jlm
zU87ZJi5Oy1Ku5P5lfvNivytysalMNZl56Zi9UQxX4jMH3E9Wh5IlSb9N/hECa8azHJN/DDAQgOc
uemKM82mbrRiIOolOnx38og9qg1x6mjuSAzFcRaai919Wa7mLya6MHehzWzS0li2zt53g2uZv8a8
qRpAyjS5a7IBy6sVpX0VHhXjehVA20shryOhxp69N+uZYFKbd/xGuz0pbvNTFnFvmKLpnRubONhF
T1dINhFyJ6nJY2mEzE+W0WtXLX97/CR/Zhbk5Qgpt98fYbhrjvlLhqCPnxqzU+sT7VyBd9DHEziB
UNEBqLjYfhoYRFU81YgHjU28D6jVftAvzqsr2AfG7CPaORpEh/u7fVkuLguuKBgapqcU4nb+LIwD
KPVjxg9UNaZYqDcYf9lZv10cbjWEQOfp5HFmfPy2RJjCRFaknMMUzS0L6ePhFJAm+J3LSZDsdhIG
pvNEfsQxIWf9vRS4GhKsTbn2siLcBOZsHbXprPz7F6bvqA12xHbtCXbRbtR8seLTJKSlhSLmXFNU
XRbwh/bztUz7su3wzUxRj0PuuKFdCBCp81oy+8D9t+go8HHtg2bwkMtMzzF+yuSVncUJ+VC3lhLz
ZnCoEByUx5Ux6wE7qOg4wbTdnias2Xz8jIBrEyTwbOZ2RIwQMNYNgyYWfGWKtA9no6JwSj2G0YYF
0jjQ+XWH7GW29BmCDsFjU3ztyDxA3N9TC7F8EXULzhpIVBIdEh6MBatr3YagQvQMRX6HmDeLIpsZ
svPYwPikaQ2KfnBxjvllDYOYsMcGLf1tJjDQMjulTFRSBHXcx+JSwGOacUxa4MeBizZ/HR/MMNph
+zSqJXfXUPZIMK5XOk0o09RYCR8yFwz1BzXvKF/pd4h/pnQqpi6JP02Ap56m9d4m2YAydoqLCDZt
lECtYwYdxSVwgVIBpDvKxJIuIINp6rY8vTLnzsMGlbXbqbOeHRpEYxW88sHebCTCEqmOeHyJTKTV
2s68r6jALEzPLUZH7yI+wOK61ZOeWUCDuDAR6OADmqudQkT7ZDRrlt3ANLBNvdfV7OYCec4Yjbwn
ja8nSm5KJvcvbQ7lg1iTj8vIxnX/71GITUQo6fvwRYgJCBEKe+XOoEsFj2To1UDDl5ve4lsjfxt6
zbbIlsJN/FEzPR8Ad4yS1fQ7cBw31GOOa3Y/VmO3+/PlbANwT/r8OY20umdluB+WX/LmeL6YWofm
N1yMi0JvHIznSntY+hD4CaWWJsLDJQ1piZu+u2DeW+efgpStspAh5iN3NRXlK5MtArKLS+hujZcZ
olja83qdqkiC0BWHKhjxlObQm1N93LIT+6RLkYFrJMXHQamdq09jdTT60RqrPlCSkWJ+9ggT/TJ7
/dtf6yA6sizah0yjywDSyEFtFYEECVkMaTdBdfIa9zO7dF8prep6FmF964lZLIcqKOVG979cdNp2
xl0TSofbFd8XsbKiFoosm7cckEARySW3OA3xCJ9mYwcT5RPyDLRHi9IO/mY8OV1XWebTKctH3Tie
X+4Y/0QeAupiOakPYvwQkVmla8+Vqru4YHNcsKnzqh7XZSv0nPFBbKJTDq822S8XVhR/CMQriNvH
PtpeCa3fmVeM2reaPyPeGZMdI4lA4E9KrmsItKCtH0vniKG3IFGdgY0+U2/r7juZcGc/aiO7XLaY
KnkxkTCxFtiANUoy9yM+WZOtezX/HigJjwkOvft0pKSgbtahlsVdzZ6BNdAm8KmghfiPQmXEbACd
OtqZo+rBugFLtqV3CNNRZxnG3oc2A1H/nxnoRlKQ5s+3+ifiLqXrVdJPXQsfdmqU+7+4RB3en7Pw
HCFFzNOz2gYGnIw09SXpYMNM6Dc9E90caW4EOqiLpnAz+YK/ssnjjg3VUq8bKrOfPHXYG0lhy6D0
uAf2VIXWDjq0H+X04lLB3oexj9Q1q3Lhs8ciLYll8Mv5+IlRRFg6+1hWjye6S3c+7ZpEeMjt5q1F
ImBrbKUuGVLX1EL1yZbdSmRXhNaIPvWd8OoGfg6s1KL/y450Ts8GQidlcltisKpEnFR4R9fQApLu
VZ+HnDvRf0tW9TMtE21QCa6q4s96YYqBqNX9DIGy/fmVZz1qxd8mbxq+fprKnBXehj0lTrdzkTQV
VB+9JfxRwFMLCrkodZBpXKdH/ITTNTr4gt1KrsxuKjwdbIZrG1FHWwQxa9vHfHFkbrrpLdUZT/Vs
feBS28VKCPn+Urk6WW++Xmhi0WHUuMH8fT5iu+9e+1DKUIvkA9f0gLkzAeYpy9T7ssQcz5ALSyzD
0zxTvmUTX/iFo+i27ggDwgNClVLn3mVDcVpelSIS7XX8huu68IBpGpxoroDX+d6mzXV0omICXWpq
xJe59aI/21YMybLKLN8sv5WZ5mtPHzHcIaa2grLbKmEl3OAtxDOsj8qoNR+AE+TxIhzi1cspMkwQ
A4uOnNmOrHFSSGAV3FoBDbSdaofaqOiIiBqIs/tUPLe5no0HAO6yLBhKar3EpaKKAyg+FhzEDWfa
hAzGR8cAY2bCbFs6B2p0VkQJb8MXMnIVJ643XUDavaxLEqT+8SqxBTC9O4SHv6XE9SYy97nGBr1H
Jo3LzWb8SZdZTM7EP/vmISXLFQrrnNVSwOZERGHo7L0Nl8lwIb4RwFgBmTnbIG4q5kLeKpZxavcz
+gaACqtXhsXFWUJ5hgyf0cTqox1yvz/FQ5tpTY9GHI7M3KnzvaTf4cXbXuPu6bSgY5izO1As3S+J
wPxPTE3XbTa0SnoPqrNrJ2YuTCmFq29BJgTrgywzM2dOc8frCpRC0avdZrfVBgZtxhP+4vtRBDeu
L23U8HZlEHVeRACdfA8BqtAGKZZdN1owEYcY4fRF6QVRnOQvFCMwaxOuY7e7RloRvs6soqEWmd0A
8dQmT5o9pF/QR2SxgfNa+Hikazz8PZQ+R5tMNrLl02MoPhmKLyuLm5TowAUmLAewK19jaPBOa2R+
aC/s0z0CK7PwKMUyqUlUpYXQxV2geKp+JRq1Gv1frzE5j0QhVTyp/If5K0ye0JkG8NRiA6Rfp/dU
VPBZYe9d4rQaJccblX1aLgKqku3wIZ/XX9m6Ag4NrRFrQwM17hUXShefGleQ7h+gqExxFzaAHX2z
MG5QFSFMq9oKExMjJY49+LbVMJ/ZPfeOPsHKKQSIvAKjNX+2KagqytDpeK5dO3VNNzaNjKL9hs78
yijAUWzM26Nt0qy5oDTHyZiVpJIx4186TJmz1zm27nNcSWY0GV8of9HiAqFbgc/Tkb+kJ7LVcM9S
5BWXzNlAZo5RplcAXyREH4Talv712tFTJz4us8kW0EEGuhWFoUZAIcK0m5XM4peHzTHFm0jknDZb
aPW+z7AyxhvFIsNGyn+njShRdIkb34QEKU+LfXDWjX4veS99VKsKG1kFQkYMb0Zh57GKUSW1FXYT
upUsfhx67iTgixnkuRECkgoo43T2FUhWELV2tnS1K2qf0aht47LPtKtafYOCkzE/pgwc1zOFAZHY
OHOx/bbgTbhnkQVN3efKojSn3zupcBCBT+Z44Xjh+CzpdGE+o7CT171XN41T/Z1iEFsrU5qWLUJj
ODI7QNqMUJ4b19FcVfvdXrjf4XmSHTkdN9pm1kbtMR7h7vvTqT4f19x9Jx85hPPaLmyvPOtrH7y+
yevhFl5nAPSzrKyhCdghrQz5ZsjtmeTZZPaFjLW514eJ+FvKUBDv0z27SLlNYMm0mcxIN+b8XCDG
LBxD/Ijmqeg0qDn/UGZns7Cpjb7Obkq6wt733zVR1b8cmDsPMtPkgNeszYkY/YIv4hSkZXtOE6/h
qm91njh9gZ2caa9gWv8gDJqgzF3mZ0XsBuLjbQF4kM6OB31vcNRFsRghpmvNZUC3GEuvenKP7PQx
E80nw9kZN5Xt/CbjspVUckRWHIjcrS1RHmnrnSVTN6cokLhX96GEMzSyA3RGDIONtcEmKNc+XSIH
fheldcVHnzx3vdXqBlr+KoCrD9/uUfJJtgz8JeYyz/nFujx3+4IXX+lTv/H/QE48u+Ve2t4WEBVh
iRRhBhJbfg6vg4+1R/Lf5C61S7EGCq35Bm0/kSodl6UXPrtCB9Ge8M8IgRWf8v/E8zAExInXJuz6
AlE2UO5EmSM6a2T2sDEqBtYenDNbGU6VEOzgibCF4I73TL6xUNvhkVCTWBNsvY0ySbI4hn5w3o1i
vrPaIepzZG5Tc2o3U2z/qmJZT1j3qu9nzoZHC1wXN8gwXeenUtoNks1JIYnKZweOMZr2yR7qSGiO
pRhrRNsW9tWzPCZQb5xGHQIRDKd+7XdqEeA9IUZvQyd06883DaRA8D+CVicp9H5kuc0twsPeZtjz
fg37OPwePLIQLxANbvF8QAiDDrAxLqTGGMhHg1C/95bal+Mz25zKstA1yw7ONwVTXCfZ5KqcrPNQ
omLcbTUD7Dy/Pkz9k7HQ+ODoWBHdpklAIiih3jewBhOlyy2dJJDsQdb84FW7uRiJ9sFnAxdNFWgb
9ieztQFjpuXQV/1FjQxnzaqiFpNH9uyXrrX4qom6QW0fl7ZQn/MNWo7WsVbbwiJyZSqSGotLh5hA
1oCL0XnDwrFXLoRLsUqP/S/PpZ8QIg94D13CQZTXRT8inUiFgzDw0Nq8n5T5V5jLMwZDqD/n4ldh
Y7lZLnrWYAuB5V7YWN4b6V8iZu0QfikHv1PxFCHLIpkCElKdvoseGEUQu7sO+IU8Nr67JcTVwMvL
p0OUqFPRBtoNNC7PKxRdjL3FtNBF5/pMGUZbPYugal6GdpLZJuHOel1d5Eb8zTyoxMohNkg7J2Mj
wrzF6SW89UbTTZe/+MAT6q54+illLl+seF/p/T5vKk7ztV3kRc6zWueFu96NdQaL7vGeZ5vpV4H/
FOYH/9rnvkLk9i6VEWN0aSg4kha6YdekRuUeX999uPIeeC+lhxgHjGM4a+7IaQkzM1l6X9oITjuI
314V/aey7Zfg5sksAuejwQhkGIa8OFRaITTLam6dmVb9EYOqcbbE1lwX9Tzvhgjjm2USxLu+htSG
wPPuI5Y9+XmoOLPnEmoS49qkfen5S/vskFYqdKvrszfuZXq6pAos7YBr5oDzsZBooXCpqjGmf5pC
3T5cyI9swEG7wvhslYEqkPgR6Yl2yH/28I+HmgkwkofROd0tzybq3roapyxdY8BbeLRoJJUtkuNp
CqmotHTFnktdVkpAKknOLva9n/HztOgPHN6ZimH0y69q0Knh2g74i4eVFT79mIW6TZ4LR03SQmqD
wahIMB1ZBvFhTyTHKDOYNFcIEFt6qMaw1bnVXvDNNLJ7pVO4R8kcGua6v1KyTjggX9W0h68I9viq
zYoY8mUM1AfgUeN7WUM6syjuZw1YPnfoR937HyoFOf6xl1vggjIMxmi91pW7nnkggXHyMbXwnLCX
QCe0OSpI43k/7yExbf+SjAga6lP2xc4y5mHnJCI8qT4jZJ1BVGMhKdjzef6gY6eUW0Sq7RytanTE
PqbJ2Pk+U4e35u2xNrXz62pKXuXcAQ7I+hXxqK3YUAUNyuCMBvzUNnZr9y592ufViQdnBlc1kKbl
2b6RmvLTCfVyQngDMojDMFodA+bvNj5drdEfMkqhyIu/+ehZEDzN2qYHThj4S2kkeoASZm7tfaA7
2UfKV0zYecetZj6kb59nPqit3cz7lT6a7IrgIWbE/vU6qQP1qOKRlh+OGCexOmTaJZ9ENQW//4gu
fKhNsvWjjJQca9Gd4NMlNp+UA6VLfRy3/g5sJfg0FRtF4V8KZB0speBi9vg1yyRF7ApwLlpW3Ivb
tBBy7V0lazLmAiyk+uYBmvF93aYrmfb5+hRXXA38UrpunKZEpkW9PRa2C0btEZ+kqYQoiPqibSGl
DYSw1MaDXuUUuG2jd/5sBuYWfwPUE9MXwbfvCcloWIVYpXr3G9GUojrAi1gXyvmFV0HoANg0tBwc
h1WCdArI281OL4JrvQ5z7NruUD583+jm57uOsXSw7c1nLOxvaNJ3bZJutdiczg/pZaZGvyl5cVKR
3DyGEdHvG+A1zssqho8cer/F3qkJCVaWIejwO+g4Yg6mOBEwJbcJxp1oPxnp/gMY8YyeWHrRy/ck
9ijlsB3BLLXp5RxPai9QCkTYAoDs6pDBoeZhAiuH3xWYdFssSNmZIXu65p6HCI1o5UmxWGA2eugr
qcDZyBXzVLg6p+ycKiKCAgAPvNfSYmYxKsh+5K6wPKbcW3/QPAkMjCexrdDtYJKti4xzStleqFjj
Meec6ivnqYE2jK9vL1wCrPnXT8+BNv1p3DI1LgATueqpypVdByuWT/mM4ufLYlTDyAj1gRhv5k55
/Q1SYXH1FStRht/qK23PD/aKv2e5PBX4SIOsiiTbDchYFTUSJeWF0zNstQhWx9vZ2MKFFSjx9j+R
todUB5yq3z2jHjlYbcoEPhpwGyPEupHMSw0xWi38/JsYmer3RRXW8af9jpx/i4VEQsBXww6QbsN9
qfc57Bif2q0GXncudCW7YH6FCQdt0DcdH/IiG640i6B5EebOmDA3gAnMYubaedL7XTtiPfWK2fNn
Bao27I31ud7kxlGt8zZKP6dnj7uvPyuRX3HcXxK82SA8TFir8hu4ESd1CMnL2euan1N4eOMA01gq
q4B8qfx0mb2Jxczxigfdy0h3eJMzEcLaPg6SAFTV9mUN5CvkHzMwiFfKyQGxAj3RWEcotPzTiL6j
/GJuTQTf5EO/pniboPry+XtFFaiV//wqLy0pLp8WGkfQTqo0QgNNvL7Y46OGTVCnJtNEDMwaq1PF
bU60c/IHxAjBk3jxki9dnwuD/q4KT9JiEx9Mvq0mumlFyikT91nkIhvqUfxlX3pOXD5pzB2vQl1e
P2qm/rqP02VQ5J6+f4tv+AiSWeG3Mxv6OaiCVd1GPHZab9MCUu37TOmZF9rwKScAW20hm/nRS1t7
JWX+HnpPxjh8XWjDQCmeEdr4pShOz6f7muLcJrg8MX+62QHJMN2Hzz12r93rOlquYNfzN3J2EcIB
RXsjsRfhl/YRPcSN1kRjsHUP7ZWl0qiG1w4O+JYDF+i+A6C1O1hmggQHuC94DdM81JFoWKDclNv2
g0ER+pgX6iF+9gRiwega36PoHGl0lBfSk8weoOqfIjaNhcx0qtzQ76MT+xNYlotpNFQUVdh0Stjr
MOehKHX3t2a6RqhtXeX8j4a+8h6CoUby8za3GAML6CgpbzZcLPBbY+v7wCefoAlNNGQ1WJ+IOXwM
tuWtVebdGOqnfJ1ii5/0+qvCW51jO4jRfUOwvJQJqlphrQJ1ggHHZJblMPV90Ump/2UsYLv3AaD1
iQ4LPzKtJ9gAv0CNJ252R4+u8wpJRy5oK2GpQbZJqaGCjiF/ny4GyNkNumb1/p0c7eiVrQbVPt4t
qo34+BbS6UHqKSeRf+9EhPCTHv313MrQVGT1ykCN1SvhspxqSGVsZIWyL/8a2mI/NnbxNnK+4O92
41dH8qYe2wMEem/r/J8KKZfh7YFsTbwMQ9vPc4eD50Qyz/zWD5dAyDJAZS0wpVF760ShyPMgXl+2
v37OIoYgWein0rCCoseNcQaaEI390BRoYCIFZ1ElegfS4Df7HGrH4Ov2xw8nT/NaRcfA/+gK3iCS
6ec1IZkJoH32dgNZvPtI6UEM+qCZdmE4Hc95aXPhoRMHj4/cq5bYZubvYx4QN1jWVtZrCcCAmW3U
AYfXIVCA0JESV5NEr5Ae/wuCo+7Ttt9xWxPPf4CtdD5bvhTmg4Q7dTnbC6XSrT6GY4Iy8VTULl3E
raMqqJdFCSu1GO6NpKhYl2Pc9vRi5GjAEQuipt40nES5GCJxbe+ckUfMQY4BHW15BENY6T8nwiMr
4vLdD4LrI4fKBQsQR/36xGM5iYTS2VKmn/Zc4QnTB998t8FxHadV3TJ0s5oA4NBlz1U/Wz53yzMQ
ZYsho5J0bi30kbzicnqy6YKo4pHBA0n8NTqWrv53pU2E7EZE1/qkQvyi/KgzZ8OVqT7k/RXs2ePx
aSGfs96LzjCtL84eKfjmkVFNjH6upm6LjBq3Vrd6h0P2ygeusVdM3qUXeHlX7YgjCgTJ3D42cfuy
Pw9aBjkxiUJDCp0vDSVsuWhJJ0pJtnIhwOTtBthMAkcUj3bRVHtB3q2r/yXoxxE2c4jku2ulhFQ0
HX/ANcbFp/5cmgTuIxbxunn4hh1X5U4IgUxGG3lX1fOBl42yJneaaQvW11JAbT6r3fsoRF4v1/xu
M4pz0/UOaoBb6F5vUYW0LTW3N/mYsOuG9uLABoSC0qwVtfYxVVG954nBSqLDa9XXFUCMx1JnLkwx
FFd//i9yiXbhlt5EMlezca4PZqdeMgGPrEvpq7cITAqWgdDEcEUfMhtz8OCgxY3Q4iO3rAtxoFzA
9rF5ihsnv6PWOTdhQAHb8MEt53+Vm2Z3EI9tFGfdUeyhNLaZ7iNgzRxFE6JVkAAvREBgGm4msZXw
FaY9vBdwtOKVYvG1mvEEQMTsyadwR08XCLgbbol/Kh11hJ4HWei/jD19T8vGikcXAZZyRtnnYa7l
eN27162y3A8wXheR4VOAPGou5Be2pzUo/bnNU2QmGcoFadIdaqxdJwM6WkarrjQwySrV4W/Oh+Ou
reyOOQF3Gqdvc7VUfsGcwafvPbHCnm2xaabiU47D40ReEbKWiR06mCRtudTIbO4zZzf9QdSkA+Sw
QxTQFsOUgldw5msfdIKKx2ZVQo3y8GOWFgUi1V3eeEODfwmUA/aaEuT+ciUSBBStgaslKbVs1vjA
8AMHP5gGqqwuJkHNAgiaCoxrLcTkp//tj7BFPriQNH4GdOwakWdxzWBCLj56ZLxlegQ+dSdk2Mod
dWJP+yj347ggJKL+3VUcWe+v4UMecyHhwi92yR8/0k09XUjUt2gZZRUW3kV8h9R6RqtaLE5dp6Wa
76y0anEnDxLOpvHAqvjtfHq+HOMmXw3itDr91L7TV3HxS5cdfh0ro2hCtZ9odVuHLPoe612bSqi3
Z8ocAQBa8cLzspmVVdwKndaPvNlPbs65kHgYk5JKtuTgDK8ijgIEnzPYeshxof+v9elHBa7R1n8p
GaroDzWC2sGczTIbkAF1120fh3V8TUPdkbDdeOpYSri1EWpDtQXkScjVF5lOm+Lu2fbcYwOgBO5r
SO3cdQzW9Icfaotg4sMy38aakGG5dhUV1oJQ7dkZEvwdmlbScxurwzYycRP7AcZWGGpsjh8zzKpl
Bw09DLvHyiwPejxtcJrQ/6zdhKYuDCtQvFXrmC/hbSQ6i6CipP4FtANDy2BapejGk4iieAoEPc/H
MIeTt8eCb+WIyv7SILfpW6k4oLdrhsz+OTUSinhTjFt9k5sFP5Qm2Q/8WZFtMyj/hJVXPonJYU6Z
EtOS6LzyhPh1sNUrRDfWvrdO75gYVaBOUKAwfUFJWRYoCeedxzSw7FTqrHkoGlpLVB3uHD7Lmnk/
QvlDA4j4hjFPfDvLKbSoVJ5o0kMZr3ACe0bXuOwQi+o7u1lXU/DPzBaqF/a05wxYVfHiMWbEYGwQ
VAMOimaqGlTwOtymxARoTrYLSDLb3sVzE8DN5e3SHla+9lEx9uWv8loHHKzVfsoTa3dPI9hduL6k
JkyOeeDuK9RIejQr7i0umWoqw+EuaJ5pGwXp7Ch/SXb8clReH3Ia1MZ9V+JbMCFXqbrhC/seTElq
xhK+HC57yeLx/9UkgCkFmo2IzCU596qK5+Yf7h8A+Ting5gT9ioNf/vW3XQ/trbkqhcRKrC9kCfK
B0k84EFsaLtc42FonpZ5S6J9B6jjxVYp4NJJs90eBh8Pm8hGlskLRgtfCR8xT+DBg82dG4TgqiH+
qBM44vDD5BZjwSpo/rG5Jc/CWe4nd/AhBUoEMh8nD25IL8A7qtoMpr0kVFB0tE0Fzyl8d7beuQ8d
TBn833gChzJqIiJTZ/XK0ulY3Zb8gseituHlLLiTvsTiCfYb4nILV1wsneG1Jva6XjAUVMxWJ94P
wMlX9YE0DN/FIwd7RcvY2I+jsfM81BVNX8n8Uj5nScsIScR5FYe1oNdQzfXJTX/RZ09yYgvdBTLJ
AYXbRKEKCHeDc14HA+ETwImGw0XCYpQrcAwo8tK91Mqul8WEKoNWUANmvY/dC0DTfjBIgmHrXMqH
mKTfVfN7HoSWtDMLQozLdw9iDiQNKiWnlB284T7JYnfa1kroO3KPkxKpM6U3InfOcNEx97a/3Pu7
PhXP6UAQSsJEIO/fHakYy6SWhftwb1PRmpV0cmEidyLj7FQpzfVAvjtnYWvaLqcRy9/nVKRH7bGx
MOx+8x1IBnJutk92++P/eYOcBPL+iBA+0IJvadMw3WeMrMQd253A1rRZEs8NLr0N6eIJQPOyjpQn
rZsvsXEGufP8TJ0BrjNVPYvXSwjc3uHO7b1FBm3tAI3ME4dKJ0IVZQYlE+ebu1XvVby6JAyI1kn8
/ka3ueWh959oI7LpXwlv50jfbxMYtFmEjdQM4xOXEAB4CmXJLvZubghxZrod9d/tdQ+c4l2BztW6
hJU7+8ELlzBluJgvsY7MtHDXRjWNEwNDv2LfKGdyA0Z9K/YI3k8ptfjz3xb4BSZQPXG6UENMaZHB
RGOKL3P8qYraiVSlthfbljbVn++mjeUQabnHyVanJDm84PmUndq6ENvVOxRRIn5RyUSmGdGvUmHV
HfvIm4mAovVB2cHr9bcyd/+iMS3wx4/l2uP3C8e0yHwat7xxr87NuypF1jMvlHDlFw8L3bBksDnJ
DzbH77lzcSYf+oULdcFwRCmuqAHCd1N+2ecfIQxZrBtKJd7eFQZXluwP7cyul6KowfUVMVXExwS6
lYoYS5l24T78YKNju0/v97X4iJIk2BQQh1GHNnMyWHiwQ4jgpp71V7Wt0lnk4bMOcND4UjqhAK30
a+emf3ZdLgRji9qXHQ47c/OhYYi3aGhzUhAYqK8u3kaZ54FZTPafp1Zr0JSjpya+8VBLUYIjWRUl
FhAKiMEXQqviiC91feqNuVkOdIu2g9hpreHSDdrKlVNfMYjRVLI8vhwW6kvP73VS86vvpIFI12u4
nhqdY/ZArD8u7VwMzJsep2yP/4YJ8xPTdGkcIUG1H+umPUpjoOnD1qqM3P5JmWfQ4Txb7qL9ZqTt
Y9wk796xKldKMk2/QYEa3rMrY12Kk+26+EJGGRZcw9RGUE3/k81k8t9ivWjov0IRpn0C8smXqEh5
T+9W2r0WMNFi6B8Y0fYIe0uyhDIqXL/Ga98UEgBjO1K9WTViF38MhpH7e7xYSt3EPJZL+wmLj9oC
mRkWQO9aThNjq+QBjBqbsjliott1s4mnrwrMrd/Z84wDOQwg8ZcGucP60AAfz3Sz0Kld/K3+c7FU
MMUDwEfgqsH0ySPM7fFgRHqNGrTQNjy11DZ1O7xEosU9ISIKFKLu/uvtlPNoFDS2XbKrW+tO6qRt
lBIdLUrU8WQ/QACy9Vo+EvCSHbxrt+2yON3YMUKvYN68BnqqUe+JHjyKV85mc7FpOxMkUjBczmGk
YvTyFADtvFug7a0IKHzrwmEtS2K4IPTsmmYpU7bw+5DqM3DozcmXOakrtPGK8vOtdJEOQc2pR5aL
gpLJVLr/Toj0SSFt28k+Z5+kx+DjQGycQOG3N64rGkpMl9BspmIFnZj9rM5ofcLD9CcfX07Gz07J
fvwX5ITSLvbJTB7kEmg7zKCHkY30xoeAOzCu9SWUthCUe0wJJFTUJqVCEp+MXX2xFRcn9WgX2n2c
sX7kdSAtD9RKN7WmB9NxT6WgRQIcFQKxBB7g8//BrGRGBlAzUlH6gWR+bcHrx+t1+iPpYyvAjyvT
CVDuO18NV3wfDSrU9HCJBKOuB2zuUtsthlcuewJSZlYkQ3T59uFlh2hLF1f8sKyXnONC9qGHV5M/
EAakoQKmA9C4A6mgNs3hrJavKVCqYshCOED8GoOoFLkHElD6axTre1NBk6I03woWDyvMWrl8l8y6
awpCLVv9s2gmmb1nDKF/nMd/Mi/ADdUMKTtwgWiiYkLChxrMIYWibw+j6tGrRw5Z2FWozcFlXba1
dsHThRcBAYA6Mj7u3mEbpRstpGoazNROLPpf5+hDIUjyciHB4obN/4aZOHL57WS1W+XfIsBZ+EhB
gzdlzjkpjmo5kmgGQh9PHIWCQIjuFLFgaRMV9qh1xD3OBSugg4sxBB88rzQesoNct0xe+j3/iyH7
7bbnbdfipxN5emtKdEMEwig19Qkl5Yru3YL85xL1q6yQkyTznZj08mOCf461BhdLja8uI9hD9PWb
uC3n57HDlFyJXAEyWgLgfxjqjf/tbA3xQD354bxaekwf5Rja6hTO3BBN2NCf6uzvRCLGI0sGqHkR
hZTJNGgT2xw4SVgeS5I3DHkCxc5Cn2O+usKA4at0URQGr6NDK84/vYUjCaWfy2kDrDVoqUrHDiY1
AKVjhHUwcSKyD5am/jHxGg0j7a3RO0/c3SYZs4uGpvs9hhZSxUvnzGy5x2N+vjpBopPvu/FQhiXX
UqjICV1r6RVJJKZQ9sCZbVA/gdkvE0UFBkvCNQsHhh6vy+kAqteqSetmkTEeQMdjSHFbh8tzilFA
szXnWcTZeAhWgmuxlD/df9daUn0dD87mss293OY+ORSoXyToMYbPFuWy3/hyFzz2i/GnhqEmxqew
WyI87PV1BnE28Pe2c9My4+1G8yJ79RAbOf9yijicb07wxJa416iEemsrciPxHTg9hEgPloNX8W3O
MDBHZQTzz4MR8S/9mVzHgkWIUJ82qob1kXtXmdNkBENmZpeuBhAPZQcA1Oq4/TMT5Mt1LrudvU49
iSB6R6+VoPQ8bA1eIMtCK1df1oteZv8Pe6Mg8yBTryRhcgweTvNp+nDs7EazUo1Eq8EwiqB750XN
NTSi3Qr1eCroVIcCFP5FD3joio7hU1v69o0AXfTP+OvztEnHxvR1LVr0/Bvvo0HLuD8M7Mwiv31Q
U9Uz1sf4ieDPWirJzr/iDfx7hGRoPoNoPXUk3n1tzgjVf/3DCDwg5wSaeazqwVL7xMj9T+fLO/c2
3+YWKKBGv4YR6ScP4ugub9Nt6amcBiVf0ApvV3KgXL31Hzw6Z1LrXIS1kZyZG4+xqneVASWjwD6U
jZwf541msAbxMUVja2EUqDmX2otdwEwGvj4P/6nCXh/tDHsd4OZBSQtpy5Uj8+uhauC9hWVaMPL6
1TAOfNJIFotN0ixt/cGtn3WB5lSBa641MVww2RAcoziLxLW7mGuEKy52llvM8HM5YhNSmpNTymq0
GXGQrLaBS1qg6oUDsIPT3qEvfH8XsqdvBfh/ZPSxNNcduPQ49gBeDNXYMjNEtoT0y9VkVacO4eil
14Q0JeVKkyZ4ukeJTS/JyNEanlNGiLt2GU9qV/aNyFqMQ1aULrMIXZHQ17q3IFkRqX6ZVON6nj4n
BoHsGYIk6OlMOmy5GChHipi9x2Fiv4Fm7JcsGvHBlAnmFjvLI8YenEqRXcIxaomRDqlyAwTTiTYA
4Pm/H9xivY8DA48lyAiXeBKeie+bzwfLLHmBNKiH711s4LXHF8ZmGEypcMYe1ZzwUd6HPrxgtr71
JLc0zVVlr0/PVr/5nJ0NrBlhAjkyghAPx79gi7SsRJoNGlojyZK92FunuFPz0ogRmfIqK4/mDzXk
E6mQyYba9UtIOEd2P+9Y9LXcRX1j0Fxqm26oKOzqoiGwDh9okKVDOWD/g7qO+G+d1sgI+8aBPRNE
hAqsduacWr182w+cwb0XdpIFq/RDxlQ0/pBuQlU3fllSeKNZfU93qRRm3EeNYwDvxHVHi+jKWtyj
eab2GmiDrA++6WygNon2duC6PZNE4pG7cNb5LWnxvLvackcAZNn/Di49+pYQn3X0OGZgbc9BSJ/q
zOCsiAc8/byaqum6miwnaCxxq1WmMtXCqe+PJ6IVlDRpVnYPh32yEGQJOvtoj+3W/d8+dWipPTMo
A94MuKHbvusgv1d/lthYlYNy6HnkN/3wDr2o0lsudaLmfe8FcuP9alitzsShl3wW3Jv5xxuwdc90
Jt2fAHDh610kVH1s9JHPyHrxviGZSVrIfSUf8MtZI1cCe+iFzn1wfRlnrkfQjKkF7FIJ8ow6Vu3k
HTFi7qrOieQrZlAwdNL/OzMCT2d01Vyzd9T5iXN0bCXQidFoNoHC0t+7YAlWRIPnugX2UnYaV3Xv
+y+wP96FCf6xb81m/vKhO1reAlcf9TjkGqGVd4NGemZ/1BonnaKBFmugu9l6b0UpQmRMTHreVkqR
xajd8cv2mKFK7NR5uzqxXrUdXrFmNGf/nhGDSjVIUAdN/2+E9QC6ksM8B9s0fWVcArSC38utswHR
Q+dqTt4OIkvzusuKtHVAdSMkPC3T15MsDKUEeMRi5CtFUoPW7K0RDkcasHiH8m5T6uGHZvDKNLDk
tcls5z3BkUEbwgV8DcIHTgL+b1BG+N/fDib4CEclrkxcjZ9uKQrJPpHKatpfFA3KLgiGRCCErtWc
nnmTomy/NCzhlCkOb7dVFbS7Yu9PCgmuXYatKsQJ9e3Nblv08kQ9FMU0McNL9gp3XzBNcea5m22o
Ds10CYxlD5DTQ5JpPLSfcOjJiYLUWKC8X0hD2h7SFni4n3jdzIay3FcIqjhchRueYso64orMmlGM
UKxi6k8LOI27h0fKXykr0IEsqoI9C1stxzR3Tbn/kopmnR3CAhDrTW2j0iKLX/ar9jAg0VcXd69q
TAVDWhfPnrkBP/g4XhY167PuiYcsf/63umcMz39SX0HtLXCCveTUwBetnpmVQ1Avr1uABU4XtM7s
jbZtjcQaDwLoienOvq5OA1gG9ZFJKH6A5/xEO+wcebknHSn9ckyK+5PTae0bZGLfeQEHgK8XHY7O
OOljHwBvr2TGpYOA9JSfUgA3VirnmEHbHR+DyKieR5b89tKp56tO01FOaNGfwnWJaDU77jxTJfik
aL5ns9TCPQInKXDQZ/TV24GSYBRlnPTcwc5qE8JUTXnzw0bvX5mynvKJop3IFmkaitTXrmkMdqjI
i78Npyy6TQQHgxhJME1gGfmdzSNQqNz9F62oIeM19xOozVIBO27grtTa7acw+LbvkubMwrz5z46r
SqRMVoJRmr4HjokFUwVIXUAUWoaJxcAUR8aNWbyP/KEJuA5JlpwksEPNZZYLDxpmsI8dXsbIpYZa
JzUQlOa0cvOsOFzJYPyOMVjEcVC5wtJ02D1HT80NTxqjCjtljAEdAc8i+hQy1nK5DShVDlanJSU1
GD+QGlxi26SMuCyRkjRak5Cfug7XOInEpIRrdxFZ8BgiVgx4UDNtvIhi+iV1XgxDCDXAvnz+XZ08
6wy397/w2VCT4xHPpY4Y7jlnIrvLqtAc+VwBAGKgFYoWL2RLVJCcO1doDGR6hKl1tkyDW4vu+5Ha
yslaP4Sy/b03JlwXgGjwQXspVBfnODnwLT0vfYd8E8ROehQGh7IyR+KRs1cMz3O7bZnNJ69ocjFZ
dwXs144KX6CLj/1AJEwG7xW9MmME0PUgdSSAroEs3laSCzz4uMoC1aDLhTsIWYP6YP2+hj31vac/
ZqzN/Xyi7hRXGSoUuNQBBMkh1jptu+ChqOT0Gv5eX9CishuuzREtBP1Q4UQLnnFXKWo3on2f4asw
WH8sY7HMgxA2eiXC9beVfLZjhgjvPSKB/pRYHwN317kHVGhzHqAOF9cjVvaSiTb6zoCHOVK2rUo3
4Z/o/RvpK+2U2ylGP//cu/19aToL/eRfjGUUlg8lUoTaMX/x/IqvhqgT4lAMrDsJOkwT8VrBU1iz
UJJW0QyBIehexWPCSV6+OCOnJ5q/detJ+wAkCxiuvwFv7qGetJr8ZzwnfIRB4/iqklnAes+JmHwA
dvEztMYwaVdMhrtj2azjaJAB2v/GsVfS1ApBN2rFsiGWrVdCae9w53z29yaTLhogacAeJ9WKT4iT
67PmLWwxxHkhGY4jEJOrkHAM2osO/vyQXNzZ6p8zfCflfzWPOO2jiuGEPAFLFMnVqwKJI3zZKnR1
jIUDkNnAxDA5FljutiXcZCUW94Mod7ETatZM5G6/ZMZph/lxt5rtgCkSGgadx3Dt2Ix1NN2gzAuF
aMisuSX88wfk1Dt3QUleueWYqG5JDaGJsjco/ntGbRoXmKpCyI8mRrBG5jMU7UUQXQI8PhL+/t3w
xNQz2du6JftM2YTwOkZbxdWmW9t9Zq2Jxi7R3ZyhC0Btzo30crcoce3Q8ix1eNcM69RBcYpq6q6h
hSHgRPheOrDFP5SCOWSfaNh1TCzjMKZIDLkO3hsa9TSrbTAYrinehzAVgzggAP+vElSEWfL2ajO6
GPyMVD9VGpmzywqg0IhwngWxO51nV5I0zp9R0ZCKyEi+jN9mzuE73E+Der3iVp50dzCbQAXJD7xK
SlrXWyKEoadg5qd0nghQUwELLnwQIM3BfWFy5SoHEiiqVEeCdA3nPrYxoEApjjTiYD9qijDqIDO/
MLZzoHxnOnDZ1xjWCKe2oYMX5w1CzI/gks6nSvpEDHrcWaJvZcisuQkKO6mtWe7CY/AG+rYt+ZqU
5yb6OsvXcwoG873RYxNmzzpXlhFzD3dT9cU+hPg1S2hMlmn4U4Y/tDetCWTx9TFvN+IpPonDhsFS
FrW/mdEkHeveQLxWx3LCXcA7KWbcyohWraGhoaK5zbvIav1WevOORZ2shDiI8l7iFM2+N2m2DT6J
eLiCwC4BumymQKBuoezPZBwydsL75+N+Yzewyi+M7oouR4hVZlLwuS62VH9HgUzHcMFo7shtSv6C
JM5ngNmo5ajp4RARhyHukeM3ZV9aNiNs+kToqofiid1syDys+YMnjD2Ibmy/scTB2xq1GuYud/b6
qj3I9pw4OuAhlQ9Tmd/2uanPYWk2mcMKPA86TspajyayBCRHV2PSJDJpjApArfyZru/UxTMspyvx
Y/MuRx0KMJse+UcTsfprhV/H8yT/mXQa5uu0Z2Dysb28azZL//e5kcM4tvXjjl2lFLFQHZFOXcuz
mwYwdp4VOSG9qlYM6m0BPAPBE/t0P1UbQA1dgJ2ByoH2flfE1379rWr5VC5OEB9sMuGzScSni4Kf
wCFSnYBP0T8iDaJVe2afQ/WoAlt2qOgInGmnkLxH0P/n986ib+ap3WKSnprpcoGEVUumTMaJ5YMA
PR1ky8e6dhhjKms49otzTO78nuScZTeGyQ0zp6ke+szTI8WL5nY3Uu0vQ6lxEMSBvvMguf9GSoqD
J6mUPR2fepYYDOV113xLpHx3lrgM0SxcvMnb0oRcGCeE2RVwLcPdnixGNMT13Jn6ZJmfuCwgBWkN
nGp9Ofm0aIA2JUO+YiV6eIJvDNaQ0zDmMYRyZICt27sRAWZaJnTmR4LRnrA5L8D25mha8h9/IUDG
icdCGl8oExx+S5NEBpC1t7eoBEPCNW4Fr+bbkesRn47FUi9xaw6LH6oUYKs2bg2Cd5464MEhEeUO
aoOGbWhX2H+i/YzED+eRjsP51XnJ4T/70DT0BS8t30SGZYCS46Mofk+hzSKSySGDKv6PwNa/3tau
Vx32ClHR0v+r9dARmOqomQCfxQTK6jd5dfUTTXnlyGD1JBLRvl3NyF7Hh3CAsHlS64smsMzKFbU5
8pG/KAmN1ujERo8hv+GZziK/5wzehtuqbm2WK0li/5Rpi+b7RYOMy2lcXzRIPl4zZpmK5RfX3emM
mQR+Pq0u5tMn9nTwHJp/CwyWKOisAwWYr9sz3f9GY6a6BB1IzlXj/VecZIqM41tLAH5pqTzvrg9Q
c4xW3T4VH9AKdNWMN5YTU7LCMdglT3VqR7HYudoNs8awjAGAWkvRqB/Top9IxjFjRv1FK1GddsEj
h63ASkXMuPvm0TYyYwyyIo1vjBaD5l/u2UajjiQwtf46iOsahVQo48ZIIpviKf9xFKcnxSt2mzUX
gaXubb+QmHvwafcCYVO6PObyRzV1ywq3aY3wNAQXS7YRqMM2JUHoi4guJ7ZAVXESWyHejGmjO2D9
mrh27ccCMFJ/bIPh6982DynCzmbyclFOo6vx4/KyRad3vGx2qfKeKydcY+PmXW5inDjH21zhziSF
8fEIH/iddEkGZqyAjQ5fr4y/R6jOwQLCO36eDk3TZlkq2a+GXkWduVvhtWMLLzhmtkjM5qVs7eq8
eNtXtDofh+voDkiiqhj/eLPSUO+vJRFuGPcK35YGXSaIexAsICoZEL4bQriWoiEivBKJUsfmbeUr
0QDzrEW3AnetrPp/QqvPOrjtLmbitjWQf0cOnxvIatHzuTIKU+kuKofralP2S4/GS2qCgvslZGhX
UnG4U6U7U6ocdk7kjwVigJhQCp56XA3NF+0QgPMqvADasDIdAYAgRoOjhtgtRqZeT2jwGX5vXFXi
Z2Le+FFV9IXPxe2oTfzdNRLBYDHihXxPjNro16aIcBvqQ7rqzeLb+0rLnOvMpaqS3kjb+F59lj+d
dxVM2Kn0Md/7GmeJrHzfGO5jEjjDy+a/yLdyuniLwkmoS0XLvhWoF51XOIYk/XnukhcuDSlPpXNy
W5bJn2GK9fNcGfz4hBzs2OVDCOm09HI41t7VtuK6qJGGr8VpZZ3URKT5Y4FOT1841WwlLcjwW/Nl
mq9F6L+jWNxn0THgCb0XLK0cr3oJUJu9iihWlsnHmMPRRfllUvWKBWuy/WPQx4o9Ihln7bkvf+ba
X8VU302O9J5Rt/PFQQEDXDxiVvfEYaBVqZn+xGepxC+UlNFdTVfD6a8EFZ3ArPqLoUVz4HLahjMb
0bAuJGgXnTUej5U269ctDOe53xLyVS6kII4I4hLTB/KCMMy51NkxJOaRJ6rNOgIbC7wtYcNltBD8
nFSluXwA0p0JXPTm00CfoRSGsFVPGyWbBnmb+eBM93cNHOPft31BTCohUquYLlZ/uRIB3ef/L1dq
9e1hf2h+S3QcVQfPMip+/oT12C608zmavQ1bga6BBEJtqKhJqQDpmkou4v0FTX3ZXlW6ozGyZrn1
eOkTDJqk7KtSwm+hgiM8+KXEMmJHRZ2eG7Cu3R22HEmpma976pa8oa4UNnveuzEOAHPmVDHWLWOX
5aGh3qie3OXHjSBiZWFaCYqjO04dXW54jKRi09G3GQHcWfpTKrfWfW/z/s8ZQ1ihTF1RHXIOoyeJ
G1S5aUUbJfztsNPsJ+wv3v8rlNdpdG9ipiturNEG3wjdAPt/YJIO1sKHmNIdrq547nwGmLYgFAg1
Ledvwq45KG3SQ/Tz06JtjyELlHNtQrWKVrEmUDCILxVht5wnI4pwiI5XVsXVaFD9DQ5qv2f0imic
b5l8C4v8zIi+Ns74Xen70BLpUOONwodHSmVbuB2+dxYCC84Y0gEYmzaebsoZVI+D94a9SmoO/ngr
iPgCqhUcQI6xUmcmNem3agb9odg5TVOeE52yiMxxkcC75HKQAJfEO9fc/X4uVouaj3nx4KwaC7VC
2LqkxX+BRMG/eTaNqdVkcdjtxWIxO5cjCKGkrzpR3GozeM6d01BG8Neb/OYtD9SNxuHW2Wyqagi3
fN1AUWKmg+SXgM4sIbaBxIdywILwrKbGewdT/FKIk3AlV+YgzpTgyWOpzbvOOoNogSohdwPTIBLz
LRARrp926iBrE09+ejtg60vnCj1XiTKKbhZ3SFRIX6BG2knByj2teBWjT+6EBJ62yaUR7RW01eEe
z4MA6fe6Lwc9z0P4fdG5syqz8HpGqVxGJYFNQac9kDs4MZFakGf1VHYKBhYqlUlC6G44c5DfAoMq
bEv6xAZAxR/XtuOm8etkagIY2z7xpGAUYdWRrFBbB1G40Yd0/b9vmBBg4yyuQEfPnT97ko70AKFA
SeLz8x8XARfkyvuY9JE+/exuG/eZbCRHSP4GrIU7BmUmAGexP00YnwlYf3SIigFKIkLwUNYCqFFb
JHR7pc5x04XsYJwp1bB4r6FFuljPaWBFGSzaWMwDmOwhd6lbCtfdXfptF+fZ+49M5JvJHZ4hg7I2
QApqVcM6BlPIlCUydvgx9CTYo64YjLLH7qciawBrCnw8LiaKAJeqR2i2fnOPIpEjaew0lme8vvHw
20ma6KhE2KZg/fzIIhhGKBK6mof81wO/ANznGuMuwb87m2Om0oc9ut8K7rMTa5TtK0TtdHwWF9SJ
5B+Fx21SMVkJbnmiyp4ac8rqlDds6IFFk96tsHpk4fu96S8iEGR1tjnhHUml1g8/wq0yqEjt3AkO
+f6aAApjtdCTBOzj1nNqQbwKAQH0U96yWN2e02x63zimmP2ytHyeeQykQRoRYrfq1+m7YiMcKoz4
Df8hnKjO/1VUUK1TJ+7UlfVZpuxwNXpOKn5//heErFKOjXbJ3ke6XowWmVAHJ+xAC6PZKReCKG0K
0vcZZF2teZGH0IHutfCsdLy2vhRN5+5vR+GoSzS6oYAAFu2duHJCJI0DYGokECIHui9M9M2Pothp
wRz+uZUd/rLvIR0r6AeufcpYlSibNa5Izc3aQsnKytypHj0jVYElPi47WHmcAjE95tXfbXYubE37
ViFCl8vWQSIOCxNlI+y6+JG4Ow7BqVaPIiN0Bvw2+DsvOOW35JvSueMxY1hybfdYxtKPFjGUGNFM
23TzrPP4fW3Ay5r+oBFU41ujRWSPegQNkE3GyOb7ojT7+t19PGRDQtFRAWux21xSssEFu6RR5j6i
oYiQ9nSc1Wp9NCNwwoa78ul+VYc3eo56/Wun7rUdByRqDR2JMkkR3nTkGqX2G7nNkEJtP0WTYIvh
aHSlBeA5SJJ87zBXGXyp7H4jPZB6W1M9JYZ1SJqhjaotMGW2mKN1hvdH0ryi7MkYs4OT/RbueQCA
424DYXOKvQ6ub4GudVlB9bOp9xrElduVKSC2IjMqItW/4xtxuMr55dAkW91QqK656FduOOGwB+TB
+63dzyIu1Qv99nf7eSa0IKVf0X8mt3kdFqkx2d4daP3mtaTtb1nZjzXie0BdRaWovA+HKhsWcldE
c+MNk+H6G0X+tm1v4DjTXtzWL9UeFFgv6jMl6B6ONLqq+awc+W2zfDo4gnwldtcd7WxOKlaXmCB9
sTpczl7PpoeoaSfXPwf8W8iS2IGPjUeg+WG47cdVJ+frQd6H2+v4l7G67BMUPZt4wCVlFuDwoQx5
abPQZ2iwQ+gIfYbia8ArCGsUdKgtfKatrwpkouUw45Ojt5wu35ddqpoon2iGZew0TdudKO2cjWli
0pv2Pv02NPOicbOYkodibCf7ogSJVOAasUmlXiyTNKgEEiRkjSJetifdn8BGZHMbzP4Lstt2aWnA
vcd+QruNJdjqWLHcV1wi2tXVz/gZXnmPRB1qAyJUGu84nFJOG/yx8R2ylfQ6YiUjXV+pJKEdeItC
NCAxPjJzNW8vqQ8E441ffGptQ4k9dJ/eaCH//tEaL3+x2XEEtYXS5HHz5LidckrtKrL+Wy9toz/n
8p/BAnVzr0/2M9MTH82TcW+CMNa6y4o7R5C0w+snTGVSWKsvim1yfKDlhlUNNmbS9LfLFTkhVoYh
hR6MhqHvo/YLKknStdPUrUYo37xaiySm0TDJwVD1KSHa5NKx8ZA7bDXKs+qQK63liuWiJgfDC6Hv
bBJrJIcJbsbG3XgHoWZ5UTkqnARSpWO9Tj15fsvpWoYI4t0LegHQCjRdj8JhDjjne3zZqwjPjVPM
PKAz+pTQqeX61E4kDWxOMX+TkETATHuCe6I+9WkfX+PtrzcnTGrbxvPFN74RPtCwBOOPbmyQ5rPG
BurkjfL1AptnsFGIdw4RfjR4ttYXDI5hn6erYSWO8KkgyCo0ut5AaI42FLi+dv1561KWOw71LZGW
j/h4EtmzMuFj9YQWs1rKv2qfGfkfodZG0QmEov9SSLJMxbt2rTRdd5R2Kr4rrgrC+zVhvQ/9MMnM
6Hmv0C1N8OWAdZ4oXTiGxMHdd/M40UX1JvXq3dHlWA43DfjKxgJB9SpSBA+Xe/Ba6CEoK5/rYlV3
gJ0y3GZUy7ceBy86j/2RjTAW1YETqudvtSrGSTf9f9PcCj8MCLg4nBvPTIHY/lHKUMEhIU1DJz8m
MMErnUIxYpIuzuFP/aQEl1TU9dF/h+pyiXDcKq/ncBbuUTUjKdsmuuwh0NLNQRAwJC7MnxtnoRVv
T/vESkGG5CaDeWvKJk58QIDXrIXPox3JL9fLXrKNMTP6EvYn1m+AYp0QJEc7PwurY0zqMQnD+HAp
T/OJsT8FozFlpW9uZZUNrj99pLL7uFOavVHjrNj79R5Hy1GXdCAnrttIDf38s45TNdgJ+A0u8rCt
11k7MTEc/g6LlW/sSxcFjxq/imhao/8tMSrJCjC4EKX06vdb+5lHQVrE+O77Cq8nPUvBvec3nVO4
XPGG8gnSsyiayUt4vxyELUoK8lOlp1tY+kcQKxyucJIAW2eBAgY85ye5cH2inAFjNXz1/vFEVbJQ
5nj7dY4q4xhJjpvOTtA49SCzEruCZPJaxdzmz8RuG/dw2s1tgQVkErPf1DXsQ0vyM5B5sZLQ27pN
vR8JF/izAcFtSXjML4N6+QajFxAPYnbQlHvUkY3wx/DpQcYRiz9CojIKeZ/00hXvbBzqBeZ9NkXx
qMvRenk9KxVIhzaw7gd0ZjmcFhLzsQRULwZh9jBvEYjgEzWIakM06xOEfQOQxAL6VN17vWmcDAb8
w4WxYT6zGFAS/RgZtfp7hqujGDkGAlrOspqaUop6GgyXGwVneTDA57aSlPHYfHboqq9M8VpNal/y
HAdp11JuibKF4m+OaTIrc71WQOn8R0OSaIt1bDswwuuJKRdsti0IvyXulPqSXeqqiAkDQ09TK39B
Xij05bFjuH1g2Pqji+l5rojPfxBi/0W9jw1SU4JZKH/ivhku73uPPMQ2z4j1uWHB5RYXUIwPPY28
kTO+MQkWcZy4q4wRrmPV55whvBO8CZLsL1nOxdTGaCF+Q1uy+jdo7T8if2Y50SmWszDxkCfP9ZEi
bJ2LjSXuyuUmQ51zhSyolN+yHLJ75eX2zPOGBAi+LSPJDGKjrturTEO2ZDPcbGBtssKjYAWLBsug
EccaopTHKEZKKpwjUzCG9KyBXkiY5p4hgSH7sXcRRx84ME7wK7xfFr8bdFufvT/UEP5U1eQB0Kdx
tzLXxsdEeYP4gKHOCIByxfvg/1DPhclvBFFupID0qrWkmDushr9qk6bBU1MJf3iNO1sunMYLLGk5
B1kBsqB0rFBrVH+2ngEZV48K8uwy6QJbuKV4aigW+tB1xLIH/jjvN3n8Je1XhOeR2wgBPTsy8BtF
vabVsmXrpOCU5UZ7eRimqZY6ivkiA0+u6d1Gk2lQTwbKepFLBe5eYRSSY1L9yzRKZLvFeSJoLgqI
tQdNj20WpHRvT0/gHU8csKtnB9kvqxEPZDhyMb3zQqFuhB5gHz0P+eBVBUYf9UgjnYCnzu3s8uNp
dnkRdkkHpT2Cv1n4B8O9U8S7IcV3omRr88lJy0jlvjpwkN75vwyadENmcuxISAy2CG87a0KUu7uZ
4o4vj9+qom7VpCNyFTobApiiFxkm6SQs4fW1/+KMXUYo32VQP1J1i0xz1b68ZQBwYcyGcQRcX0f0
FSczEpv9cKFgr++QQF/FXPfNkJHHChO8ZfCL/oM5fDFFHDJ/4NU5dDKM4/U2rVMMvgfDaaKBzstV
OOl4pstfGkVYhnr13ZXjHK2kD3n2j412vnXPAh+fYx708Rz9NZpSUBKDfOMEKiMVCrzlcH3WzH3n
e/miPAUp6MoDjKeFZFTIZAkpaMVtyymQL6qMdFiiMmc81rkWGO+Ra9CPlR6V4HpSvr4o0x1KcVu2
ORQoaYHCkZ4fN7JVKoQZrAvsTpiy9MqAeEgklAEWqGdPg/QPTVpPKwb5qw3KamLaQ3xbegL1U2BG
tqAs9XcviojVJeaKa5DHuPCtf4JZV2ugvwUhyrN0lOFqfgfpETHUwgiqKBzG5rueoqN/KCQw55V1
Z6xWA38wL4E4sjCcQK6Hzfb5GvWpB2g+1brUGc9UvqfVug+tMz6kFx+ABxmtxPVvPTz8GZalEdJo
FcFchdJKXf6Ub4NEE4KVf3OeCHQjAPShEr3/6IaHXSGlPg6SLtxyk2+WxmtEea5uQPhrOIT4o7rS
5ngfw71a8uHX3fo75Fm4FEykzel2tyDzkFrl3//CiJHVjitAtBRGML9vUpsnTlF5u2LxC7icPONk
36jnuVTm6Smqshx/unFBQcvBHM5g+laRo9mneE1EKJt6tmFvhhzU11vMSRzgW34Jia2QdsAkpNDE
a/+4KNH8FiB9+wF45/DDzPPbEHjCsybrRhu1nylQfX5jOdLXo5eqORB05qED6LawdyKKOZF9oOlL
BElwG5od4iKqrOmvwEl4oKm4ebMy8p+tcbhSKqrwSZDQMPOyDiP5gny7YEzYT/illB6PgwKPmlpj
QyZ+AyvCQ5YXNYURMGfNgBQamX494PCLEVzpTx2ukZka1vxBvSw2qG3CTbeD4L6xh4a5rG1TdoE9
Wbz2T4BNhUZTvwbn5WAv9HyE5NQQBUnON0eqEFKf5gSXQ7akNdTrlLZPkwD1zOC/yKUHHPihlh7E
5OfgAyaxVdeFyh+4Hcm8BKwdxsqGFoYqVqs8EnNzkvzyAPu25vmNjhbxz/L0g+l41Ydyc1OKOnvj
j/ZRYlH67wEeSYZjQojDDeXi9jrgi3IZpIdaGYsjwftl77kwW8mI4bn59mUs8NZycuzMTDlIBarg
t5xdQxKz6Fa4qPYfgaHAjFfskKk3rgcpprzD43ypGSr4m3kEZ1u+ZTFSv4G/ZT7Bpyr2nah6dmKE
N4Ei/3tsHzK/9Vppg9zHCoA92dW2KQrpy2ee/QgFdvjEDSQPZ8fA4A4Zu/yKjPHkz6hp8WkyDG/+
9+tvpIa3q11diasVDuPezVto0gXfWfmqTWQL9EHdz5S4zOXiF0hpDVmAxGbV0eCfNzYgG3olHvOS
aFDXbNhEx93tWicBD9JpMQJMzrf/HGDmz50k7IQu8J8/ZUHJ6X/s5qQ7dxvy8WcJzMcFGCKawm88
ZEPSqwLClBXtmi+fYJ4iJu3mRVaod/dwyTXLm9jSxcLCe5Cap5QkQETgKIYhPQq5OvN5nlvM36wl
bgLJdVfzfzkV8/OnJwKqD3qNM9zyCJ0s7Q21UFcuHBrQjLS/V7YCzQw20uFSBQB7tV6x64zWdlb2
Bl3lxpB8pCDrz+IMJvMkEstetACj4ScU3hTV94yHE89RvtPrGDdmUPzx7Au2iI0vXdmf4kVGubSL
gRkDg+KvsjO2+suKfXMhS1Y5DmBhOcfPkZVC9WMVH1UH8hEjC92DIeIIBhXm4WKA42gz9BIdiqFe
lJiUSkUCYew6rXOAv7XQK3GUbe47Ubi56YVNCHbqvcwV3OsatoBUEXDDpLjU+KuZSJI8e+r1vQr7
I4UqPk4AVP7akaMsuwhkR8vE1fTbEd6/HeDqxJOjkdV4TFKOPY2bej1nBx2zx11zS/DXYl0yV3Ih
/h12um84R6GO0is6htMm9Ow1sYJ8TbKcMVdnpFsknhfRH5CJD09BHqPpxqxOvl/jfu/CstKW9rAy
4eyty/NNzkqnZQaz5FPDgSQKN4nkEtAldJfKemjEXGDXB91zXlmD1U32fkumg9vWhEIZv/lVV4nD
5mN1ZPBgqFKWnhZkihbOfIu8e35zs3A5HiGxtnw8uikm5v3kvij6zLSlzPsRKB4V6t67BoCu+WtZ
sN55NCPooN9aZSOEKcdKwkLlkZUR0AwffDw07xwDDp+D3tkRuDEzL5fN7DVGH/gtBkoQDYaHrd2q
wnPO90Kyet8jrp56t2IdiPTMefx36TH6vxe1EKsY3b4dXfi5BMxVt1lj3NHymuGxwBikuXtYzgGJ
6t7Shjm+THhRQjqZo7BgOWorNhY7fPjYlIOpV1BM+dj6weZjGgySTPVQOHTZ3qPF1PtxHZ4aPExg
IsemjuVceTQDUaMSHZqIeSu/v52VresBMuWg/TCchCvgCLikrTN1Zd6rLh5d6Ujp2rARGvDbUDA+
IFcDfaRG3tgGgI6cpQfSQKMDXIF6PgCm4EAIZEGzKFe9QpFzABUNglDDDkAX0GFvcTvJ+9UooY/c
HKWvzgJkWxYGoqdw6epnsneQaPpbeBEYyhVwU+J4glJPeehN1t6EHjny0AbWHtfyJXoGnuRkKRtJ
HLr1cRo6oENFhZszeq3oL7iDAGY+9evdqOKvRaBK6pM4p9aM0AUYPAZrnAp6UccoOce4MtIndc0u
RTW8E2wpto8gp1kUroh2PakVdYU/XtkuqvvToz2JR5Cg7TDCY/vrnGODrySzSO0/V84cYrPAaPwr
foHeptJJILPOQlD78/bJUL3MSH9l8OA+W6I2+VjynuPJkwhrWWm9r+DOAlIeP4Y7/vPPO/NMFbew
CZwWV84RzbTIjjE8q997teNnXqAjEVKhs52DKD4xoWQuaI8ViDS5ih/iAembmIraIu0q/Yl4Xw16
nMQyhh+y3HC8BTZ2iYgAZrSvQTTeXyUF5+goByCUsIUBF8+0/GdDdQvhM7vyGN3E13ISGoF0u0Zs
5VLaMSmhirDx1JuS/XyEBBYd255og0sV4wOXGea7/VuSqAIzYr9/ypH4FX3Tp6OxtV50eTfpDuux
dCrzWchN0dc9Ab0Fj+SX5sLiFySmhQxjJlgho2cP5oFl/D0sE48RxQR4Fz7UBnFytKcx+HxXDFPm
IxZhNuC6Avo72CwhbyWq1vrXgILOf1hCUNfO/yxbjHxncGOlRn55TwM8o53vG3CSmzTIAyuMquKE
eZ/1YaM+OS82weysq8B+G3Ahg5EG5bjdzRQkjVFiA977OqxxxrHn5J8sFPlJbY5g/P17+8u36Ewm
4yytq8eXuevB5l+PC7EUN70u7Zc3gDlLT1Ff5sLxtjOuzhZ762AIr83PdHUzGN0932L0vI7l/Zqg
aqOJh4WQeFT9lQpuLzgoZwc43qijC7B9LLt349MblhuvvGHFAIbq8ADHNUgO2vA3sRq1g6/o6sJs
hLeKnlvoDZgKRYKF4pNInwCjgDfVsNsJuFTM0YLq2lTMsLmAUkl0gHedvpblhJ0fKn9bi3Wrlk3f
0MJpxNQ1b9ttwyeMzNfPz8S0enSBrr9lfVHHVPaP9P7Zbm3EKZ2f1BGqXRwdtvW22KpLdtSvRF5x
whRPzhgZrjbATkH7yczVEuBVk1W3JrskBYDOd8Me1OHI6sUgRSGX6/mGXc3ZKRRkWNVvHBquOEXH
Tny3BLhwbdFoW7EgATZ5AKvex/Y7yIL+V+ohXizprTb4XWDfN5ajeMcYyhKwaOo0dd+vDinTXt7D
pDKGWm4LgBoxFIITkuMVDQxZT9l+gH5HeFFxzlAkSYZ9gvLg56c6Zqq86z8NZ4wwZuRRmXCGuRX8
0P1A0yPR6cWVqEuwIThmBYDyJG9OvC3zFwys86P+3l9LJePHIR5UzuLZF/HmslRgHx8yiA1NFluy
0IA8a4R+sw7lHFpsfv9YG4qN+HQ+BxLjqUv6FCebU+3zWOWigVZPgKcCCP7ilEJ6ZxC7EivFAtBw
HluG2msYBER6pBP7ioJmThE6kNkR9nJUVRboyqLIPUTQGeOwEdMIQZS8+ZAlel99ne9DMf1WNAAq
Jq4fOwI4pRFSLNlDgXMlyO1zgsCanZ7CxhMb+XYwtZrbZGoqtCde8wKc7e5kxyJKwYSxuBUphsuK
2a5vHZDuBGFGjrX7uJTqM6tZl9HU4LidXl+lCvaCu8fKWcmvbjb8OCA06V20IddAk0QBgCDFHJcP
04CPcNQJqEnjz4JilOdGq3VCZ2swanKohkktIZJTjRY3xSlzfNxZqmb8SxiUa2cSkmUbGbUBT/QW
JTB+69aJk39iNxO1ipUZiD0i/J9LvFEKYIDaY0/b397C6aVP8XohDKKcbSBuDWfvmqPjgP7hgT/S
SrqEQyDy/0JB4CMfW9+9uf407I3cbO8HEAnNurYFlxgt2b5fplOSxnW/7hYqqeIv94K6X18n+o96
hLlJUT1r/6n8l/S2IJrmn9tAi4uka9Nxv1lopuNtxE1TB+aEVfZtY4ebZWKIVLbbGkSpjBj1XqY0
6z/+LSn9KSMPkJBxfpbLkmZQ4aF5/fS1ymdXdCaBw/IiWdRMnTvVFoje67XeFkG+j/fZF+C3DMMS
tqpITZ/zlv1MT+VBcD4UxYlxP0vGInOYbI829Oh+KtMjrxiqUtl01ac1X7X93HPXmucBKHXHkMli
xOqBIHqEwYavRyJiHVTOWYeB7tY8kXwN7/m/mR1oMPX0LbZvEWw/UoYkmZDHa+iOs0wlSkH5TSlG
dPAyErQC9CeUSEr+JoRw1v4TTokNCJWZ781Wt71Vs4M4oHsK6CPEgCkPC+hdt2M8eplkOd+0cj00
CI8DLb7R7Nfwd1l4cnBgbF8PwmHWFq9XYo/Co0vrbFTP9NvLE0rn2/5BggNnahVSI4azqTzNN9I+
+aR8EMXGw0fZsh7Shc06T8Wf+VFqIQdc07utGI6H0ZYi2mDVCx3gBMx6hFUExXF4VY4pWWIfxmim
j+7jsoUer4zuaRhkqZG5lfJEMTEq7iA8IkteFXHF1RnC7tc9i4+KK7sKY+F7/DjMf8SjoLrEJ2Ea
QS1WzA/rSfJJYXrp9kpb/7WWYAuROrmz4PaLNCuOxL4yMjvVOzLPOGEDBw3ZNMR518eZAM0wQ1oN
cnAYlttnJf5czlGuXmlNpmwDFu0kkb9V5mR9HVyrfgeYn0/8Ns7kAUXn3b97wJMzW0YXXnIt8XQE
4bOlv1RAR7Mk/jWWmTtY/lscAn75znhVpLi3qULxdpQgd+VrvWD17xsuQrQRv0DnHQhnVSRfSIig
qQTRxhrDXXq4M3ORkjsUztdzR/xOhin/c4q3l5sdYqFJYbT/pMSqz4QsVZ8b9G6eK4VlSiRUKKk2
KeCCQGe/grQeU1HzvgIjin5DWp4Ay1mdgTi8GoWAkIJ9HSVLlbWfbNdI54RxBdOlnY7nm93AklMj
6B/lULjdhRO3MiwnakgXtlX+tdsZ9fFikZNz2XW2HDXa82jeBvfl6BccpQwoxTUk92svbnldiPW0
jbev+5hu47o1dvHVGn4N5hXEp9i+4t9SHdhPQEdSHhOsT13b/e90KHWUdp4JF3SlnARIjo6kFl4F
0ZpRKmAlGiRGWEcsWZc7JpE5rwH9BRXtPXZRcXQ4arsSTCjlS7NCCH89e76MsC3ZlHMsSkl1A2xb
vhvcllXhEge7TViFnwGlTuMEM5u8yyWeCS+CGAUWzPSMg/Pz5n43zm6xZxTlSSXHWLz1wREa+Na2
ezr3wXAiVh3eF5fYNZ9v05xBg/dk1ETuA5bMFjdlyazlhlj9ud+JijZesE22FRd0HWndvgerqset
gpIJemT8+U/3+BF9T7I8dlAmqcMLHlBrEeJ0vehGiPUIoPgCK6MLz2zuCrM9UQNjXcTpQJ5vDHwn
AGH6EijvtNw2CtavGRhdIyiiwrem8NRR+MiGzdI/RmtyT7FIKmH5rJmQbG23VBBGumap3H1Fjo+G
f8Y2NkNsLEJYAKChhjklwtpcCdKHq7HXDTplAsLdIQpDsAcodVaq9y2xzABo0Bt15U2QM2g9jVjb
wsWdNuqSvQcdnCI/qlAmyNaezA7IWphh+HRJkkJnorx+VqTouuDrReoa18txBhA1+hyIIYhxvrKF
4PvjoDbHUwNiC3iabibDm7tz5HAmbvhWy8+kvVaMzlqQfgrWbvC6ZIJbUDdevUKWthskL4JmwT4h
Th8TfT1l1/zYxy39AbTRKBY7GazwjNgIkR5rrIztUaFec0MZ51CshuzYjwpCpziFAHDsj6IslIlg
VeN1mcVbkoZihf3EzSiKbP9k7i53iN9aRpjvdsWDNc1MYMd/1ZAHdeVI0D1a4pcEV5x/5aReNc1X
uND46EP//JLyhKnkVyU8G+LVZZ5KtujRiNtFfQz077pCYkJsA2cXDQYA6Ldt2I6zqnDtppYZa+kB
6sHeTgMrRBbWxfOvqftDx1SNo+trcPf1+d1WOe/YakFM+vl+Nne83vziurS1to0aGmSoIdxuR4VU
+BXriCc0ViIPo6jYO4VklHRbPAG8KMmOev8NBnJVb9K01TxxozHMfl5RwG1b6zn2SgkyYEPta5vE
WXRNArXTmBNcYLrKiLS74YFdF5oQQHHn/nYyW63iY7t0+BxV3CMS0cm6wozrrlaucRKtejmluXii
wJlIiCxTCUd1fhNCEkutiUVYHlbxgs5YJ3V8x2tBJw7eLD699WSLoeqOaYi36T9coVRIj9Cclrpj
5aBvmZxXSlq9nAAFLdjvT1VdKwdYp4rTPuP4aU6SVWJjT4Qdj0KRtaAtC67xA9Y/HiTQQkcgSaup
V5AN6xWU6O/vUeqYL/EPo6TNhAVCcfPER3D6Rr2PGe6HjalDsxrhMcXWtDI40yBCMhMDtTEJMOfF
BhggfE1qtrf0rTIDgHQfUX1y3SCk5iJbd6Hnf9pF/KuUdejUifJ4m8T1ExLt8IN+8IzOCA1zNX9y
SBUVNGeyuKozZpffT4/yoeoiWyJDd+2CVz85ISWXiauu2bv42wGTQ8f8g0vX9bcA6qVrgwMQ8Jxt
QPeqANjxEpyDu1jgjDT8P0JFEmiuTmvf4Fpt1UlM1f5irgfTp5AZt5CqbdVMhi4+MAfSeByRsSQ1
JHRwk+f77QvAe9rRlMmrSWr2FSxrgrZCO4TMaCwb4xE0Knml++dtGgeoU01vl/8xjnKIrFYJFnQ0
p6ik/USeTv7ikXRs6eLpsplTPwAWu0Nh2Jsx8HvvGTUAas+Czyd7hxzW9MnkknS6AsG6k3simjv2
Od6HbB88Y//IdUOM8SKOcmVB2rk7zCpEYVxgxEJmatzV1/qHVjFAN1gNKi16+UzYmBo7EvXKaAjz
FkldtHszEqqJJNULF6DFUdtX3ajsd8bmP/r5nL7PH8CqFKZ5meABC2aHoyBxhF0NgW0LgL7tTYJd
mMzxb3KZYG9lmZJl/BSALKyyVpxGztY7uOF2As3gip+zmtBQg6JGll+6UVcOV5oJRiMGuHNMIsmu
/3bIqzn2d27ocQkcoPS1nbRWOuLZbt1Z3fwaEXlojdku1MMPNrg1aWXT9xB2lJfW+gbMZUFKcqpn
13MpKQT7k860hQMFVBdve8HzlfnNwsLr/W2nIT0CQlcGhB+tDAi9hJ0MayYz9owDwxNypurBY0/i
BjlkC1UBSl5GSNvtynSKSVtga34cuuZmcheMKHQ3ujvQ0jK4IJsX5HcD/tRfSalMgGV51MnwPN9P
vm98I6iBrh/krIzsGfp0PBj7jsfNO7Vz/OThD/OINIlbpUrHgyzSq5ShMluDkaA4BHnyBq8JfYqZ
kg0+lWrywYfBYHBWO7mvDWXPe2J8iHr1WBVYVwr5ZVAjKEKfqolCxI9VrM++iDA8zTO0+6k+/61E
aqrDKfSkSVqAwTjB2XzVzI5v2eRGtqaaNIgJMGJyd9ob1x1gRIhK+D5qIK5camp4bi6INqZGkud9
NMwO/4GR0peXLtVOCy4VtautCtM3UFOYy1ZDLJR5GczI+1BT1nBHWsHlC9LXjLFcqi9ic+CxMzSe
fatjrmOEgCGwfxLITzk0hpWXWw6RDqTtDAm3n5N/EsxzkyGscYlLKmX3R5wGG0YR0a4F7Ajd2fgY
pwHuX+HmcrQvwvYlhWMUOaXs4SRKdpy0xliNidOIieg95jDfEMUu9dFx/uWX4locJVhZGgGXyP6b
Uu/hmwgJkXWIiqxMSwx0J8VK1lOywC0DbYAMZae0Z9MEJkVVcYgXQqpIxDo6czlVG7h10OjLmyQi
xgeewd7Vrqpn6gNgFhNAhA032Hj8iMRP4dR66vPQvREVkCdgZ2nnVGH9PN0v6FytIjXBqGDFzBFo
28euScM2pg2ibBB1i8HfIMtYAud9fSIOzzLrNjb/RrVWBN9dsliqbrGDnUD6IMjQLPzkBbQsjoca
IOLp/vn8sg3b9OAdwLXpr28V0Vivrx5s/rRIIuv68+eYCvpCiHzgb9ssWkfQwYxUg9vV1f1LagII
YsU+t2aCT7Y8yy+07oameYWq9k0HeEH5JYCFVpvI33vGB7K4QR7dS27JXjdKGEBy+sRhXkx6dSFj
JxpewIfHNXka6qcJvCNx/rNdnWfPuQINCf9TthGzfGrdFK0F48ean3eSPb7y6FgDb1/rp832sIEy
hSD+nzG/9e382HjqYb2vHUae2debS/RtEAVu+gx0RcAnUuumol+dQq3c+fx+2Igl81/TgIvY/cLC
nrTmA9aLiNNP5tdzu0BX0OBwDb+YEThVtZWScgmXki3+CQsC4dny37Kzmq6sV/hU9lzwVfEXqcyM
jvsUD2k0pbIExhXyT5kmoKoO5XMMblDMoqtorEtBgH0vZTjILyYyBQa9l6S4PB6qjUYYDLTHJoJa
WX08AZq7/F2p6q8Z5gJHceGOrlGZIjsBv2nlAISYJKs6YDdrcKTTybBVtWsNaOKwXyx6eYffamKO
/szzizx6DDtuHnZGRKGw0JVWamwwUowLdi7TI72tzqHKwtuW3129/Mf+UrMsZoddjxtzKvPO1KJc
riHPVTPYhvpgPz+Kb7kYXdeX73nSMr02iHBeNis0xFMUW67tI22zK8tTwYJNTEuKY7o35j3j+Zyv
+8EQFmcXP3QXMMLriRuSJlV7mVGhvdqVmnRiVkDjh/oP8SVeMmZdInFFmjY4dzoQBcj5nFOqvZlx
C99f5WOKo1TrV9D77QLvzQRVtU2ninyB6DRHSmT0fVAlk2y/5CxrigYj95HvKuwXxMXck7F0f9iR
OYDppSvnJWw6QYkBCYoHZMYfk5043l5p6fjMks36XsHQtfHvw8oti7eq/Qxjz6YnUn2kmmZ3l9bB
YzGBEZXLSSwuA+JlT6orBIpcD+Hgghjhm/PsVbb2b78Q2Uo2kFjsB+P5UPQ4V6sO1b5TxLI2078T
eOJhzykfHstiLWy1BJNKk245XGCLirf19+V52ihydhP0oYVudiCDq6zZuHoltIDGliThePxWeSwn
P6Pp/NYen+OyZGX/yL480D1AQLJkuiqa32YFciIUiUpBf6gM1TyVrG4kwvHg8Rvb/wHMIPpGy7Be
O7fEBbHo69UT5o4osVeQnZbtmgul6ZkJUQYdSfVUqRqV2Qdk1Z+nbzLP/ZJyq4L5V4+QztGcyzL7
p88O9t+1iF6V4uL+ExyoH2560ib45gozaLxY6tolbFTJmucYY05msjlQwB3MRQP8RyM+XKcIApt2
NiNUlCp2dKjWSwAolaHr4S2hnbgIh1S95jgte8w/KoZSn0TjAK0GST8VOjs6V3jxw2zGUjJmoqAb
8vVTGoMgoRgYeuvdKIb6kvIzMBiwqWzLOZ3uIQBl/hRkzOUIOsOxO2fXX3ipPGQNn9fUABgkeQ4d
UsOK3vpRAj6WoWZms1LQU18ax9MiMGMRg2QUAszZBH+dVgvlRqtnj9vH4rOSFAOIE6M9ssilD8lH
MDnPnueFunmi9h1Dr2JgtYVjMqOiGmksmy9sRVsVQmO4QdVLSCWZuKbWM0Dyi/049HKSSp5Xg8AG
DmhPL9AXDIYsvbsSXQlivs65UrCiAl0houkre0eyZYVNwybRLuGsLn9BG3Ad0jPPfKpwBvxn2agd
R7s2e6pMXu6aFnDkg94I34S1r2ZaZxSiDn0bCexUC6KrhXiUmn10K2Ga0BUQi28+WXZTvbPTk9cK
xeELTLFY61pItd88rHF9wf5pC5ePxI0YBz+48DlPthcgUmdBLSQDHOd3RzEsMsx42uxRUuCRUCyl
VhCU6rJaT7IOVeN7sYQsyMYKMW1zDMJeierHhXIXdAkDmtcHl125sLk2nd+cCNfSBF27c1T1S1/R
DItVRE9sElJbkt1Yk8XECy6ajoDCE67ZELcBzgsm7vedBPprjUionoN1acFqxNVlpqJGb6G5/oGw
B76NsMncMr/Xa9klreF1y/xkZty6c8cO1aqvOfmmko1GXJRW7452+6GpVdKOs5I6NoS/ell3u2bK
r3ybQGAQGFylTfek7uPzvJwCJmHfKNx+grYnu/YCSjzDKyaFvuzQUjjVaTfjclyfyzRWu4X4hzhB
VfyyhwcWVKAk/RSi3D41VbFZb4bKi/eP3BNd4cK8paDZ6byNuDZvxmCuU/URm0wLT7W0wtYUr9U8
k1n7qGpotdMBicDG3ZO6/o9obDpVTg9rJiNW/OCF1m5Yy2f4tc4hKwGxQd9CStrcpS1JUJCbRpQ5
C3ZkJIVKRfRfjbxSgokRdH8s2wZ9ojrXeBb/v3g+JvWPyhMMSGuBcQGM2BPna5b9gfvMOjyhkmt2
0KUXr+dxF/thw3T6NBXl5LM6xmBLQnnj0AfQOGmZNlZWPQDyYmm+OlUxQvzSelN/WFu9Q1LnzwBd
So7wqwgG24DLZeOxl20vRe1QzyvLGgdxa6ZLWrmfa5FUWSyRHbjKbkC9/WgFYkJkTsZlB+Ff/Zsf
mve255u3EHcZQ4l8Agpc7w3EuPX4qhXJga1+XYYhplWybukCxOK9YBEp2Nt5Ddh4HG3ca4I3gPLE
+UPH3krLy/m9S+rW7XB+OEWusJDEpb+k494SMGkemudr5YaArn3aPt4VNne3eP1GgOKSfY9IlMwf
HIvv2uVGy84JI690IB7exU/6yQs9SbGwIHtM3xwvZqyBECrHfDdJHqdMCoXIq85udvO+WbppdFQT
QdpHU7qzF5WNZSQWFA5KGyvAwIGgEgQtl4pakjgWSNtOYhNNFJBnnVK0jEORxYtmzyVWJ3ODMWpc
gmDYKiu5+jKpFL6wbvm1fjFoXPzMFtV6bIL/G/O/1Wligt2nESXw1EmKm8zx5oQZ0Ve/gHXa176d
K8gnoqInSZ5TzAMecJ01uHtVPRI/Jf/92qMGbEFkoj0kd9oKFBj3e/kCjGs6bQOgJH1vOHqn/03L
MhTnlbedZxQRcoLeu6a1r3N272H+HU80u7nGudChdgeNolamKVWtOZB78VCO/jdkin9RAwbnFo1v
1TSwkUE3rAxXWrASpZedVNvcd0qxtAEf2yH7A+bHUK39uJLyTvK7Zf8Nbnn62kfDxBTIiADdPjQQ
6zmjkC+0Y0+HWk6VM38bBLzu45ob8gPGwt9CejTlW1smgiO5eompLLpaYLkpp6Kj+f/6aei1a35G
xgJaTNSHnrmlUJb3rr4wcHsh3orrPeUqDovZQqLtehtKIhOvD+NEfUROPDQEggNt2aeV89EpcFPe
jKJ9WanSZPZ3nV70WAFLnpm4C/1kuy/d4LUSw8Qm+B0w2cTjlBZXvnSqMp/mlmJYjdtq83Rgnvvs
PkIPP8DmCqOUx78/91UlT0JhBrI0T8qCsOATom711tdWExkrtGRLwMV6LrflAkMoGNRMMolZ1PYM
5PYhqydqKe6KyTNcNCkcMgIMBaLAW4NSAftNi7FjvzLw+iHHmiBLUv8LWBpmUtogwmSkT0MqFf1G
V9zDmeCDObFnpap3j0RGRZuiDDmIR8aOMvfxb+7bDKaOcMqicOjSzqx9vIV5JHVKJxrb7mLlOzDI
QiknTMjTkpp2USQqsxTcQ2qMmzLP2L6nIuEBo+Mdif93ClSzDJfkiiHnpij016y8Dd8zTcQkkz50
3IbCu8jP8jg1E2cqIzjpapnwkUQyUe/RLKJf0lMAEzEs5fMFeHuaoLFhv8YN9lwBNZfDnm6I2rrT
n3zyW1xm1gSg2z3SptjdVZm7fkgwB5aKXRWHc153r8A98Bu0kwBTiI5iz2AQTbGn0RLbWuqPsgDy
ZQRAnl6ByoqAiXcrQqh4RnkCged3X0Rb0TL0ptuHcfcFWei5FTREn3OyoR/xqVAiNociEjd4q6t9
m7YaH1iZ15z/qhNDWHnpfCqwTHmz8kSCUV6LmpsRjWEZtssxZCnxIaKxer2EcLiJ2iIpoWVAHMNm
yOiG/ks/ovTX6yKajEIvHiKnYy2GX6KoI1Qg5kPaYFYmtng6ZhFfCIloYmiG2yVbiWnVFMW4sNqe
Xz/lLrPsVfKJcFfB32YelRBNPFWJbOXt01k/8H89mhkyksUllRkMT/Yrx7+KzXhThFoBR+rNMMj3
lq5wRvacRn9cleyIsMUwdLkqslb1ovZMiEn5+hDHf5uoXdyzljIoIyIRKy+/aw0gYAxy51cNdwk4
iyRiqNI2rWAqO9MSW5h0xTf13kRZFHthVt4HJNf3qxZTUOYUTScEIrzC8X5vkoYpt4NerKQo9oVA
pa/itOO5eize/LESOpWmoxTn+3Qb02jvcJ7T1SEzHNjQjJHvGNtsjmkiojzYvnzxjBXbrIeYtYsc
XW/D3OuRKd2jc8ecZR3rEatRSbmZKgxtHUgEcyyAQr6zC/fU6/Bp9uIKA4e61EL0ueVE7i010nRl
scV3DCueuxZBVjvX7ymCngxwIIyAoiHNB1yWylLckwzkbNeHNLXIQnxf4pKLHeCYlpRBA1zUJQwR
LedaOHHhIiJ/KLkVYdEoD8sCb9zh5tBVxvWeExtG+QHWeUmzHus3XLtKezDchDDZiUwctmx9lFDS
+QXQ+wdri6Z+8YeSuDwBFqiyN3xglrJzWEhYSZ8Ax5JHmghX6GFjFTQvLl1rveNcWjbgvoGakwVv
njh2lERYvdUg0NOzuHGywEha+f6pBs/DT66SiHiDy9seMVI61PbVKWfG1bNv5M3zq2xq1812pGsM
bwG19dRgXlboYLmPj2iox/hNIe8wYzwmW/zZ6lIW9njVat3cHoCv2Xi99c1CORvkBY2ZkwYBHSx/
GavANfxs2uSCmW+8zmuFOs3PfK7GHc8bvTiM89AKi7uheu+tBb+fCBkIJaXim4bldEJBrTFOhynZ
yBdQjpNDhnw77E4YXqZpo2gJqXDhXd/BP7JCLP/WuG7fWn/FHW7AQvSpbo+0uXLeXN7UpPv+CTf8
exBhiQOiR/U5yj9MnWYOVTrh5rQT+L1Wthb2czhMvzPBxg0+FAsKnxzxvbCFFjkpZaSElAPNMesI
PJci+aHrsFvWLHZW4RKfv0oGeLs+Ff90uPPec5gUkoe/uyW9qjBtZImaduxQXCzeRrFE3hxsoJVo
N7Da4SCkDPsb3BHqRGCLFz/CFyO5DJx4p9syod7XQW5dJD7pdBXiimuGRKD+IT9wFyz76S5ge7KO
+GxitK8esqFJMNGnrfvxatB4tRYw5K7NipamUdjJJ4Se4ByBHRY6mDT6XVIM3AQFySf0KxMHexpz
JScuiG9L8atp+wX35Po15z1pucKcS/M2eHtSuvX9wP3/lcRbvaOeeXuUNMdDS5n1ow7ZRrOoxe98
gf6LuEes6wmuJj6U+UG90nDc2TFsGrH04E8UJZLzdrw2EAdt/kPSxEJLMjOQRqf1gGO325zN5jzp
7wvYw27II3rOyoJRft9gTPJ303a4rRiMgaJ39yzcXppiAKbbiGQGrQ7OFqkneq6JXx4yqivfGkec
BQXGv1YdrlFxetx+1IXoQCd0QCbYwZp59pHYWPznkCeHW7crEdOmOVCddkjOI9EYTN8nwG1KQLmF
PG2+nk6S7LGsCruPzYExubkFuy/pk+SNf722UPAHvz/wsQibJ4woGhuCkyLbKh8lfV6uGCOii91Y
ECSLt5CQxN3Txwui+NI453KZwrT0EjLTo+BroyZli4+eEmHD/Mnog0n5KMLkCFnopqtf2DMV/X1D
2AnuUVRYPIvEWFc2bbZ7SvsfHHg52ut4hdH0Qty7ODsPIL1ztAlr0Q56kRlmlXGeKzAlzHtZIWVD
ODso31XOYiolcay3DkPxj6cyneJ0pXmbux7CWEwa/fRZbtOt5VLihpo9tUGtu/ud+stc+V/VtWZH
bOjIRGmKiC67uX/3EDWOu+riqJnyyZItST1UvF6RGeAGSE8FsB074Wu4ba6gQD4Mo4I9d7XOJ3Y5
lHJHml6hZlMpwSVaqoI4uFSHQN26gVO05k4MVt7uWwAxsjIxhvdUJi4VWTsDeuvp+oZ36k6PBLs6
KJ3J6UbJAsP1gx2oIhg+Ph758kH9uOd1OH1V9p2yRDezSOG8Dz27Pqs8cE56WrpqasDVjibtfWK3
bYpVRLctn/PDH44SX0THUxoq00SPOgN8QT0qDD2mFJosA6AdD5CcKOCUNHLxMvMJei+CCw995Oaf
g01wf6mx45KzwKI+jTJxKkLOBxGZbVeep3TKGoS8PjNixh9cE3kkXjK5G9Zu1uSbw4bgx8GJ/2bK
5JMT4IpgIMJGEdys/7mGt09H4tXMQH7LKgGUYBlvoynBX+QsRGAGfVNZM8ycIPfiGP3tKusl9lHc
/X7wrAf6KPlOoAzWaHuSGca8Z1oHa+VRdVW+TpPxB0YkMNLwncMqo3Ih3ClHAGXwzm2LQfh7aln7
hR9QL2yVo6QTILLMWVP2okYAL1m4GAeS5oAYbMlwzyEaf7emYEF5AIug1bYEoBYV5P6a0mk2wf9J
c2g1E5Ra8ozGCF8dVkSDseKoATstWcB26D6S+cNmcZqldpJZJx2147HW/mD+uTqAyJSdItxhsL8r
G7ZlcADT5edL92gWPG0EedhPtvFnuK8K4X2l1bcNF244/xTmiwq4rNbx2WmxCNLXD0JfGvDTurhs
kExhBvd+et34ISlXMQB9uLkUUQP8gk8WqisDkwf2s7BCO3JDBp2AXka//qI7IplOqgsgIAggH8Kb
oj+TsP1JvaMLH1nmgcFpW+ZfipkETRKWRygulD+qpfxOiWdAhCYoo7RiWRAahPQDEoylpvmq+Qie
a64Ibuuazea273KFx8YVHVy+0D4MIDQe6O5nJSlXsX5SDg/FNO9jf/fQEwaB4D0xmtA5zAseIAU8
jnF8UFYvxxhKzSXAtJP1lifCAAYnadVGsUf246wAUlDchh0N8AZl4X4tVe8NqC0cCtEPYN0k5B4n
xZfaJ1LJdR3FDkMxTv8nZgoR1cJUmQ53TQDseUsL/EufV8ppgV8HNtpgPwuhSK1yMHhAS+2/ScV5
mZwiZxHxdiID+X4zX95ebkWeSJYgE8wKhN2ej2lmjeM5YY4vPYEQ9NUnnRiZy/q3tiMude1jzSdL
azUDI8eDkxNu5YtHG8DvrB0o7b0gMSZ9jFmy3j+dxAMYH9ineS+RkV9lsoqTeLI2wCTmo2Z9zbFt
pYKy7c/PGA1umqtsESqsivhH4cpQWaulPNwM60Xy+QpUBKe58mApLjmIDPBoLE6EKOjGGFXjTMyA
uSAhYkdRvuRuyNcFRlkz1xevyWWsHkQECm3fh0pwOC8+O6Spl/+ga2jR3e6/Tx46hTobBqnEvSFi
HaRAAXXEFAEdYFS8t9b9u2wmeIN6Ycl41j34R54L25hRJmAPnBiZzyD4jxOXjUGbVdb6aegA75Ct
JG6HBEia9iGQ7o6LH6Bpxwo0XU1j1C6VYchUz2o89zIdkjroE3spMaC5yEgvqbyeVMR2IMQ70sNb
jYOLrCJPPhU+ain9//qYge4WjAgsgbNIELYlLnAyOgZSs7dHu2zcIJI69b0e8GwzTDJExz0DNoZr
JQLv7BBeHZpml6skY0quOi0RrPYOjyS5/JE/1J7OmZHbkuBB2eIl8nhDxxwZuJnT1/koaA8JCTxj
MhsHltdbe3c+7SshiDmahkfjerjRf1pp0MpItTZ9W9RZzTsb/e+xmG7smpgXoilBck5LaAlg/sIY
zvw84MHwE9Hgjn5oYxyGy9GyqSANt9AB+FMjEEbTsG4+2rO/SZEMzfcff/Mwy9A3YzLYQuydo6Sp
mjWEMZgBx2dAlXDtH5Jn1mC7GvPSjLCaNmXPSYmj8mlu674XMau24O+K62SjqM31R9hVSmGvgFRm
77NHiNFpdqBrAWGxGhB+GaI9g23uuSLqxXYgPHsnGByUt2Y5TmZlj4hW9C7QDS1PZC9cqon/DAZc
eWb8O0WTmEd9Iq09ohwLSdM2blciDHcUdgjK/4ZCtOWzp8snQBPJUsyFIw9DCRPvCBn7DYHB4RoA
hz8NDXCdWLJ8t+l/HnHIL3dE09MjYeuxl0hGNiZ2LbVqY6a7mi/oII0vVq+t4OBiXmvsgloGfdPF
sIOULdJOtclwgNe1EYaWSqiRMpj8JLtLmXczR9QvmSxjJ1jv5O18E0ir38BVJpdY4Zhxy+CIzmOI
Fc4YAksVwCtXprW4TO91apP9nRHp+csLEK3HW0qZ4+LF/eaiNca7cltsbKyR0YDkGOOiAhNmmh7E
+RdKj+avYGNusPiCKgoTldgCW9JO5DskTzxUAv1sHTEB12SZeqVhBBnZojfCeaG9/rCBtJ/OFv0M
fLGWoIBKJzuD1Lh0awD0e22lAnjXW4hL+sA3ogsZGV+hhi9ovfvzgVZr0QQzO6CeCHqYiwuu9MJS
8fCqfBgrzzZQ7fehwo5xGLjZ2/XbeTgQbjRqfo8Vl7iiWaxhuooSA4ocblojNXi85s8hm6ChQb3y
EM88r4m3bwmbCMxbfQcKc7mY8qQ2axULT6v+dNHx7SfTHZHAV7j5mmq/UZKjqOgcIZNY3Q2XnYq7
2R6fblE9qLFOfU+Di7NSA0+TpNTrKUKB7aq8y2xHc5W6ksc7T0wKDTMCabllBusxbrwMYipFYKcP
wdrRHVbRHiOigTlYHVwgAiYGsFOZT8QE9EKRtboQ3g+2S3AfiNtquE/7ZuEKQroBerBGn/X8G+3B
qQL5+K39FrIhRv2fbr5tk3hRlDNvzlOBahd3KH8MtvILdRVEUb1/Bl0TSl9V0qUdABG4V1Ceghp2
MxSlG5eys0ybFSHRcMYZ7ZidgKns3Fity2jXNfBzLRnT3gae2UbrM8FNMCZ4oXR4aZ+962FIB+kg
vYDMGC7bmlMvvWR0YiCumDQ1m70uAU3zMKcNbSoCBnfgpJb0V+6TPlcqiKJc1QZKFYiawAynbErE
XjmQKQBxfe3nA0ULfBoDkYB6fK8uEN/K3pPDFAKnxu8foPSXvw4Bp3B7jMR5sxaN4w0lKvXxJfC9
PMkj161D3txf1oDsUMDzeTL6t0BhZTLYAAMD0t8oRUsfBVe1Y/dh/9XFgDOu4PJ3BE35/kEg1hRw
Hn+DPAw/qJdl+HvhdayNyR4/QY9TjTP2zb/zhnrV90AsVChbmfPrhRc+kdGm3DVWfYQ4iNSm2Qon
/KvtrSopOINsnU/omKwVXhPb9Aszd4HY7YzmIkIN6wmkdas/zdwesbEoLsUWZ+KhHZEXKzUQLArb
uZWkpQFPp2RGCLXN8Cr+PpwqjxM26/ccbaMbxR7iYPj9IfjZay0PBKhbw+eLqJTvesDGjeKbSs14
KZs5rbeRrjP8UzsmDphe7BfL1QNRwXr1HL8hHbNmUXP0vzlDr2tNtr1Vz7GtMlK6uwy7Ie1SXeT2
L93hIcwfpitvpYdXliTldl/N+52QHqBpGmrdOzFItrEFdyK+/BrTEqz7wGABOuNSNk8wCVCjIOVz
dlQjEPwfU1aMO18cWVleQJOOOUmaAHZ/XX7ji/RfeIyQq/vV4Vhw1feQtjHf/cgjxD0aPMiQnZ0Y
IvSMrONl97cWhbwlJDMnzUUSBC1U3ndw4q+ckUIn1jshgIGSc2+LYMGVevdN8VIC+p3GUO000i65
SprUWrcwsLnqXMpTLUljJ+jSJQYEEW6i4C1JJZ05JJmLmOtKQq3N+LjEGDSqrSP4tihCIRxjmC2+
obwYn+vFNMGTI8t9+bT1ik3tnxSFpdb0VabpO8a2TXJrhSaCW63/uAnHdInomX1UhTEI9wmDhpz+
/AcxEkx4pKWmsEaLPNJagpdo1nnERGuwg6xC7n554OWX4BtwkRBsLmo6ZgTFw8M/yy0dscWZsPGD
0OdK5vBdbu0FDpPP9jL2n0Er/P+U3M/8evRtkH4gw2FGCnEm3VVvh18YmQ2O6a8e3IdVT17X0QDg
OMH1Xzfpndp+n1KqiMi5GsV/zyfYYPxvmsk58KXl2ntQG85AcxevjMkhxr+RmI7prMVc6iAIHtrG
XQRphb7VYyQaDV+vCikqad/fotdUSp/Nscwo8x5jVMKp3wn+0J84gTYIcnrOa80acVf4kWdz3RwJ
tFlgqE/21MNOyMhyz+AJzu07QAuYnEKcgzSVN+sejNX0e57AuJHDP1Scoe7oYoWjtRcPvKx2zGEj
E/qJDJEfnYkkkrkhSfszqng8TqSycQzmXTnxMukaOlGC2iPWNwTTn4pfVW00whX7QydzQ1lYQ/Fv
vB/XYNhRjHhiY5VqvL4EjLrm2gZqyjkW/LH12ZRsuT0i6w67U3A0VbHrlI5yPlOEN0NWYFopGOdu
VEtCra0Kc7SCfIfLJxPnjPwqaimf49CYO9fdZ/S5gdOy24ueEpKpPi3HQEn06B9AcwPo0L3oNWyx
UFJisRhBHWOVNlJQ/5GxKXAD2Iegl9t2unuHMlrQCY6z5CyXgctiljFdx0DTVMO971Hdvz9hGG3p
2NenVDfuxYSKEhRKd43d9kpSAGP9K+mKgMaeU08+LrZS0Bl5LCD06CVS4ZSJsVDYECFmC9AsWOvi
XB+GXqs9+1nVLdvD6RXB6SPSUePuTpwoyn+n+dSE2aZ2Kcm4FoJPaZz4ORt4nombkQpNOxolyd95
AaeyhZygVErlg2n378ycDIoh0kJL1AijWg467betfFQtmpjBfPi7Hfg9HwyzAMe3xOeTjErTz460
GD6tG7ebwzbAC4/yoTfxNOc+FRSc2vWnj9zBbc/9kirmI1iR+XFLMlV7dbulXiVUa/TVoK3PKCeA
pBKv+04l4xkOJHWoeLulLG9w7fzHhdTdcTUjbQv70CgziixKJedxtNzmr7aPJXIFJqIh3nLTHOxH
Ad3iMs4RTuTJaJUGPtRkLEnyb9PhIRT+RTF6S/0dpbmTbDsdu8BVyyQt8tjh4rpp6UGciLHgYRqJ
+UQQiOfVW56VhlRjbHCrZsx7vSwm6UcZpoYJaYUvoPM9QT2iQF9lSpCm1TOfqfl4juNtOCoBqQsc
s/P3b7jWHvqac/Ss6V73IGHq6YM+QJzse2MnDNpnCyTPtHw8Dl1bTZNEO8iXcA8KzqWd9sm4VeRv
ALwzzsC6i02D11lJQztkqrpd+gbi4CXTYvsrjN8Sja+XFOh6QiKuVMOIdcaOTjOsKa8+pIvPsN/X
G37qtfSSW32QFQ79gpoyiU7uhPhB4pCbDGzYEFsOq7343cdW0cW7oFQNCib97YQxhcYFyNpXNrQ5
Z5VwPfDwscszHOtF1kmema/dDpA85aqcFVafKw1jnjRzjhWOYQtebmmmLZ6tyigTXJTBfyPd2nz+
rooV/naBxv7pC0JKxMnEBe2ipJlUsZmgHhFWHamatdRGJpSK5wuGTuk97JMkfOFiAsnGxOq9BcEL
b7yT3cXeX47MPFInr8NSen+W7MPjIrKTV1ggwRISX3szhWmku/T3IUDNE6mqnh/8qu/s/SOy68/E
sKKZ/zkoQgVHXZUDHDklYtibZMfeQ2iI7kY+8aoPvz3iJcTpT5r67oygbNLgOa0s2q5esYrV8dF6
EOOySkaVG9hR5IqPnEx+VVE3jyy1KG7WLCH5jPz3P7n6DIX1MTMHFUCDk1Gq4b31uzrEptZHEaK+
e8YEa0aK+Mh71mAQjbZeekMgFek9rZkUZaLQvwUmbESlTnw7uLKg6b1XvqASxf5j6hLr5kRZlvMQ
IZ4kmKx6NYMpbQGiMjEKHkcQ0zauQ/bgHvs9H3LFwx+q7TvH4X/i1WdqTjnLMnPORbef1Qbx07A1
6aQDE9sP3aMRrxlKVxWSBB5EEdmW23iu7GHUpIXY4j29+lGAf9OecrJHDD6jh98bKGpvYXaKYDBV
gvVfk207HQMR0dMQQCyQ+Eyq8EfQW/sGxOvZLJOMVfT0v5V+gFPUJ0io6DyrZhFm/RG/BUnNBld9
jzn7aSHvaHVZooydGKX8GZzdsFs4EIQZpKEHajXUsn9AlZAPynvDfd18/FoQqi6mW7bv+cxTnTHb
BhMKRh1JDLnNUawdz4hGjbf3z3VPT59KsJxKdHULHGrzT7ghOWVlb/MFgeUPcyE5SP9ZAbnMJG5t
azDYVjDT3OsZEQap1zAfNRrbR+Jy6hMfC/FO7ucTr1XBb13jYc6fQ9nA2V49Ak3GVlMVW+P8TCYa
EPy+7vvLt6mlDp5e28PZDn/1Ehc2eORYsq9i3mcZoxDZOxkIHQJ5MQYV940MhH1r6+iwE5kXcTcS
GFo91fhhLFHhIKaFqNaFxfIwjrt8i3C/j0asCDv6XkwXQ2i4wIJUM2gUPNhv+PLoO0wo+HtdKoli
gfDW7GIh+rqgdYMQrZ96W5xDCJkRpcQ5IQ7plH0w556ho3mLL3QwRKEz65PbD5rT9kvH2dfcle/K
ztuNsz4ZvHYOABc2KEyT0avh/U13FxSjRXbfbEd8EcAoGrkxsjlpMwUpux14nrSZHVm3dsYiAQv8
0AakKtiztGLLrkcVasDgW3pY8gj6vU5tr72qn8DMto0A8Uw2OG8U3Xn5JzsnuNqofgfHf6pVJQnp
eaIPmPDp7cKWL8bwqqV/KTBU3cUvrB/2iQAp/k1yRxCtqPuJ+So1FeEUWXyUw2Rlu2CKYr4kgAcJ
dAG6O5V+yqg0yrmodybkfkbFYmDjHccW+bCKckEO2VD6PHpROdm5ADKmIPqipJJPA0L8nlmRAx/E
0K09E/Q1URitzvKPPap/Sw+dLfI42U5FOdWzxX2bhQo2RYebeFNlJTFVHEggLdUucFw0rSQ3ycGI
3kp44ZRB2shySc6idJ4vz0PN4EyGCH0AWnFcorrhQlwxuVd9uGICxzXvwdx1VHrqYvJvQ94gWkiE
4mH2QJyVIWoLcusgRzNHAOXaB3cl6+J/doQGWd1BGDc72yJIBTqugxucOfrAg3lIGL7hwzzEkx3P
L8zwg69kvylMtVDRFUG9+au6yHpBciNpgXbyzPqDZK2eGJ5xAYM3qB1u61pmSH23Zt7CX/PvLdMp
gci0qgUA5xHv2yujXpoSvHl/JEcnuBgDWUaQJH146cCILniXN6A7zeSyYNT4DYbaGBjwcvstoJNE
P2xKzQkgbLfptk402P4TLrmZDunjNX0yx1pJEk4HAdOP8xYZ2bG6WT2rqmoaKsHfY/PbPien11aL
hdM6WnGdiI27xmcAqtH65KiN1lQBKsOPaqYzeclFYZuhmuDjCLYCX01YjzQppD5GhhckNw31mVI0
xZOwVQgBDjJ4A8oW2maTfb3RIlVYnlUbgzU0s87662zPvTxzW/wa7NI2I6XITd9ZGZ3efuR8ik66
inxag+JHjhOjWo4As5fIG6u9PaCoocRGr9P21h+2ccKSf/OcZrsq7OO8RzNAG6O3ZHSrU5jkM1pm
7aTQfHRUzVTkuypwFeQMsTatKerD9PW0oo1+8zuVrrv6hdn/IYepkorlC7U7PmzxhkgzVBeeKqA+
tXffZI11y1JJo/h5+7YPfP1BLcOhz2Fqn8PutdHJj4Knqc/PY1zqL8pS3APQz4ab87QuWfDrlR9u
+k4QqAyE9Ht95HrzTWLBe2Eukp+CdBkCloXcOKJ3eHx//LNSjwgCWgE6Kh5oxBAvdzcm4yfCl+uh
O/o17jlAmEax5hsE8xAg69DBJijYctwjsvHNL1h+04S4+FX8tpV2IjLR3cHpkeqvrBrgWHaRyw1H
po+XaegsVcqheWuZPiiEQKx1zagzMt2/d9c8NRQJBO9SCD9A4MQgT55SEdrd989OfdEWaCt0GTSZ
FOU1dJfPptsk53aBO6t+6P/SVtfni51uZr/snP57VnpLB2UeouFQOoHJ/N51MyoD6mbCeefCArzV
nd5SzwSSpFb1TFK19aXqHx/+g1TM+fzHVsSfIdMY1cBmtLNaOuBaKbkMAb6oFtOJnefPe3Bxp2wX
1iB9TRaEUIw0gh3rEv6MHCcaXXnIOhrrzRiDWazzlUcmwTfApUf/NpXP84Xwfsejt4bCQKAqYBGh
3aSmBQjwxGM7Q6bH6n79D/y22b71qtLabbBGuDWlcji+yezS4k6Y96TAAxL84F1KUoC9x/O6jDn5
7zgn90qWDwfeGJ+C2905bu721l8Wj82zb9mnrE+uzxiolpnDmjffeIsEIZy0DOgy1EsRuSxdSl7k
s05tOPjd0vKU0VhsiGhKKmj8XiK2APc1q1MUUXhX6z5RfaR19ZEv0aNDDTUn8dzc2yCNERBCyY88
W3gEgBIuB5WAEeTAVBVRPOblZ6ueOOC73hH+QgL5608ox1fxmGwNOKrCTtB10UEa+c+cU0Q7gwX8
bxFNzJ4IqhOWZZXT8wG9rEIm21vZZaNwqNPHDuRPtopU8p+r8BQfilxWl30L1/RzLJzMYX81tyED
e4jKynhCPR7SzPPISiBfSj9RF0FGPT2ONxkpEF8OTHGVafszJbzQ9CRuRaWjSnM3t5ldUqJTcASg
thfshiW4CICgSbPW376Hk+fRRKj9LRjQxCSlaXTBGzJCGDTpAquj6gK3mxtQvH09hHCc7tr5EXUP
GKels7E4r39KFOnSa+F49qMbLbLEh9m0eQwSGsJxqbSobh/wg7EWd2I+RnpGOWj8wOARiyH4dIP9
Ido4SY98P6j6LP9+jLTSPdmEgJzfAm2y5kgObo8YGQK3MmVoF/1ZX+AZSH9SRs1pz5sz5bm9Z/Pg
Jjt5fMJmkYhLLnH4YKtxkzxdvKLJSw8+J6CCOTVaVn1zkaItCpwKblwYNqSI3dB6MFRcFQzkrlQ/
ZC7eOCG83eiiALOpaALKAaDN3iuBJ98OdhRr3TwDvjFEL+OzNUDkahum7FRddzCGsRJhJJ2ZrIox
ga2d4rUuTPEI+6Ph8bX6O3TuxBqnOkJGIQb+khiAAUloxHy+TDlfAB+kZJEfFcwauq/f/uXY+7e+
oyyZDeJBBPlQt4j4LNpixeHbYrO4LC4xmzZMgGRQ7euv+tVCuxjOIw0qUBGtSbDZlc/M0fwm88OM
9qwrQEvlMChRPyUCKVKe05SFeUBfEfxtuQvyNVvUrK0lZPKHeMvqFIEOKinlDd9vLvtqA5kNgcJR
aQtAAFKADu6dzZndAr7p6XCFqKfC5IT9+zpEj6OTH802SOk9SJ5pWO4H7RdANGeXHnTxh3/5/+tm
dRun34TSadfcHKEIMRzR7/569wa6qLg4cKZIwQRXuJvJhAa+qttSCBXBOujxDe/NPmmAMzwJ85zj
e1EFe0zG34RLPUZ56t8EGOauhuSN5M5up9RFASS6GkTWNK9sY8tP810LZrKGZzUfc4jhLbZZryhj
vI8T0RczbAdVkdBMnOA0VW16rXBJGoyjBZM2j2EY5+W/QEnIgWAGcjH9YpOzgrZipxuHd1+O08By
5dXRWHWZrCXfZ8mqYT08j3/s36RI2iePbTQX9YG/nHKSYjkBfjlkYUcMaSS7qLvmZu54yci1i/tb
uj3t2W2cppMLJ26DdiwvwkufuzVsNoZvekhXGOk4i+3vNLWrXWszbL6aIc7bPfc7v+4Uq9xC0AdE
RgJAGIp8i/u2knhxZpy7YKoZHasUoCXZ+IQWcc2nK+JViIhlgPJqmAOW5zpkZmtnE9vhNqBtVAzt
M2zNGMVMNRNif2KE6EOvlOvXGIrWGPAfOF97tgkipKV0sfXcmpXug9Xmg4h9KIswamo2KIEom0cE
SE+4DxuRVQdl3947/8u8J5nZmSx9IATiCWpr88dH12LUXE4pFzrs5gnjNQPA/rrYNDH9HWfR7nRB
PSWOSmmgZITNtM9uhz/HimpuomW/gCVoLiIu/kyHNvT0cEusqO5/Epen9hze3eLGFmEwAZxaE42q
Uye2O3M5KFj2Zic/Z7MtNjY9NyiIrVZmdzABZyZIMxGCJgdk2UEcKZ9RlrutaBdreXASIvmqgKUM
y2tk4fOqHY5xK3TXSmCmhOHaoP4KN7ViLhQoc4/qhMF6Pabm2XhBN7ZoDySjufjvfUUFMiNSz3Vd
xUarc7qRBLs1HQa7nUmcj/cibz1TYxJrtbjLrTvSKkCLNOuW9IKnBS57UqDUdsCYxcQBz6uX5Dwv
fXkj5ly725TogxWJHfgS6tdJHrotcCObmcf5xUL/3S3RBnHCJnikPBuUUkw+VTVwQFAf1bJgUakv
qMLXym1kVQDdHGD1Gi0a8LrX+gGoC3/72DHnLV27uXFqgK8kDX5EQbSoZNp1HTHSuJZC7hThE0Wy
MkefgYmfv1CVZLDJDj+fgML2CAVEpHshv4eJLNw7nlqWoMVnDYiLFa+P3ED5HuQ8zJN+px1eTRDO
I6SkewX/vZc3D6BKMaHXtRubpM7EBlpSu1ssUGKtnOQh9CWtT/jr9SbO9dxzTYgoqlQv3WKZwCUv
xA/Ue89AKFnaNnccYulbC6qCJFJ0wsNGhK/QpCGamZexvSkqHXHdI9hzKdr2ntlagDp4WgkEdW/C
Gygk7eghVmyOVGptTBG0fZLcwh6/jKl4IwURsgjnj3w5Vow9SLBfKlB0gw6Z8THIKsZKE/WUUGTX
rhi7fzN6ksFXr9MetOgsvv49ZHMzdf6YTJqlcwe6DAyKbHEPULXW9LcKazLzhouOxJPb98xwGM2O
9lN0nQjh9nGfTlU8p9f3BKAYyGeI1KVNhyUnP+pF8Y1aUEg1dNay9xPwrN/nhPatcBrQO51I6hXz
yr4UyOpLzlhuj4g9hxEGVUpnfDvt3WYXbqabFihfJAaVKbKpfdV6YiP9JSDCmX8X1IriSL74p9mf
5lz6hPZygcwg60U2JyCRmljckH9IWhe0UQjaxMI8yluOjZNU9qtcUZIqSBIxYECnMr67pFGaVMWb
isCek9LSyyTqtSIM26KqHLJuxxL7ueR7mI1uvfUVpe6Mc3ZvGovYWssfEdhjoiU5uYnOLjJ/Z2EF
34l9/CFxzE6+6a8ADmDFifG9eRNFnLhsJi2pvVAg2tqCvL02w9lrG/kPH0U6bI7jMwRihqoYfrj4
QdCEpVtQC+fl9eseDICoTUdbUrFfHcOBmxKYz8U2CDJzBA1os8U6LvgcdYY8gJMhSz3kzm/yqs3g
VHuVncMEfL8G8FUpGJNY777euIL+snBg6T15V0CwvyW98f5hsTgP2g0hYVWrQEMg7uQ+KSh+P/uY
rJJOpXAmSvuafuoM+wwMf/m+l31js7PKg/n+N4vuNzMJCsRBseTZsdkdAART70d317ZCdifTY/3U
yHag2wyEO2obx27Vc1uyZDhZKsiyFC/jbq5wbKh0452WeFbWMGLo1QS6sas7Y/Qm6Zw8N5QAMkVK
5KDsSWH6cZ3jKs6FIEwB/imM+u/UUHbuwSCsT5J9aR6VCLCZsc+7581HdMsKGbiB/A3Tqm7w4smZ
9nCUgB1ExrQpjGXyex6SFjYn8t/LedVtYeSfkpnWP3+9F5IMW7lF8cGr90dJWxt/4J2PkYJjIQG9
pa4XJhMhbaKrb8Cl6Rfz2VgR9X14Ef5b+10Q5cLSahelbrgMhf7b4shNj8pziXaHtO+Ufh67nhGP
P22U3WKAh7u45JShhReIUlBartlbKMSlojg/cKEfnZ+iK87Eull2yGMhnqeHbfR28I7T7h+lYyY9
ras0n3IKuAUmDy2nwraIdkLGzF8VqXqn43bN2iTv4cezBo9UMK7pkmCMV+Lcm0/ocH9YhbeS3eBC
DRvM9ZXfb+dSobmBE2ycxyicwn3ebsBNvsmpKxvy9k25glMF2z0Bwrs0y75mb25Nn7Y+700eEvfa
gLx/EvfBBVY+D3CapSaze1IOpfTFNg5ooxis2sqTkI8kCz/vs9YRDWHa/AGTW2bHU9ugD1+Musqf
ueSuabrhLZQRLq1i2G6DN7Y1bAAtT0PMm6Kt0LPq3fg8uBKVQo6BX8znZP6SQYj6UXALsCifof8q
GgN2obiUAOzHD2PgJxtXa8dJMwAbYes8xISdU/6CBSzd6SDtjlvBHecBR65QD2nOtcoA5tOc2RLU
Zg+rmZmOzICByQjw5gwYElkttej4RbRuxx5BlqETRmCXfHY85EZQf2HCfIimkhlMvLL0e8yG1ysj
FmyJy1USEf60Hr22dxKBvOnrIj70eTLuTjzjiYXBYdXFvTB8VDk4biDUDNdoLLrtffUX0oZ7mpvO
kVgIA3dNmZUNkqNLjfpsF6fy8iSzQe6OcRuqKJD65ur1brBoT72sABZU2s4At3hDAtltkMOYznKV
hr63lOCpR9BV5bBQLC7L6AalRR0uv/+EOIcUJv0Pm1hP3u6MTiFWqCbLBjNCFoVUBYSINKulNgs9
zm6nwwapIQrTUIWI7ksPIGlYJ8A0EUcB7KL+Ns1aIg0Zcet0VB2iTq1RdISA8etCA9jtPOHPI3ng
BUyqNGpTdFSxrtK6ygwCKb12DTKBHhGQPOQzjK3mzHoPs/JYvwLttuzvMDDTWGmzq66xk3K3Kk8/
YDdSSlm3s23SSE8uRrGI1Wyd3xVIWZ5miI1W3Y5Y63R2ggGcRI2oqKiyjP74jE+9luT5en/gjXtC
xz32W2r2nW0/deoe9Vr2r1thI06RL+wBYTrowFLtch56FvLEXPkW5/mrQHEH3xYWUP1oKH8CCnZj
EFsGM8JDZQXu4AEYrktXydSwi8UiKfPFxsGRnpPjm2FS5EFg2/PPjNEWYQZK202Skc2Wz8tPGWbf
GQOtk4Wksurp+vpx+a4YqTImwr5NKwKrH5daiMx8yNfFRibAMFxxVHmHSG0QLGUr5zCGD9BVQvll
PPv1mBT926ZdDrxRt6MEohI+jaIngzRuxJ5toJotQY1YIQYsNa/IfATXnnDt6BnWL9wKxkZoGOqd
ECR3z+fW6blLHGPdZEX2dkmcmoaMjHPZ0S0SWT1S7aztjONgEzijhRbt+c5BMHbm0GqO0n1cdfGJ
O19Kfp/VVKLc/lVf37UPH6+gVEXdfiKwDKhms2MxlLPfsnm//FqnV7l0mrsb8IeqbZft5ewOGYHc
L/Avty7Bl8C/RjW8X2YMK8yU65E9qWcWRbQxE2jBNADswG7JnHN5dc7yCWMnNIMc5iZIOW02EXCQ
+RYWv0mMFHuHX434xIz5X7VvnFa6pSRaCI0FX6ABDWJ+DNObyN2zN6keDUulVCLdgYgzPOuELzgs
VddbjnK6lr2lAvn9r+F77kCaUIqGiXKKhWcxsX+xHGggnrP170eDcYBnsGO4PMe6Skbaa/ST+NTd
bUllSedH+cJFTD5INyDTI06MesHLzF2o0h3XJsKSFlaHXEB+nS84iz9wtpIbrAdvYAUOolTW085d
K1JBTZNEhDYCIOj7CfoVruc7YLFBPVy970u+0O4ojd7639hDaLvbHezKZVCjI+oXCC1Jv1MwMUwA
eQwENFUxzJ1I+4DtjPFLbd3CDueepYdGvYHiY/ZAU5x5+EUpyg3/IhT+6kTd8azcyr5uyRF0bhZW
OtNAkkcazQjh2bIeHTeJiSurIm9s6E7SYGatyzRGo7ieGin7+G66GyKVVDvsEK5NIUveUKB8FoUO
m91wMAfNv2JljerUQS6lnrFCNLmlJd9fpMqviIos5BveJSXeU5/Pxp6sIP+TiHAKqdw1tvQtbZ9/
icHvx3D1G5xx9SsRNUSHoCc6Ovy2vfbVPeqUedtneSouBdwwsZSrOiCYczHl9RH0Utvx4Hn/MwGV
Xccpo9mUHBzh7bgl3O+rawo4jCTND1RXnZXmSoXBpnsIqo5YB+OVZic76de2qE458Au4NVCsyrxd
Ft6/46Tj0Q9GlXRm+/lE1fYUpV6s3AusW0bLTsf+kKnzem/8m30sevkeNU9tQvMYH7p93ZzzyHrL
DOe0B/7sULehPCHvYuXgHnwdTb0tU0EZlUnAlcNNj/XwQjZGSUnj63d4Z6tQ+oaqlgXEmaM6GVYU
UjBP7HYMTtlDdn38Fggy9OknGqNujJvmvf+bZS8zE0jUedeNAEmySK/pbkkFLBxRQ5YgLIgIvsqc
RlD5SUwiHeyUuGU+S7cBEJI8KWDNw7fXVZl/MBYvkt7pjDU78KOjmRrjnrwQk9r4n24R9lpDMiVc
CS2SBCogk+UEDORdY7wQdrU43DxKWYEPC/kaaFK/BXnOb/YSeAaiocmPw5p+w+HvhpWqbu44pc3D
bHG/UiwFLpMbnKUXJ452TI+SGbDqrtX7S7wRCCIXVKDhME3n8JX/ss+FwueHWmVN5A4jG8aHumgZ
EhmWt2QSCIrE+RBDMH6Czx75VyQbalhpA4InLQWXKf+QItC8VA95ilb+OrM2D8A0c9OFKPc4pDo7
5sfDiDXnEbEwJv8pszP7R4QBdUHADdLBZcL0MSHG0EVJr2vfkfuq46fpz7sTz0/IB8412A5+4nTu
ta+lPjPBctSF5nfd5Br+5KHKv5HyJqiIlbJaOUunXdrIm6gqjpkLs251LUoRpocnGfYLWhWcfzTv
p+yi19B53RVYubFvDoo9dxVtK19i/V2z6KfGc84nOR9iC1EogmoqjAvFFdhuX9l6nairMK0qs4ma
SVB/IPVnRgZz+8HlUe1hzFXwQNsZt/8qkThyCUHzjx1y3M/6sxZd8cT1GSmWZO8Ojyg6Al4Nj+Iz
RseFaMgD8WBCF402cPxU0yuA+bSn75+B2cLbI8Hl4uo9FR8j6AIy0wm7hls0yW8f7jFwf3utxU+p
b0IYzsFfefM8Og+mYBgvDTrbJBAUssYKOmDp/GJf9uemDs9CFksmwTyJ33nwwrdLOo1SMLRiyk1d
ZMW8P3ThlV8vmNLgalL/AMUrV66/nNSwjDykJTqtiECcjtVq6S8HuAvzRl6nUbK7bi/xsbn8T7LK
5zWaFHTpg3GtL6UoNlkJVZnhSGjsL7tQc3/MU6DSqErCfULY15ojwPcaH790Y2rU9nBwNJ0ouvpB
0rAhF4q4G54IJ7J/Pd0sEyjBd7oc1RcPH9IIl0Nym9jxVxZdg4GSXs8OVIsLB9n/Rq/aZIe5U4OF
jKcs9HA7nTnokS6cjinHaGvdk2fnY/JY9OL8/fNoibjscaFnC0FQs+goSFb6wJKGNFUCWDwiV1jf
jz/1Fvu1eEXrkFNo2JgVuzHssyz3xryxyp7HqOZT3epkCBuVghZG3d8VUndZqFL39DBQ9abekx4x
zM6VxPc96spuxAzV8jbcNdeA3l0fZT02zcLw+PElxJQTGN6bUJvmGxhpoC/zrzEA/wmvMcD2TbgK
fFytg92A+uqzyscIVpBiQc6IGSlgcGU7uYV5Z41ATI7SNaFUzWDrc21RDMEBn4wcubxB157cPJJ/
uggkZGPlFlLDp/hUzUjnoH3leKNNzNNrZxueKskyQiTk966uZuUltfCZt76QhFrS0ut2P9aIfA5u
GogDVBYyg6cz9GUERvs/XPFIlOl3fXGZDNSWzUn9eTzM0YuetT+hFTdj8RHQ5m2TyKcD1VnDvxZR
J9AV3gQ7c/HGRhA4fkp3GvHfzMQRMvDZsJVy00rjujLVoMNzVGNI6KtaV65rsGSQCGgoTdOmJS3h
x5p5cK0f9ciVEdUDubcqDfgDRZSEZiFUJPcJ07QHYgsHZMLpeXB1DsE6KG8OnMdJaI56n+Jj/W8H
EFBD63tRJfKBno23nNLYCMCObhdDEG+h3XgLzfu81sR8E/yeS3w44N2iKtzCKD5XLDi/2GI451Hx
nMf/pkLMKDlhfbwLQe943l57XxjAvz5E3og3ktbSwXTwGGpc8CXlGpilpzzAIs5xfcSaCPsG2bgW
Trq3GmUXyy+tJV5IrCeRbtbajcdnbqpfe6ADCfbL/UjsDEUPRQ35UWlBupaN+8WfkgXDIxFPfzoo
9/HyVwTXZYl0Zu/otufcqM/EVgUoihoDoip1Wbjs7Y1fJVOsgNimoznKRL8PDoRB+VVmLNuApV9b
6tC2XUPI63Z83WLmIOvASmc6cJ7EMlS3DPrs1B0UZA425rHagzbeX/awt+4Ukw4eVVMlP/9lQmiD
4ygKGVfa8hsM5liwiCNTe21hFRbbCNMxl+apN9I3Vent1bzmJ6W8nTmjXxtTXQQqEpQ85JuCWmFv
BmIdNeNhAwMVgqKk/k2w+GeFwN/Nd9pTv3iAgnWmluYIXWM66FCWZnrj4NT3KEqdAJdTwpBRvwng
0rwHwhtG26m7ZtXqHVErzrdg1AUR7U0oQWD4uWAa6nbB457wvsE4TLEwdZx4CS8Fv1MsB1PnhUqZ
7t3W4RHgdTFK56mkzaRJHTS1FYIau5TdGwNM4+2pLAbFsgzP8KnTLlO0v1xVmqiD69z09ojnfvaO
+twDK820Rh8Kln1OxYtunZiv5LLthjAwLswkDML98Mop855J9gz6GqaAe+/f0ujfjikxzK2R3Gb1
q2wFfg0ZydNy7sw21dsWm2PSv3O2eGoSW2yINjPvumt1pUM3waC4Wh0lJ0JSLRhTynY5+FyWjR4R
WNfa405fj4+/2eopXMBIxyqLEkHOBuSpX88XbAnqyrx5sd9k7YZoQ5bdO26x+KD7ZAIS0vsxDLjv
2MQez7Xx/LVlX7NmM3cxay2ydxBSzAxpZwAaO0DaJKo1RCYEjfDRuKkMBley9fqNCpUWEk5fQygt
dwGppV0nS4zeAaBxN0UrUcBj6lufuyi/fGWv+EGoCgzJ7ifNVzffOSScTVfPpyPGg+b8EIE1H+J4
JwSwlfeu0Ly1y4e4kYQXlW9Dy0bckYKBe05QRaXijlr0njQ5XNPvUQwSe84heRzu9jVfkABRTBGK
TzdtrKOg3Xkt2Ryulcghnxqp3n1lEpNg1n0EZkHphZkZ0OV/baQQre0nOdns8uIWvy1ESeGpplAr
rDIwlllRpmh1sSo+wdhgGY9885CtTOHOv8Kvfz29HOqBk9s6knjwVz8sm53kP3eo80TkRZLHpM/J
CSmcxsBvpuW8t7bTQhfD9QCnRnRt4C29yKa0w66nBf4IFk7fziJBjKp+5YSNzz9g2i3Fp4SKaPAr
DHa8l9L5kiWOcuYpzjEA0Tm8MM918jCGDRG5ARJ3A0StLNo3VUkR9zWfP9IycN6pjB141dh5yxDa
5djwUi+dhmZDiK9go+UuP59bWeo+G54thUfUl4MhJphB0ZCexW8Rz+H/mJ+IN1Z1ps8R/x1kLPeU
9hmnL16KrBN27RH/8u7/7ehGvIic53g98Pcrssm8bcL9pKY9GMjA6ofTPpCPCzFcuOSdw4/XIBUP
C/uOrgrwp9t0H1aCc3mvjx4v93s/lEaYRz4RT2j32EEswIXzxCqMZo+rfqeoDTJ57w36NsQNdp3Q
JcsVfpvQOS7qu3VVwPmA1I996ZCDxgts+N7ii8RQyMfbvp/JQFsr6EMRTXZUhoW6JZiUxeqDre4o
4hwvDhoW0CmBbKQwryjDbaf0H9UbNDR36lWnNWWKyRuuuoY/AqQMHeQgIcGHe0vFMPIbUUdxNexF
i4kphG2sgF6PLjjwHTAH68A8q8FkwMXwmCjBt4MPydybGpbZdkAfJR0VE/ZKfgwLnopz7XoY9vGl
XfOx42bJZ8AhHvvd8+1oRVkC/Xy18CyLOmfse2GOtvG7+fUTT+dMUbtsvMRWlbw3goAU/ZWoid+u
sCFd185ZTjjzj3zJpZYlM47D6D3v0JRq7QGYL7NslfeBOa5zS9k+9NxKj2u1T3qK5M4HXP/QgQmC
ChNcakQFxYk62STEUCy84tg0HAbZrA0361Om/Ttm1NdmlLhiL52+664m21xX7WFKNem/h4igf/Jj
0dhmxsRVDdjYKTUNmjTvpcZ3y+l9oPeBqqPhRs69HivHNfdKbQedONM0Tfx0h4TBL0e3CPznbzlG
uB9T5J14PwbHQ+NXwWUP9BaI4zaMmjM4B3keVjkIDVZVKsXhsYXq9ChzZO0N1mRDk0DPpYR8Q05O
gh1Nn4LPBEag7cidFB834Frb3KKDn3lT8/yMDmOE7dDtR7T64wKdhE7sENCG47QW0tKKHxcjqtpv
H8ixuEYItPp6AyCt01fjevF2JHB9h/2k3w1eFESIR3E3XWbHnj0My10Jx2GQYM8G/KcUvgI8quWh
hRTsDply9JqLp3p6q6JcJ1XxZxEtv3NmHBOf6Cx+9nbw6sG+ZLjExsj8rG8bFTFWPp2bAsfyT4eV
wZvfLVQ+yw5yaEYb9uE70AtmvW50V+CVrSjJw3K3yVf4rywlwQAPK8yoS5EhDjXphzdFr+xYfPBJ
4G12cUxE+yD5OkiskPSjFlK6338dlMJ6yjjl2ga5TRfQUd98O4O6wwimtL3xDaDvvMHQIu2wMnKM
UPfkZ2p6cB+2OITiMo35S0iGi+K/DwPMCakfVvxvSeQMJpIuk+xVAbTBWO73c+GqL14TwZt47CrF
MEJnZLg/LGQlvzixqbFK6qYsbz19IkOkI2ZO7vbHeqY2Z2o2/q1PsW3M5NPP0vnHAWe8QCw/I88N
y7tIZEAp9W+RRjZUP2MK5eGyEfA7FARwAxEVo5xVLaFP+Awd5LOuCeG1hETO/aoD9SlvyuljR/lu
1SqdmsfYIKpcQty8+EXRPSjxLjPAHuz3tLEG7RkLCKJ73GAGG/rF3lQHi2yws5/xSeHEJvTDY4iJ
LlQXNT4lZt7gnG3EK2ZbsXzMGnNAuxjBWWInUBAXerveYhHukWqYRaANPRBOmeQtHQwyNtsFaO19
Svbg7euvW/T+Zz7GjkD6adJKvlsJvlN/js5tVorOV11t4ezqR4wIhQxQ+C8IixC10j5jOt4K00xO
twCwKfZ0766aRF3UDfcoXFmdW2mAnNbYpBd13fgHADN9zsAndJGAYfybkmFcDMK2/mw1GAeZPO7C
sfOWTu39tzG9XHSk/NcTNG8JsSO4d7U1rObs0yY3gFKrKJyedVcyxXbfz7fki+pzvnxtCWHz7ufF
2Wi3tba4hFX2u17maqzmmimHmXlo6b4J9uUJpDV8TIZJtSTuLVyAW+xi9PQvQJ1Vdfr1emD3c5XY
Y3KVx3G3CthIu9fwrLIA2LlUVJCkhG1w1IGQlFJZssI/np7b4kcXrNUOTGeVF9KpELXreEu5V3a2
+TNWchioiuKBgjOhkxMRPK+wAUfZ4oRe1r7TyIHNwQp7KCaJwOjwUL+cZtoQTq/tMgyVPxnAjqXM
7uHDQSYczkisTAuXEmMPAAqfGnfifM/jwgkgBjIIxQYXnmNuvjz0eGMw2EnC8UOACRuMGkP7h69p
Asp1g/J0rC89Xfrm75tuXceOr4k2K6GEPHCYKzNIoAg7jNfmVDBf5034PTdLdT+zSQye/NYE8aku
ILJ5z9zepiLmSMwS8NbHgLyLa1h0Bn8pjPdvB7Qvz3g/ZfCOWnaRZrdh15XaBL/6hXVbnl1GzdGP
nbR2Awt/cfBvsAknw2SzQrOVsDsiWpCxSG1hr2Ka4t7b6y6HAlRWl5/LDO5ltuSKk4XRvVZZUyE2
p1BvGhKn8wnqiqDWBD/xc4VCV0i9hEOiKo5BH85ev3Wyf6TaJdNB7o/zMnKxE1OGCoupI4Na4Ceb
7teljc+g3f81E+XKyeOViLePyR/E4qERyAv7U4oPXkZFyokJG93/2coKm6AVegtSCRJu96eKVgZq
K1Yx8K/LzQd0+oVoq0WGGtum423cUJpK8xvpaj4I6SpPmKsXY0KEGawRFxBfjkUefrYX+eCgh1w4
anCZsdw9gnCBAv0lybw4Qns6jdc2Rqj6DKKEkIllisC1m4RD/5A04d76fcdG/yeKHfNV9AahkUnw
aBjP0B5Yu/0toZ7bnMkWBZLNKvT++416fT7URqb71UP5VDMMLIXf+bbUmePfCAiSm3BxfaM8EM2g
sXGbWL3mwz+pz+S+AIhBXiHXnVPQ47RoSmxiMJb5wu/mxg2sKQDcEc86sdFe7mj1RKypqS6VjD5C
nSFI82HODcdmt27k0y68DwnECvxiPI58P/oRAEblEfA0yMlmybufo3uniCxt3Qdev4OZRBIjZoIL
pgOVCV4sypQuYmpi5fubWORV03XK2t5Ytn6LNmCIMM0zOumDJ/ve98kByN0XYWEmDwl8Zw/zpkQF
Kyzq5U6SKD/ySpPe5NiLv9mfwl6hVcNFTTHHLeVsnZ5MMJJw47ah+ATyFzPZPjO7LfBL+qnTo78U
fC4nyt/AnX340nx4bUFkOHxMC7oR/kymlE7KqsROsVntNWBEbQhcFWI8wY97MRUyfd3elQ9+qY9D
NKKKJDsdwgvPy4anB+A0waUCS3473LZcYgaFZup0ybs/Res3gj/6bEn4nabMeKctWh1rUa6h9t1K
+t7Gof70N3FadKvEOZyoTfSmZGY++LCcEwwoU40CTEwgC5ctTVzW1TO0+7eN1DFzRQKMzrX874ea
q8KHu3bhHS+13Ao0i3SGfHvkjVA1S3wTv+v8wHZGJr3MBBgLJNHTqDl0oCxW/CpOgTJQWmq2pu5t
nAnvalzSkjXBlFa1igfXAP0WAB/NctCId94grxHrwORxpTmizbAivmA5ooNY1mqWlXmB/BuRzqM0
YkfTENb99jOEbi5lCmGaTA2H4GloAQutN++H5IRAO2bqw0D/ZbSZLz2doWZsafPhLyC3mW1Xnx3n
+olasQmWB4Le8Dfck1rGoQ49FQE/8HhfHYSdnsJ71/kdn2ZBbwJlL1bmMjmRGjKZggW+ijnS7akr
BFdJ7HofXzEz3QUi+8cKVhjA+/usHDo7VddL+v2NwSZIqNRjvg779FgzEtAfm9EVF84mW93xWQuq
fX0TgMWjnhJkc4WH+Ogww4hRaKkGErzUQTGKxp12PRfh5AZTsyPHfKf07ClPFSkI+0iW+/5TXkrY
1VKaYc1U4SPMVyoGNTbFr4c1NdvAjZBBdBJxEKodMuQrkYeqGoNGcXeImvYfFxR2pweTUwpHHZkM
a6ChCP+CwFOOBQtgj9sVFspmcY8Ct/IEUGNQSn9ZMopl4A52iir9kL1Ezp1nk6r9GPaOlAQl3JLA
hoCwNMYWX6LS1XyDTV4nyfR1jiIOnkUKaYfRzJF4Un9CXsaV48NyVExEOqfeEfwe2d8BOhwmEhDi
dfVATBy3lWp1m7a/KT0A22z/f4B4CeZYQR/VNr6sKtmPJHMBiLYtPDZmc/Wo+zb7c10ZKkFIqY2g
7STxSfky5P2DDqjOdyAJbi8AbJjnZuJIHrqUZlb9Z+Yks3vh4Bvi/LoNXM8J38FWFtmVBrXJ3uJG
3At5iDzLXtc/vUzpttkg8kARb/GugyOx1HK/fAFBGHqcNPj0ILH33s7v5bGRBAJ805cPW8EgLtgU
lN7DSfpk8oGA4EAhz/3HN4ESbptg12NbPpzAmAslp3PV0GE7gDHIkPOZXOSLgNjtYJf70pBgeCcg
hV01YeihhRiI8Qds6mWTtoP5RUNycDq4yoUykVnccLWLejZCmDwJU13O7PGSYcz5UToHruVMgBIV
HPobhSOzXu14yFOtbzwkk+KfphuqAfIhpGbhPNLTNltpwe2li3xztJSQeWgmdS4NDPt7+pNBTIod
zL4dRb/33rN+TLBPJ9EAEEiAJGNIkZNOrER3TKwBn/JcuO/TtVrdeJzleVCjWkpGrUTg3XcsYUpY
IwgndaAySCvPiLkbpjoEidxjZt9isoM7rvRpEmrYT3LH8MpDe1JXXZSjX4X/q9mhsYgjsJN4G+HK
OvFRFC3pg9d+t1Lc9fhicAaXXnSvkpbeZT6usKv0cwQaNZ54IHDbOCRt+JJLM6o+Y/cOvx3g92/+
fgDYRKQrf5W3NktrMeJ3QEcDdG4JoVSTDjZPzusyObndlohGBX9FJ8i4Ag1K9iPw9dcTrPxT4Ddj
xOakkIcOCc4MBxd9fnU/DRIllL9kaQcZbjpSH9ndXoscB8GKW9BFPYNJql3pA3DRds14GbZdiZw3
Bvy6MafbmN3SZ7ahwp8Twy/nAFRiDC4I8Otm644smFJyC7VHzBO2hdATFw35bFvlWBy+nLJslLIu
klwxiGMq8470oH5nC/Vw45IRcE2M6DVmonuW0Tp3c819CklZdtHq+goDSoRt+xCxffeJZaxxaQls
qaTteO7yb20DH1T8gGGQnNXpO30f9nrj2ygzctLZdhaJdL7TctsCSnLxRVVYWspuRM3xs5a2NwNL
0tLAT1iEOskvhYCoIFgcWq7BQsquBMaKOYWvfsAYMG6C4iSg2osyv9uJN5Hc5LlRp2JxCqf1e0jF
YECZb0ESJNssGd6q6/UXLBpwcAyx8smct96pUgocag1plcDt90N+IkWnMoEAbx9IdNlTzA/jLeh4
bA60y9EcxMlGd0xbbpXsj9+FsynZGCJqabW3+QAXafx5mJ9zGUhcWpluZoA8k3S5kSVscn+UAy5u
ZntdEzWa+kAaQezgj/Q88jbonBBSl1HdQjz70CtyyH69dZpt8LeZuWOLDp9kUkbghC7bwfcdUM3r
wOhQBAxBzlfV/ZYqkV8qXsZk9psMNoRVfR8f8k8GqlVVHkudkeLg3sKpOKKh4LJWJKymTujuAEp1
dY4IgcwrW3kBIcw5A3Mk4GoTtDxNjd9mxLArzOTGBS+XU3NPt0RH4x9gk55tENZSEOm1AVmtqcz+
/vAm8sdh2d3+84GLeLu/s3hVM1wybFreQXRHNKX4j9AlotAvB8aaZ5lBBTLToCG5kH5/rFk3AI6t
gsAEEmLWMa2RrIAOijkQN7tZUvr62c6ZUYntHmKa8QrKlFuZ0nsjHnZscW19CUjGyjljmXSwT/E9
Y3rah9B0EZMHxmhyKNsF3Fm6uoUYb9Q4dL0svoqIJdG12uUNTTVNXiuPNAMOlwUq2iBJU8M7/mv/
Trdg80N0wHpLwaWw5sgF8S38KrttZ/B2L0q/iD3i+BV79Xf/1dX129jfN6YTjleViN2JY+iJrjRe
WqLPAmgYMZS5z/4Hmzl4i72+/m+lNnbonphIS43KguaUwNvFSWcpVS+fHa4VVgAO+oYt+0H6vnzw
TrHz4Ityq3PPXVblKex2GSjP0FrPlD3bETXlvumiWKQBN21ExyjOJrOvkMejefPa5TVLc3KurHLY
SpHfIuRAtZhuU1T5C4v0Xz2MVxX/cK3INTGQ0vaZiyMdURsOvA4PUJCRNBaohWb9Bt6+nonbHFYl
dh7bvfFHvDVXIwSl24tV3HueF/she1uTImm7+0G/R9ktbDpy0JHExWJZ99l9ktlNdfCmnymyYkiF
Zmyeq1Uri3NM0qioYn6oU1aGBFSAb/6pAHr9E06zIEk9WagMcTV4n4Lu95m3DQ3sz7Guj3f2ZmtY
6kt5WDipkq70Ef02G2Yag/Tk+gYhHGTVKLTHFLPzS6qg7a24Kqojn4RKCyzxTk5Z17B0xcKRy+O7
K5Dyz5kkvAQe3GNKRKTFNJGkfz5Bdg+T/9FrfL5OZs5fbl1ZWZmIu32HLm6sjZZsCrLauQxbdHMW
i6cBDQzsKJ7nUnP75dh0GHFpZOt5i8R/AK/4E7XN2X2QgzXpwPHUa/ewQW8pHeVoN2cft3REhmRP
2TKgSBCixmThvE9HlyVFXor8dcP2QqmMmKbq7UwAh4OgHJpwaPsBZL77YsKkzhUEPjhvSURzvXYP
YfHyFctXZ6CflJKaVOil9MLXywr5tXg4v20QmQ5Z3kAWhIZj5tqehNuU4G3u5tM9t+hzTYibRZZR
DBsW08Fhu0Smlw2M82GREiWOJR/DoUYmB5nXORTgTD7Xd4tSp5ZFiDDm3HNDW+zcPNQd6prPrdLd
5EzAeJajHOytlxITimqQshZOajaCiCWn2II493snvXvHHHWNEyNu034kLEjbcxLiHw/sQrsey2lK
ANNlbOzrNQeGCqB94J3riyDevKRfzx5VwYf0G7NgWZ6JsbmFRpI914YQI/cHEwa6ueZuU51BESYj
a0/ratO7wnONy8Qe2cZQWrJwAHIbP2zaB/fsGTXf0D4aC3qKHYafrmatDmntr8rIgXeUB5ifqdSY
AElVGibj3NUgvp8FA4hnqHK6LRSwtNAJSYe6kiEwHZYXvvifuaZ03gZW4cxo0sO16kEQXqc5kmog
Z5gGyAC5RaeLQVf/1JoeKcmGYUgDjyZF4sbUhCBE+XTYckLM7Y1agXYzvX+BGIeS8FUCZbTYDzR5
mKbmDLr2byjqFx6nOAhRmUlNkB9gC39FNN12Y7scxqWvydjKtsbF8k2dY2xAtcHuquJa3T5cKD0/
IftyZXQZFYYTx1kQp9Vk4HZiZRcuBMzazFsg6708XQDkFmpQ14Oqx8+A4AStmr18JdtMxbn4YEbC
epThat55HJoh0P2L6hGLxAN/hcELGz3uOU7OxfAUxnJISsArh0gfycfk2ZpzXO8QlZFJaeXhMD67
kacfdNRPA/LakvW+usyP6o2qojF0HgD9SmZW/E4gPerggehk3TsBGOlEvgANwyl7GAu7glhfCHlL
7GcnH3petnfGK/Z3LLPRXMXAVka+QafjnSIM7vbWWaVUgPWG37mgf1f2U7CHx7T4NlTH0IXz1hZS
+Jqi1I0ZzSt/L2uTJJBSRykMkP0vU3yyHe7xUe+taMM1U4xjRhaKHehgbroJHq8acNRovKxR7Gv7
GVy3Gaw3tYm9XUtfvbLHFklWa2sflcpAnEKdcTnd4AzIhD9RSFwfPym4Akm3i6sV46FVaNPTTT+M
Df/JCjxmtR1Lw6X5i0AB/NXWLqGpla3d+b/MRJ6J/0TGJGkYi5K4WOVw1SMW5BgPkXd1t7BSMzpC
yoDpVB1r8SEDgXOYd5wiYlVWl49wAcFzp5JqRBhFu30pQ2tLOC8s0TB8YAu4n9zWCa/1hAwe4U/v
y+6JkGET4fY+pEd+k/cf0FHAneWrFHBtFP4mgaiNND5YfwOGGmeu9sN9HNB8vV2foYQXOO1d3OuX
v3O8MZfK7ARnJX4vEurxkA/3hOsPOk9sNJ/oxXLMsesMIRJOTz3nILPHw2vCuVxAgpDjZjVzq8mw
zBwt04Z31LYYNkE0tt749YCrAqsVBQvyBjthi1TTzJUUwDv2m2kTFO0kTymf9iwVrpFjipyLKuto
1nRTCtlDUMtLbHxWpQInZpIwPxktt9vb9a5MIITiZeqAtEOa6MhUJJ3PySXjvH19XxRhnJ3nFNP2
pcLlKLONLMSlHHbaf6TkM8+uxmFZMUQEGtooHQszJ/+1FO/Dz+Ps1OlkUIX+/dpQnzid7my3UDhs
RoAC7O16cDB+5haXXqUXnlz7muqAbfxtl4msrhcaAMeA7H9j76ckEzRMic0XuWXvNoFmoqtSaCDz
yNCtjtS5c9GsU7yWr9FsBdrKyoTLP1tZ+pDs5Prg3IZSwtoeMd+QkrNG4hlCCmLVQBC6VROlicS8
AdPWrBKTwWTyPSZ1GZ13Q/9/14n7v0EpdTcityVqqURmq0gNcY1Bs9aAWYugGoDZPQcD5E01Dhks
m/oZXIhMUmNcsx+/2nRw6gYwwTa7twXt6ZPBmPETap4u8lsVX7VHMpDWRP1ZTLO/UWMVnK3fwUwA
/y2XC7Usxmz6S94EBBQ3NYo7AaH+hvP7ZB+nrC0ixExi2OeeOjN0TGrg9wvXPnv0ev5GgU2ViYSL
YysJ7iC05CNquYZMVgKTqHJyHlzeN+fxdU5x/zlpmWg+MAOXwdNR85Zwc1NnPTjmRontoMvAhwIr
Y6w41gDrPC8XePrmXypnR4bQtiVR0iGjP105y7cUoaVrn/LBGyhU/tebbhzotF5v4XA5C5V3zHXa
hFpuEbZCvpkKmbiUoEBooIGtZkE6yycXsZVHUeVB73sgNd8fI6CE5Ceaem870apg+RkR8Fni/MQv
gkB1FtQ/V+dXi8osADWO1zY15VFHuWyhsEskokNkQE+PoISV/TZBfPwEUiba90Q+k5w67jKrMAvT
BDIx0njE+Sf7sqfZj9jKMsoYbInp6OhGbT2NAJHt3+0GHJtacDgLqLDur7iDmX99hE2NcKAqwJ7X
pzeOJKRp54+U8pYOckKj7kyTU95tC6KlTT0diccA9VuYjOIuzz9PGHgXRWZTfsEnTSqT4WG0nPiN
muu/CeqcL0TVhWBYR8lIqfmIop0pG2INO8rTJqqs4G6dZ5eUSejnAgD8lqGuQMFYp+3hfGCFNdZQ
EANckznjUmTA8pPVK5j0JZvj7OS86OD34OmsXlQGGQ67FZn8Fari5QZ5BckNsksXVRgO5BHAxuI3
cenlIoDfAYDhMUiYt0/lgfcA+83kda4mxHsYR9Hw5qzZwaYsX8/UPE4+HOdxNIJjv3j7ckta8Aps
BrnAyN0kGGrk0HHO0YMAP2bZalEF28wtcxG8jpRX8o0ASiXWc7/s97e8KRGlhnEFLZzUMWj+M0YO
anJbcC6i+LFbQT7u2Pni0J52vMPU7oTjwLWhL7UlM4iK4I3GrQKLggFVo7nCOyhOesb2hw1zBwIv
eZPuUQuwi3y3L/Iy+ls3tdv82DgK+l4oMrJa0Jt+5UdWGQGwJuPITYiPxyxIJIV7I/NMld/ulaIA
C9mS/Q0AvjcacqUSry5ML7etL3dwsgRHSDdChi01b6zgSbi7OdIMKkQPhNt7p9U4v5HMc9wGDBxk
s5yXBbNsjJKxH5prLD2Z/vFp7F/mWdt4hGHOMGv0OvllAswxM967AcyVRUQf2NR+omvNSOM5k3Ws
bGhMsoNKTsbAmW26gBNfCFlQqyAIOrT1B1lbA22gIjwqhDgy3Cnh/uoJ57x9QkEH+FzTN51xkYoE
23PDTmr/gV1ZFZzqBHV6AkTpSY/XSpRHaPYIvgbkriUwyTGr9zFfNxgOtE9QciKIMEzvvgUJv19X
BdFh8N0TqzKp1Olo3R0NCuX7KKbKiOgNn1fVTWGEelj6npdeghm0nidhBDWMdKF14ou3PdXShj05
n7WnBuQDwUnMWK6qZrnd7WAN/8zvMGWnL3aIlArdSRxQyXMUw7dyIV5yAre5DbNJngWmz032vpsm
DCjLu8wXpLQonpiauEhbViilM3jAeLoHB9KdRxiLSEl1/1VvJKGKQAh+3f4NcrTN2HzLvlFKrB+Y
lVXdKEB+2qd7fz1KjMZqMoWk5dLMQyQwWjhMBydhxlvZDfyOaZrVmBXeJ/2TKNAMPJ6HcEzdBMh7
OCfCe7p/VfrLAXU=
`pragma protect end_protected


endmodule
