// =============================================================================
// Copyright 2016 Amazon.com, Inc. or its affiliates.
// All Rights Reserved Worldwide.
// Amazon Confidential information
// Restricted NDA Material
// =============================================================================
`define CL_NAME cl_simple
`define FPGA_LESS_RST
`define NO_XDMA

