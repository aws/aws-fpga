`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinx_2014_03", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
L/yhz0ZaRTYSpXjqwG9WZJBcOtq0XmLNTysRJQNVJOgGahEtCh7NqY/+u0QRj3WUWPxL1Ufw+Xw5
NqE0PHyDMWFotRkhe0af3hx/a34zIQ6g75B385s9iGUuYZYC6UQan9sYZwYXpwVkdVdI22CrhTAl
LvFUwyGerelX64yLQzFs/NJPYMpy5ITtBf+pCd+M5fWjiNywyUOWMT9z8MasSVfEuQyYPQGvug87
6UCVuh12SomKw68/lmzFenOgsqLpLO1fHoyUHLb/+KGHa1u5tdvG48b8rhDqXDCFZeDSagApvVdx
IieEy6yu8bHXe2eLIsJ8vGKNEiL44Ar3tKmDqA==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
IO0R5hnfUS844IJXrVorlwHRxUCTNuIyB8wzYVPcSVE9edF0LQMfJnHgHROF2kluEihoBDcwlY9t
mdw8Qh/4Z/UvrDywX8/ggcsrZdTSUKv1Jbuu4MlmoQfzWf8Dbc5vcHblk72bdleDjSA8ZWnSwwyl
mmWBtBmBWG9flsDfOkM=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
FygEYR40xD0CeRZXKFznTtGndvjNK8SxO44X11RQHwrkKIgg+8nm5febWYKzHLOtEYRf7UAnU3kv
mCdlEA3i2q+tO+IptJBZbpE9yy6mU9ou2sLRKe1BXgA4ycNxgL0fLAzrfeiyYaO6qb1Paxw8O31Y
MMqr9zt1mQSzRySht1Q=

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2624)
`pragma protect data_block
8T7qo6/JeJv1i6lNrYI9A3nuNoyit4DOCT0JpK5hXJKINE1qXGitcBWBzDa0igX9QOCejcaWSRey
s8zYCCyYUPuqhLpDQWxLr9cM56mkLX7qFtIPZM3YXuYniIyz3a7WnmcjI5JGhgAPM0Lb/E1XbPk8
CVUhwGPdGkDatt9QdbUE1JfcRnqKZ+GYF50qyCBT7fnZP+D19S1sZGRCTtFQ4gL75sYNUvPi3nsb
emjst1P0i791xWl/Ru/KvSV75uGBBIVemV7Dm3/DKU4ciKnSXzYGIXRp/+bjISr1fhc066xvinQZ
hTnUEU++ot45iwPGtVnUt1BcoNZYggyc+xiX9xTj2V3N1IrdkME0rCNGRiSQZmnhYngLPSvUVzGN
geYgVxTRx8MDcMMxErKo6pg2pUSzG3owrPF1/t2mWtnJogWwkIB1acy8tdIdOB7KX0ImdNhpwNEL
dzKw1okQw7lWPerW8/BY4izvx2dQ2i3R9GtXGIDG9MTZRcGaB8KbAss/dP1LO68V9z4ZjGzU9dLl
6qkgf+B/Cs1cqmmGjGpHG3ELhDLcSTf/E3T8F52XvGawiCo+7MhWqguFfVIHI6DSfh6joyyjrTJD
NXI+kTeR1H5K4GI4fnkMBKnXMMUyfiKC30+FtkGnBZI6PZV4BnCGkK6pXSj0+02cAiWlIrKUBphx
erkjhckMSuYV7RXzHiR38A0vW8xTRqk240X1i4KMcGpu9JanzEi1V4/01EvFYXzD9obs+3mUGXxJ
ZecX+QZu5Me/ee6hmG/xA1vqa5luTxjFiEsegXiLX4gON9MrgHk5mulXAN7qt+DpYvDQMaBdYkks
8aP1OGaO11wV4TMC72HIiFhOjxKPN4JtfTmF0u7hksKEGSmN0FdD6SDJsLKcWa1zKT8Nk39NvD+Y
29vg7jDsQV/OtQfCKM7+emIFpdUCAiOTXU3qR/qy8TnFa5HXyZvax9eVCEe3JuVnS/LaHJ56OWnh
DJh8UhCnGww0WRe4xZJvkSggct382DgbOqloHDk7ilYPCGOYZYXH7PzWCgrTFcOEWKoAionpmNcv
znzO+pFQtZ13Xz5PaXnEUq3w/OmqkOdo0XZmMT6CHDCNeq7ji1iG/zoL6STVBXaOff1DyERclbCh
6ujxgh7TJ8ou2LqhYmbHTPRs5ToQrovJVdwGdqeFOdFC+yfcurgQ2rLEB9EIjCZeXp5AxYxHj1JR
8AgOfPBsYBNQSIEi3QK47jeSFNs+h84glC9ve7MxQu+LA2Ja3WABiUO35JRw4ykDmoihIUBTU/LZ
9ZWjB+lgqWkMcs7KM0u3UEYw+P1byhQpmtfAay5jBZPjcSzgJPYzxhx4SANRuL//YO+GGHi8FasW
fpGIdMsAqPh8/XFfE/4at7IWAX4NLh/RT1mxqxL7gSXnGHcwFAB+cYK8WTD/IcBwIg94nLXKw7sY
2EFD0BiIrCoepJqDXrq7bJwtq+37/TlEKMC89neoOnYUQ9s5ZmdmDyexp/9UvxLY6psbCadSR3+X
azX+YGpXeaSt9tkqT0OzCO8+B3j8mFWYtty3pGyxMHf7sk0kfaKMAYAAZAn7/JIYdN0cfzlquKpe
vVRtbtuZmtSOUelKYnyfA1iL6gW3pBeI3YjwfYfUaP0yL5NA2vkhviDlOCJmyGJyedcQMvcd8QDb
JrNKBw7q3wVfC1cJs+79LDO3jISDBC8HiWx808C16CdQsSsHVuzROpU0BdND0PvOu9HcykXyblAJ
P2+1M1EvS1alGjNkuh+s+WUPulz7GycetUSV4ga5u2c64Rf6HYCUykC2C9G0abUMI7deHeFJq8Rb
xnbpgMVflIpIjxOerLQ1xacOnDmUw7gilMaj8vqWiIfYpV4vjNbFtJ5nvoEzcdF3rxIj5l8m6unS
Uz+Ud2UmT6nvTi5kjRnYbrzOPgbZws2W2mwgs9LsyF13Y8dooB0IXaTJ6vjHSXSTdsIIAc0NnIf5
dpHJWSUqcGaUY6l2xr+1KQ8zkeXToGcp0Pz1Gdc5re9XAwEmznJRY9cxiDV2YsWs+otK0dpNPdk1
pS69HZv8qWdTo6c6ojKeEU6o3eY55wt3OoH2AMKMb/kHXTsecrOvLd2Rv6f/PVjNy2yV1GyYaEGF
u1LnRX/PP+BUbyYsswx8RXGGOTfdd0fpIEO54H3gbpgb8xJqncahF9RSXzTvk55bl8d4zYZZLJoO
DinznL0CKdy+hN1JpH1LXCjJ3AucciXFPru0+CI3VmhGOjnaaQdcARQoh3jhjpjaWetuTAPWUUdk
P/iAlvxnhettjBV7hk4Rfx1tMjaQXzAWsF2Wv5pFteGvsaSd6ZSyA5fvbNpIR6Uo/o/MAnMH51Ar
EygKwDHjZwqLyyoqpT9YXmIEiBwN1r9KE6MZAhbC+ObPUAIcPgUrNP06uBvyEsNu+S3Sq7/55Ahb
xi+cywAxa0SVlS4Ra5382jbgwrfew0pnFNniuZkxY+a3tE8UWi3huO/QkzHr3cwCyYkZvGaElijy
q15S2qJxudnzLPJiSLT77IPC8UqE8UVnEIGEsPm77DA6SrWPaEFPMKe5PgGar01VIaARhKXci+y0
/RKybOmIM7abyWtmqXlmysZPBQtDaJQaK+rEQACXwCiuQIGJZ8KSdjFWk8+feX4zdvGBdFKwh9Ua
mnQ/Ss3dRKcqPk5bAxHvZGdywckq9NX3guHGH3FXYSQ1hIEKUJuwSkS8PTNQlcVXyV9roFmCvApc
FJ1kWSRxqnROl7nWZiPXM1VJ4+YDaI9M8H1nQvMyFAxi87tJ9yj8rPb/AfUia4QkcqaU0OJfjXE7
0xHkxlP/78uX1IT46GTk9RSeuLeFseuNxdD30IDmZSsF4DYPBwuK0sUwUVs5oO6irbBT1rGKPZDR
gTlQmfOn2w4vu7x5FlQwCeCY0qc0ob0W19i+42dXpTU0hOWZma1m1vxsBzH2wE5F0XF3KD1Ve+OV
GgB505cAv0RihmilRx9cr9s4MAn5o8GsHnXR/JMc9FNSJlJGm3okwHbRZS1afAIrggnq8Z+gKiy5
Q+zdVDQFfQuEl8rVeDVr2iwQKQ1Zu36l7fnFMZ2AhnJ5obQ/kj29Ekn949QjBP5jQ5JNw+LYi6XD
1t4taW9T66WeBPWXAL2OdjlAmnfynWZVdCIoVmR3VYOQq4XcPpwwslehqgEg9JgCtbkKZrVhKyKN
WcLRnQizxIdXOWLXJlMrJD5pECk83n669bQIMl+g5KokNeAw3npj9rb35sNyg0+If5Zl0tEv2pNl
3Qa3pThXnLHzT0yml4DqKf5U3Cnxg2qwVsezB+XW7zbt/F/JHaaJtsSdeq3BlFelkTnVN2kLA7h2
X2Y3vjnUd6Jrtfic3wGHHikWsn3DIJnQzLuqDSvxppMWcjSNFa9f/ZGDu6flel5gSQRnzYOKptbx
M6rFzTHGEkr6mCvetdhC0lS0A6oZmyw/jUyFC4/HjXr+FvLzotw4AGVJ24aaeVGerOGJ7zhjfvTj
B2g=
`pragma protect end_protected
